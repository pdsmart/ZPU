-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use pkgs.config_pkg.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8a",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"88",
           281 => x"00",
           282 => x"70",
           283 => x"8b",
           284 => x"70",
           285 => x"0c",
           286 => x"88",
           287 => x"99",
           288 => x"02",
           289 => x"3d",
           290 => x"94",
           291 => x"08",
           292 => x"88",
           293 => x"82",
           294 => x"08",
           295 => x"54",
           296 => x"94",
           297 => x"08",
           298 => x"fd",
           299 => x"53",
           300 => x"05",
           301 => x"08",
           302 => x"51",
           303 => x"88",
           304 => x"0c",
           305 => x"0d",
           306 => x"94",
           307 => x"0c",
           308 => x"80",
           309 => x"fc",
           310 => x"08",
           311 => x"80",
           312 => x"94",
           313 => x"08",
           314 => x"88",
           315 => x"0b",
           316 => x"05",
           317 => x"fc",
           318 => x"38",
           319 => x"08",
           320 => x"94",
           321 => x"08",
           322 => x"05",
           323 => x"8c",
           324 => x"25",
           325 => x"08",
           326 => x"30",
           327 => x"05",
           328 => x"94",
           329 => x"0c",
           330 => x"05",
           331 => x"81",
           332 => x"f0",
           333 => x"08",
           334 => x"94",
           335 => x"0c",
           336 => x"08",
           337 => x"52",
           338 => x"05",
           339 => x"a7",
           340 => x"70",
           341 => x"05",
           342 => x"08",
           343 => x"80",
           344 => x"94",
           345 => x"08",
           346 => x"f8",
           347 => x"08",
           348 => x"70",
           349 => x"89",
           350 => x"0c",
           351 => x"02",
           352 => x"3d",
           353 => x"94",
           354 => x"0c",
           355 => x"05",
           356 => x"93",
           357 => x"88",
           358 => x"94",
           359 => x"0c",
           360 => x"08",
           361 => x"94",
           362 => x"08",
           363 => x"38",
           364 => x"05",
           365 => x"08",
           366 => x"81",
           367 => x"8c",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"08",
           372 => x"54",
           373 => x"05",
           374 => x"8c",
           375 => x"f8",
           376 => x"94",
           377 => x"0c",
           378 => x"05",
           379 => x"0c",
           380 => x"0d",
           381 => x"94",
           382 => x"0c",
           383 => x"81",
           384 => x"fc",
           385 => x"0b",
           386 => x"05",
           387 => x"8c",
           388 => x"08",
           389 => x"27",
           390 => x"08",
           391 => x"80",
           392 => x"80",
           393 => x"8c",
           394 => x"99",
           395 => x"8c",
           396 => x"94",
           397 => x"0c",
           398 => x"05",
           399 => x"08",
           400 => x"c9",
           401 => x"fc",
           402 => x"2e",
           403 => x"94",
           404 => x"08",
           405 => x"05",
           406 => x"38",
           407 => x"05",
           408 => x"8c",
           409 => x"94",
           410 => x"0c",
           411 => x"05",
           412 => x"fc",
           413 => x"94",
           414 => x"0c",
           415 => x"05",
           416 => x"94",
           417 => x"0c",
           418 => x"05",
           419 => x"94",
           420 => x"0c",
           421 => x"94",
           422 => x"08",
           423 => x"38",
           424 => x"05",
           425 => x"08",
           426 => x"51",
           427 => x"08",
           428 => x"70",
           429 => x"05",
           430 => x"08",
           431 => x"88",
           432 => x"0d",
           433 => x"ff",
           434 => x"88",
           435 => x"92",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"8c",
           441 => x"06",
           442 => x"80",
           443 => x"87",
           444 => x"08",
           445 => x"38",
           446 => x"8c",
           447 => x"80",
           448 => x"93",
           449 => x"98",
           450 => x"70",
           451 => x"38",
           452 => x"0b",
           453 => x"0b",
           454 => x"a8",
           455 => x"83",
           456 => x"fa",
           457 => x"7b",
           458 => x"56",
           459 => x"0b",
           460 => x"33",
           461 => x"55",
           462 => x"75",
           463 => x"06",
           464 => x"85",
           465 => x"98",
           466 => x"87",
           467 => x"0c",
           468 => x"c0",
           469 => x"87",
           470 => x"08",
           471 => x"70",
           472 => x"52",
           473 => x"2e",
           474 => x"c0",
           475 => x"70",
           476 => x"76",
           477 => x"53",
           478 => x"2e",
           479 => x"80",
           480 => x"71",
           481 => x"05",
           482 => x"14",
           483 => x"55",
           484 => x"51",
           485 => x"8b",
           486 => x"98",
           487 => x"70",
           488 => x"87",
           489 => x"08",
           490 => x"38",
           491 => x"c0",
           492 => x"87",
           493 => x"08",
           494 => x"51",
           495 => x"38",
           496 => x"80",
           497 => x"52",
           498 => x"09",
           499 => x"38",
           500 => x"8c",
           501 => x"72",
           502 => x"06",
           503 => x"52",
           504 => x"88",
           505 => x"fe",
           506 => x"81",
           507 => x"33",
           508 => x"07",
           509 => x"51",
           510 => x"04",
           511 => x"75",
           512 => x"82",
           513 => x"90",
           514 => x"2b",
           515 => x"33",
           516 => x"88",
           517 => x"71",
           518 => x"52",
           519 => x"54",
           520 => x"0d",
           521 => x"0d",
           522 => x"0b",
           523 => x"57",
           524 => x"27",
           525 => x"76",
           526 => x"27",
           527 => x"75",
           528 => x"82",
           529 => x"74",
           530 => x"38",
           531 => x"74",
           532 => x"83",
           533 => x"76",
           534 => x"17",
           535 => x"88",
           536 => x"55",
           537 => x"88",
           538 => x"74",
           539 => x"3f",
           540 => x"ff",
           541 => x"ad",
           542 => x"76",
           543 => x"fc",
           544 => x"87",
           545 => x"08",
           546 => x"3d",
           547 => x"fd",
           548 => x"08",
           549 => x"51",
           550 => x"88",
           551 => x"06",
           552 => x"81",
           553 => x"0c",
           554 => x"04",
           555 => x"0b",
           556 => x"ac",
           557 => x"88",
           558 => x"05",
           559 => x"80",
           560 => x"27",
           561 => x"14",
           562 => x"29",
           563 => x"05",
           564 => x"88",
           565 => x"0d",
           566 => x"0d",
           567 => x"0b",
           568 => x"9f",
           569 => x"33",
           570 => x"71",
           571 => x"81",
           572 => x"94",
           573 => x"ef",
           574 => x"90",
           575 => x"14",
           576 => x"3f",
           577 => x"ff",
           578 => x"07",
           579 => x"3d",
           580 => x"3d",
           581 => x"0b",
           582 => x"08",
           583 => x"75",
           584 => x"08",
           585 => x"2e",
           586 => x"14",
           587 => x"85",
           588 => x"b0",
           589 => x"38",
           590 => x"71",
           591 => x"81",
           592 => x"90",
           593 => x"72",
           594 => x"72",
           595 => x"38",
           596 => x"d8",
           597 => x"52",
           598 => x"14",
           599 => x"90",
           600 => x"52",
           601 => x"86",
           602 => x"fa",
           603 => x"0b",
           604 => x"ac",
           605 => x"81",
           606 => x"ff",
           607 => x"54",
           608 => x"80",
           609 => x"90",
           610 => x"72",
           611 => x"52",
           612 => x"73",
           613 => x"71",
           614 => x"81",
           615 => x"0c",
           616 => x"53",
           617 => x"83",
           618 => x"22",
           619 => x"76",
           620 => x"b5",
           621 => x"33",
           622 => x"84",
           623 => x"71",
           624 => x"51",
           625 => x"81",
           626 => x"08",
           627 => x"83",
           628 => x"88",
           629 => x"96",
           630 => x"8c",
           631 => x"08",
           632 => x"3f",
           633 => x"16",
           634 => x"23",
           635 => x"88",
           636 => x"0d",
           637 => x"0d",
           638 => x"58",
           639 => x"33",
           640 => x"2e",
           641 => x"88",
           642 => x"70",
           643 => x"39",
           644 => x"56",
           645 => x"2e",
           646 => x"84",
           647 => x"43",
           648 => x"1d",
           649 => x"33",
           650 => x"9f",
           651 => x"7b",
           652 => x"3f",
           653 => x"80",
           654 => x"d3",
           655 => x"84",
           656 => x"58",
           657 => x"55",
           658 => x"81",
           659 => x"ff",
           660 => x"ff",
           661 => x"06",
           662 => x"70",
           663 => x"7f",
           664 => x"7a",
           665 => x"81",
           666 => x"13",
           667 => x"af",
           668 => x"a0",
           669 => x"80",
           670 => x"51",
           671 => x"5d",
           672 => x"80",
           673 => x"ae",
           674 => x"06",
           675 => x"55",
           676 => x"75",
           677 => x"80",
           678 => x"79",
           679 => x"30",
           680 => x"70",
           681 => x"07",
           682 => x"51",
           683 => x"75",
           684 => x"58",
           685 => x"ab",
           686 => x"19",
           687 => x"06",
           688 => x"5a",
           689 => x"75",
           690 => x"39",
           691 => x"0c",
           692 => x"a0",
           693 => x"81",
           694 => x"1a",
           695 => x"fc",
           696 => x"08",
           697 => x"a0",
           698 => x"70",
           699 => x"e0",
           700 => x"90",
           701 => x"7c",
           702 => x"3f",
           703 => x"88",
           704 => x"38",
           705 => x"74",
           706 => x"ee",
           707 => x"33",
           708 => x"70",
           709 => x"56",
           710 => x"38",
           711 => x"1e",
           712 => x"59",
           713 => x"ff",
           714 => x"ff",
           715 => x"79",
           716 => x"5b",
           717 => x"81",
           718 => x"71",
           719 => x"56",
           720 => x"2e",
           721 => x"39",
           722 => x"92",
           723 => x"fc",
           724 => x"8e",
           725 => x"56",
           726 => x"38",
           727 => x"56",
           728 => x"8b",
           729 => x"55",
           730 => x"8b",
           731 => x"84",
           732 => x"06",
           733 => x"74",
           734 => x"56",
           735 => x"56",
           736 => x"51",
           737 => x"88",
           738 => x"0c",
           739 => x"75",
           740 => x"3d",
           741 => x"3d",
           742 => x"59",
           743 => x"83",
           744 => x"52",
           745 => x"fb",
           746 => x"88",
           747 => x"38",
           748 => x"b3",
           749 => x"83",
           750 => x"55",
           751 => x"82",
           752 => x"09",
           753 => x"ce",
           754 => x"b6",
           755 => x"76",
           756 => x"3f",
           757 => x"88",
           758 => x"76",
           759 => x"3f",
           760 => x"ff",
           761 => x"74",
           762 => x"2e",
           763 => x"54",
           764 => x"77",
           765 => x"f6",
           766 => x"08",
           767 => x"94",
           768 => x"f7",
           769 => x"08",
           770 => x"06",
           771 => x"82",
           772 => x"38",
           773 => x"88",
           774 => x"0d",
           775 => x"0d",
           776 => x"0b",
           777 => x"9f",
           778 => x"9b",
           779 => x"81",
           780 => x"56",
           781 => x"38",
           782 => x"8d",
           783 => x"57",
           784 => x"3f",
           785 => x"ff",
           786 => x"81",
           787 => x"06",
           788 => x"54",
           789 => x"74",
           790 => x"f5",
           791 => x"08",
           792 => x"3d",
           793 => x"80",
           794 => x"95",
           795 => x"51",
           796 => x"88",
           797 => x"53",
           798 => x"fe",
           799 => x"08",
           800 => x"57",
           801 => x"09",
           802 => x"38",
           803 => x"99",
           804 => x"2e",
           805 => x"56",
           806 => x"a4",
           807 => x"79",
           808 => x"f4",
           809 => x"56",
           810 => x"fd",
           811 => x"e5",
           812 => x"b3",
           813 => x"83",
           814 => x"58",
           815 => x"95",
           816 => x"51",
           817 => x"88",
           818 => x"af",
           819 => x"71",
           820 => x"05",
           821 => x"54",
           822 => x"f6",
           823 => x"08",
           824 => x"06",
           825 => x"1a",
           826 => x"33",
           827 => x"95",
           828 => x"51",
           829 => x"88",
           830 => x"23",
           831 => x"05",
           832 => x"3f",
           833 => x"ff",
           834 => x"75",
           835 => x"3d",
           836 => x"f5",
           837 => x"08",
           838 => x"f5",
           839 => x"08",
           840 => x"06",
           841 => x"79",
           842 => x"22",
           843 => x"82",
           844 => x"72",
           845 => x"59",
           846 => x"ee",
           847 => x"08",
           848 => x"88",
           849 => x"08",
           850 => x"56",
           851 => x"df",
           852 => x"38",
           853 => x"ff",
           854 => x"85",
           855 => x"89",
           856 => x"76",
           857 => x"c1",
           858 => x"34",
           859 => x"09",
           860 => x"38",
           861 => x"05",
           862 => x"3f",
           863 => x"1a",
           864 => x"8c",
           865 => x"90",
           866 => x"83",
           867 => x"8c",
           868 => x"71",
           869 => x"94",
           870 => x"80",
           871 => x"34",
           872 => x"0b",
           873 => x"80",
           874 => x"0c",
           875 => x"04",
           876 => x"0b",
           877 => x"ac",
           878 => x"54",
           879 => x"80",
           880 => x"0b",
           881 => x"98",
           882 => x"45",
           883 => x"3d",
           884 => x"ec",
           885 => x"9d",
           886 => x"54",
           887 => x"c0",
           888 => x"33",
           889 => x"2e",
           890 => x"a7",
           891 => x"84",
           892 => x"06",
           893 => x"73",
           894 => x"38",
           895 => x"39",
           896 => x"d5",
           897 => x"a0",
           898 => x"3d",
           899 => x"f3",
           900 => x"08",
           901 => x"73",
           902 => x"81",
           903 => x"34",
           904 => x"98",
           905 => x"f6",
           906 => x"7f",
           907 => x"0b",
           908 => x"59",
           909 => x"80",
           910 => x"57",
           911 => x"81",
           912 => x"16",
           913 => x"55",
           914 => x"80",
           915 => x"38",
           916 => x"81",
           917 => x"39",
           918 => x"17",
           919 => x"81",
           920 => x"16",
           921 => x"08",
           922 => x"78",
           923 => x"74",
           924 => x"2e",
           925 => x"98",
           926 => x"83",
           927 => x"57",
           928 => x"38",
           929 => x"ff",
           930 => x"2a",
           931 => x"ff",
           932 => x"79",
           933 => x"87",
           934 => x"08",
           935 => x"a4",
           936 => x"f3",
           937 => x"08",
           938 => x"27",
           939 => x"74",
           940 => x"a4",
           941 => x"f3",
           942 => x"08",
           943 => x"80",
           944 => x"38",
           945 => x"a8",
           946 => x"16",
           947 => x"06",
           948 => x"31",
           949 => x"75",
           950 => x"77",
           951 => x"98",
           952 => x"ff",
           953 => x"16",
           954 => x"51",
           955 => x"88",
           956 => x"38",
           957 => x"15",
           958 => x"77",
           959 => x"08",
           960 => x"58",
           961 => x"fe",
           962 => x"19",
           963 => x"39",
           964 => x"88",
           965 => x"0d",
           966 => x"0d",
           967 => x"e4",
           968 => x"94",
           969 => x"90",
           970 => x"87",
           971 => x"0c",
           972 => x"0b",
           973 => x"84",
           974 => x"83",
           975 => x"94",
           976 => x"b0",
           977 => x"3f",
           978 => x"38",
           979 => x"fc",
           980 => x"08",
           981 => x"80",
           982 => x"87",
           983 => x"0c",
           984 => x"fc",
           985 => x"80",
           986 => x"fd",
           987 => x"08",
           988 => x"54",
           989 => x"86",
           990 => x"55",
           991 => x"80",
           992 => x"80",
           993 => x"00",
           994 => x"ff",
           995 => x"ff",
           996 => x"ff",
           997 => x"00",
           998 => x"54",
           999 => x"59",
          1000 => x"4d",
          1001 => x"00",
          1002 => x"00",
          2048 => x"c4",
          2049 => x"0b",
          2050 => x"04",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"c4",
          2057 => x"0b",
          2058 => x"04",
          2059 => x"c4",
          2060 => x"0b",
          2061 => x"04",
          2062 => x"c4",
          2063 => x"0b",
          2064 => x"04",
          2065 => x"c4",
          2066 => x"0b",
          2067 => x"04",
          2068 => x"c4",
          2069 => x"0b",
          2070 => x"04",
          2071 => x"c5",
          2072 => x"0b",
          2073 => x"04",
          2074 => x"c5",
          2075 => x"0b",
          2076 => x"04",
          2077 => x"c5",
          2078 => x"0b",
          2079 => x"04",
          2080 => x"c5",
          2081 => x"0b",
          2082 => x"04",
          2083 => x"c6",
          2084 => x"0b",
          2085 => x"04",
          2086 => x"c6",
          2087 => x"0b",
          2088 => x"04",
          2089 => x"c6",
          2090 => x"0b",
          2091 => x"04",
          2092 => x"c6",
          2093 => x"0b",
          2094 => x"04",
          2095 => x"c7",
          2096 => x"0b",
          2097 => x"04",
          2098 => x"c7",
          2099 => x"0b",
          2100 => x"04",
          2101 => x"c7",
          2102 => x"0b",
          2103 => x"04",
          2104 => x"c7",
          2105 => x"0b",
          2106 => x"04",
          2107 => x"c8",
          2108 => x"0b",
          2109 => x"04",
          2110 => x"c8",
          2111 => x"0b",
          2112 => x"04",
          2113 => x"c8",
          2114 => x"0b",
          2115 => x"04",
          2116 => x"c8",
          2117 => x"0b",
          2118 => x"04",
          2119 => x"c9",
          2120 => x"0b",
          2121 => x"04",
          2122 => x"c9",
          2123 => x"0b",
          2124 => x"04",
          2125 => x"c9",
          2126 => x"0b",
          2127 => x"04",
          2128 => x"c9",
          2129 => x"0b",
          2130 => x"04",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"d4",
          2178 => x"80",
          2179 => x"d4",
          2180 => x"90",
          2181 => x"d4",
          2182 => x"c0",
          2183 => x"d4",
          2184 => x"90",
          2185 => x"d4",
          2186 => x"85",
          2187 => x"d4",
          2188 => x"90",
          2189 => x"d4",
          2190 => x"a3",
          2191 => x"d4",
          2192 => x"90",
          2193 => x"d4",
          2194 => x"f7",
          2195 => x"d4",
          2196 => x"90",
          2197 => x"d4",
          2198 => x"8b",
          2199 => x"d4",
          2200 => x"90",
          2201 => x"d4",
          2202 => x"c4",
          2203 => x"d4",
          2204 => x"90",
          2205 => x"d4",
          2206 => x"a8",
          2207 => x"d4",
          2208 => x"90",
          2209 => x"d4",
          2210 => x"be",
          2211 => x"d4",
          2212 => x"90",
          2213 => x"d4",
          2214 => x"9d",
          2215 => x"d4",
          2216 => x"90",
          2217 => x"d4",
          2218 => x"b3",
          2219 => x"d4",
          2220 => x"90",
          2221 => x"d4",
          2222 => x"d7",
          2223 => x"d4",
          2224 => x"90",
          2225 => x"d4",
          2226 => x"80",
          2227 => x"d4",
          2228 => x"90",
          2229 => x"d4",
          2230 => x"ce",
          2231 => x"d4",
          2232 => x"90",
          2233 => x"d4",
          2234 => x"d8",
          2235 => x"d4",
          2236 => x"90",
          2237 => x"d4",
          2238 => x"90",
          2239 => x"d4",
          2240 => x"90",
          2241 => x"d4",
          2242 => x"ea",
          2243 => x"d4",
          2244 => x"90",
          2245 => x"d4",
          2246 => x"f2",
          2247 => x"d4",
          2248 => x"90",
          2249 => x"d4",
          2250 => x"e9",
          2251 => x"d4",
          2252 => x"90",
          2253 => x"d4",
          2254 => x"f8",
          2255 => x"d4",
          2256 => x"90",
          2257 => x"d4",
          2258 => x"df",
          2259 => x"d4",
          2260 => x"90",
          2261 => x"d4",
          2262 => x"92",
          2263 => x"d4",
          2264 => x"90",
          2265 => x"d4",
          2266 => x"86",
          2267 => x"d4",
          2268 => x"90",
          2269 => x"d4",
          2270 => x"9a",
          2271 => x"d4",
          2272 => x"90",
          2273 => x"d4",
          2274 => x"bd",
          2275 => x"d4",
          2276 => x"90",
          2277 => x"d4",
          2278 => x"e1",
          2279 => x"d4",
          2280 => x"90",
          2281 => x"d4",
          2282 => x"8a",
          2283 => x"d4",
          2284 => x"90",
          2285 => x"d4",
          2286 => x"9a",
          2287 => x"d4",
          2288 => x"90",
          2289 => x"d4",
          2290 => x"92",
          2291 => x"d4",
          2292 => x"90",
          2293 => x"d4",
          2294 => x"f3",
          2295 => x"d4",
          2296 => x"90",
          2297 => x"d4",
          2298 => x"80",
          2299 => x"d4",
          2300 => x"90",
          2301 => x"d4",
          2302 => x"f7",
          2303 => x"d4",
          2304 => x"90",
          2305 => x"d4",
          2306 => x"fd",
          2307 => x"d4",
          2308 => x"90",
          2309 => x"d4",
          2310 => x"c9",
          2311 => x"d4",
          2312 => x"90",
          2313 => x"d4",
          2314 => x"a2",
          2315 => x"d4",
          2316 => x"90",
          2317 => x"d4",
          2318 => x"cc",
          2319 => x"d4",
          2320 => x"90",
          2321 => x"d4",
          2322 => x"da",
          2323 => x"d4",
          2324 => x"90",
          2325 => x"d4",
          2326 => x"f6",
          2327 => x"d4",
          2328 => x"90",
          2329 => x"d4",
          2330 => x"81",
          2331 => x"d4",
          2332 => x"90",
          2333 => x"d4",
          2334 => x"ee",
          2335 => x"d4",
          2336 => x"90",
          2337 => x"d4",
          2338 => x"83",
          2339 => x"d4",
          2340 => x"90",
          2341 => x"d4",
          2342 => x"df",
          2343 => x"d4",
          2344 => x"90",
          2345 => x"d4",
          2346 => x"fe",
          2347 => x"d4",
          2348 => x"90",
          2349 => x"d4",
          2350 => x"d7",
          2351 => x"d4",
          2352 => x"90",
          2353 => x"d4",
          2354 => x"b1",
          2355 => x"d4",
          2356 => x"90",
          2357 => x"d4",
          2358 => x"81",
          2359 => x"d4",
          2360 => x"90",
          2361 => x"d4",
          2362 => x"e6",
          2363 => x"d4",
          2364 => x"90",
          2365 => x"d4",
          2366 => x"f3",
          2367 => x"d4",
          2368 => x"90",
          2369 => x"d4",
          2370 => x"dd",
          2371 => x"d4",
          2372 => x"90",
          2373 => x"c8",
          2374 => x"cc",
          2375 => x"80",
          2376 => x"05",
          2377 => x"0b",
          2378 => x"04",
          2379 => x"51",
          2380 => x"04",
          2381 => x"93",
          2382 => x"82",
          2383 => x"fd",
          2384 => x"53",
          2385 => x"08",
          2386 => x"52",
          2387 => x"08",
          2388 => x"51",
          2389 => x"82",
          2390 => x"70",
          2391 => x"0c",
          2392 => x"0d",
          2393 => x"0c",
          2394 => x"d4",
          2395 => x"93",
          2396 => x"3d",
          2397 => x"82",
          2398 => x"8c",
          2399 => x"82",
          2400 => x"88",
          2401 => x"93",
          2402 => x"c8",
          2403 => x"93",
          2404 => x"85",
          2405 => x"93",
          2406 => x"82",
          2407 => x"02",
          2408 => x"0c",
          2409 => x"81",
          2410 => x"d4",
          2411 => x"0c",
          2412 => x"93",
          2413 => x"05",
          2414 => x"d4",
          2415 => x"08",
          2416 => x"08",
          2417 => x"27",
          2418 => x"93",
          2419 => x"05",
          2420 => x"ae",
          2421 => x"82",
          2422 => x"8c",
          2423 => x"a2",
          2424 => x"d4",
          2425 => x"08",
          2426 => x"d4",
          2427 => x"0c",
          2428 => x"08",
          2429 => x"10",
          2430 => x"08",
          2431 => x"ff",
          2432 => x"93",
          2433 => x"05",
          2434 => x"80",
          2435 => x"93",
          2436 => x"05",
          2437 => x"d4",
          2438 => x"08",
          2439 => x"82",
          2440 => x"88",
          2441 => x"93",
          2442 => x"05",
          2443 => x"93",
          2444 => x"05",
          2445 => x"d4",
          2446 => x"08",
          2447 => x"08",
          2448 => x"07",
          2449 => x"08",
          2450 => x"82",
          2451 => x"fc",
          2452 => x"2a",
          2453 => x"08",
          2454 => x"82",
          2455 => x"8c",
          2456 => x"2a",
          2457 => x"08",
          2458 => x"ff",
          2459 => x"93",
          2460 => x"05",
          2461 => x"93",
          2462 => x"d4",
          2463 => x"08",
          2464 => x"d4",
          2465 => x"0c",
          2466 => x"82",
          2467 => x"f8",
          2468 => x"82",
          2469 => x"f4",
          2470 => x"82",
          2471 => x"f4",
          2472 => x"93",
          2473 => x"3d",
          2474 => x"d4",
          2475 => x"3d",
          2476 => x"71",
          2477 => x"9f",
          2478 => x"55",
          2479 => x"72",
          2480 => x"74",
          2481 => x"70",
          2482 => x"38",
          2483 => x"71",
          2484 => x"38",
          2485 => x"81",
          2486 => x"ff",
          2487 => x"ff",
          2488 => x"06",
          2489 => x"82",
          2490 => x"86",
          2491 => x"74",
          2492 => x"75",
          2493 => x"90",
          2494 => x"54",
          2495 => x"27",
          2496 => x"71",
          2497 => x"53",
          2498 => x"70",
          2499 => x"0c",
          2500 => x"84",
          2501 => x"72",
          2502 => x"05",
          2503 => x"12",
          2504 => x"26",
          2505 => x"72",
          2506 => x"72",
          2507 => x"05",
          2508 => x"12",
          2509 => x"26",
          2510 => x"53",
          2511 => x"fb",
          2512 => x"79",
          2513 => x"83",
          2514 => x"52",
          2515 => x"71",
          2516 => x"54",
          2517 => x"73",
          2518 => x"c6",
          2519 => x"54",
          2520 => x"70",
          2521 => x"52",
          2522 => x"2e",
          2523 => x"33",
          2524 => x"2e",
          2525 => x"95",
          2526 => x"81",
          2527 => x"70",
          2528 => x"54",
          2529 => x"70",
          2530 => x"33",
          2531 => x"ff",
          2532 => x"ff",
          2533 => x"31",
          2534 => x"0c",
          2535 => x"3d",
          2536 => x"09",
          2537 => x"fd",
          2538 => x"70",
          2539 => x"81",
          2540 => x"51",
          2541 => x"38",
          2542 => x"16",
          2543 => x"56",
          2544 => x"08",
          2545 => x"73",
          2546 => x"ff",
          2547 => x"0b",
          2548 => x"0c",
          2549 => x"04",
          2550 => x"80",
          2551 => x"71",
          2552 => x"87",
          2553 => x"93",
          2554 => x"ff",
          2555 => x"81",
          2556 => x"83",
          2557 => x"38",
          2558 => x"c8",
          2559 => x"0d",
          2560 => x"0d",
          2561 => x"70",
          2562 => x"73",
          2563 => x"cd",
          2564 => x"51",
          2565 => x"09",
          2566 => x"38",
          2567 => x"33",
          2568 => x"a0",
          2569 => x"73",
          2570 => x"81",
          2571 => x"72",
          2572 => x"70",
          2573 => x"38",
          2574 => x"30",
          2575 => x"74",
          2576 => x"70",
          2577 => x"33",
          2578 => x"2e",
          2579 => x"88",
          2580 => x"70",
          2581 => x"34",
          2582 => x"73",
          2583 => x"93",
          2584 => x"3d",
          2585 => x"3d",
          2586 => x"72",
          2587 => x"91",
          2588 => x"fc",
          2589 => x"51",
          2590 => x"82",
          2591 => x"85",
          2592 => x"83",
          2593 => x"72",
          2594 => x"0c",
          2595 => x"04",
          2596 => x"7d",
          2597 => x"ff",
          2598 => x"81",
          2599 => x"26",
          2600 => x"83",
          2601 => x"05",
          2602 => x"79",
          2603 => x"b1",
          2604 => x"33",
          2605 => x"79",
          2606 => x"a5",
          2607 => x"33",
          2608 => x"79",
          2609 => x"99",
          2610 => x"33",
          2611 => x"79",
          2612 => x"8d",
          2613 => x"22",
          2614 => x"79",
          2615 => x"81",
          2616 => x"1c",
          2617 => x"5b",
          2618 => x"26",
          2619 => x"8a",
          2620 => x"88",
          2621 => x"86",
          2622 => x"85",
          2623 => x"84",
          2624 => x"83",
          2625 => x"82",
          2626 => x"7b",
          2627 => x"f6",
          2628 => x"89",
          2629 => x"98",
          2630 => x"7b",
          2631 => x"87",
          2632 => x"0c",
          2633 => x"87",
          2634 => x"0c",
          2635 => x"87",
          2636 => x"0c",
          2637 => x"87",
          2638 => x"0c",
          2639 => x"87",
          2640 => x"0c",
          2641 => x"87",
          2642 => x"0c",
          2643 => x"87",
          2644 => x"0c",
          2645 => x"87",
          2646 => x"0c",
          2647 => x"80",
          2648 => x"93",
          2649 => x"3d",
          2650 => x"3d",
          2651 => x"87",
          2652 => x"5c",
          2653 => x"87",
          2654 => x"08",
          2655 => x"23",
          2656 => x"b8",
          2657 => x"82",
          2658 => x"c0",
          2659 => x"5b",
          2660 => x"34",
          2661 => x"b0",
          2662 => x"84",
          2663 => x"c0",
          2664 => x"5b",
          2665 => x"34",
          2666 => x"a8",
          2667 => x"86",
          2668 => x"c0",
          2669 => x"5b",
          2670 => x"23",
          2671 => x"a0",
          2672 => x"8a",
          2673 => x"7c",
          2674 => x"22",
          2675 => x"22",
          2676 => x"33",
          2677 => x"33",
          2678 => x"33",
          2679 => x"33",
          2680 => x"33",
          2681 => x"52",
          2682 => x"51",
          2683 => x"8d",
          2684 => x"80",
          2685 => x"8b",
          2686 => x"30",
          2687 => x"51",
          2688 => x"0b",
          2689 => x"c0",
          2690 => x"0d",
          2691 => x"0d",
          2692 => x"82",
          2693 => x"54",
          2694 => x"94",
          2695 => x"80",
          2696 => x"87",
          2697 => x"51",
          2698 => x"96",
          2699 => x"06",
          2700 => x"70",
          2701 => x"38",
          2702 => x"70",
          2703 => x"51",
          2704 => x"71",
          2705 => x"32",
          2706 => x"51",
          2707 => x"2e",
          2708 => x"93",
          2709 => x"06",
          2710 => x"ff",
          2711 => x"0b",
          2712 => x"33",
          2713 => x"94",
          2714 => x"80",
          2715 => x"87",
          2716 => x"52",
          2717 => x"73",
          2718 => x"0c",
          2719 => x"04",
          2720 => x"02",
          2721 => x"0b",
          2722 => x"c0",
          2723 => x"87",
          2724 => x"51",
          2725 => x"86",
          2726 => x"94",
          2727 => x"08",
          2728 => x"70",
          2729 => x"52",
          2730 => x"2e",
          2731 => x"91",
          2732 => x"06",
          2733 => x"d7",
          2734 => x"2a",
          2735 => x"81",
          2736 => x"70",
          2737 => x"38",
          2738 => x"70",
          2739 => x"51",
          2740 => x"38",
          2741 => x"8b",
          2742 => x"87",
          2743 => x"52",
          2744 => x"86",
          2745 => x"94",
          2746 => x"72",
          2747 => x"0d",
          2748 => x"0d",
          2749 => x"74",
          2750 => x"70",
          2751 => x"f7",
          2752 => x"81",
          2753 => x"0b",
          2754 => x"c0",
          2755 => x"87",
          2756 => x"51",
          2757 => x"86",
          2758 => x"94",
          2759 => x"08",
          2760 => x"70",
          2761 => x"52",
          2762 => x"2e",
          2763 => x"91",
          2764 => x"06",
          2765 => x"d7",
          2766 => x"2a",
          2767 => x"81",
          2768 => x"70",
          2769 => x"38",
          2770 => x"70",
          2771 => x"51",
          2772 => x"38",
          2773 => x"8b",
          2774 => x"87",
          2775 => x"52",
          2776 => x"86",
          2777 => x"94",
          2778 => x"72",
          2779 => x"74",
          2780 => x"70",
          2781 => x"75",
          2782 => x"0c",
          2783 => x"04",
          2784 => x"0b",
          2785 => x"c0",
          2786 => x"c0",
          2787 => x"71",
          2788 => x"38",
          2789 => x"94",
          2790 => x"70",
          2791 => x"81",
          2792 => x"51",
          2793 => x"e2",
          2794 => x"82",
          2795 => x"51",
          2796 => x"80",
          2797 => x"2e",
          2798 => x"c0",
          2799 => x"71",
          2800 => x"ff",
          2801 => x"c8",
          2802 => x"3d",
          2803 => x"3d",
          2804 => x"82",
          2805 => x"51",
          2806 => x"84",
          2807 => x"2e",
          2808 => x"c0",
          2809 => x"71",
          2810 => x"2a",
          2811 => x"51",
          2812 => x"52",
          2813 => x"a2",
          2814 => x"82",
          2815 => x"51",
          2816 => x"80",
          2817 => x"2e",
          2818 => x"c0",
          2819 => x"71",
          2820 => x"2b",
          2821 => x"51",
          2822 => x"82",
          2823 => x"83",
          2824 => x"fd",
          2825 => x"c0",
          2826 => x"08",
          2827 => x"8a",
          2828 => x"53",
          2829 => x"83",
          2830 => x"8b",
          2831 => x"c0",
          2832 => x"71",
          2833 => x"87",
          2834 => x"08",
          2835 => x"88",
          2836 => x"9e",
          2837 => x"0c",
          2838 => x"87",
          2839 => x"08",
          2840 => x"90",
          2841 => x"9e",
          2842 => x"0c",
          2843 => x"87",
          2844 => x"08",
          2845 => x"98",
          2846 => x"9e",
          2847 => x"0c",
          2848 => x"87",
          2849 => x"08",
          2850 => x"a0",
          2851 => x"9e",
          2852 => x"0c",
          2853 => x"52",
          2854 => x"13",
          2855 => x"87",
          2856 => x"08",
          2857 => x"81",
          2858 => x"34",
          2859 => x"80",
          2860 => x"9e",
          2861 => x"a0",
          2862 => x"52",
          2863 => x"2e",
          2864 => x"53",
          2865 => x"80",
          2866 => x"9e",
          2867 => x"81",
          2868 => x"51",
          2869 => x"80",
          2870 => x"81",
          2871 => x"8b",
          2872 => x"0b",
          2873 => x"88",
          2874 => x"c0",
          2875 => x"52",
          2876 => x"2e",
          2877 => x"52",
          2878 => x"f3",
          2879 => x"87",
          2880 => x"08",
          2881 => x"06",
          2882 => x"70",
          2883 => x"38",
          2884 => x"82",
          2885 => x"80",
          2886 => x"9e",
          2887 => x"88",
          2888 => x"52",
          2889 => x"2e",
          2890 => x"52",
          2891 => x"f5",
          2892 => x"87",
          2893 => x"08",
          2894 => x"06",
          2895 => x"70",
          2896 => x"38",
          2897 => x"82",
          2898 => x"80",
          2899 => x"9e",
          2900 => x"82",
          2901 => x"52",
          2902 => x"2e",
          2903 => x"52",
          2904 => x"f7",
          2905 => x"87",
          2906 => x"08",
          2907 => x"06",
          2908 => x"70",
          2909 => x"38",
          2910 => x"82",
          2911 => x"82",
          2912 => x"87",
          2913 => x"70",
          2914 => x"e0",
          2915 => x"2c",
          2916 => x"53",
          2917 => x"81",
          2918 => x"71",
          2919 => x"08",
          2920 => x"51",
          2921 => x"80",
          2922 => x"81",
          2923 => x"34",
          2924 => x"c0",
          2925 => x"70",
          2926 => x"52",
          2927 => x"2e",
          2928 => x"52",
          2929 => x"fb",
          2930 => x"9e",
          2931 => x"87",
          2932 => x"70",
          2933 => x"34",
          2934 => x"04",
          2935 => x"81",
          2936 => x"84",
          2937 => x"8b",
          2938 => x"73",
          2939 => x"38",
          2940 => x"51",
          2941 => x"81",
          2942 => x"84",
          2943 => x"8b",
          2944 => x"55",
          2945 => x"2e",
          2946 => x"15",
          2947 => x"8b",
          2948 => x"81",
          2949 => x"8a",
          2950 => x"8b",
          2951 => x"55",
          2952 => x"2e",
          2953 => x"15",
          2954 => x"15",
          2955 => x"f7",
          2956 => x"e9",
          2957 => x"f3",
          2958 => x"55",
          2959 => x"81",
          2960 => x"73",
          2961 => x"38",
          2962 => x"70",
          2963 => x"11",
          2964 => x"81",
          2965 => x"89",
          2966 => x"8b",
          2967 => x"73",
          2968 => x"38",
          2969 => x"51",
          2970 => x"82",
          2971 => x"54",
          2972 => x"88",
          2973 => x"fc",
          2974 => x"3f",
          2975 => x"33",
          2976 => x"2e",
          2977 => x"f8",
          2978 => x"97",
          2979 => x"f8",
          2980 => x"55",
          2981 => x"8c",
          2982 => x"33",
          2983 => x"94",
          2984 => x"3f",
          2985 => x"33",
          2986 => x"2e",
          2987 => x"f8",
          2988 => x"ef",
          2989 => x"fb",
          2990 => x"55",
          2991 => x"8c",
          2992 => x"33",
          2993 => x"d0",
          2994 => x"3f",
          2995 => x"51",
          2996 => x"82",
          2997 => x"70",
          2998 => x"52",
          2999 => x"f8",
          3000 => x"55",
          3001 => x"73",
          3002 => x"f9",
          3003 => x"ad",
          3004 => x"08",
          3005 => x"c8",
          3006 => x"3f",
          3007 => x"52",
          3008 => x"51",
          3009 => x"90",
          3010 => x"81",
          3011 => x"88",
          3012 => x"3d",
          3013 => x"3d",
          3014 => x"05",
          3015 => x"85",
          3016 => x"71",
          3017 => x"0b",
          3018 => x"05",
          3019 => x"04",
          3020 => x"51",
          3021 => x"ac",
          3022 => x"c8",
          3023 => x"3f",
          3024 => x"fa",
          3025 => x"a9",
          3026 => x"81",
          3027 => x"f7",
          3028 => x"39",
          3029 => x"51",
          3030 => x"88",
          3031 => x"e4",
          3032 => x"3f",
          3033 => x"04",
          3034 => x"0c",
          3035 => x"87",
          3036 => x"0c",
          3037 => x"0d",
          3038 => x"84",
          3039 => x"52",
          3040 => x"70",
          3041 => x"82",
          3042 => x"72",
          3043 => x"0d",
          3044 => x"0d",
          3045 => x"84",
          3046 => x"8c",
          3047 => x"80",
          3048 => x"09",
          3049 => x"80",
          3050 => x"82",
          3051 => x"73",
          3052 => x"3d",
          3053 => x"8c",
          3054 => x"c0",
          3055 => x"04",
          3056 => x"02",
          3057 => x"53",
          3058 => x"09",
          3059 => x"38",
          3060 => x"3f",
          3061 => x"08",
          3062 => x"38",
          3063 => x"08",
          3064 => x"34",
          3065 => x"08",
          3066 => x"93",
          3067 => x"39",
          3068 => x"08",
          3069 => x"38",
          3070 => x"93",
          3071 => x"71",
          3072 => x"0d",
          3073 => x"0d",
          3074 => x"33",
          3075 => x"08",
          3076 => x"d8",
          3077 => x"ff",
          3078 => x"82",
          3079 => x"84",
          3080 => x"fe",
          3081 => x"70",
          3082 => x"71",
          3083 => x"38",
          3084 => x"05",
          3085 => x"ff",
          3086 => x"33",
          3087 => x"38",
          3088 => x"04",
          3089 => x"76",
          3090 => x"08",
          3091 => x"d8",
          3092 => x"54",
          3093 => x"80",
          3094 => x"72",
          3095 => x"54",
          3096 => x"dc",
          3097 => x"52",
          3098 => x"73",
          3099 => x"0c",
          3100 => x"04",
          3101 => x"66",
          3102 => x"78",
          3103 => x"5a",
          3104 => x"80",
          3105 => x"38",
          3106 => x"88",
          3107 => x"fe",
          3108 => x"39",
          3109 => x"70",
          3110 => x"33",
          3111 => x"75",
          3112 => x"81",
          3113 => x"81",
          3114 => x"05",
          3115 => x"5d",
          3116 => x"ad",
          3117 => x"06",
          3118 => x"79",
          3119 => x"5b",
          3120 => x"75",
          3121 => x"81",
          3122 => x"7b",
          3123 => x"08",
          3124 => x"05",
          3125 => x"5c",
          3126 => x"39",
          3127 => x"72",
          3128 => x"38",
          3129 => x"16",
          3130 => x"70",
          3131 => x"33",
          3132 => x"57",
          3133 => x"27",
          3134 => x"80",
          3135 => x"30",
          3136 => x"80",
          3137 => x"cc",
          3138 => x"70",
          3139 => x"25",
          3140 => x"59",
          3141 => x"54",
          3142 => x"8c",
          3143 => x"07",
          3144 => x"05",
          3145 => x"5d",
          3146 => x"83",
          3147 => x"55",
          3148 => x"27",
          3149 => x"16",
          3150 => x"06",
          3151 => x"be",
          3152 => x"96",
          3153 => x"38",
          3154 => x"81",
          3155 => x"53",
          3156 => x"7b",
          3157 => x"08",
          3158 => x"80",
          3159 => x"54",
          3160 => x"8d",
          3161 => x"70",
          3162 => x"51",
          3163 => x"f5",
          3164 => x"2a",
          3165 => x"51",
          3166 => x"38",
          3167 => x"55",
          3168 => x"27",
          3169 => x"81",
          3170 => x"56",
          3171 => x"b0",
          3172 => x"38",
          3173 => x"55",
          3174 => x"26",
          3175 => x"51",
          3176 => x"73",
          3177 => x"53",
          3178 => x"fd",
          3179 => x"51",
          3180 => x"73",
          3181 => x"53",
          3182 => x"f2",
          3183 => x"39",
          3184 => x"83",
          3185 => x"5d",
          3186 => x"3f",
          3187 => x"82",
          3188 => x"88",
          3189 => x"8a",
          3190 => x"90",
          3191 => x"75",
          3192 => x"3f",
          3193 => x"7c",
          3194 => x"81",
          3195 => x"72",
          3196 => x"38",
          3197 => x"71",
          3198 => x"53",
          3199 => x"80",
          3200 => x"81",
          3201 => x"7b",
          3202 => x"08",
          3203 => x"89",
          3204 => x"1d",
          3205 => x"5d",
          3206 => x"c4",
          3207 => x"70",
          3208 => x"25",
          3209 => x"24",
          3210 => x"55",
          3211 => x"2e",
          3212 => x"30",
          3213 => x"5e",
          3214 => x"7a",
          3215 => x"e6",
          3216 => x"93",
          3217 => x"ff",
          3218 => x"77",
          3219 => x"e6",
          3220 => x"c8",
          3221 => x"75",
          3222 => x"74",
          3223 => x"81",
          3224 => x"54",
          3225 => x"f8",
          3226 => x"87",
          3227 => x"ff",
          3228 => x"96",
          3229 => x"e0",
          3230 => x"54",
          3231 => x"34",
          3232 => x"30",
          3233 => x"9f",
          3234 => x"74",
          3235 => x"51",
          3236 => x"ff",
          3237 => x"84",
          3238 => x"06",
          3239 => x"80",
          3240 => x"96",
          3241 => x"e0",
          3242 => x"73",
          3243 => x"58",
          3244 => x"06",
          3245 => x"55",
          3246 => x"a0",
          3247 => x"2a",
          3248 => x"51",
          3249 => x"38",
          3250 => x"55",
          3251 => x"27",
          3252 => x"81",
          3253 => x"56",
          3254 => x"e4",
          3255 => x"38",
          3256 => x"55",
          3257 => x"26",
          3258 => x"18",
          3259 => x"05",
          3260 => x"53",
          3261 => x"c8",
          3262 => x"38",
          3263 => x"55",
          3264 => x"27",
          3265 => x"a0",
          3266 => x"3f",
          3267 => x"55",
          3268 => x"26",
          3269 => x"e3",
          3270 => x"0d",
          3271 => x"0d",
          3272 => x"70",
          3273 => x"08",
          3274 => x"51",
          3275 => x"85",
          3276 => x"fe",
          3277 => x"82",
          3278 => x"85",
          3279 => x"52",
          3280 => x"b0",
          3281 => x"e0",
          3282 => x"73",
          3283 => x"82",
          3284 => x"84",
          3285 => x"fd",
          3286 => x"93",
          3287 => x"82",
          3288 => x"87",
          3289 => x"53",
          3290 => x"fa",
          3291 => x"82",
          3292 => x"85",
          3293 => x"fa",
          3294 => x"7a",
          3295 => x"53",
          3296 => x"08",
          3297 => x"fa",
          3298 => x"73",
          3299 => x"39",
          3300 => x"93",
          3301 => x"71",
          3302 => x"c8",
          3303 => x"06",
          3304 => x"2e",
          3305 => x"8d",
          3306 => x"38",
          3307 => x"70",
          3308 => x"70",
          3309 => x"2a",
          3310 => x"06",
          3311 => x"53",
          3312 => x"8e",
          3313 => x"74",
          3314 => x"52",
          3315 => x"3f",
          3316 => x"74",
          3317 => x"38",
          3318 => x"74",
          3319 => x"b2",
          3320 => x"52",
          3321 => x"81",
          3322 => x"ff",
          3323 => x"f7",
          3324 => x"9e",
          3325 => x"52",
          3326 => x"8a",
          3327 => x"3f",
          3328 => x"82",
          3329 => x"88",
          3330 => x"fe",
          3331 => x"93",
          3332 => x"82",
          3333 => x"77",
          3334 => x"53",
          3335 => x"72",
          3336 => x"0c",
          3337 => x"04",
          3338 => x"7a",
          3339 => x"80",
          3340 => x"75",
          3341 => x"56",
          3342 => x"a0",
          3343 => x"06",
          3344 => x"08",
          3345 => x"0c",
          3346 => x"33",
          3347 => x"a0",
          3348 => x"73",
          3349 => x"81",
          3350 => x"81",
          3351 => x"76",
          3352 => x"70",
          3353 => x"58",
          3354 => x"09",
          3355 => x"d3",
          3356 => x"81",
          3357 => x"74",
          3358 => x"55",
          3359 => x"e2",
          3360 => x"73",
          3361 => x"09",
          3362 => x"38",
          3363 => x"14",
          3364 => x"08",
          3365 => x"54",
          3366 => x"39",
          3367 => x"81",
          3368 => x"75",
          3369 => x"56",
          3370 => x"39",
          3371 => x"74",
          3372 => x"38",
          3373 => x"80",
          3374 => x"89",
          3375 => x"38",
          3376 => x"d0",
          3377 => x"56",
          3378 => x"80",
          3379 => x"39",
          3380 => x"e1",
          3381 => x"80",
          3382 => x"57",
          3383 => x"74",
          3384 => x"38",
          3385 => x"27",
          3386 => x"14",
          3387 => x"06",
          3388 => x"14",
          3389 => x"06",
          3390 => x"74",
          3391 => x"f9",
          3392 => x"ff",
          3393 => x"89",
          3394 => x"38",
          3395 => x"c5",
          3396 => x"29",
          3397 => x"81",
          3398 => x"75",
          3399 => x"56",
          3400 => x"a0",
          3401 => x"38",
          3402 => x"84",
          3403 => x"56",
          3404 => x"81",
          3405 => x"93",
          3406 => x"3d",
          3407 => x"3d",
          3408 => x"5a",
          3409 => x"7a",
          3410 => x"70",
          3411 => x"58",
          3412 => x"09",
          3413 => x"38",
          3414 => x"05",
          3415 => x"08",
          3416 => x"53",
          3417 => x"f0",
          3418 => x"2e",
          3419 => x"8e",
          3420 => x"08",
          3421 => x"75",
          3422 => x"56",
          3423 => x"b0",
          3424 => x"06",
          3425 => x"74",
          3426 => x"75",
          3427 => x"70",
          3428 => x"73",
          3429 => x"9a",
          3430 => x"f8",
          3431 => x"06",
          3432 => x"0b",
          3433 => x"0c",
          3434 => x"33",
          3435 => x"80",
          3436 => x"75",
          3437 => x"76",
          3438 => x"70",
          3439 => x"57",
          3440 => x"56",
          3441 => x"81",
          3442 => x"14",
          3443 => x"88",
          3444 => x"27",
          3445 => x"f3",
          3446 => x"53",
          3447 => x"89",
          3448 => x"38",
          3449 => x"56",
          3450 => x"80",
          3451 => x"39",
          3452 => x"56",
          3453 => x"80",
          3454 => x"e0",
          3455 => x"38",
          3456 => x"81",
          3457 => x"53",
          3458 => x"81",
          3459 => x"53",
          3460 => x"8e",
          3461 => x"70",
          3462 => x"55",
          3463 => x"27",
          3464 => x"77",
          3465 => x"76",
          3466 => x"75",
          3467 => x"76",
          3468 => x"70",
          3469 => x"56",
          3470 => x"ff",
          3471 => x"80",
          3472 => x"75",
          3473 => x"79",
          3474 => x"75",
          3475 => x"0c",
          3476 => x"04",
          3477 => x"02",
          3478 => x"51",
          3479 => x"72",
          3480 => x"82",
          3481 => x"33",
          3482 => x"93",
          3483 => x"3d",
          3484 => x"3d",
          3485 => x"05",
          3486 => x"05",
          3487 => x"55",
          3488 => x"72",
          3489 => x"ed",
          3490 => x"29",
          3491 => x"8c",
          3492 => x"52",
          3493 => x"84",
          3494 => x"52",
          3495 => x"72",
          3496 => x"c0",
          3497 => x"51",
          3498 => x"85",
          3499 => x"98",
          3500 => x"52",
          3501 => x"8c",
          3502 => x"70",
          3503 => x"51",
          3504 => x"87",
          3505 => x"51",
          3506 => x"72",
          3507 => x"c0",
          3508 => x"70",
          3509 => x"80",
          3510 => x"71",
          3511 => x"c0",
          3512 => x"51",
          3513 => x"87",
          3514 => x"8c",
          3515 => x"82",
          3516 => x"33",
          3517 => x"93",
          3518 => x"3d",
          3519 => x"3d",
          3520 => x"65",
          3521 => x"80",
          3522 => x"56",
          3523 => x"83",
          3524 => x"fe",
          3525 => x"93",
          3526 => x"06",
          3527 => x"71",
          3528 => x"80",
          3529 => x"87",
          3530 => x"73",
          3531 => x"c0",
          3532 => x"87",
          3533 => x"12",
          3534 => x"57",
          3535 => x"76",
          3536 => x"92",
          3537 => x"71",
          3538 => x"75",
          3539 => x"70",
          3540 => x"81",
          3541 => x"54",
          3542 => x"8e",
          3543 => x"52",
          3544 => x"81",
          3545 => x"81",
          3546 => x"a2",
          3547 => x"80",
          3548 => x"75",
          3549 => x"d5",
          3550 => x"52",
          3551 => x"87",
          3552 => x"80",
          3553 => x"81",
          3554 => x"c0",
          3555 => x"53",
          3556 => x"82",
          3557 => x"71",
          3558 => x"1b",
          3559 => x"84",
          3560 => x"1e",
          3561 => x"06",
          3562 => x"7a",
          3563 => x"38",
          3564 => x"80",
          3565 => x"87",
          3566 => x"26",
          3567 => x"73",
          3568 => x"06",
          3569 => x"2e",
          3570 => x"52",
          3571 => x"82",
          3572 => x"90",
          3573 => x"f3",
          3574 => x"62",
          3575 => x"05",
          3576 => x"56",
          3577 => x"83",
          3578 => x"fc",
          3579 => x"93",
          3580 => x"06",
          3581 => x"71",
          3582 => x"80",
          3583 => x"98",
          3584 => x"2b",
          3585 => x"8c",
          3586 => x"92",
          3587 => x"41",
          3588 => x"56",
          3589 => x"87",
          3590 => x"19",
          3591 => x"52",
          3592 => x"80",
          3593 => x"70",
          3594 => x"81",
          3595 => x"54",
          3596 => x"8c",
          3597 => x"81",
          3598 => x"78",
          3599 => x"53",
          3600 => x"70",
          3601 => x"52",
          3602 => x"87",
          3603 => x"52",
          3604 => x"75",
          3605 => x"80",
          3606 => x"72",
          3607 => x"99",
          3608 => x"0c",
          3609 => x"8c",
          3610 => x"08",
          3611 => x"51",
          3612 => x"38",
          3613 => x"8d",
          3614 => x"70",
          3615 => x"84",
          3616 => x"5d",
          3617 => x"2e",
          3618 => x"fc",
          3619 => x"52",
          3620 => x"7d",
          3621 => x"fc",
          3622 => x"80",
          3623 => x"71",
          3624 => x"38",
          3625 => x"54",
          3626 => x"c8",
          3627 => x"0d",
          3628 => x"0d",
          3629 => x"05",
          3630 => x"02",
          3631 => x"05",
          3632 => x"55",
          3633 => x"8c",
          3634 => x"c8",
          3635 => x"52",
          3636 => x"bc",
          3637 => x"72",
          3638 => x"38",
          3639 => x"88",
          3640 => x"2e",
          3641 => x"39",
          3642 => x"9a",
          3643 => x"74",
          3644 => x"c0",
          3645 => x"70",
          3646 => x"94",
          3647 => x"0a",
          3648 => x"54",
          3649 => x"80",
          3650 => x"54",
          3651 => x"54",
          3652 => x"c8",
          3653 => x"0d",
          3654 => x"0d",
          3655 => x"81",
          3656 => x"88",
          3657 => x"82",
          3658 => x"52",
          3659 => x"3d",
          3660 => x"3d",
          3661 => x"11",
          3662 => x"33",
          3663 => x"71",
          3664 => x"81",
          3665 => x"07",
          3666 => x"88",
          3667 => x"93",
          3668 => x"54",
          3669 => x"85",
          3670 => x"ff",
          3671 => x"02",
          3672 => x"05",
          3673 => x"70",
          3674 => x"05",
          3675 => x"88",
          3676 => x"72",
          3677 => x"0d",
          3678 => x"0d",
          3679 => x"52",
          3680 => x"81",
          3681 => x"70",
          3682 => x"70",
          3683 => x"05",
          3684 => x"88",
          3685 => x"72",
          3686 => x"54",
          3687 => x"2a",
          3688 => x"34",
          3689 => x"04",
          3690 => x"76",
          3691 => x"54",
          3692 => x"2e",
          3693 => x"70",
          3694 => x"33",
          3695 => x"05",
          3696 => x"11",
          3697 => x"38",
          3698 => x"04",
          3699 => x"75",
          3700 => x"52",
          3701 => x"70",
          3702 => x"34",
          3703 => x"70",
          3704 => x"3d",
          3705 => x"3d",
          3706 => x"79",
          3707 => x"74",
          3708 => x"56",
          3709 => x"81",
          3710 => x"71",
          3711 => x"16",
          3712 => x"52",
          3713 => x"86",
          3714 => x"2e",
          3715 => x"82",
          3716 => x"86",
          3717 => x"fe",
          3718 => x"76",
          3719 => x"54",
          3720 => x"2e",
          3721 => x"73",
          3722 => x"81",
          3723 => x"52",
          3724 => x"2e",
          3725 => x"73",
          3726 => x"06",
          3727 => x"33",
          3728 => x"0c",
          3729 => x"04",
          3730 => x"93",
          3731 => x"80",
          3732 => x"c8",
          3733 => x"3d",
          3734 => x"80",
          3735 => x"33",
          3736 => x"78",
          3737 => x"38",
          3738 => x"16",
          3739 => x"16",
          3740 => x"17",
          3741 => x"fa",
          3742 => x"93",
          3743 => x"2e",
          3744 => x"b8",
          3745 => x"c8",
          3746 => x"34",
          3747 => x"a4",
          3748 => x"55",
          3749 => x"08",
          3750 => x"82",
          3751 => x"74",
          3752 => x"81",
          3753 => x"81",
          3754 => x"08",
          3755 => x"05",
          3756 => x"81",
          3757 => x"fa",
          3758 => x"39",
          3759 => x"82",
          3760 => x"89",
          3761 => x"fa",
          3762 => x"7a",
          3763 => x"56",
          3764 => x"75",
          3765 => x"76",
          3766 => x"3f",
          3767 => x"08",
          3768 => x"c8",
          3769 => x"81",
          3770 => x"b4",
          3771 => x"17",
          3772 => x"8a",
          3773 => x"c8",
          3774 => x"85",
          3775 => x"81",
          3776 => x"18",
          3777 => x"93",
          3778 => x"3d",
          3779 => x"3d",
          3780 => x"52",
          3781 => x"3f",
          3782 => x"08",
          3783 => x"c8",
          3784 => x"38",
          3785 => x"74",
          3786 => x"81",
          3787 => x"38",
          3788 => x"59",
          3789 => x"09",
          3790 => x"e3",
          3791 => x"53",
          3792 => x"08",
          3793 => x"70",
          3794 => x"80",
          3795 => x"d5",
          3796 => x"17",
          3797 => x"3f",
          3798 => x"a4",
          3799 => x"51",
          3800 => x"86",
          3801 => x"f2",
          3802 => x"17",
          3803 => x"3f",
          3804 => x"52",
          3805 => x"51",
          3806 => x"8c",
          3807 => x"84",
          3808 => x"fb",
          3809 => x"17",
          3810 => x"70",
          3811 => x"79",
          3812 => x"52",
          3813 => x"51",
          3814 => x"77",
          3815 => x"80",
          3816 => x"81",
          3817 => x"fa",
          3818 => x"93",
          3819 => x"2e",
          3820 => x"58",
          3821 => x"c8",
          3822 => x"0d",
          3823 => x"0d",
          3824 => x"98",
          3825 => x"05",
          3826 => x"80",
          3827 => x"27",
          3828 => x"14",
          3829 => x"29",
          3830 => x"05",
          3831 => x"82",
          3832 => x"87",
          3833 => x"f9",
          3834 => x"7a",
          3835 => x"54",
          3836 => x"27",
          3837 => x"14",
          3838 => x"86",
          3839 => x"81",
          3840 => x"74",
          3841 => x"72",
          3842 => x"f5",
          3843 => x"24",
          3844 => x"81",
          3845 => x"81",
          3846 => x"83",
          3847 => x"38",
          3848 => x"74",
          3849 => x"70",
          3850 => x"16",
          3851 => x"74",
          3852 => x"93",
          3853 => x"c8",
          3854 => x"38",
          3855 => x"06",
          3856 => x"33",
          3857 => x"89",
          3858 => x"08",
          3859 => x"54",
          3860 => x"fc",
          3861 => x"93",
          3862 => x"fe",
          3863 => x"ff",
          3864 => x"11",
          3865 => x"2b",
          3866 => x"81",
          3867 => x"2a",
          3868 => x"51",
          3869 => x"e2",
          3870 => x"ff",
          3871 => x"da",
          3872 => x"2a",
          3873 => x"05",
          3874 => x"fc",
          3875 => x"93",
          3876 => x"c6",
          3877 => x"83",
          3878 => x"05",
          3879 => x"f8",
          3880 => x"93",
          3881 => x"ff",
          3882 => x"ae",
          3883 => x"2a",
          3884 => x"05",
          3885 => x"fc",
          3886 => x"93",
          3887 => x"38",
          3888 => x"83",
          3889 => x"05",
          3890 => x"f8",
          3891 => x"93",
          3892 => x"0a",
          3893 => x"39",
          3894 => x"82",
          3895 => x"89",
          3896 => x"f7",
          3897 => x"7d",
          3898 => x"55",
          3899 => x"74",
          3900 => x"38",
          3901 => x"08",
          3902 => x"38",
          3903 => x"72",
          3904 => x"a8",
          3905 => x"24",
          3906 => x"81",
          3907 => x"82",
          3908 => x"83",
          3909 => x"38",
          3910 => x"73",
          3911 => x"70",
          3912 => x"17",
          3913 => x"75",
          3914 => x"9b",
          3915 => x"c8",
          3916 => x"93",
          3917 => x"ea",
          3918 => x"ff",
          3919 => x"11",
          3920 => x"81",
          3921 => x"51",
          3922 => x"72",
          3923 => x"38",
          3924 => x"9f",
          3925 => x"33",
          3926 => x"07",
          3927 => x"78",
          3928 => x"83",
          3929 => x"89",
          3930 => x"08",
          3931 => x"51",
          3932 => x"82",
          3933 => x"57",
          3934 => x"08",
          3935 => x"78",
          3936 => x"15",
          3937 => x"81",
          3938 => x"2a",
          3939 => x"58",
          3940 => x"75",
          3941 => x"33",
          3942 => x"76",
          3943 => x"07",
          3944 => x"34",
          3945 => x"16",
          3946 => x"39",
          3947 => x"a4",
          3948 => x"52",
          3949 => x"8f",
          3950 => x"c8",
          3951 => x"93",
          3952 => x"de",
          3953 => x"ff",
          3954 => x"73",
          3955 => x"06",
          3956 => x"05",
          3957 => x"3f",
          3958 => x"16",
          3959 => x"39",
          3960 => x"a4",
          3961 => x"52",
          3962 => x"db",
          3963 => x"c8",
          3964 => x"93",
          3965 => x"38",
          3966 => x"06",
          3967 => x"83",
          3968 => x"11",
          3969 => x"54",
          3970 => x"f6",
          3971 => x"93",
          3972 => x"0a",
          3973 => x"52",
          3974 => x"dd",
          3975 => x"83",
          3976 => x"82",
          3977 => x"8b",
          3978 => x"f9",
          3979 => x"7b",
          3980 => x"58",
          3981 => x"81",
          3982 => x"38",
          3983 => x"74",
          3984 => x"82",
          3985 => x"39",
          3986 => x"aa",
          3987 => x"75",
          3988 => x"fd",
          3989 => x"93",
          3990 => x"82",
          3991 => x"80",
          3992 => x"39",
          3993 => x"ed",
          3994 => x"80",
          3995 => x"93",
          3996 => x"80",
          3997 => x"52",
          3998 => x"eb",
          3999 => x"c8",
          4000 => x"93",
          4001 => x"2e",
          4002 => x"82",
          4003 => x"81",
          4004 => x"82",
          4005 => x"ff",
          4006 => x"80",
          4007 => x"74",
          4008 => x"3f",
          4009 => x"08",
          4010 => x"15",
          4011 => x"54",
          4012 => x"74",
          4013 => x"90",
          4014 => x"05",
          4015 => x"84",
          4016 => x"07",
          4017 => x"16",
          4018 => x"98",
          4019 => x"26",
          4020 => x"80",
          4021 => x"93",
          4022 => x"3d",
          4023 => x"3d",
          4024 => x"71",
          4025 => x"5c",
          4026 => x"8c",
          4027 => x"77",
          4028 => x"38",
          4029 => x"78",
          4030 => x"81",
          4031 => x"7a",
          4032 => x"f9",
          4033 => x"55",
          4034 => x"c8",
          4035 => x"e9",
          4036 => x"c8",
          4037 => x"93",
          4038 => x"2e",
          4039 => x"82",
          4040 => x"55",
          4041 => x"82",
          4042 => x"26",
          4043 => x"7a",
          4044 => x"90",
          4045 => x"2e",
          4046 => x"80",
          4047 => x"2e",
          4048 => x"80",
          4049 => x"1b",
          4050 => x"08",
          4051 => x"38",
          4052 => x"52",
          4053 => x"8f",
          4054 => x"c8",
          4055 => x"5a",
          4056 => x"08",
          4057 => x"81",
          4058 => x"82",
          4059 => x"5a",
          4060 => x"70",
          4061 => x"07",
          4062 => x"7d",
          4063 => x"51",
          4064 => x"73",
          4065 => x"75",
          4066 => x"38",
          4067 => x"56",
          4068 => x"8a",
          4069 => x"1a",
          4070 => x"38",
          4071 => x"57",
          4072 => x"38",
          4073 => x"17",
          4074 => x"08",
          4075 => x"38",
          4076 => x"78",
          4077 => x"38",
          4078 => x"51",
          4079 => x"82",
          4080 => x"56",
          4081 => x"08",
          4082 => x"38",
          4083 => x"93",
          4084 => x"2e",
          4085 => x"86",
          4086 => x"c8",
          4087 => x"ff",
          4088 => x"70",
          4089 => x"25",
          4090 => x"51",
          4091 => x"73",
          4092 => x"76",
          4093 => x"81",
          4094 => x"38",
          4095 => x"f9",
          4096 => x"76",
          4097 => x"f9",
          4098 => x"93",
          4099 => x"93",
          4100 => x"70",
          4101 => x"08",
          4102 => x"7d",
          4103 => x"07",
          4104 => x"06",
          4105 => x"56",
          4106 => x"2e",
          4107 => x"53",
          4108 => x"51",
          4109 => x"82",
          4110 => x"56",
          4111 => x"76",
          4112 => x"98",
          4113 => x"05",
          4114 => x"08",
          4115 => x"38",
          4116 => x"ff",
          4117 => x"0c",
          4118 => x"81",
          4119 => x"84",
          4120 => x"39",
          4121 => x"81",
          4122 => x"89",
          4123 => x"89",
          4124 => x"85",
          4125 => x"76",
          4126 => x"93",
          4127 => x"3d",
          4128 => x"3d",
          4129 => x"52",
          4130 => x"3f",
          4131 => x"93",
          4132 => x"db",
          4133 => x"76",
          4134 => x"3f",
          4135 => x"08",
          4136 => x"08",
          4137 => x"5a",
          4138 => x"80",
          4139 => x"70",
          4140 => x"98",
          4141 => x"81",
          4142 => x"84",
          4143 => x"56",
          4144 => x"55",
          4145 => x"97",
          4146 => x"75",
          4147 => x"52",
          4148 => x"51",
          4149 => x"82",
          4150 => x"80",
          4151 => x"80",
          4152 => x"22",
          4153 => x"76",
          4154 => x"81",
          4155 => x"74",
          4156 => x"0c",
          4157 => x"04",
          4158 => x"7a",
          4159 => x"58",
          4160 => x"f0",
          4161 => x"8a",
          4162 => x"06",
          4163 => x"2e",
          4164 => x"58",
          4165 => x"74",
          4166 => x"88",
          4167 => x"73",
          4168 => x"33",
          4169 => x"27",
          4170 => x"16",
          4171 => x"9b",
          4172 => x"2a",
          4173 => x"88",
          4174 => x"58",
          4175 => x"81",
          4176 => x"16",
          4177 => x"0c",
          4178 => x"8a",
          4179 => x"89",
          4180 => x"72",
          4181 => x"38",
          4182 => x"51",
          4183 => x"82",
          4184 => x"54",
          4185 => x"08",
          4186 => x"38",
          4187 => x"93",
          4188 => x"8b",
          4189 => x"08",
          4190 => x"08",
          4191 => x"82",
          4192 => x"39",
          4193 => x"55",
          4194 => x"cc",
          4195 => x"75",
          4196 => x"3f",
          4197 => x"08",
          4198 => x"73",
          4199 => x"82",
          4200 => x"08",
          4201 => x"38",
          4202 => x"58",
          4203 => x"89",
          4204 => x"08",
          4205 => x"0c",
          4206 => x"06",
          4207 => x"9c",
          4208 => x"58",
          4209 => x"c8",
          4210 => x"0d",
          4211 => x"0d",
          4212 => x"08",
          4213 => x"a0",
          4214 => x"59",
          4215 => x"0a",
          4216 => x"38",
          4217 => x"16",
          4218 => x"98",
          4219 => x"2e",
          4220 => x"75",
          4221 => x"54",
          4222 => x"38",
          4223 => x"81",
          4224 => x"0c",
          4225 => x"98",
          4226 => x"2a",
          4227 => x"59",
          4228 => x"26",
          4229 => x"73",
          4230 => x"84",
          4231 => x"39",
          4232 => x"ff",
          4233 => x"2a",
          4234 => x"72",
          4235 => x"94",
          4236 => x"74",
          4237 => x"3f",
          4238 => x"08",
          4239 => x"81",
          4240 => x"c8",
          4241 => x"84",
          4242 => x"82",
          4243 => x"ff",
          4244 => x"38",
          4245 => x"82",
          4246 => x"26",
          4247 => x"77",
          4248 => x"98",
          4249 => x"53",
          4250 => x"94",
          4251 => x"74",
          4252 => x"3f",
          4253 => x"08",
          4254 => x"82",
          4255 => x"80",
          4256 => x"38",
          4257 => x"93",
          4258 => x"2e",
          4259 => x"53",
          4260 => x"08",
          4261 => x"38",
          4262 => x"08",
          4263 => x"fb",
          4264 => x"53",
          4265 => x"08",
          4266 => x"94",
          4267 => x"52",
          4268 => x"89",
          4269 => x"c8",
          4270 => x"0c",
          4271 => x"0c",
          4272 => x"06",
          4273 => x"9c",
          4274 => x"53",
          4275 => x"c8",
          4276 => x"0d",
          4277 => x"0d",
          4278 => x"08",
          4279 => x"80",
          4280 => x"fc",
          4281 => x"93",
          4282 => x"82",
          4283 => x"80",
          4284 => x"93",
          4285 => x"98",
          4286 => x"77",
          4287 => x"3f",
          4288 => x"08",
          4289 => x"c8",
          4290 => x"38",
          4291 => x"08",
          4292 => x"70",
          4293 => x"55",
          4294 => x"2e",
          4295 => x"83",
          4296 => x"72",
          4297 => x"25",
          4298 => x"53",
          4299 => x"8b",
          4300 => x"57",
          4301 => x"9a",
          4302 => x"80",
          4303 => x"75",
          4304 => x"3f",
          4305 => x"08",
          4306 => x"c8",
          4307 => x"ff",
          4308 => x"84",
          4309 => x"06",
          4310 => x"54",
          4311 => x"c8",
          4312 => x"0d",
          4313 => x"0d",
          4314 => x"52",
          4315 => x"3f",
          4316 => x"08",
          4317 => x"06",
          4318 => x"51",
          4319 => x"83",
          4320 => x"06",
          4321 => x"14",
          4322 => x"3f",
          4323 => x"08",
          4324 => x"07",
          4325 => x"93",
          4326 => x"3d",
          4327 => x"3d",
          4328 => x"70",
          4329 => x"06",
          4330 => x"53",
          4331 => x"ab",
          4332 => x"33",
          4333 => x"83",
          4334 => x"06",
          4335 => x"90",
          4336 => x"15",
          4337 => x"3f",
          4338 => x"04",
          4339 => x"7b",
          4340 => x"84",
          4341 => x"58",
          4342 => x"80",
          4343 => x"38",
          4344 => x"52",
          4345 => x"df",
          4346 => x"c8",
          4347 => x"93",
          4348 => x"f1",
          4349 => x"08",
          4350 => x"53",
          4351 => x"84",
          4352 => x"39",
          4353 => x"8b",
          4354 => x"bf",
          4355 => x"ff",
          4356 => x"51",
          4357 => x"17",
          4358 => x"e5",
          4359 => x"76",
          4360 => x"30",
          4361 => x"9f",
          4362 => x"55",
          4363 => x"80",
          4364 => x"76",
          4365 => x"38",
          4366 => x"06",
          4367 => x"88",
          4368 => x"06",
          4369 => x"54",
          4370 => x"99",
          4371 => x"75",
          4372 => x"3f",
          4373 => x"08",
          4374 => x"c8",
          4375 => x"98",
          4376 => x"fc",
          4377 => x"2e",
          4378 => x"0b",
          4379 => x"77",
          4380 => x"0c",
          4381 => x"04",
          4382 => x"7a",
          4383 => x"56",
          4384 => x"51",
          4385 => x"82",
          4386 => x"54",
          4387 => x"08",
          4388 => x"86",
          4389 => x"80",
          4390 => x"16",
          4391 => x"51",
          4392 => x"82",
          4393 => x"57",
          4394 => x"08",
          4395 => x"9c",
          4396 => x"33",
          4397 => x"80",
          4398 => x"9c",
          4399 => x"11",
          4400 => x"55",
          4401 => x"17",
          4402 => x"33",
          4403 => x"70",
          4404 => x"55",
          4405 => x"38",
          4406 => x"16",
          4407 => x"ea",
          4408 => x"93",
          4409 => x"2e",
          4410 => x"52",
          4411 => x"dd",
          4412 => x"c8",
          4413 => x"93",
          4414 => x"2e",
          4415 => x"76",
          4416 => x"93",
          4417 => x"3d",
          4418 => x"3d",
          4419 => x"08",
          4420 => x"52",
          4421 => x"bd",
          4422 => x"c8",
          4423 => x"93",
          4424 => x"38",
          4425 => x"52",
          4426 => x"9b",
          4427 => x"c8",
          4428 => x"93",
          4429 => x"38",
          4430 => x"93",
          4431 => x"9c",
          4432 => x"e9",
          4433 => x"53",
          4434 => x"9c",
          4435 => x"e8",
          4436 => x"0b",
          4437 => x"74",
          4438 => x"0c",
          4439 => x"04",
          4440 => x"76",
          4441 => x"12",
          4442 => x"53",
          4443 => x"d7",
          4444 => x"c8",
          4445 => x"93",
          4446 => x"38",
          4447 => x"53",
          4448 => x"81",
          4449 => x"34",
          4450 => x"c8",
          4451 => x"0d",
          4452 => x"0d",
          4453 => x"57",
          4454 => x"17",
          4455 => x"08",
          4456 => x"89",
          4457 => x"55",
          4458 => x"08",
          4459 => x"81",
          4460 => x"52",
          4461 => x"ad",
          4462 => x"2e",
          4463 => x"84",
          4464 => x"53",
          4465 => x"09",
          4466 => x"38",
          4467 => x"05",
          4468 => x"81",
          4469 => x"15",
          4470 => x"88",
          4471 => x"81",
          4472 => x"15",
          4473 => x"27",
          4474 => x"15",
          4475 => x"80",
          4476 => x"34",
          4477 => x"52",
          4478 => x"88",
          4479 => x"17",
          4480 => x"51",
          4481 => x"82",
          4482 => x"76",
          4483 => x"08",
          4484 => x"e6",
          4485 => x"93",
          4486 => x"17",
          4487 => x"08",
          4488 => x"e5",
          4489 => x"93",
          4490 => x"17",
          4491 => x"0d",
          4492 => x"0d",
          4493 => x"7f",
          4494 => x"5a",
          4495 => x"a0",
          4496 => x"e7",
          4497 => x"70",
          4498 => x"79",
          4499 => x"73",
          4500 => x"81",
          4501 => x"38",
          4502 => x"33",
          4503 => x"ae",
          4504 => x"70",
          4505 => x"82",
          4506 => x"51",
          4507 => x"54",
          4508 => x"7a",
          4509 => x"74",
          4510 => x"58",
          4511 => x"af",
          4512 => x"77",
          4513 => x"70",
          4514 => x"06",
          4515 => x"51",
          4516 => x"74",
          4517 => x"38",
          4518 => x"a0",
          4519 => x"38",
          4520 => x"0c",
          4521 => x"76",
          4522 => x"a0",
          4523 => x"1c",
          4524 => x"82",
          4525 => x"17",
          4526 => x"19",
          4527 => x"a0",
          4528 => x"8c",
          4529 => x"32",
          4530 => x"80",
          4531 => x"30",
          4532 => x"71",
          4533 => x"53",
          4534 => x"55",
          4535 => x"b5",
          4536 => x"81",
          4537 => x"77",
          4538 => x"51",
          4539 => x"af",
          4540 => x"06",
          4541 => x"5a",
          4542 => x"70",
          4543 => x"55",
          4544 => x"2e",
          4545 => x"83",
          4546 => x"79",
          4547 => x"73",
          4548 => x"bc",
          4549 => x"32",
          4550 => x"80",
          4551 => x"27",
          4552 => x"54",
          4553 => x"a2",
          4554 => x"32",
          4555 => x"ae",
          4556 => x"72",
          4557 => x"9f",
          4558 => x"51",
          4559 => x"74",
          4560 => x"88",
          4561 => x"fe",
          4562 => x"98",
          4563 => x"80",
          4564 => x"75",
          4565 => x"81",
          4566 => x"33",
          4567 => x"51",
          4568 => x"82",
          4569 => x"80",
          4570 => x"78",
          4571 => x"81",
          4572 => x"59",
          4573 => x"d7",
          4574 => x"c8",
          4575 => x"89",
          4576 => x"54",
          4577 => x"86",
          4578 => x"80",
          4579 => x"18",
          4580 => x"34",
          4581 => x"11",
          4582 => x"74",
          4583 => x"58",
          4584 => x"75",
          4585 => x"f0",
          4586 => x"3f",
          4587 => x"08",
          4588 => x"ff",
          4589 => x"73",
          4590 => x"38",
          4591 => x"81",
          4592 => x"54",
          4593 => x"75",
          4594 => x"18",
          4595 => x"39",
          4596 => x"0c",
          4597 => x"80",
          4598 => x"7a",
          4599 => x"81",
          4600 => x"81",
          4601 => x"85",
          4602 => x"54",
          4603 => x"8d",
          4604 => x"86",
          4605 => x"86",
          4606 => x"80",
          4607 => x"1c",
          4608 => x"73",
          4609 => x"0c",
          4610 => x"04",
          4611 => x"78",
          4612 => x"56",
          4613 => x"33",
          4614 => x"72",
          4615 => x"38",
          4616 => x"7a",
          4617 => x"54",
          4618 => x"dc",
          4619 => x"81",
          4620 => x"06",
          4621 => x"2e",
          4622 => x"17",
          4623 => x"0c",
          4624 => x"1a",
          4625 => x"70",
          4626 => x"55",
          4627 => x"09",
          4628 => x"38",
          4629 => x"7a",
          4630 => x"54",
          4631 => x"dc",
          4632 => x"06",
          4633 => x"54",
          4634 => x"53",
          4635 => x"80",
          4636 => x"0c",
          4637 => x"51",
          4638 => x"26",
          4639 => x"80",
          4640 => x"34",
          4641 => x"51",
          4642 => x"82",
          4643 => x"55",
          4644 => x"85",
          4645 => x"39",
          4646 => x"05",
          4647 => x"fb",
          4648 => x"93",
          4649 => x"82",
          4650 => x"81",
          4651 => x"51",
          4652 => x"82",
          4653 => x"ab",
          4654 => x"55",
          4655 => x"08",
          4656 => x"c2",
          4657 => x"c8",
          4658 => x"09",
          4659 => x"ec",
          4660 => x"2a",
          4661 => x"51",
          4662 => x"2e",
          4663 => x"82",
          4664 => x"06",
          4665 => x"80",
          4666 => x"38",
          4667 => x"ab",
          4668 => x"55",
          4669 => x"73",
          4670 => x"81",
          4671 => x"72",
          4672 => x"55",
          4673 => x"82",
          4674 => x"06",
          4675 => x"ac",
          4676 => x"33",
          4677 => x"70",
          4678 => x"54",
          4679 => x"2e",
          4680 => x"90",
          4681 => x"ff",
          4682 => x"05",
          4683 => x"f4",
          4684 => x"93",
          4685 => x"17",
          4686 => x"39",
          4687 => x"c8",
          4688 => x"0d",
          4689 => x"0d",
          4690 => x"79",
          4691 => x"54",
          4692 => x"74",
          4693 => x"d0",
          4694 => x"81",
          4695 => x"70",
          4696 => x"30",
          4697 => x"71",
          4698 => x"51",
          4699 => x"70",
          4700 => x"ba",
          4701 => x"06",
          4702 => x"74",
          4703 => x"52",
          4704 => x"26",
          4705 => x"15",
          4706 => x"06",
          4707 => x"59",
          4708 => x"2e",
          4709 => x"80",
          4710 => x"e8",
          4711 => x"10",
          4712 => x"08",
          4713 => x"57",
          4714 => x"81",
          4715 => x"75",
          4716 => x"57",
          4717 => x"12",
          4718 => x"70",
          4719 => x"38",
          4720 => x"81",
          4721 => x"51",
          4722 => x"51",
          4723 => x"89",
          4724 => x"70",
          4725 => x"54",
          4726 => x"74",
          4727 => x"30",
          4728 => x"80",
          4729 => x"2a",
          4730 => x"53",
          4731 => x"b9",
          4732 => x"75",
          4733 => x"30",
          4734 => x"9f",
          4735 => x"2a",
          4736 => x"53",
          4737 => x"2e",
          4738 => x"18",
          4739 => x"25",
          4740 => x"8b",
          4741 => x"24",
          4742 => x"77",
          4743 => x"79",
          4744 => x"82",
          4745 => x"51",
          4746 => x"c8",
          4747 => x"0d",
          4748 => x"0d",
          4749 => x"0b",
          4750 => x"ff",
          4751 => x"0c",
          4752 => x"51",
          4753 => x"84",
          4754 => x"c8",
          4755 => x"38",
          4756 => x"51",
          4757 => x"82",
          4758 => x"83",
          4759 => x"54",
          4760 => x"82",
          4761 => x"09",
          4762 => x"e7",
          4763 => x"b4",
          4764 => x"55",
          4765 => x"2e",
          4766 => x"83",
          4767 => x"73",
          4768 => x"70",
          4769 => x"25",
          4770 => x"51",
          4771 => x"38",
          4772 => x"54",
          4773 => x"2e",
          4774 => x"b5",
          4775 => x"81",
          4776 => x"80",
          4777 => x"de",
          4778 => x"93",
          4779 => x"82",
          4780 => x"80",
          4781 => x"85",
          4782 => x"84",
          4783 => x"16",
          4784 => x"3f",
          4785 => x"08",
          4786 => x"c8",
          4787 => x"83",
          4788 => x"74",
          4789 => x"0c",
          4790 => x"04",
          4791 => x"60",
          4792 => x"80",
          4793 => x"58",
          4794 => x"0c",
          4795 => x"d5",
          4796 => x"c8",
          4797 => x"56",
          4798 => x"93",
          4799 => x"87",
          4800 => x"93",
          4801 => x"10",
          4802 => x"05",
          4803 => x"53",
          4804 => x"80",
          4805 => x"38",
          4806 => x"76",
          4807 => x"75",
          4808 => x"72",
          4809 => x"38",
          4810 => x"51",
          4811 => x"82",
          4812 => x"81",
          4813 => x"81",
          4814 => x"72",
          4815 => x"80",
          4816 => x"73",
          4817 => x"81",
          4818 => x"8a",
          4819 => x"cf",
          4820 => x"86",
          4821 => x"75",
          4822 => x"16",
          4823 => x"81",
          4824 => x"d6",
          4825 => x"93",
          4826 => x"ff",
          4827 => x"06",
          4828 => x"56",
          4829 => x"38",
          4830 => x"8f",
          4831 => x"2a",
          4832 => x"51",
          4833 => x"72",
          4834 => x"80",
          4835 => x"52",
          4836 => x"3f",
          4837 => x"08",
          4838 => x"57",
          4839 => x"09",
          4840 => x"e4",
          4841 => x"73",
          4842 => x"90",
          4843 => x"10",
          4844 => x"83",
          4845 => x"55",
          4846 => x"57",
          4847 => x"8d",
          4848 => x"16",
          4849 => x"3f",
          4850 => x"08",
          4851 => x"0c",
          4852 => x"83",
          4853 => x"38",
          4854 => x"3d",
          4855 => x"05",
          4856 => x"5b",
          4857 => x"79",
          4858 => x"38",
          4859 => x"51",
          4860 => x"82",
          4861 => x"81",
          4862 => x"81",
          4863 => x"38",
          4864 => x"83",
          4865 => x"38",
          4866 => x"84",
          4867 => x"38",
          4868 => x"81",
          4869 => x"38",
          4870 => x"d9",
          4871 => x"93",
          4872 => x"ff",
          4873 => x"8d",
          4874 => x"80",
          4875 => x"06",
          4876 => x"80",
          4877 => x"d9",
          4878 => x"93",
          4879 => x"ff",
          4880 => x"73",
          4881 => x"d8",
          4882 => x"e6",
          4883 => x"c8",
          4884 => x"9c",
          4885 => x"c4",
          4886 => x"16",
          4887 => x"15",
          4888 => x"53",
          4889 => x"81",
          4890 => x"38",
          4891 => x"74",
          4892 => x"c1",
          4893 => x"55",
          4894 => x"16",
          4895 => x"ff",
          4896 => x"72",
          4897 => x"38",
          4898 => x"06",
          4899 => x"2e",
          4900 => x"56",
          4901 => x"80",
          4902 => x"d8",
          4903 => x"93",
          4904 => x"16",
          4905 => x"c8",
          4906 => x"ff",
          4907 => x"53",
          4908 => x"83",
          4909 => x"c7",
          4910 => x"dd",
          4911 => x"c8",
          4912 => x"ff",
          4913 => x"8d",
          4914 => x"15",
          4915 => x"3f",
          4916 => x"08",
          4917 => x"15",
          4918 => x"3f",
          4919 => x"08",
          4920 => x"06",
          4921 => x"78",
          4922 => x"b3",
          4923 => x"22",
          4924 => x"84",
          4925 => x"56",
          4926 => x"73",
          4927 => x"38",
          4928 => x"52",
          4929 => x"51",
          4930 => x"3f",
          4931 => x"08",
          4932 => x"82",
          4933 => x"80",
          4934 => x"38",
          4935 => x"93",
          4936 => x"ff",
          4937 => x"26",
          4938 => x"57",
          4939 => x"f5",
          4940 => x"82",
          4941 => x"f5",
          4942 => x"81",
          4943 => x"76",
          4944 => x"db",
          4945 => x"98",
          4946 => x"a0",
          4947 => x"19",
          4948 => x"77",
          4949 => x"0c",
          4950 => x"09",
          4951 => x"38",
          4952 => x"51",
          4953 => x"82",
          4954 => x"83",
          4955 => x"53",
          4956 => x"82",
          4957 => x"15",
          4958 => x"56",
          4959 => x"38",
          4960 => x"51",
          4961 => x"82",
          4962 => x"a8",
          4963 => x"15",
          4964 => x"53",
          4965 => x"15",
          4966 => x"56",
          4967 => x"81",
          4968 => x"15",
          4969 => x"16",
          4970 => x"2e",
          4971 => x"88",
          4972 => x"08",
          4973 => x"39",
          4974 => x"10",
          4975 => x"05",
          4976 => x"98",
          4977 => x"06",
          4978 => x"83",
          4979 => x"2a",
          4980 => x"72",
          4981 => x"26",
          4982 => x"ff",
          4983 => x"0c",
          4984 => x"16",
          4985 => x"0b",
          4986 => x"76",
          4987 => x"81",
          4988 => x"38",
          4989 => x"51",
          4990 => x"82",
          4991 => x"83",
          4992 => x"53",
          4993 => x"09",
          4994 => x"f9",
          4995 => x"52",
          4996 => x"b3",
          4997 => x"c8",
          4998 => x"38",
          4999 => x"08",
          5000 => x"84",
          5001 => x"d5",
          5002 => x"93",
          5003 => x"ff",
          5004 => x"72",
          5005 => x"2e",
          5006 => x"80",
          5007 => x"15",
          5008 => x"3f",
          5009 => x"08",
          5010 => x"a4",
          5011 => x"81",
          5012 => x"84",
          5013 => x"d5",
          5014 => x"93",
          5015 => x"8a",
          5016 => x"2e",
          5017 => x"9d",
          5018 => x"15",
          5019 => x"3f",
          5020 => x"08",
          5021 => x"84",
          5022 => x"d5",
          5023 => x"93",
          5024 => x"16",
          5025 => x"34",
          5026 => x"22",
          5027 => x"72",
          5028 => x"23",
          5029 => x"23",
          5030 => x"16",
          5031 => x"75",
          5032 => x"0c",
          5033 => x"04",
          5034 => x"77",
          5035 => x"73",
          5036 => x"38",
          5037 => x"2e",
          5038 => x"08",
          5039 => x"53",
          5040 => x"a4",
          5041 => x"22",
          5042 => x"57",
          5043 => x"2e",
          5044 => x"94",
          5045 => x"33",
          5046 => x"3f",
          5047 => x"08",
          5048 => x"71",
          5049 => x"55",
          5050 => x"73",
          5051 => x"06",
          5052 => x"08",
          5053 => x"71",
          5054 => x"82",
          5055 => x"87",
          5056 => x"fa",
          5057 => x"ab",
          5058 => x"58",
          5059 => x"05",
          5060 => x"b1",
          5061 => x"c8",
          5062 => x"54",
          5063 => x"93",
          5064 => x"80",
          5065 => x"93",
          5066 => x"10",
          5067 => x"05",
          5068 => x"54",
          5069 => x"84",
          5070 => x"34",
          5071 => x"86",
          5072 => x"80",
          5073 => x"10",
          5074 => x"e4",
          5075 => x"0c",
          5076 => x"75",
          5077 => x"38",
          5078 => x"3d",
          5079 => x"05",
          5080 => x"3f",
          5081 => x"08",
          5082 => x"93",
          5083 => x"3d",
          5084 => x"3d",
          5085 => x"84",
          5086 => x"05",
          5087 => x"89",
          5088 => x"2e",
          5089 => x"76",
          5090 => x"54",
          5091 => x"05",
          5092 => x"84",
          5093 => x"f6",
          5094 => x"93",
          5095 => x"82",
          5096 => x"84",
          5097 => x"5c",
          5098 => x"3d",
          5099 => x"f0",
          5100 => x"93",
          5101 => x"82",
          5102 => x"92",
          5103 => x"d7",
          5104 => x"98",
          5105 => x"74",
          5106 => x"38",
          5107 => x"9c",
          5108 => x"80",
          5109 => x"38",
          5110 => x"9c",
          5111 => x"2e",
          5112 => x"8e",
          5113 => x"d4",
          5114 => x"9e",
          5115 => x"c8",
          5116 => x"88",
          5117 => x"39",
          5118 => x"33",
          5119 => x"74",
          5120 => x"38",
          5121 => x"39",
          5122 => x"70",
          5123 => x"55",
          5124 => x"83",
          5125 => x"75",
          5126 => x"76",
          5127 => x"81",
          5128 => x"74",
          5129 => x"a7",
          5130 => x"7a",
          5131 => x"3f",
          5132 => x"08",
          5133 => x"b2",
          5134 => x"8e",
          5135 => x"b9",
          5136 => x"a0",
          5137 => x"34",
          5138 => x"52",
          5139 => x"ce",
          5140 => x"62",
          5141 => x"d2",
          5142 => x"55",
          5143 => x"16",
          5144 => x"2e",
          5145 => x"7a",
          5146 => x"77",
          5147 => x"99",
          5148 => x"53",
          5149 => x"b3",
          5150 => x"c8",
          5151 => x"93",
          5152 => x"e6",
          5153 => x"7a",
          5154 => x"3f",
          5155 => x"08",
          5156 => x"8c",
          5157 => x"56",
          5158 => x"82",
          5159 => x"b2",
          5160 => x"84",
          5161 => x"06",
          5162 => x"74",
          5163 => x"38",
          5164 => x"39",
          5165 => x"70",
          5166 => x"55",
          5167 => x"8f",
          5168 => x"05",
          5169 => x"55",
          5170 => x"83",
          5171 => x"75",
          5172 => x"76",
          5173 => x"81",
          5174 => x"74",
          5175 => x"38",
          5176 => x"07",
          5177 => x"11",
          5178 => x"0c",
          5179 => x"0c",
          5180 => x"f6",
          5181 => x"74",
          5182 => x"3f",
          5183 => x"08",
          5184 => x"62",
          5185 => x"d0",
          5186 => x"93",
          5187 => x"19",
          5188 => x"0c",
          5189 => x"84",
          5190 => x"90",
          5191 => x"91",
          5192 => x"9c",
          5193 => x"94",
          5194 => x"80",
          5195 => x"a8",
          5196 => x"98",
          5197 => x"2a",
          5198 => x"51",
          5199 => x"2e",
          5200 => x"8c",
          5201 => x"2e",
          5202 => x"8c",
          5203 => x"19",
          5204 => x"11",
          5205 => x"2b",
          5206 => x"8c",
          5207 => x"5a",
          5208 => x"a5",
          5209 => x"77",
          5210 => x"3f",
          5211 => x"08",
          5212 => x"c8",
          5213 => x"83",
          5214 => x"76",
          5215 => x"81",
          5216 => x"81",
          5217 => x"31",
          5218 => x"70",
          5219 => x"25",
          5220 => x"26",
          5221 => x"55",
          5222 => x"76",
          5223 => x"75",
          5224 => x"78",
          5225 => x"55",
          5226 => x"b9",
          5227 => x"7a",
          5228 => x"3f",
          5229 => x"08",
          5230 => x"56",
          5231 => x"89",
          5232 => x"c8",
          5233 => x"9c",
          5234 => x"81",
          5235 => x"a8",
          5236 => x"81",
          5237 => x"55",
          5238 => x"82",
          5239 => x"80",
          5240 => x"81",
          5241 => x"2e",
          5242 => x"78",
          5243 => x"74",
          5244 => x"0c",
          5245 => x"04",
          5246 => x"7f",
          5247 => x"5f",
          5248 => x"80",
          5249 => x"3d",
          5250 => x"76",
          5251 => x"3f",
          5252 => x"08",
          5253 => x"c8",
          5254 => x"91",
          5255 => x"74",
          5256 => x"38",
          5257 => x"ae",
          5258 => x"33",
          5259 => x"87",
          5260 => x"2e",
          5261 => x"bd",
          5262 => x"91",
          5263 => x"56",
          5264 => x"81",
          5265 => x"34",
          5266 => x"8a",
          5267 => x"91",
          5268 => x"56",
          5269 => x"81",
          5270 => x"34",
          5271 => x"f6",
          5272 => x"91",
          5273 => x"56",
          5274 => x"81",
          5275 => x"34",
          5276 => x"e2",
          5277 => x"08",
          5278 => x"31",
          5279 => x"27",
          5280 => x"59",
          5281 => x"82",
          5282 => x"17",
          5283 => x"ff",
          5284 => x"74",
          5285 => x"7d",
          5286 => x"ff",
          5287 => x"2a",
          5288 => x"7a",
          5289 => x"87",
          5290 => x"08",
          5291 => x"98",
          5292 => x"76",
          5293 => x"3f",
          5294 => x"08",
          5295 => x"27",
          5296 => x"74",
          5297 => x"fb",
          5298 => x"18",
          5299 => x"08",
          5300 => x"d1",
          5301 => x"93",
          5302 => x"2e",
          5303 => x"82",
          5304 => x"1b",
          5305 => x"5b",
          5306 => x"2e",
          5307 => x"79",
          5308 => x"11",
          5309 => x"56",
          5310 => x"85",
          5311 => x"31",
          5312 => x"77",
          5313 => x"7d",
          5314 => x"52",
          5315 => x"3f",
          5316 => x"08",
          5317 => x"90",
          5318 => x"98",
          5319 => x"74",
          5320 => x"38",
          5321 => x"78",
          5322 => x"7a",
          5323 => x"84",
          5324 => x"17",
          5325 => x"80",
          5326 => x"cc",
          5327 => x"89",
          5328 => x"f9",
          5329 => x"08",
          5330 => x"c9",
          5331 => x"33",
          5332 => x"56",
          5333 => x"25",
          5334 => x"54",
          5335 => x"53",
          5336 => x"7d",
          5337 => x"52",
          5338 => x"3f",
          5339 => x"08",
          5340 => x"90",
          5341 => x"ff",
          5342 => x"90",
          5343 => x"54",
          5344 => x"17",
          5345 => x"11",
          5346 => x"c6",
          5347 => x"93",
          5348 => x"d7",
          5349 => x"18",
          5350 => x"08",
          5351 => x"84",
          5352 => x"57",
          5353 => x"27",
          5354 => x"56",
          5355 => x"17",
          5356 => x"06",
          5357 => x"52",
          5358 => x"ec",
          5359 => x"31",
          5360 => x"7e",
          5361 => x"94",
          5362 => x"94",
          5363 => x"59",
          5364 => x"38",
          5365 => x"82",
          5366 => x"8f",
          5367 => x"f3",
          5368 => x"62",
          5369 => x"5f",
          5370 => x"7d",
          5371 => x"fc",
          5372 => x"51",
          5373 => x"82",
          5374 => x"55",
          5375 => x"08",
          5376 => x"17",
          5377 => x"80",
          5378 => x"74",
          5379 => x"39",
          5380 => x"70",
          5381 => x"81",
          5382 => x"56",
          5383 => x"80",
          5384 => x"38",
          5385 => x"0b",
          5386 => x"82",
          5387 => x"39",
          5388 => x"18",
          5389 => x"83",
          5390 => x"0b",
          5391 => x"81",
          5392 => x"39",
          5393 => x"18",
          5394 => x"83",
          5395 => x"0b",
          5396 => x"81",
          5397 => x"39",
          5398 => x"18",
          5399 => x"83",
          5400 => x"17",
          5401 => x"74",
          5402 => x"27",
          5403 => x"17",
          5404 => x"78",
          5405 => x"8c",
          5406 => x"08",
          5407 => x"06",
          5408 => x"82",
          5409 => x"8a",
          5410 => x"05",
          5411 => x"06",
          5412 => x"80",
          5413 => x"96",
          5414 => x"08",
          5415 => x"38",
          5416 => x"51",
          5417 => x"82",
          5418 => x"55",
          5419 => x"17",
          5420 => x"51",
          5421 => x"82",
          5422 => x"55",
          5423 => x"82",
          5424 => x"81",
          5425 => x"38",
          5426 => x"fe",
          5427 => x"98",
          5428 => x"17",
          5429 => x"74",
          5430 => x"90",
          5431 => x"98",
          5432 => x"74",
          5433 => x"38",
          5434 => x"17",
          5435 => x"17",
          5436 => x"11",
          5437 => x"c5",
          5438 => x"93",
          5439 => x"ba",
          5440 => x"33",
          5441 => x"55",
          5442 => x"34",
          5443 => x"52",
          5444 => x"a9",
          5445 => x"c8",
          5446 => x"fe",
          5447 => x"93",
          5448 => x"79",
          5449 => x"58",
          5450 => x"80",
          5451 => x"1b",
          5452 => x"22",
          5453 => x"74",
          5454 => x"38",
          5455 => x"5a",
          5456 => x"53",
          5457 => x"81",
          5458 => x"55",
          5459 => x"82",
          5460 => x"fd",
          5461 => x"17",
          5462 => x"55",
          5463 => x"9b",
          5464 => x"53",
          5465 => x"29",
          5466 => x"17",
          5467 => x"3f",
          5468 => x"80",
          5469 => x"74",
          5470 => x"79",
          5471 => x"80",
          5472 => x"17",
          5473 => x"a1",
          5474 => x"08",
          5475 => x"27",
          5476 => x"54",
          5477 => x"17",
          5478 => x"11",
          5479 => x"c2",
          5480 => x"93",
          5481 => x"b0",
          5482 => x"18",
          5483 => x"08",
          5484 => x"84",
          5485 => x"57",
          5486 => x"27",
          5487 => x"56",
          5488 => x"52",
          5489 => x"83",
          5490 => x"a8",
          5491 => x"d8",
          5492 => x"33",
          5493 => x"55",
          5494 => x"34",
          5495 => x"7d",
          5496 => x"0c",
          5497 => x"19",
          5498 => x"94",
          5499 => x"1a",
          5500 => x"5d",
          5501 => x"27",
          5502 => x"55",
          5503 => x"0c",
          5504 => x"38",
          5505 => x"80",
          5506 => x"74",
          5507 => x"80",
          5508 => x"93",
          5509 => x"3d",
          5510 => x"3d",
          5511 => x"3d",
          5512 => x"70",
          5513 => x"80",
          5514 => x"c8",
          5515 => x"93",
          5516 => x"aa",
          5517 => x"33",
          5518 => x"70",
          5519 => x"56",
          5520 => x"2e",
          5521 => x"75",
          5522 => x"74",
          5523 => x"38",
          5524 => x"18",
          5525 => x"18",
          5526 => x"11",
          5527 => x"c2",
          5528 => x"55",
          5529 => x"08",
          5530 => x"90",
          5531 => x"ff",
          5532 => x"90",
          5533 => x"18",
          5534 => x"51",
          5535 => x"82",
          5536 => x"57",
          5537 => x"08",
          5538 => x"a4",
          5539 => x"11",
          5540 => x"56",
          5541 => x"17",
          5542 => x"08",
          5543 => x"77",
          5544 => x"fa",
          5545 => x"08",
          5546 => x"51",
          5547 => x"82",
          5548 => x"52",
          5549 => x"c5",
          5550 => x"52",
          5551 => x"c5",
          5552 => x"55",
          5553 => x"16",
          5554 => x"c8",
          5555 => x"93",
          5556 => x"19",
          5557 => x"06",
          5558 => x"90",
          5559 => x"55",
          5560 => x"c8",
          5561 => x"0d",
          5562 => x"0d",
          5563 => x"54",
          5564 => x"82",
          5565 => x"53",
          5566 => x"08",
          5567 => x"3d",
          5568 => x"73",
          5569 => x"3f",
          5570 => x"08",
          5571 => x"c8",
          5572 => x"82",
          5573 => x"74",
          5574 => x"93",
          5575 => x"3d",
          5576 => x"3d",
          5577 => x"51",
          5578 => x"8b",
          5579 => x"82",
          5580 => x"24",
          5581 => x"93",
          5582 => x"93",
          5583 => x"53",
          5584 => x"c8",
          5585 => x"0d",
          5586 => x"0d",
          5587 => x"3d",
          5588 => x"94",
          5589 => x"84",
          5590 => x"c8",
          5591 => x"93",
          5592 => x"df",
          5593 => x"63",
          5594 => x"d4",
          5595 => x"9c",
          5596 => x"c8",
          5597 => x"93",
          5598 => x"38",
          5599 => x"05",
          5600 => x"2b",
          5601 => x"80",
          5602 => x"76",
          5603 => x"0c",
          5604 => x"02",
          5605 => x"70",
          5606 => x"81",
          5607 => x"56",
          5608 => x"93",
          5609 => x"53",
          5610 => x"d7",
          5611 => x"93",
          5612 => x"15",
          5613 => x"85",
          5614 => x"2e",
          5615 => x"83",
          5616 => x"74",
          5617 => x"0c",
          5618 => x"04",
          5619 => x"a3",
          5620 => x"3d",
          5621 => x"80",
          5622 => x"53",
          5623 => x"b8",
          5624 => x"3d",
          5625 => x"3f",
          5626 => x"08",
          5627 => x"c8",
          5628 => x"38",
          5629 => x"7f",
          5630 => x"4a",
          5631 => x"59",
          5632 => x"81",
          5633 => x"3d",
          5634 => x"40",
          5635 => x"52",
          5636 => x"e4",
          5637 => x"c8",
          5638 => x"93",
          5639 => x"de",
          5640 => x"7e",
          5641 => x"3f",
          5642 => x"08",
          5643 => x"c8",
          5644 => x"38",
          5645 => x"51",
          5646 => x"82",
          5647 => x"48",
          5648 => x"51",
          5649 => x"82",
          5650 => x"57",
          5651 => x"08",
          5652 => x"7c",
          5653 => x"73",
          5654 => x"3f",
          5655 => x"08",
          5656 => x"c8",
          5657 => x"6c",
          5658 => x"d5",
          5659 => x"93",
          5660 => x"2e",
          5661 => x"52",
          5662 => x"d1",
          5663 => x"c8",
          5664 => x"93",
          5665 => x"2e",
          5666 => x"84",
          5667 => x"06",
          5668 => x"57",
          5669 => x"38",
          5670 => x"bc",
          5671 => x"05",
          5672 => x"3f",
          5673 => x"70",
          5674 => x"11",
          5675 => x"57",
          5676 => x"80",
          5677 => x"81",
          5678 => x"81",
          5679 => x"55",
          5680 => x"38",
          5681 => x"78",
          5682 => x"38",
          5683 => x"39",
          5684 => x"99",
          5685 => x"ff",
          5686 => x"08",
          5687 => x"70",
          5688 => x"56",
          5689 => x"33",
          5690 => x"eb",
          5691 => x"a3",
          5692 => x"55",
          5693 => x"34",
          5694 => x"fe",
          5695 => x"81",
          5696 => x"7c",
          5697 => x"06",
          5698 => x"19",
          5699 => x"11",
          5700 => x"74",
          5701 => x"82",
          5702 => x"70",
          5703 => x"fb",
          5704 => x"08",
          5705 => x"52",
          5706 => x"58",
          5707 => x"8d",
          5708 => x"70",
          5709 => x"51",
          5710 => x"f5",
          5711 => x"54",
          5712 => x"a5",
          5713 => x"77",
          5714 => x"38",
          5715 => x"73",
          5716 => x"81",
          5717 => x"81",
          5718 => x"78",
          5719 => x"ba",
          5720 => x"05",
          5721 => x"18",
          5722 => x"38",
          5723 => x"96",
          5724 => x"08",
          5725 => x"5a",
          5726 => x"7a",
          5727 => x"5c",
          5728 => x"26",
          5729 => x"7a",
          5730 => x"93",
          5731 => x"3d",
          5732 => x"3d",
          5733 => x"90",
          5734 => x"54",
          5735 => x"57",
          5736 => x"82",
          5737 => x"5a",
          5738 => x"08",
          5739 => x"17",
          5740 => x"80",
          5741 => x"79",
          5742 => x"39",
          5743 => x"78",
          5744 => x"90",
          5745 => x"81",
          5746 => x"06",
          5747 => x"74",
          5748 => x"17",
          5749 => x"17",
          5750 => x"70",
          5751 => x"5b",
          5752 => x"82",
          5753 => x"8a",
          5754 => x"89",
          5755 => x"55",
          5756 => x"b6",
          5757 => x"ff",
          5758 => x"96",
          5759 => x"93",
          5760 => x"17",
          5761 => x"53",
          5762 => x"96",
          5763 => x"93",
          5764 => x"26",
          5765 => x"30",
          5766 => x"18",
          5767 => x"18",
          5768 => x"18",
          5769 => x"80",
          5770 => x"17",
          5771 => x"be",
          5772 => x"76",
          5773 => x"3f",
          5774 => x"08",
          5775 => x"c8",
          5776 => x"09",
          5777 => x"38",
          5778 => x"18",
          5779 => x"82",
          5780 => x"93",
          5781 => x"2e",
          5782 => x"8b",
          5783 => x"91",
          5784 => x"55",
          5785 => x"82",
          5786 => x"88",
          5787 => x"98",
          5788 => x"80",
          5789 => x"38",
          5790 => x"80",
          5791 => x"79",
          5792 => x"08",
          5793 => x"0c",
          5794 => x"70",
          5795 => x"81",
          5796 => x"5d",
          5797 => x"2e",
          5798 => x"52",
          5799 => x"be",
          5800 => x"c8",
          5801 => x"93",
          5802 => x"38",
          5803 => x"08",
          5804 => x"75",
          5805 => x"c2",
          5806 => x"93",
          5807 => x"75",
          5808 => x"e1",
          5809 => x"27",
          5810 => x"55",
          5811 => x"76",
          5812 => x"82",
          5813 => x"34",
          5814 => x"d8",
          5815 => x"18",
          5816 => x"26",
          5817 => x"94",
          5818 => x"94",
          5819 => x"83",
          5820 => x"74",
          5821 => x"38",
          5822 => x"51",
          5823 => x"82",
          5824 => x"8b",
          5825 => x"91",
          5826 => x"55",
          5827 => x"77",
          5828 => x"93",
          5829 => x"5b",
          5830 => x"94",
          5831 => x"92",
          5832 => x"08",
          5833 => x"90",
          5834 => x"c0",
          5835 => x"90",
          5836 => x"17",
          5837 => x"06",
          5838 => x"2e",
          5839 => x"9c",
          5840 => x"2e",
          5841 => x"90",
          5842 => x"98",
          5843 => x"74",
          5844 => x"38",
          5845 => x"17",
          5846 => x"17",
          5847 => x"11",
          5848 => x"ff",
          5849 => x"82",
          5850 => x"80",
          5851 => x"81",
          5852 => x"34",
          5853 => x"39",
          5854 => x"80",
          5855 => x"74",
          5856 => x"81",
          5857 => x"a8",
          5858 => x"81",
          5859 => x"55",
          5860 => x"3f",
          5861 => x"08",
          5862 => x"38",
          5863 => x"18",
          5864 => x"90",
          5865 => x"91",
          5866 => x"55",
          5867 => x"9c",
          5868 => x"55",
          5869 => x"c8",
          5870 => x"0d",
          5871 => x"0d",
          5872 => x"54",
          5873 => x"81",
          5874 => x"53",
          5875 => x"05",
          5876 => x"84",
          5877 => x"84",
          5878 => x"c8",
          5879 => x"93",
          5880 => x"ef",
          5881 => x"0c",
          5882 => x"51",
          5883 => x"82",
          5884 => x"55",
          5885 => x"08",
          5886 => x"ab",
          5887 => x"98",
          5888 => x"80",
          5889 => x"38",
          5890 => x"70",
          5891 => x"81",
          5892 => x"57",
          5893 => x"93",
          5894 => x"08",
          5895 => x"ce",
          5896 => x"93",
          5897 => x"17",
          5898 => x"85",
          5899 => x"38",
          5900 => x"14",
          5901 => x"23",
          5902 => x"51",
          5903 => x"82",
          5904 => x"55",
          5905 => x"09",
          5906 => x"38",
          5907 => x"80",
          5908 => x"80",
          5909 => x"54",
          5910 => x"c8",
          5911 => x"0d",
          5912 => x"0d",
          5913 => x"fc",
          5914 => x"52",
          5915 => x"3f",
          5916 => x"08",
          5917 => x"c8",
          5918 => x"82",
          5919 => x"74",
          5920 => x"93",
          5921 => x"3d",
          5922 => x"3d",
          5923 => x"89",
          5924 => x"54",
          5925 => x"54",
          5926 => x"82",
          5927 => x"53",
          5928 => x"08",
          5929 => x"74",
          5930 => x"93",
          5931 => x"73",
          5932 => x"3f",
          5933 => x"08",
          5934 => x"80",
          5935 => x"ce",
          5936 => x"93",
          5937 => x"82",
          5938 => x"84",
          5939 => x"06",
          5940 => x"53",
          5941 => x"74",
          5942 => x"d1",
          5943 => x"52",
          5944 => x"e9",
          5945 => x"c8",
          5946 => x"93",
          5947 => x"2e",
          5948 => x"83",
          5949 => x"72",
          5950 => x"0c",
          5951 => x"04",
          5952 => x"64",
          5953 => x"88",
          5954 => x"95",
          5955 => x"db",
          5956 => x"93",
          5957 => x"82",
          5958 => x"b5",
          5959 => x"73",
          5960 => x"3f",
          5961 => x"08",
          5962 => x"c8",
          5963 => x"02",
          5964 => x"33",
          5965 => x"55",
          5966 => x"25",
          5967 => x"55",
          5968 => x"80",
          5969 => x"75",
          5970 => x"d4",
          5971 => x"c1",
          5972 => x"93",
          5973 => x"3d",
          5974 => x"3d",
          5975 => x"55",
          5976 => x"90",
          5977 => x"52",
          5978 => x"da",
          5979 => x"93",
          5980 => x"82",
          5981 => x"82",
          5982 => x"74",
          5983 => x"98",
          5984 => x"05",
          5985 => x"15",
          5986 => x"93",
          5987 => x"08",
          5988 => x"e9",
          5989 => x"81",
          5990 => x"59",
          5991 => x"80",
          5992 => x"56",
          5993 => x"81",
          5994 => x"06",
          5995 => x"82",
          5996 => x"75",
          5997 => x"f0",
          5998 => x"bc",
          5999 => x"93",
          6000 => x"2e",
          6001 => x"93",
          6002 => x"2e",
          6003 => x"93",
          6004 => x"70",
          6005 => x"08",
          6006 => x"78",
          6007 => x"7d",
          6008 => x"54",
          6009 => x"76",
          6010 => x"80",
          6011 => x"98",
          6012 => x"12",
          6013 => x"54",
          6014 => x"98",
          6015 => x"81",
          6016 => x"58",
          6017 => x"3f",
          6018 => x"08",
          6019 => x"c8",
          6020 => x"38",
          6021 => x"51",
          6022 => x"2e",
          6023 => x"a0",
          6024 => x"b4",
          6025 => x"b5",
          6026 => x"93",
          6027 => x"ff",
          6028 => x"30",
          6029 => x"19",
          6030 => x"59",
          6031 => x"39",
          6032 => x"05",
          6033 => x"ea",
          6034 => x"c8",
          6035 => x"06",
          6036 => x"80",
          6037 => x"18",
          6038 => x"54",
          6039 => x"06",
          6040 => x"55",
          6041 => x"38",
          6042 => x"7a",
          6043 => x"0c",
          6044 => x"11",
          6045 => x"55",
          6046 => x"16",
          6047 => x"93",
          6048 => x"3d",
          6049 => x"3d",
          6050 => x"3d",
          6051 => x"70",
          6052 => x"94",
          6053 => x"c8",
          6054 => x"93",
          6055 => x"38",
          6056 => x"57",
          6057 => x"86",
          6058 => x"81",
          6059 => x"18",
          6060 => x"2a",
          6061 => x"51",
          6062 => x"56",
          6063 => x"81",
          6064 => x"18",
          6065 => x"08",
          6066 => x"38",
          6067 => x"9a",
          6068 => x"88",
          6069 => x"77",
          6070 => x"cf",
          6071 => x"c8",
          6072 => x"0b",
          6073 => x"80",
          6074 => x"18",
          6075 => x"51",
          6076 => x"3f",
          6077 => x"08",
          6078 => x"08",
          6079 => x"30",
          6080 => x"80",
          6081 => x"58",
          6082 => x"c8",
          6083 => x"09",
          6084 => x"38",
          6085 => x"9b",
          6086 => x"75",
          6087 => x"27",
          6088 => x"18",
          6089 => x"52",
          6090 => x"bd",
          6091 => x"93",
          6092 => x"94",
          6093 => x"19",
          6094 => x"33",
          6095 => x"55",
          6096 => x"34",
          6097 => x"74",
          6098 => x"74",
          6099 => x"38",
          6100 => x"18",
          6101 => x"18",
          6102 => x"11",
          6103 => x"ff",
          6104 => x"82",
          6105 => x"80",
          6106 => x"81",
          6107 => x"90",
          6108 => x"ff",
          6109 => x"90",
          6110 => x"80",
          6111 => x"76",
          6112 => x"76",
          6113 => x"76",
          6114 => x"93",
          6115 => x"3d",
          6116 => x"3d",
          6117 => x"8c",
          6118 => x"d5",
          6119 => x"9f",
          6120 => x"05",
          6121 => x"51",
          6122 => x"82",
          6123 => x"56",
          6124 => x"08",
          6125 => x"81",
          6126 => x"ff",
          6127 => x"77",
          6128 => x"9f",
          6129 => x"51",
          6130 => x"82",
          6131 => x"81",
          6132 => x"56",
          6133 => x"3f",
          6134 => x"38",
          6135 => x"05",
          6136 => x"2a",
          6137 => x"51",
          6138 => x"80",
          6139 => x"86",
          6140 => x"95",
          6141 => x"98",
          6142 => x"f5",
          6143 => x"f7",
          6144 => x"98",
          6145 => x"73",
          6146 => x"38",
          6147 => x"39",
          6148 => x"05",
          6149 => x"54",
          6150 => x"83",
          6151 => x"75",
          6152 => x"6a",
          6153 => x"c6",
          6154 => x"93",
          6155 => x"84",
          6156 => x"05",
          6157 => x"2a",
          6158 => x"51",
          6159 => x"73",
          6160 => x"e5",
          6161 => x"9c",
          6162 => x"a5",
          6163 => x"55",
          6164 => x"08",
          6165 => x"d1",
          6166 => x"a0",
          6167 => x"91",
          6168 => x"76",
          6169 => x"a4",
          6170 => x"85",
          6171 => x"89",
          6172 => x"54",
          6173 => x"82",
          6174 => x"56",
          6175 => x"08",
          6176 => x"82",
          6177 => x"52",
          6178 => x"c0",
          6179 => x"c8",
          6180 => x"93",
          6181 => x"38",
          6182 => x"84",
          6183 => x"70",
          6184 => x"2c",
          6185 => x"56",
          6186 => x"dd",
          6187 => x"a8",
          6188 => x"bd",
          6189 => x"d4",
          6190 => x"a4",
          6191 => x"c8",
          6192 => x"c8",
          6193 => x"82",
          6194 => x"07",
          6195 => x"30",
          6196 => x"9f",
          6197 => x"52",
          6198 => x"56",
          6199 => x"9b",
          6200 => x"ac",
          6201 => x"89",
          6202 => x"76",
          6203 => x"d4",
          6204 => x"ba",
          6205 => x"93",
          6206 => x"75",
          6207 => x"51",
          6208 => x"3f",
          6209 => x"08",
          6210 => x"b0",
          6211 => x"e1",
          6212 => x"93",
          6213 => x"3d",
          6214 => x"3d",
          6215 => x"98",
          6216 => x"52",
          6217 => x"d3",
          6218 => x"93",
          6219 => x"82",
          6220 => x"82",
          6221 => x"5d",
          6222 => x"3d",
          6223 => x"cd",
          6224 => x"93",
          6225 => x"82",
          6226 => x"83",
          6227 => x"74",
          6228 => x"81",
          6229 => x"38",
          6230 => x"05",
          6231 => x"2a",
          6232 => x"51",
          6233 => x"80",
          6234 => x"86",
          6235 => x"2e",
          6236 => x"81",
          6237 => x"59",
          6238 => x"3d",
          6239 => x"ff",
          6240 => x"82",
          6241 => x"56",
          6242 => x"93",
          6243 => x"2e",
          6244 => x"83",
          6245 => x"75",
          6246 => x"81",
          6247 => x"82",
          6248 => x"2e",
          6249 => x"83",
          6250 => x"82",
          6251 => x"57",
          6252 => x"38",
          6253 => x"51",
          6254 => x"3f",
          6255 => x"08",
          6256 => x"c8",
          6257 => x"38",
          6258 => x"52",
          6259 => x"ff",
          6260 => x"77",
          6261 => x"b4",
          6262 => x"54",
          6263 => x"15",
          6264 => x"80",
          6265 => x"ff",
          6266 => x"75",
          6267 => x"52",
          6268 => x"aa",
          6269 => x"b4",
          6270 => x"d4",
          6271 => x"af",
          6272 => x"54",
          6273 => x"d5",
          6274 => x"53",
          6275 => x"52",
          6276 => x"8a",
          6277 => x"81",
          6278 => x"34",
          6279 => x"05",
          6280 => x"3f",
          6281 => x"08",
          6282 => x"c8",
          6283 => x"76",
          6284 => x"05",
          6285 => x"c1",
          6286 => x"63",
          6287 => x"c2",
          6288 => x"54",
          6289 => x"15",
          6290 => x"81",
          6291 => x"34",
          6292 => x"b1",
          6293 => x"93",
          6294 => x"8e",
          6295 => x"75",
          6296 => x"c4",
          6297 => x"b7",
          6298 => x"82",
          6299 => x"98",
          6300 => x"db",
          6301 => x"3d",
          6302 => x"cd",
          6303 => x"53",
          6304 => x"84",
          6305 => x"3d",
          6306 => x"3f",
          6307 => x"08",
          6308 => x"c8",
          6309 => x"38",
          6310 => x"3d",
          6311 => x"3d",
          6312 => x"ca",
          6313 => x"93",
          6314 => x"82",
          6315 => x"82",
          6316 => x"81",
          6317 => x"81",
          6318 => x"73",
          6319 => x"38",
          6320 => x"82",
          6321 => x"53",
          6322 => x"52",
          6323 => x"88",
          6324 => x"ad",
          6325 => x"53",
          6326 => x"05",
          6327 => x"70",
          6328 => x"ad",
          6329 => x"3d",
          6330 => x"51",
          6331 => x"82",
          6332 => x"55",
          6333 => x"08",
          6334 => x"6e",
          6335 => x"06",
          6336 => x"55",
          6337 => x"08",
          6338 => x"88",
          6339 => x"2e",
          6340 => x"81",
          6341 => x"3d",
          6342 => x"51",
          6343 => x"82",
          6344 => x"55",
          6345 => x"08",
          6346 => x"67",
          6347 => x"a7",
          6348 => x"05",
          6349 => x"51",
          6350 => x"3f",
          6351 => x"33",
          6352 => x"8b",
          6353 => x"84",
          6354 => x"06",
          6355 => x"73",
          6356 => x"a0",
          6357 => x"8b",
          6358 => x"54",
          6359 => x"15",
          6360 => x"33",
          6361 => x"70",
          6362 => x"55",
          6363 => x"2e",
          6364 => x"6d",
          6365 => x"d5",
          6366 => x"77",
          6367 => x"e5",
          6368 => x"c8",
          6369 => x"51",
          6370 => x"3f",
          6371 => x"93",
          6372 => x"2e",
          6373 => x"93",
          6374 => x"77",
          6375 => x"a7",
          6376 => x"c8",
          6377 => x"19",
          6378 => x"93",
          6379 => x"38",
          6380 => x"54",
          6381 => x"09",
          6382 => x"38",
          6383 => x"52",
          6384 => x"bf",
          6385 => x"54",
          6386 => x"15",
          6387 => x"38",
          6388 => x"05",
          6389 => x"3f",
          6390 => x"08",
          6391 => x"c8",
          6392 => x"77",
          6393 => x"a6",
          6394 => x"c8",
          6395 => x"82",
          6396 => x"a7",
          6397 => x"ed",
          6398 => x"80",
          6399 => x"02",
          6400 => x"df",
          6401 => x"57",
          6402 => x"3d",
          6403 => x"96",
          6404 => x"c8",
          6405 => x"c8",
          6406 => x"93",
          6407 => x"d4",
          6408 => x"65",
          6409 => x"d4",
          6410 => x"e0",
          6411 => x"c8",
          6412 => x"93",
          6413 => x"38",
          6414 => x"05",
          6415 => x"06",
          6416 => x"2e",
          6417 => x"55",
          6418 => x"75",
          6419 => x"71",
          6420 => x"33",
          6421 => x"74",
          6422 => x"57",
          6423 => x"8b",
          6424 => x"54",
          6425 => x"15",
          6426 => x"ff",
          6427 => x"82",
          6428 => x"55",
          6429 => x"c8",
          6430 => x"0d",
          6431 => x"0d",
          6432 => x"53",
          6433 => x"05",
          6434 => x"51",
          6435 => x"82",
          6436 => x"55",
          6437 => x"08",
          6438 => x"77",
          6439 => x"94",
          6440 => x"51",
          6441 => x"82",
          6442 => x"55",
          6443 => x"08",
          6444 => x"80",
          6445 => x"81",
          6446 => x"73",
          6447 => x"38",
          6448 => x"a9",
          6449 => x"22",
          6450 => x"70",
          6451 => x"07",
          6452 => x"7f",
          6453 => x"ff",
          6454 => x"77",
          6455 => x"83",
          6456 => x"51",
          6457 => x"3f",
          6458 => x"08",
          6459 => x"93",
          6460 => x"3d",
          6461 => x"3d",
          6462 => x"5c",
          6463 => x"98",
          6464 => x"52",
          6465 => x"cb",
          6466 => x"93",
          6467 => x"93",
          6468 => x"70",
          6469 => x"08",
          6470 => x"7b",
          6471 => x"07",
          6472 => x"06",
          6473 => x"56",
          6474 => x"2e",
          6475 => x"7b",
          6476 => x"80",
          6477 => x"70",
          6478 => x"b7",
          6479 => x"93",
          6480 => x"82",
          6481 => x"80",
          6482 => x"52",
          6483 => x"bc",
          6484 => x"93",
          6485 => x"82",
          6486 => x"bb",
          6487 => x"c8",
          6488 => x"c8",
          6489 => x"58",
          6490 => x"81",
          6491 => x"56",
          6492 => x"33",
          6493 => x"18",
          6494 => x"27",
          6495 => x"19",
          6496 => x"34",
          6497 => x"8f",
          6498 => x"79",
          6499 => x"51",
          6500 => x"a0",
          6501 => x"75",
          6502 => x"81",
          6503 => x"80",
          6504 => x"56",
          6505 => x"77",
          6506 => x"7c",
          6507 => x"07",
          6508 => x"06",
          6509 => x"55",
          6510 => x"bc",
          6511 => x"11",
          6512 => x"ff",
          6513 => x"82",
          6514 => x"56",
          6515 => x"08",
          6516 => x"70",
          6517 => x"80",
          6518 => x"83",
          6519 => x"80",
          6520 => x"84",
          6521 => x"a7",
          6522 => x"b4",
          6523 => x"a6",
          6524 => x"93",
          6525 => x"0c",
          6526 => x"c8",
          6527 => x"0d",
          6528 => x"0d",
          6529 => x"3d",
          6530 => x"52",
          6531 => x"c9",
          6532 => x"93",
          6533 => x"82",
          6534 => x"83",
          6535 => x"53",
          6536 => x"3d",
          6537 => x"51",
          6538 => x"3f",
          6539 => x"71",
          6540 => x"55",
          6541 => x"27",
          6542 => x"74",
          6543 => x"05",
          6544 => x"ff",
          6545 => x"ff",
          6546 => x"82",
          6547 => x"80",
          6548 => x"6a",
          6549 => x"53",
          6550 => x"a7",
          6551 => x"93",
          6552 => x"2e",
          6553 => x"88",
          6554 => x"6b",
          6555 => x"56",
          6556 => x"56",
          6557 => x"54",
          6558 => x"8a",
          6559 => x"70",
          6560 => x"06",
          6561 => x"ff",
          6562 => x"38",
          6563 => x"16",
          6564 => x"80",
          6565 => x"75",
          6566 => x"f8",
          6567 => x"f7",
          6568 => x"c8",
          6569 => x"81",
          6570 => x"88",
          6571 => x"26",
          6572 => x"39",
          6573 => x"86",
          6574 => x"82",
          6575 => x"ff",
          6576 => x"38",
          6577 => x"05",
          6578 => x"76",
          6579 => x"55",
          6580 => x"81",
          6581 => x"3d",
          6582 => x"bc",
          6583 => x"74",
          6584 => x"6b",
          6585 => x"56",
          6586 => x"26",
          6587 => x"89",
          6588 => x"86",
          6589 => x"e5",
          6590 => x"38",
          6591 => x"a8",
          6592 => x"05",
          6593 => x"70",
          6594 => x"56",
          6595 => x"2e",
          6596 => x"94",
          6597 => x"57",
          6598 => x"8c",
          6599 => x"70",
          6600 => x"73",
          6601 => x"38",
          6602 => x"41",
          6603 => x"3d",
          6604 => x"ff",
          6605 => x"82",
          6606 => x"54",
          6607 => x"08",
          6608 => x"81",
          6609 => x"ff",
          6610 => x"82",
          6611 => x"54",
          6612 => x"08",
          6613 => x"80",
          6614 => x"8b",
          6615 => x"ff",
          6616 => x"65",
          6617 => x"c0",
          6618 => x"65",
          6619 => x"34",
          6620 => x"0b",
          6621 => x"77",
          6622 => x"92",
          6623 => x"c8",
          6624 => x"df",
          6625 => x"c8",
          6626 => x"09",
          6627 => x"d3",
          6628 => x"76",
          6629 => x"cb",
          6630 => x"9a",
          6631 => x"51",
          6632 => x"3f",
          6633 => x"08",
          6634 => x"c8",
          6635 => x"a0",
          6636 => x"c8",
          6637 => x"51",
          6638 => x"3f",
          6639 => x"0b",
          6640 => x"8b",
          6641 => x"ff",
          6642 => x"65",
          6643 => x"d8",
          6644 => x"81",
          6645 => x"34",
          6646 => x"a6",
          6647 => x"93",
          6648 => x"73",
          6649 => x"93",
          6650 => x"3d",
          6651 => x"3d",
          6652 => x"02",
          6653 => x"cf",
          6654 => x"3d",
          6655 => x"72",
          6656 => x"58",
          6657 => x"82",
          6658 => x"57",
          6659 => x"08",
          6660 => x"18",
          6661 => x"80",
          6662 => x"76",
          6663 => x"39",
          6664 => x"95",
          6665 => x"08",
          6666 => x"18",
          6667 => x"2a",
          6668 => x"51",
          6669 => x"90",
          6670 => x"82",
          6671 => x"57",
          6672 => x"81",
          6673 => x"39",
          6674 => x"22",
          6675 => x"70",
          6676 => x"58",
          6677 => x"f9",
          6678 => x"16",
          6679 => x"30",
          6680 => x"9f",
          6681 => x"c8",
          6682 => x"8c",
          6683 => x"52",
          6684 => x"80",
          6685 => x"27",
          6686 => x"14",
          6687 => x"83",
          6688 => x"78",
          6689 => x"80",
          6690 => x"77",
          6691 => x"d7",
          6692 => x"c8",
          6693 => x"61",
          6694 => x"98",
          6695 => x"26",
          6696 => x"55",
          6697 => x"ff",
          6698 => x"ff",
          6699 => x"38",
          6700 => x"81",
          6701 => x"7e",
          6702 => x"85",
          6703 => x"80",
          6704 => x"2e",
          6705 => x"c1",
          6706 => x"76",
          6707 => x"7b",
          6708 => x"38",
          6709 => x"55",
          6710 => x"b3",
          6711 => x"54",
          6712 => x"09",
          6713 => x"38",
          6714 => x"53",
          6715 => x"51",
          6716 => x"3f",
          6717 => x"08",
          6718 => x"c8",
          6719 => x"74",
          6720 => x"18",
          6721 => x"75",
          6722 => x"39",
          6723 => x"76",
          6724 => x"7f",
          6725 => x"0c",
          6726 => x"2e",
          6727 => x"88",
          6728 => x"8c",
          6729 => x"18",
          6730 => x"07",
          6731 => x"19",
          6732 => x"11",
          6733 => x"55",
          6734 => x"08",
          6735 => x"38",
          6736 => x"7e",
          6737 => x"0c",
          6738 => x"33",
          6739 => x"55",
          6740 => x"34",
          6741 => x"82",
          6742 => x"91",
          6743 => x"ea",
          6744 => x"02",
          6745 => x"e7",
          6746 => x"3d",
          6747 => x"ff",
          6748 => x"82",
          6749 => x"56",
          6750 => x"0b",
          6751 => x"08",
          6752 => x"38",
          6753 => x"08",
          6754 => x"93",
          6755 => x"74",
          6756 => x"87",
          6757 => x"55",
          6758 => x"75",
          6759 => x"5a",
          6760 => x"51",
          6761 => x"3f",
          6762 => x"08",
          6763 => x"70",
          6764 => x"56",
          6765 => x"8c",
          6766 => x"82",
          6767 => x"06",
          6768 => x"57",
          6769 => x"38",
          6770 => x"05",
          6771 => x"79",
          6772 => x"dd",
          6773 => x"c8",
          6774 => x"66",
          6775 => x"38",
          6776 => x"80",
          6777 => x"66",
          6778 => x"06",
          6779 => x"2e",
          6780 => x"47",
          6781 => x"77",
          6782 => x"38",
          6783 => x"92",
          6784 => x"80",
          6785 => x"38",
          6786 => x"06",
          6787 => x"2e",
          6788 => x"57",
          6789 => x"7d",
          6790 => x"fe",
          6791 => x"82",
          6792 => x"6c",
          6793 => x"53",
          6794 => x"f6",
          6795 => x"93",
          6796 => x"82",
          6797 => x"29",
          6798 => x"62",
          6799 => x"82",
          6800 => x"30",
          6801 => x"c8",
          6802 => x"25",
          6803 => x"59",
          6804 => x"41",
          6805 => x"8a",
          6806 => x"3d",
          6807 => x"81",
          6808 => x"ff",
          6809 => x"81",
          6810 => x"c8",
          6811 => x"38",
          6812 => x"70",
          6813 => x"55",
          6814 => x"64",
          6815 => x"06",
          6816 => x"44",
          6817 => x"66",
          6818 => x"38",
          6819 => x"46",
          6820 => x"ff",
          6821 => x"bc",
          6822 => x"77",
          6823 => x"8a",
          6824 => x"81",
          6825 => x"06",
          6826 => x"80",
          6827 => x"7c",
          6828 => x"74",
          6829 => x"38",
          6830 => x"55",
          6831 => x"83",
          6832 => x"7c",
          6833 => x"93",
          6834 => x"74",
          6835 => x"84",
          6836 => x"61",
          6837 => x"81",
          6838 => x"38",
          6839 => x"65",
          6840 => x"5c",
          6841 => x"81",
          6842 => x"71",
          6843 => x"56",
          6844 => x"2e",
          6845 => x"77",
          6846 => x"81",
          6847 => x"71",
          6848 => x"22",
          6849 => x"5b",
          6850 => x"86",
          6851 => x"27",
          6852 => x"52",
          6853 => x"f4",
          6854 => x"93",
          6855 => x"93",
          6856 => x"10",
          6857 => x"87",
          6858 => x"fe",
          6859 => x"82",
          6860 => x"5c",
          6861 => x"0b",
          6862 => x"17",
          6863 => x"ff",
          6864 => x"27",
          6865 => x"8e",
          6866 => x"39",
          6867 => x"65",
          6868 => x"5c",
          6869 => x"81",
          6870 => x"71",
          6871 => x"56",
          6872 => x"2e",
          6873 => x"77",
          6874 => x"81",
          6875 => x"71",
          6876 => x"22",
          6877 => x"5b",
          6878 => x"86",
          6879 => x"27",
          6880 => x"52",
          6881 => x"f3",
          6882 => x"93",
          6883 => x"84",
          6884 => x"93",
          6885 => x"f5",
          6886 => x"81",
          6887 => x"c8",
          6888 => x"11",
          6889 => x"83",
          6890 => x"42",
          6891 => x"1e",
          6892 => x"fe",
          6893 => x"82",
          6894 => x"5c",
          6895 => x"5b",
          6896 => x"51",
          6897 => x"3f",
          6898 => x"08",
          6899 => x"06",
          6900 => x"7c",
          6901 => x"68",
          6902 => x"69",
          6903 => x"06",
          6904 => x"58",
          6905 => x"61",
          6906 => x"81",
          6907 => x"76",
          6908 => x"41",
          6909 => x"76",
          6910 => x"90",
          6911 => x"65",
          6912 => x"74",
          6913 => x"be",
          6914 => x"31",
          6915 => x"53",
          6916 => x"52",
          6917 => x"9e",
          6918 => x"c8",
          6919 => x"83",
          6920 => x"06",
          6921 => x"93",
          6922 => x"ff",
          6923 => x"38",
          6924 => x"78",
          6925 => x"77",
          6926 => x"8e",
          6927 => x"39",
          6928 => x"09",
          6929 => x"d3",
          6930 => x"f5",
          6931 => x"38",
          6932 => x"78",
          6933 => x"80",
          6934 => x"38",
          6935 => x"f1",
          6936 => x"2a",
          6937 => x"74",
          6938 => x"38",
          6939 => x"e1",
          6940 => x"38",
          6941 => x"81",
          6942 => x"fc",
          6943 => x"57",
          6944 => x"75",
          6945 => x"93",
          6946 => x"38",
          6947 => x"81",
          6948 => x"fc",
          6949 => x"57",
          6950 => x"80",
          6951 => x"2e",
          6952 => x"83",
          6953 => x"75",
          6954 => x"75",
          6955 => x"57",
          6956 => x"38",
          6957 => x"52",
          6958 => x"9a",
          6959 => x"53",
          6960 => x"52",
          6961 => x"99",
          6962 => x"52",
          6963 => x"ff",
          6964 => x"78",
          6965 => x"34",
          6966 => x"ff",
          6967 => x"1f",
          6968 => x"f7",
          6969 => x"90",
          6970 => x"83",
          6971 => x"70",
          6972 => x"80",
          6973 => x"55",
          6974 => x"ff",
          6975 => x"65",
          6976 => x"26",
          6977 => x"80",
          6978 => x"52",
          6979 => x"ff",
          6980 => x"8a",
          6981 => x"a0",
          6982 => x"98",
          6983 => x"7f",
          6984 => x"bf",
          6985 => x"51",
          6986 => x"3f",
          6987 => x"9a",
          6988 => x"98",
          6989 => x"52",
          6990 => x"ff",
          6991 => x"61",
          6992 => x"81",
          6993 => x"38",
          6994 => x"0a",
          6995 => x"1f",
          6996 => x"a5",
          6997 => x"a4",
          6998 => x"98",
          6999 => x"52",
          7000 => x"ff",
          7001 => x"81",
          7002 => x"51",
          7003 => x"3f",
          7004 => x"1f",
          7005 => x"e3",
          7006 => x"7f",
          7007 => x"34",
          7008 => x"c2",
          7009 => x"53",
          7010 => x"52",
          7011 => x"51",
          7012 => x"3f",
          7013 => x"88",
          7014 => x"a7",
          7015 => x"97",
          7016 => x"83",
          7017 => x"52",
          7018 => x"ff",
          7019 => x"ff",
          7020 => x"05",
          7021 => x"a6",
          7022 => x"53",
          7023 => x"52",
          7024 => x"ff",
          7025 => x"82",
          7026 => x"83",
          7027 => x"ff",
          7028 => x"81",
          7029 => x"7e",
          7030 => x"ff",
          7031 => x"81",
          7032 => x"c8",
          7033 => x"38",
          7034 => x"09",
          7035 => x"f0",
          7036 => x"63",
          7037 => x"7e",
          7038 => x"ff",
          7039 => x"7d",
          7040 => x"7e",
          7041 => x"c4",
          7042 => x"85",
          7043 => x"7e",
          7044 => x"e5",
          7045 => x"85",
          7046 => x"83",
          7047 => x"ff",
          7048 => x"ff",
          7049 => x"e8",
          7050 => x"96",
          7051 => x"52",
          7052 => x"51",
          7053 => x"3f",
          7054 => x"52",
          7055 => x"51",
          7056 => x"3f",
          7057 => x"87",
          7058 => x"52",
          7059 => x"93",
          7060 => x"54",
          7061 => x"53",
          7062 => x"51",
          7063 => x"3f",
          7064 => x"52",
          7065 => x"96",
          7066 => x"56",
          7067 => x"83",
          7068 => x"06",
          7069 => x"52",
          7070 => x"95",
          7071 => x"52",
          7072 => x"ff",
          7073 => x"f0",
          7074 => x"1f",
          7075 => x"e9",
          7076 => x"87",
          7077 => x"55",
          7078 => x"83",
          7079 => x"74",
          7080 => x"ff",
          7081 => x"7b",
          7082 => x"74",
          7083 => x"38",
          7084 => x"54",
          7085 => x"52",
          7086 => x"92",
          7087 => x"93",
          7088 => x"86",
          7089 => x"80",
          7090 => x"ff",
          7091 => x"76",
          7092 => x"31",
          7093 => x"d1",
          7094 => x"5b",
          7095 => x"ff",
          7096 => x"55",
          7097 => x"83",
          7098 => x"60",
          7099 => x"26",
          7100 => x"57",
          7101 => x"53",
          7102 => x"51",
          7103 => x"3f",
          7104 => x"08",
          7105 => x"76",
          7106 => x"31",
          7107 => x"db",
          7108 => x"61",
          7109 => x"38",
          7110 => x"83",
          7111 => x"8a",
          7112 => x"61",
          7113 => x"38",
          7114 => x"83",
          7115 => x"58",
          7116 => x"38",
          7117 => x"52",
          7118 => x"95",
          7119 => x"d4",
          7120 => x"fe",
          7121 => x"94",
          7122 => x"be",
          7123 => x"76",
          7124 => x"81",
          7125 => x"0b",
          7126 => x"77",
          7127 => x"76",
          7128 => x"63",
          7129 => x"80",
          7130 => x"76",
          7131 => x"c6",
          7132 => x"85",
          7133 => x"93",
          7134 => x"2a",
          7135 => x"74",
          7136 => x"82",
          7137 => x"87",
          7138 => x"52",
          7139 => x"51",
          7140 => x"3f",
          7141 => x"ca",
          7142 => x"93",
          7143 => x"54",
          7144 => x"52",
          7145 => x"90",
          7146 => x"57",
          7147 => x"08",
          7148 => x"53",
          7149 => x"51",
          7150 => x"3f",
          7151 => x"93",
          7152 => x"38",
          7153 => x"57",
          7154 => x"57",
          7155 => x"57",
          7156 => x"57",
          7157 => x"c8",
          7158 => x"0d",
          7159 => x"0d",
          7160 => x"93",
          7161 => x"38",
          7162 => x"81",
          7163 => x"52",
          7164 => x"82",
          7165 => x"ff",
          7166 => x"81",
          7167 => x"82",
          7168 => x"80",
          7169 => x"c9",
          7170 => x"98",
          7171 => x"93",
          7172 => x"39",
          7173 => x"51",
          7174 => x"3f",
          7175 => x"82",
          7176 => x"fe",
          7177 => x"81",
          7178 => x"82",
          7179 => x"ff",
          7180 => x"9d",
          7181 => x"e0",
          7182 => x"e7",
          7183 => x"39",
          7184 => x"51",
          7185 => x"3f",
          7186 => x"82",
          7187 => x"fe",
          7188 => x"80",
          7189 => x"83",
          7190 => x"ff",
          7191 => x"f1",
          7192 => x"b8",
          7193 => x"bb",
          7194 => x"39",
          7195 => x"51",
          7196 => x"3f",
          7197 => x"82",
          7198 => x"fe",
          7199 => x"80",
          7200 => x"84",
          7201 => x"ff",
          7202 => x"c5",
          7203 => x"a8",
          7204 => x"8f",
          7205 => x"82",
          7206 => x"fe",
          7207 => x"b1",
          7208 => x"dc",
          7209 => x"fb",
          7210 => x"82",
          7211 => x"fe",
          7212 => x"9d",
          7213 => x"8c",
          7214 => x"e7",
          7215 => x"82",
          7216 => x"fe",
          7217 => x"89",
          7218 => x"b0",
          7219 => x"d3",
          7220 => x"0d",
          7221 => x"0d",
          7222 => x"56",
          7223 => x"26",
          7224 => x"52",
          7225 => x"29",
          7226 => x"ca",
          7227 => x"c8",
          7228 => x"39",
          7229 => x"74",
          7230 => x"ba",
          7231 => x"c8",
          7232 => x"51",
          7233 => x"3f",
          7234 => x"08",
          7235 => x"79",
          7236 => x"82",
          7237 => x"ff",
          7238 => x"87",
          7239 => x"fe",
          7240 => x"81",
          7241 => x"81",
          7242 => x"02",
          7243 => x"e3",
          7244 => x"73",
          7245 => x"07",
          7246 => x"ff",
          7247 => x"54",
          7248 => x"57",
          7249 => x"75",
          7250 => x"81",
          7251 => x"81",
          7252 => x"d8",
          7253 => x"bc",
          7254 => x"93",
          7255 => x"82",
          7256 => x"bb",
          7257 => x"c8",
          7258 => x"98",
          7259 => x"93",
          7260 => x"81",
          7261 => x"d4",
          7262 => x"84",
          7263 => x"52",
          7264 => x"51",
          7265 => x"82",
          7266 => x"58",
          7267 => x"08",
          7268 => x"80",
          7269 => x"7a",
          7270 => x"58",
          7271 => x"81",
          7272 => x"d8",
          7273 => x"c1",
          7274 => x"70",
          7275 => x"25",
          7276 => x"9f",
          7277 => x"51",
          7278 => x"74",
          7279 => x"38",
          7280 => x"53",
          7281 => x"88",
          7282 => x"51",
          7283 => x"77",
          7284 => x"93",
          7285 => x"96",
          7286 => x"f8",
          7287 => x"b7",
          7288 => x"ff",
          7289 => x"80",
          7290 => x"7a",
          7291 => x"3f",
          7292 => x"08",
          7293 => x"80",
          7294 => x"76",
          7295 => x"38",
          7296 => x"55",
          7297 => x"93",
          7298 => x"52",
          7299 => x"2d",
          7300 => x"08",
          7301 => x"75",
          7302 => x"93",
          7303 => x"3d",
          7304 => x"3d",
          7305 => x"05",
          7306 => x"ec",
          7307 => x"f4",
          7308 => x"81",
          7309 => x"8b",
          7310 => x"52",
          7311 => x"d6",
          7312 => x"80",
          7313 => x"8c",
          7314 => x"33",
          7315 => x"94",
          7316 => x"c9",
          7317 => x"2e",
          7318 => x"f6",
          7319 => x"3d",
          7320 => x"3d",
          7321 => x"96",
          7322 => x"fe",
          7323 => x"81",
          7324 => x"ff",
          7325 => x"b0",
          7326 => x"f5",
          7327 => x"fe",
          7328 => x"72",
          7329 => x"81",
          7330 => x"71",
          7331 => x"38",
          7332 => x"ee",
          7333 => x"86",
          7334 => x"f0",
          7335 => x"51",
          7336 => x"3f",
          7337 => x"70",
          7338 => x"52",
          7339 => x"95",
          7340 => x"fe",
          7341 => x"82",
          7342 => x"fe",
          7343 => x"80",
          7344 => x"af",
          7345 => x"2a",
          7346 => x"51",
          7347 => x"2e",
          7348 => x"51",
          7349 => x"3f",
          7350 => x"51",
          7351 => x"3f",
          7352 => x"ee",
          7353 => x"84",
          7354 => x"06",
          7355 => x"80",
          7356 => x"81",
          7357 => x"fb",
          7358 => x"84",
          7359 => x"f1",
          7360 => x"fe",
          7361 => x"72",
          7362 => x"81",
          7363 => x"71",
          7364 => x"38",
          7365 => x"ed",
          7366 => x"87",
          7367 => x"ef",
          7368 => x"51",
          7369 => x"3f",
          7370 => x"70",
          7371 => x"52",
          7372 => x"95",
          7373 => x"fe",
          7374 => x"82",
          7375 => x"fe",
          7376 => x"80",
          7377 => x"ab",
          7378 => x"2a",
          7379 => x"51",
          7380 => x"2e",
          7381 => x"51",
          7382 => x"3f",
          7383 => x"51",
          7384 => x"3f",
          7385 => x"ed",
          7386 => x"88",
          7387 => x"06",
          7388 => x"80",
          7389 => x"81",
          7390 => x"f7",
          7391 => x"d4",
          7392 => x"ed",
          7393 => x"fe",
          7394 => x"fe",
          7395 => x"84",
          7396 => x"fa",
          7397 => x"70",
          7398 => x"56",
          7399 => x"2e",
          7400 => x"8e",
          7401 => x"0c",
          7402 => x"53",
          7403 => x"81",
          7404 => x"75",
          7405 => x"72",
          7406 => x"38",
          7407 => x"30",
          7408 => x"75",
          7409 => x"72",
          7410 => x"33",
          7411 => x"2e",
          7412 => x"88",
          7413 => x"70",
          7414 => x"34",
          7415 => x"90",
          7416 => x"88",
          7417 => x"53",
          7418 => x"54",
          7419 => x"3f",
          7420 => x"08",
          7421 => x"14",
          7422 => x"81",
          7423 => x"38",
          7424 => x"81",
          7425 => x"53",
          7426 => x"d2",
          7427 => x"72",
          7428 => x"0c",
          7429 => x"04",
          7430 => x"80",
          7431 => x"c8",
          7432 => x"5d",
          7433 => x"5a",
          7434 => x"51",
          7435 => x"3f",
          7436 => x"08",
          7437 => x"59",
          7438 => x"09",
          7439 => x"38",
          7440 => x"52",
          7441 => x"52",
          7442 => x"e7",
          7443 => x"78",
          7444 => x"1b",
          7445 => x"ab",
          7446 => x"c8",
          7447 => x"80",
          7448 => x"82",
          7449 => x"fe",
          7450 => x"85",
          7451 => x"5e",
          7452 => x"d0",
          7453 => x"ab",
          7454 => x"70",
          7455 => x"f8",
          7456 => x"80",
          7457 => x"fe",
          7458 => x"79",
          7459 => x"fe",
          7460 => x"b4",
          7461 => x"05",
          7462 => x"3f",
          7463 => x"08",
          7464 => x"90",
          7465 => x"78",
          7466 => x"85",
          7467 => x"10",
          7468 => x"88",
          7469 => x"08",
          7470 => x"fe",
          7471 => x"fe",
          7472 => x"fe",
          7473 => x"82",
          7474 => x"8c",
          7475 => x"d4",
          7476 => x"c9",
          7477 => x"39",
          7478 => x"f0",
          7479 => x"f8",
          7480 => x"fe",
          7481 => x"93",
          7482 => x"2e",
          7483 => x"60",
          7484 => x"80",
          7485 => x"05",
          7486 => x"80",
          7487 => x"51",
          7488 => x"3f",
          7489 => x"08",
          7490 => x"59",
          7491 => x"82",
          7492 => x"fe",
          7493 => x"81",
          7494 => x"39",
          7495 => x"51",
          7496 => x"3f",
          7497 => x"b4",
          7498 => x"11",
          7499 => x"05",
          7500 => x"f4",
          7501 => x"c8",
          7502 => x"fe",
          7503 => x"53",
          7504 => x"80",
          7505 => x"51",
          7506 => x"3f",
          7507 => x"08",
          7508 => x"8c",
          7509 => x"c5",
          7510 => x"39",
          7511 => x"f4",
          7512 => x"f8",
          7513 => x"fd",
          7514 => x"93",
          7515 => x"2e",
          7516 => x"89",
          7517 => x"38",
          7518 => x"f0",
          7519 => x"f8",
          7520 => x"fd",
          7521 => x"93",
          7522 => x"38",
          7523 => x"08",
          7524 => x"82",
          7525 => x"96",
          7526 => x"59",
          7527 => x"3f",
          7528 => x"33",
          7529 => x"60",
          7530 => x"82",
          7531 => x"51",
          7532 => x"3f",
          7533 => x"08",
          7534 => x"38",
          7535 => x"08",
          7536 => x"3f",
          7537 => x"82",
          7538 => x"fe",
          7539 => x"81",
          7540 => x"39",
          7541 => x"f8",
          7542 => x"e4",
          7543 => x"93",
          7544 => x"3d",
          7545 => x"52",
          7546 => x"fa",
          7547 => x"82",
          7548 => x"52",
          7549 => x"a7",
          7550 => x"c8",
          7551 => x"fc",
          7552 => x"93",
          7553 => x"f3",
          7554 => x"e5",
          7555 => x"fe",
          7556 => x"fe",
          7557 => x"82",
          7558 => x"b5",
          7559 => x"05",
          7560 => x"e4",
          7561 => x"93",
          7562 => x"3d",
          7563 => x"52",
          7564 => x"b2",
          7565 => x"c8",
          7566 => x"fe",
          7567 => x"59",
          7568 => x"3f",
          7569 => x"58",
          7570 => x"57",
          7571 => x"55",
          7572 => x"08",
          7573 => x"54",
          7574 => x"52",
          7575 => x"fb",
          7576 => x"c8",
          7577 => x"fc",
          7578 => x"93",
          7579 => x"f2",
          7580 => x"fd",
          7581 => x"98",
          7582 => x"a7",
          7583 => x"fe",
          7584 => x"fb",
          7585 => x"89",
          7586 => x"f3",
          7587 => x"51",
          7588 => x"3f",
          7589 => x"84",
          7590 => x"87",
          7591 => x"0c",
          7592 => x"0b",
          7593 => x"94",
          7594 => x"c8",
          7595 => x"f3",
          7596 => x"39",
          7597 => x"51",
          7598 => x"3f",
          7599 => x"0b",
          7600 => x"84",
          7601 => x"83",
          7602 => x"94",
          7603 => x"a1",
          7604 => x"fe",
          7605 => x"fe",
          7606 => x"fe",
          7607 => x"82",
          7608 => x"80",
          7609 => x"38",
          7610 => x"89",
          7611 => x"f8",
          7612 => x"59",
          7613 => x"3d",
          7614 => x"53",
          7615 => x"51",
          7616 => x"3f",
          7617 => x"08",
          7618 => x"e5",
          7619 => x"82",
          7620 => x"fe",
          7621 => x"60",
          7622 => x"82",
          7623 => x"5e",
          7624 => x"08",
          7625 => x"c9",
          7626 => x"c8",
          7627 => x"8a",
          7628 => x"f7",
          7629 => x"b9",
          7630 => x"c4",
          7631 => x"e3",
          7632 => x"bc",
          7633 => x"39",
          7634 => x"51",
          7635 => x"3f",
          7636 => x"a0",
          7637 => x"84",
          7638 => x"39",
          7639 => x"51",
          7640 => x"2e",
          7641 => x"7c",
          7642 => x"78",
          7643 => x"cb",
          7644 => x"fe",
          7645 => x"fe",
          7646 => x"82",
          7647 => x"82",
          7648 => x"55",
          7649 => x"54",
          7650 => x"8a",
          7651 => x"3d",
          7652 => x"fe",
          7653 => x"82",
          7654 => x"82",
          7655 => x"80",
          7656 => x"05",
          7657 => x"80",
          7658 => x"80",
          7659 => x"80",
          7660 => x"f4",
          7661 => x"93",
          7662 => x"7c",
          7663 => x"81",
          7664 => x"78",
          7665 => x"ff",
          7666 => x"06",
          7667 => x"82",
          7668 => x"fe",
          7669 => x"f9",
          7670 => x"3d",
          7671 => x"82",
          7672 => x"9b",
          7673 => x"0b",
          7674 => x"8c",
          7675 => x"86",
          7676 => x"c0",
          7677 => x"8c",
          7678 => x"87",
          7679 => x"0c",
          7680 => x"0b",
          7681 => x"94",
          7682 => x"8d",
          7683 => x"d8",
          7684 => x"80",
          7685 => x"dc",
          7686 => x"87",
          7687 => x"cd",
          7688 => x"9c",
          7689 => x"c9",
          7690 => x"a8",
          7691 => x"f3",
          7692 => x"e2",
          7693 => x"b0",
          7694 => x"f3",
          7695 => x"d8",
          7696 => x"00",
          7697 => x"5d",
          7698 => x"30",
          7699 => x"39",
          7700 => x"42",
          7701 => x"4b",
          7702 => x"54",
          7703 => x"cf",
          7704 => x"c0",
          7705 => x"d7",
          7706 => x"df",
          7707 => x"df",
          7708 => x"df",
          7709 => x"df",
          7710 => x"df",
          7711 => x"df",
          7712 => x"df",
          7713 => x"df",
          7714 => x"df",
          7715 => x"df",
          7716 => x"d3",
          7717 => x"df",
          7718 => x"df",
          7719 => x"df",
          7720 => x"53",
          7721 => x"df",
          7722 => x"d7",
          7723 => x"df",
          7724 => x"df",
          7725 => x"db",
          7726 => x"bf",
          7727 => x"f3",
          7728 => x"fe",
          7729 => x"09",
          7730 => x"14",
          7731 => x"1f",
          7732 => x"2a",
          7733 => x"35",
          7734 => x"40",
          7735 => x"4b",
          7736 => x"56",
          7737 => x"61",
          7738 => x"6c",
          7739 => x"77",
          7740 => x"82",
          7741 => x"8d",
          7742 => x"97",
          7743 => x"a1",
          7744 => x"ab",
          7745 => x"b5",
          7746 => x"71",
          7747 => x"5c",
          7748 => x"b9",
          7749 => x"5c",
          7750 => x"27",
          7751 => x"5c",
          7752 => x"5c",
          7753 => x"5c",
          7754 => x"5c",
          7755 => x"5c",
          7756 => x"5c",
          7757 => x"5c",
          7758 => x"5c",
          7759 => x"5c",
          7760 => x"5c",
          7761 => x"5c",
          7762 => x"5c",
          7763 => x"5c",
          7764 => x"5c",
          7765 => x"5c",
          7766 => x"5c",
          7767 => x"5c",
          7768 => x"5c",
          7769 => x"5c",
          7770 => x"5c",
          7771 => x"5c",
          7772 => x"5c",
          7773 => x"5c",
          7774 => x"5c",
          7775 => x"5c",
          7776 => x"5c",
          7777 => x"5c",
          7778 => x"5c",
          7779 => x"5c",
          7780 => x"5c",
          7781 => x"5c",
          7782 => x"5c",
          7783 => x"5c",
          7784 => x"5c",
          7785 => x"5c",
          7786 => x"5c",
          7787 => x"5c",
          7788 => x"5c",
          7789 => x"d4",
          7790 => x"5c",
          7791 => x"5c",
          7792 => x"5c",
          7793 => x"5c",
          7794 => x"0d",
          7795 => x"5c",
          7796 => x"5c",
          7797 => x"5c",
          7798 => x"5c",
          7799 => x"5c",
          7800 => x"5c",
          7801 => x"5c",
          7802 => x"5c",
          7803 => x"5c",
          7804 => x"5c",
          7805 => x"5c",
          7806 => x"5c",
          7807 => x"5c",
          7808 => x"5c",
          7809 => x"5c",
          7810 => x"5c",
          7811 => x"5c",
          7812 => x"5c",
          7813 => x"5c",
          7814 => x"5c",
          7815 => x"5c",
          7816 => x"5c",
          7817 => x"5c",
          7818 => x"5c",
          7819 => x"5c",
          7820 => x"5c",
          7821 => x"5c",
          7822 => x"5c",
          7823 => x"5c",
          7824 => x"5c",
          7825 => x"5c",
          7826 => x"75",
          7827 => x"86",
          7828 => x"5c",
          7829 => x"5c",
          7830 => x"97",
          7831 => x"b4",
          7832 => x"5c",
          7833 => x"5c",
          7834 => x"5c",
          7835 => x"5c",
          7836 => x"5c",
          7837 => x"5c",
          7838 => x"5c",
          7839 => x"5c",
          7840 => x"5c",
          7841 => x"5c",
          7842 => x"5c",
          7843 => x"5c",
          7844 => x"5c",
          7845 => x"5c",
          7846 => x"5c",
          7847 => x"5c",
          7848 => x"5c",
          7849 => x"5c",
          7850 => x"5c",
          7851 => x"5c",
          7852 => x"5c",
          7853 => x"5c",
          7854 => x"5c",
          7855 => x"5c",
          7856 => x"5c",
          7857 => x"5c",
          7858 => x"5c",
          7859 => x"5c",
          7860 => x"5c",
          7861 => x"5c",
          7862 => x"5c",
          7863 => x"5c",
          7864 => x"5c",
          7865 => x"5c",
          7866 => x"d1",
          7867 => x"f6",
          7868 => x"5c",
          7869 => x"5c",
          7870 => x"5c",
          7871 => x"5c",
          7872 => x"5c",
          7873 => x"5c",
          7874 => x"5c",
          7875 => x"5c",
          7876 => x"39",
          7877 => x"48",
          7878 => x"5c",
          7879 => x"55",
          7880 => x"5c",
          7881 => x"71",
          7882 => x"25",
          7883 => x"64",
          7884 => x"3a",
          7885 => x"25",
          7886 => x"64",
          7887 => x"00",
          7888 => x"20",
          7889 => x"66",
          7890 => x"72",
          7891 => x"6f",
          7892 => x"00",
          7893 => x"72",
          7894 => x"53",
          7895 => x"63",
          7896 => x"69",
          7897 => x"00",
          7898 => x"65",
          7899 => x"65",
          7900 => x"6d",
          7901 => x"6d",
          7902 => x"65",
          7903 => x"00",
          7904 => x"20",
          7905 => x"4e",
          7906 => x"41",
          7907 => x"53",
          7908 => x"74",
          7909 => x"38",
          7910 => x"53",
          7911 => x"3d",
          7912 => x"58",
          7913 => x"00",
          7914 => x"20",
          7915 => x"4d",
          7916 => x"74",
          7917 => x"3d",
          7918 => x"58",
          7919 => x"69",
          7920 => x"25",
          7921 => x"29",
          7922 => x"00",
          7923 => x"20",
          7924 => x"20",
          7925 => x"61",
          7926 => x"25",
          7927 => x"2c",
          7928 => x"7a",
          7929 => x"30",
          7930 => x"2e",
          7931 => x"00",
          7932 => x"20",
          7933 => x"54",
          7934 => x"00",
          7935 => x"20",
          7936 => x"0a",
          7937 => x"00",
          7938 => x"20",
          7939 => x"0a",
          7940 => x"00",
          7941 => x"20",
          7942 => x"43",
          7943 => x"20",
          7944 => x"76",
          7945 => x"73",
          7946 => x"32",
          7947 => x"0a",
          7948 => x"00",
          7949 => x"20",
          7950 => x"45",
          7951 => x"50",
          7952 => x"4f",
          7953 => x"4f",
          7954 => x"52",
          7955 => x"00",
          7956 => x"20",
          7957 => x"45",
          7958 => x"28",
          7959 => x"65",
          7960 => x"25",
          7961 => x"29",
          7962 => x"00",
          7963 => x"72",
          7964 => x"65",
          7965 => x"00",
          7966 => x"20",
          7967 => x"20",
          7968 => x"65",
          7969 => x"65",
          7970 => x"72",
          7971 => x"64",
          7972 => x"73",
          7973 => x"25",
          7974 => x"0a",
          7975 => x"00",
          7976 => x"20",
          7977 => x"20",
          7978 => x"6f",
          7979 => x"53",
          7980 => x"74",
          7981 => x"64",
          7982 => x"73",
          7983 => x"25",
          7984 => x"0a",
          7985 => x"00",
          7986 => x"20",
          7987 => x"63",
          7988 => x"74",
          7989 => x"20",
          7990 => x"72",
          7991 => x"20",
          7992 => x"20",
          7993 => x"25",
          7994 => x"0a",
          7995 => x"00",
          7996 => x"20",
          7997 => x"20",
          7998 => x"20",
          7999 => x"20",
          8000 => x"20",
          8001 => x"20",
          8002 => x"20",
          8003 => x"25",
          8004 => x"0a",
          8005 => x"00",
          8006 => x"20",
          8007 => x"74",
          8008 => x"43",
          8009 => x"6b",
          8010 => x"65",
          8011 => x"20",
          8012 => x"20",
          8013 => x"25",
          8014 => x"0a",
          8015 => x"00",
          8016 => x"6c",
          8017 => x"00",
          8018 => x"69",
          8019 => x"00",
          8020 => x"78",
          8021 => x"00",
          8022 => x"00",
          8023 => x"6d",
          8024 => x"00",
          8025 => x"6e",
          8026 => x"00",
          8027 => x"00",
          8028 => x"2c",
          8029 => x"3d",
          8030 => x"5d",
          8031 => x"00",
          8032 => x"00",
          8033 => x"33",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"00",
          8045 => x"4d",
          8046 => x"53",
          8047 => x"00",
          8048 => x"4e",
          8049 => x"20",
          8050 => x"46",
          8051 => x"32",
          8052 => x"00",
          8053 => x"4e",
          8054 => x"20",
          8055 => x"46",
          8056 => x"20",
          8057 => x"00",
          8058 => x"6c",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"41",
          8063 => x"80",
          8064 => x"49",
          8065 => x"8f",
          8066 => x"4f",
          8067 => x"55",
          8068 => x"9b",
          8069 => x"9f",
          8070 => x"55",
          8071 => x"a7",
          8072 => x"ab",
          8073 => x"af",
          8074 => x"b3",
          8075 => x"b7",
          8076 => x"bb",
          8077 => x"bf",
          8078 => x"c3",
          8079 => x"c7",
          8080 => x"cb",
          8081 => x"cf",
          8082 => x"d3",
          8083 => x"d7",
          8084 => x"db",
          8085 => x"df",
          8086 => x"e3",
          8087 => x"e7",
          8088 => x"eb",
          8089 => x"ef",
          8090 => x"f3",
          8091 => x"f7",
          8092 => x"fb",
          8093 => x"ff",
          8094 => x"3b",
          8095 => x"2f",
          8096 => x"3a",
          8097 => x"7c",
          8098 => x"00",
          8099 => x"04",
          8100 => x"40",
          8101 => x"00",
          8102 => x"00",
          8103 => x"02",
          8104 => x"08",
          8105 => x"20",
          8106 => x"00",
          8107 => x"31",
          8108 => x"00",
          8109 => x"31",
          8110 => x"00",
          8111 => x"41",
          8112 => x"00",
          8113 => x"4b",
          8114 => x"20",
          8115 => x"54",
          8116 => x"53",
          8117 => x"00",
          8118 => x"4b",
          8119 => x"46",
          8120 => x"20",
          8121 => x"54",
          8122 => x"53",
          8123 => x"00",
          8124 => x"45",
          8125 => x"54",
          8126 => x"43",
          8127 => x"52",
          8128 => x"00",
          8129 => x"4f",
          8130 => x"00",
          8131 => x"44",
          8132 => x"45",
          8133 => x"00",
          8134 => x"54",
          8135 => x"00",
          8136 => x"43",
          8137 => x"4f",
          8138 => x"00",
          8139 => x"43",
          8140 => x"4d",
          8141 => x"44",
          8142 => x"00",
          8143 => x"6d",
          8144 => x"00",
          8145 => x"69",
          8146 => x"00",
          8147 => x"61",
          8148 => x"00",
          8149 => x"63",
          8150 => x"00",
          8151 => x"6d",
          8152 => x"00",
          8153 => x"69",
          8154 => x"00",
          8155 => x"61",
          8156 => x"00",
          8157 => x"69",
          8158 => x"00",
          8159 => x"6c",
          8160 => x"00",
          8161 => x"6e",
          8162 => x"00",
          8163 => x"69",
          8164 => x"00",
          8165 => x"65",
          8166 => x"00",
          8167 => x"6f",
          8168 => x"00",
          8169 => x"65",
          8170 => x"00",
          8171 => x"61",
          8172 => x"00",
          8173 => x"73",
          8174 => x"74",
          8175 => x"00",
          8176 => x"69",
          8177 => x"00",
          8178 => x"75",
          8179 => x"00",
          8180 => x"6c",
          8181 => x"00",
          8182 => x"74",
          8183 => x"00",
          8184 => x"6d",
          8185 => x"00",
          8186 => x"6e",
          8187 => x"00",
          8188 => x"6c",
          8189 => x"00",
          8190 => x"64",
          8191 => x"00",
          8192 => x"61",
          8193 => x"00",
          8194 => x"72",
          8195 => x"00",
          8196 => x"74",
          8197 => x"00",
          8198 => x"00",
          8199 => x"6e",
          8200 => x"00",
          8201 => x"72",
          8202 => x"00",
          8203 => x"61",
          8204 => x"00",
          8205 => x"65",
          8206 => x"00",
          8207 => x"76",
          8208 => x"00",
          8209 => x"6d",
          8210 => x"00",
          8211 => x"00",
          8212 => x"69",
          8213 => x"00",
          8214 => x"6f",
          8215 => x"72",
          8216 => x"00",
          8217 => x"62",
          8218 => x"00",
          8219 => x"66",
          8220 => x"00",
          8221 => x"72",
          8222 => x"00",
          8223 => x"6d",
          8224 => x"00",
          8225 => x"00",
          8226 => x"00",
          8227 => x"00",
          8228 => x"00",
          8229 => x"00",
          8230 => x"00",
          8231 => x"00",
          8232 => x"00",
          8233 => x"00",
          8234 => x"79",
          8235 => x"00",
          8236 => x"65",
          8237 => x"6b",
          8238 => x"00",
          8239 => x"6c",
          8240 => x"00",
          8241 => x"00",
          8242 => x"74",
          8243 => x"00",
          8244 => x"65",
          8245 => x"00",
          8246 => x"70",
          8247 => x"00",
          8248 => x"6f",
          8249 => x"00",
          8250 => x"65",
          8251 => x"00",
          8252 => x"74",
          8253 => x"00",
          8254 => x"6b",
          8255 => x"72",
          8256 => x"00",
          8257 => x"65",
          8258 => x"6c",
          8259 => x"72",
          8260 => x"0a",
          8261 => x"00",
          8262 => x"6b",
          8263 => x"74",
          8264 => x"61",
          8265 => x"0a",
          8266 => x"00",
          8267 => x"66",
          8268 => x"20",
          8269 => x"6e",
          8270 => x"00",
          8271 => x"70",
          8272 => x"20",
          8273 => x"6e",
          8274 => x"00",
          8275 => x"61",
          8276 => x"20",
          8277 => x"65",
          8278 => x"65",
          8279 => x"00",
          8280 => x"65",
          8281 => x"64",
          8282 => x"65",
          8283 => x"00",
          8284 => x"65",
          8285 => x"72",
          8286 => x"79",
          8287 => x"69",
          8288 => x"2e",
          8289 => x"00",
          8290 => x"65",
          8291 => x"6e",
          8292 => x"20",
          8293 => x"61",
          8294 => x"2e",
          8295 => x"00",
          8296 => x"69",
          8297 => x"72",
          8298 => x"20",
          8299 => x"74",
          8300 => x"65",
          8301 => x"00",
          8302 => x"76",
          8303 => x"75",
          8304 => x"72",
          8305 => x"20",
          8306 => x"61",
          8307 => x"2e",
          8308 => x"00",
          8309 => x"6b",
          8310 => x"74",
          8311 => x"61",
          8312 => x"64",
          8313 => x"00",
          8314 => x"63",
          8315 => x"61",
          8316 => x"6c",
          8317 => x"69",
          8318 => x"79",
          8319 => x"6d",
          8320 => x"75",
          8321 => x"6f",
          8322 => x"69",
          8323 => x"0a",
          8324 => x"00",
          8325 => x"6d",
          8326 => x"61",
          8327 => x"74",
          8328 => x"0a",
          8329 => x"00",
          8330 => x"65",
          8331 => x"2c",
          8332 => x"65",
          8333 => x"69",
          8334 => x"63",
          8335 => x"65",
          8336 => x"64",
          8337 => x"00",
          8338 => x"65",
          8339 => x"20",
          8340 => x"6b",
          8341 => x"0a",
          8342 => x"00",
          8343 => x"75",
          8344 => x"63",
          8345 => x"74",
          8346 => x"6d",
          8347 => x"2e",
          8348 => x"00",
          8349 => x"20",
          8350 => x"79",
          8351 => x"65",
          8352 => x"69",
          8353 => x"2e",
          8354 => x"00",
          8355 => x"61",
          8356 => x"65",
          8357 => x"69",
          8358 => x"72",
          8359 => x"74",
          8360 => x"00",
          8361 => x"63",
          8362 => x"2e",
          8363 => x"00",
          8364 => x"6e",
          8365 => x"20",
          8366 => x"6f",
          8367 => x"00",
          8368 => x"75",
          8369 => x"74",
          8370 => x"25",
          8371 => x"74",
          8372 => x"75",
          8373 => x"74",
          8374 => x"73",
          8375 => x"0a",
          8376 => x"00",
          8377 => x"64",
          8378 => x"00",
          8379 => x"54",
          8380 => x"00",
          8381 => x"20",
          8382 => x"28",
          8383 => x"00",
          8384 => x"30",
          8385 => x"30",
          8386 => x"00",
          8387 => x"33",
          8388 => x"00",
          8389 => x"55",
          8390 => x"65",
          8391 => x"30",
          8392 => x"20",
          8393 => x"25",
          8394 => x"2a",
          8395 => x"00",
          8396 => x"54",
          8397 => x"6e",
          8398 => x"72",
          8399 => x"20",
          8400 => x"64",
          8401 => x"0a",
          8402 => x"00",
          8403 => x"65",
          8404 => x"6e",
          8405 => x"72",
          8406 => x"0a",
          8407 => x"00",
          8408 => x"20",
          8409 => x"65",
          8410 => x"70",
          8411 => x"00",
          8412 => x"54",
          8413 => x"44",
          8414 => x"74",
          8415 => x"75",
          8416 => x"00",
          8417 => x"54",
          8418 => x"52",
          8419 => x"74",
          8420 => x"75",
          8421 => x"00",
          8422 => x"54",
          8423 => x"58",
          8424 => x"74",
          8425 => x"75",
          8426 => x"00",
          8427 => x"54",
          8428 => x"58",
          8429 => x"74",
          8430 => x"75",
          8431 => x"00",
          8432 => x"54",
          8433 => x"58",
          8434 => x"74",
          8435 => x"75",
          8436 => x"00",
          8437 => x"54",
          8438 => x"58",
          8439 => x"74",
          8440 => x"75",
          8441 => x"00",
          8442 => x"74",
          8443 => x"20",
          8444 => x"74",
          8445 => x"72",
          8446 => x"0a",
          8447 => x"00",
          8448 => x"62",
          8449 => x"67",
          8450 => x"6d",
          8451 => x"2e",
          8452 => x"00",
          8453 => x"00",
          8454 => x"6c",
          8455 => x"74",
          8456 => x"6e",
          8457 => x"61",
          8458 => x"65",
          8459 => x"20",
          8460 => x"64",
          8461 => x"20",
          8462 => x"61",
          8463 => x"69",
          8464 => x"20",
          8465 => x"75",
          8466 => x"79",
          8467 => x"00",
          8468 => x"00",
          8469 => x"20",
          8470 => x"6b",
          8471 => x"21",
          8472 => x"00",
          8473 => x"74",
          8474 => x"69",
          8475 => x"2e",
          8476 => x"00",
          8477 => x"6c",
          8478 => x"74",
          8479 => x"6e",
          8480 => x"61",
          8481 => x"65",
          8482 => x"00",
          8483 => x"25",
          8484 => x"00",
          8485 => x"00",
          8486 => x"61",
          8487 => x"6e",
          8488 => x"6e",
          8489 => x"72",
          8490 => x"73",
          8491 => x"00",
          8492 => x"62",
          8493 => x"67",
          8494 => x"74",
          8495 => x"75",
          8496 => x"0a",
          8497 => x"00",
          8498 => x"61",
          8499 => x"64",
          8500 => x"72",
          8501 => x"69",
          8502 => x"00",
          8503 => x"62",
          8504 => x"67",
          8505 => x"72",
          8506 => x"69",
          8507 => x"00",
          8508 => x"63",
          8509 => x"6e",
          8510 => x"6f",
          8511 => x"40",
          8512 => x"38",
          8513 => x"2e",
          8514 => x"00",
          8515 => x"6c",
          8516 => x"20",
          8517 => x"65",
          8518 => x"25",
          8519 => x"20",
          8520 => x"0a",
          8521 => x"00",
          8522 => x"6c",
          8523 => x"74",
          8524 => x"65",
          8525 => x"6f",
          8526 => x"28",
          8527 => x"2e",
          8528 => x"00",
          8529 => x"74",
          8530 => x"69",
          8531 => x"61",
          8532 => x"69",
          8533 => x"69",
          8534 => x"2e",
          8535 => x"00",
          8536 => x"64",
          8537 => x"62",
          8538 => x"69",
          8539 => x"2e",
          8540 => x"00",
          8541 => x"00",
          8542 => x"00",
          8543 => x"5c",
          8544 => x"25",
          8545 => x"73",
          8546 => x"00",
          8547 => x"20",
          8548 => x"6d",
          8549 => x"2e",
          8550 => x"00",
          8551 => x"6e",
          8552 => x"2e",
          8553 => x"00",
          8554 => x"62",
          8555 => x"67",
          8556 => x"74",
          8557 => x"75",
          8558 => x"2e",
          8559 => x"00",
          8560 => x"00",
          8561 => x"00",
          8562 => x"ff",
          8563 => x"00",
          8564 => x"ff",
          8565 => x"00",
          8566 => x"ff",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"00",
          8572 => x"01",
          8573 => x"01",
          8574 => x"01",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"3c",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"44",
          8583 => x"00",
          8584 => x"00",
          8585 => x"00",
          8586 => x"4c",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"54",
          8591 => x"00",
          8592 => x"00",
          8593 => x"00",
          8594 => x"5c",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"64",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"6c",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"74",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"7c",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"84",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"8c",
          8619 => x"00",
          8620 => x"00",
          8621 => x"00",
          8622 => x"94",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"9c",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"a4",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"ac",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"b4",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"c0",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"c8",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"d0",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"d8",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"e0",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"e8",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"f0",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"f8",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"08",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"10",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"18",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"1c",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"24",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"2c",
          8699 => x"00",
          8700 => x"00",
          8701 => x"00",
          8702 => x"34",
          8703 => x"00",
          8704 => x"00",
          8705 => x"00",
          8706 => x"3c",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"44",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"4c",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"50",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"58",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"64",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"6c",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"74",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"7c",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"84",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"88",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"8c",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"90",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"94",
          8759 => x"00",
          8760 => x"00",
          8761 => x"00",
          8762 => x"98",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"9c",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"a0",
          8771 => x"00",
          8772 => x"00",
          8773 => x"00",
          8774 => x"a4",
          8775 => x"00",
          8776 => x"00",
          8777 => x"00",
          8778 => x"a8",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"b0",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"bc",
          8787 => x"00",
          8788 => x"00",
          8789 => x"00",
          8790 => x"c4",
          8791 => x"00",
          8792 => x"00",
          8793 => x"00",
          8794 => x"c8",
          8795 => x"00",
          8796 => x"00",
          8797 => x"00",
          8798 => x"d0",
          8799 => x"00",
          8800 => x"00",
          8801 => x"00",
          8802 => x"d8",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"e0",
          8807 => x"00",
          8808 => x"00",
          8809 => x"00",
          8810 => x"e8",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"f0",
          8815 => x"00",
          8816 => x"00",
          8817 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"00",
           281 => x"00",
           282 => x"ac",
           283 => x"27",
           284 => x"71",
           285 => x"53",
           286 => x"04",
           287 => x"9e",
           288 => x"08",
           289 => x"fd",
           290 => x"53",
           291 => x"05",
           292 => x"08",
           293 => x"51",
           294 => x"88",
           295 => x"0c",
           296 => x"0d",
           297 => x"94",
           298 => x"0c",
           299 => x"81",
           300 => x"8c",
           301 => x"94",
           302 => x"08",
           303 => x"3f",
           304 => x"88",
           305 => x"3d",
           306 => x"04",
           307 => x"94",
           308 => x"0d",
           309 => x"08",
           310 => x"94",
           311 => x"08",
           312 => x"38",
           313 => x"05",
           314 => x"08",
           315 => x"80",
           316 => x"f4",
           317 => x"08",
           318 => x"88",
           319 => x"94",
           320 => x"0c",
           321 => x"05",
           322 => x"fc",
           323 => x"08",
           324 => x"80",
           325 => x"94",
           326 => x"08",
           327 => x"8c",
           328 => x"0b",
           329 => x"05",
           330 => x"fc",
           331 => x"38",
           332 => x"08",
           333 => x"94",
           334 => x"08",
           335 => x"05",
           336 => x"94",
           337 => x"08",
           338 => x"88",
           339 => x"81",
           340 => x"08",
           341 => x"f8",
           342 => x"94",
           343 => x"08",
           344 => x"38",
           345 => x"05",
           346 => x"08",
           347 => x"94",
           348 => x"08",
           349 => x"54",
           350 => x"94",
           351 => x"08",
           352 => x"fb",
           353 => x"0b",
           354 => x"05",
           355 => x"88",
           356 => x"25",
           357 => x"08",
           358 => x"30",
           359 => x"05",
           360 => x"94",
           361 => x"0c",
           362 => x"05",
           363 => x"8c",
           364 => x"8c",
           365 => x"94",
           366 => x"0c",
           367 => x"08",
           368 => x"52",
           369 => x"05",
           370 => x"3f",
           371 => x"94",
           372 => x"0c",
           373 => x"fc",
           374 => x"2e",
           375 => x"08",
           376 => x"30",
           377 => x"05",
           378 => x"f8",
           379 => x"88",
           380 => x"3d",
           381 => x"04",
           382 => x"94",
           383 => x"0d",
           384 => x"08",
           385 => x"80",
           386 => x"f8",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"94",
           391 => x"08",
           392 => x"38",
           393 => x"08",
           394 => x"24",
           395 => x"08",
           396 => x"10",
           397 => x"05",
           398 => x"fc",
           399 => x"94",
           400 => x"0c",
           401 => x"08",
           402 => x"80",
           403 => x"38",
           404 => x"05",
           405 => x"88",
           406 => x"a1",
           407 => x"88",
           408 => x"08",
           409 => x"31",
           410 => x"05",
           411 => x"f8",
           412 => x"08",
           413 => x"07",
           414 => x"05",
           415 => x"fc",
           416 => x"2a",
           417 => x"05",
           418 => x"8c",
           419 => x"2a",
           420 => x"05",
           421 => x"39",
           422 => x"05",
           423 => x"8f",
           424 => x"88",
           425 => x"94",
           426 => x"0c",
           427 => x"94",
           428 => x"08",
           429 => x"f4",
           430 => x"94",
           431 => x"08",
           432 => x"3d",
           433 => x"04",
           434 => x"81",
           435 => x"c0",
           436 => x"81",
           437 => x"92",
           438 => x"0b",
           439 => x"8c",
           440 => x"92",
           441 => x"82",
           442 => x"70",
           443 => x"38",
           444 => x"8c",
           445 => x"e9",
           446 => x"92",
           447 => x"80",
           448 => x"71",
           449 => x"c0",
           450 => x"51",
           451 => x"88",
           452 => x"0b",
           453 => x"34",
           454 => x"9f",
           455 => x"0c",
           456 => x"04",
           457 => x"78",
           458 => x"58",
           459 => x"0b",
           460 => x"a8",
           461 => x"52",
           462 => x"70",
           463 => x"81",
           464 => x"38",
           465 => x"c0",
           466 => x"79",
           467 => x"80",
           468 => x"87",
           469 => x"0c",
           470 => x"8c",
           471 => x"2a",
           472 => x"51",
           473 => x"80",
           474 => x"87",
           475 => x"08",
           476 => x"06",
           477 => x"52",
           478 => x"80",
           479 => x"70",
           480 => x"38",
           481 => x"81",
           482 => x"ff",
           483 => x"15",
           484 => x"06",
           485 => x"2e",
           486 => x"c0",
           487 => x"51",
           488 => x"38",
           489 => x"8c",
           490 => x"95",
           491 => x"87",
           492 => x"0c",
           493 => x"8c",
           494 => x"06",
           495 => x"f4",
           496 => x"fc",
           497 => x"52",
           498 => x"2e",
           499 => x"8f",
           500 => x"98",
           501 => x"70",
           502 => x"81",
           503 => x"81",
           504 => x"0c",
           505 => x"04",
           506 => x"74",
           507 => x"71",
           508 => x"2b",
           509 => x"53",
           510 => x"0d",
           511 => x"0d",
           512 => x"33",
           513 => x"71",
           514 => x"88",
           515 => x"14",
           516 => x"07",
           517 => x"33",
           518 => x"0c",
           519 => x"56",
           520 => x"3d",
           521 => x"3d",
           522 => x"0b",
           523 => x"08",
           524 => x"77",
           525 => x"38",
           526 => x"08",
           527 => x"38",
           528 => x"74",
           529 => x"38",
           530 => x"ae",
           531 => x"39",
           532 => x"10",
           533 => x"53",
           534 => x"8c",
           535 => x"52",
           536 => x"52",
           537 => x"3f",
           538 => x"38",
           539 => x"f8",
           540 => x"83",
           541 => x"55",
           542 => x"54",
           543 => x"83",
           544 => x"76",
           545 => x"17",
           546 => x"88",
           547 => x"55",
           548 => x"88",
           549 => x"74",
           550 => x"3f",
           551 => x"0a",
           552 => x"39",
           553 => x"88",
           554 => x"0d",
           555 => x"0d",
           556 => x"9f",
           557 => x"19",
           558 => x"fe",
           559 => x"54",
           560 => x"73",
           561 => x"82",
           562 => x"71",
           563 => x"08",
           564 => x"75",
           565 => x"3d",
           566 => x"3d",
           567 => x"80",
           568 => x"0b",
           569 => x"70",
           570 => x"53",
           571 => x"09",
           572 => x"38",
           573 => x"fd",
           574 => x"08",
           575 => x"9a",
           576 => x"e4",
           577 => x"83",
           578 => x"73",
           579 => x"85",
           580 => x"fc",
           581 => x"0b",
           582 => x"ac",
           583 => x"80",
           584 => x"15",
           585 => x"81",
           586 => x"88",
           587 => x"26",
           588 => x"52",
           589 => x"90",
           590 => x"52",
           591 => x"09",
           592 => x"38",
           593 => x"53",
           594 => x"0c",
           595 => x"8b",
           596 => x"fe",
           597 => x"08",
           598 => x"90",
           599 => x"71",
           600 => x"80",
           601 => x"0c",
           602 => x"04",
           603 => x"78",
           604 => x"9f",
           605 => x"22",
           606 => x"83",
           607 => x"57",
           608 => x"73",
           609 => x"38",
           610 => x"53",
           611 => x"83",
           612 => x"39",
           613 => x"52",
           614 => x"38",
           615 => x"16",
           616 => x"08",
           617 => x"38",
           618 => x"17",
           619 => x"73",
           620 => x"38",
           621 => x"16",
           622 => x"74",
           623 => x"52",
           624 => x"72",
           625 => x"3f",
           626 => x"88",
           627 => x"38",
           628 => x"08",
           629 => x"27",
           630 => x"08",
           631 => x"88",
           632 => x"c9",
           633 => x"90",
           634 => x"75",
           635 => x"71",
           636 => x"3d",
           637 => x"3d",
           638 => x"64",
           639 => x"75",
           640 => x"a0",
           641 => x"06",
           642 => x"16",
           643 => x"ef",
           644 => x"33",
           645 => x"af",
           646 => x"06",
           647 => x"16",
           648 => x"88",
           649 => x"70",
           650 => x"74",
           651 => x"38",
           652 => x"df",
           653 => x"56",
           654 => x"82",
           655 => x"3d",
           656 => x"70",
           657 => x"8a",
           658 => x"70",
           659 => x"34",
           660 => x"74",
           661 => x"81",
           662 => x"80",
           663 => x"88",
           664 => x"5a",
           665 => x"70",
           666 => x"60",
           667 => x"70",
           668 => x"30",
           669 => x"71",
           670 => x"51",
           671 => x"53",
           672 => x"74",
           673 => x"76",
           674 => x"81",
           675 => x"81",
           676 => x"27",
           677 => x"74",
           678 => x"38",
           679 => x"70",
           680 => x"32",
           681 => x"73",
           682 => x"53",
           683 => x"56",
           684 => x"88",
           685 => x"ff",
           686 => x"81",
           687 => x"ff",
           688 => x"53",
           689 => x"76",
           690 => x"98",
           691 => x"7f",
           692 => x"76",
           693 => x"38",
           694 => x"8b",
           695 => x"51",
           696 => x"88",
           697 => x"38",
           698 => x"22",
           699 => x"83",
           700 => x"55",
           701 => x"52",
           702 => x"a8",
           703 => x"57",
           704 => x"fb",
           705 => x"55",
           706 => x"80",
           707 => x"1d",
           708 => x"2a",
           709 => x"51",
           710 => x"b2",
           711 => x"84",
           712 => x"08",
           713 => x"58",
           714 => x"77",
           715 => x"38",
           716 => x"05",
           717 => x"70",
           718 => x"33",
           719 => x"52",
           720 => x"80",
           721 => x"86",
           722 => x"2e",
           723 => x"51",
           724 => x"ff",
           725 => x"08",
           726 => x"b4",
           727 => x"76",
           728 => x"08",
           729 => x"51",
           730 => x"38",
           731 => x"70",
           732 => x"81",
           733 => x"56",
           734 => x"83",
           735 => x"81",
           736 => x"7c",
           737 => x"3f",
           738 => x"1d",
           739 => x"39",
           740 => x"90",
           741 => x"f9",
           742 => x"7b",
           743 => x"54",
           744 => x"77",
           745 => x"f6",
           746 => x"56",
           747 => x"e7",
           748 => x"f8",
           749 => x"08",
           750 => x"06",
           751 => x"74",
           752 => x"2e",
           753 => x"80",
           754 => x"54",
           755 => x"52",
           756 => x"d0",
           757 => x"56",
           758 => x"38",
           759 => x"88",
           760 => x"83",
           761 => x"55",
           762 => x"c6",
           763 => x"82",
           764 => x"53",
           765 => x"51",
           766 => x"88",
           767 => x"08",
           768 => x"51",
           769 => x"88",
           770 => x"ff",
           771 => x"81",
           772 => x"83",
           773 => x"75",
           774 => x"3d",
           775 => x"3d",
           776 => x"80",
           777 => x"0b",
           778 => x"f5",
           779 => x"08",
           780 => x"82",
           781 => x"f2",
           782 => x"53",
           783 => x"53",
           784 => x"d3",
           785 => x"81",
           786 => x"76",
           787 => x"81",
           788 => x"90",
           789 => x"53",
           790 => x"51",
           791 => x"88",
           792 => x"8d",
           793 => x"74",
           794 => x"38",
           795 => x"05",
           796 => x"3f",
           797 => x"08",
           798 => x"5a",
           799 => x"88",
           800 => x"06",
           801 => x"2e",
           802 => x"86",
           803 => x"82",
           804 => x"80",
           805 => x"86",
           806 => x"39",
           807 => x"53",
           808 => x"51",
           809 => x"81",
           810 => x"81",
           811 => x"3d",
           812 => x"f6",
           813 => x"08",
           814 => x"06",
           815 => x"38",
           816 => x"05",
           817 => x"3f",
           818 => x"02",
           819 => x"78",
           820 => x"88",
           821 => x"70",
           822 => x"5b",
           823 => x"88",
           824 => x"ff",
           825 => x"8c",
           826 => x"3d",
           827 => x"34",
           828 => x"05",
           829 => x"3f",
           830 => x"1a",
           831 => x"e2",
           832 => x"e4",
           833 => x"83",
           834 => x"56",
           835 => x"95",
           836 => x"51",
           837 => x"88",
           838 => x"51",
           839 => x"88",
           840 => x"ff",
           841 => x"31",
           842 => x"1b",
           843 => x"2a",
           844 => x"56",
           845 => x"55",
           846 => x"55",
           847 => x"88",
           848 => x"70",
           849 => x"88",
           850 => x"05",
           851 => x"83",
           852 => x"83",
           853 => x"83",
           854 => x"27",
           855 => x"57",
           856 => x"56",
           857 => x"80",
           858 => x"79",
           859 => x"2e",
           860 => x"90",
           861 => x"fb",
           862 => x"81",
           863 => x"90",
           864 => x"39",
           865 => x"18",
           866 => x"79",
           867 => x"06",
           868 => x"19",
           869 => x"05",
           870 => x"55",
           871 => x"1a",
           872 => x"0b",
           873 => x"0c",
           874 => x"88",
           875 => x"0d",
           876 => x"0d",
           877 => x"9f",
           878 => x"85",
           879 => x"2e",
           880 => x"80",
           881 => x"34",
           882 => x"11",
           883 => x"89",
           884 => x"57",
           885 => x"f8",
           886 => x"08",
           887 => x"80",
           888 => x"3d",
           889 => x"80",
           890 => x"02",
           891 => x"70",
           892 => x"81",
           893 => x"57",
           894 => x"85",
           895 => x"a1",
           896 => x"f5",
           897 => x"08",
           898 => x"98",
           899 => x"51",
           900 => x"88",
           901 => x"0c",
           902 => x"0c",
           903 => x"16",
           904 => x"0c",
           905 => x"04",
           906 => x"7d",
           907 => x"0b",
           908 => x"08",
           909 => x"58",
           910 => x"85",
           911 => x"2e",
           912 => x"81",
           913 => x"06",
           914 => x"74",
           915 => x"c3",
           916 => x"74",
           917 => x"86",
           918 => x"81",
           919 => x"57",
           920 => x"9c",
           921 => x"17",
           922 => x"74",
           923 => x"38",
           924 => x"80",
           925 => x"38",
           926 => x"70",
           927 => x"56",
           928 => x"c7",
           929 => x"33",
           930 => x"89",
           931 => x"81",
           932 => x"55",
           933 => x"76",
           934 => x"16",
           935 => x"39",
           936 => x"51",
           937 => x"88",
           938 => x"75",
           939 => x"38",
           940 => x"0c",
           941 => x"51",
           942 => x"88",
           943 => x"08",
           944 => x"8f",
           945 => x"1a",
           946 => x"98",
           947 => x"ff",
           948 => x"71",
           949 => x"77",
           950 => x"38",
           951 => x"54",
           952 => x"83",
           953 => x"a8",
           954 => x"78",
           955 => x"3f",
           956 => x"e5",
           957 => x"08",
           958 => x"0c",
           959 => x"7b",
           960 => x"0c",
           961 => x"2e",
           962 => x"74",
           963 => x"e2",
           964 => x"76",
           965 => x"3d",
           966 => x"3d",
           967 => x"86",
           968 => x"c0",
           969 => x"9b",
           970 => x"0b",
           971 => x"9c",
           972 => x"83",
           973 => x"94",
           974 => x"80",
           975 => x"c0",
           976 => x"9f",
           977 => x"d6",
           978 => x"b8",
           979 => x"51",
           980 => x"88",
           981 => x"a0",
           982 => x"08",
           983 => x"88",
           984 => x"3d",
           985 => x"84",
           986 => x"51",
           987 => x"88",
           988 => x"75",
           989 => x"2e",
           990 => x"15",
           991 => x"a0",
           992 => x"04",
           993 => x"39",
           994 => x"ff",
           995 => x"ff",
           996 => x"00",
           997 => x"ff",
           998 => x"4f",
           999 => x"4e",
          1000 => x"4f",
          1001 => x"00",
          1002 => x"00",
          2048 => x"80",
          2049 => x"0b",
          2050 => x"95",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"80",
          2057 => x"0b",
          2058 => x"85",
          2059 => x"80",
          2060 => x"0b",
          2061 => x"a5",
          2062 => x"80",
          2063 => x"0b",
          2064 => x"c5",
          2065 => x"80",
          2066 => x"0b",
          2067 => x"e5",
          2068 => x"80",
          2069 => x"0b",
          2070 => x"85",
          2071 => x"80",
          2072 => x"0b",
          2073 => x"a5",
          2074 => x"80",
          2075 => x"0b",
          2076 => x"c5",
          2077 => x"80",
          2078 => x"0b",
          2079 => x"e5",
          2080 => x"80",
          2081 => x"0b",
          2082 => x"85",
          2083 => x"80",
          2084 => x"0b",
          2085 => x"a5",
          2086 => x"80",
          2087 => x"0b",
          2088 => x"c5",
          2089 => x"80",
          2090 => x"0b",
          2091 => x"e5",
          2092 => x"80",
          2093 => x"0b",
          2094 => x"85",
          2095 => x"80",
          2096 => x"0b",
          2097 => x"a5",
          2098 => x"80",
          2099 => x"0b",
          2100 => x"c5",
          2101 => x"80",
          2102 => x"0b",
          2103 => x"e5",
          2104 => x"80",
          2105 => x"0b",
          2106 => x"85",
          2107 => x"80",
          2108 => x"0b",
          2109 => x"a5",
          2110 => x"80",
          2111 => x"0b",
          2112 => x"c5",
          2113 => x"80",
          2114 => x"0b",
          2115 => x"e5",
          2116 => x"80",
          2117 => x"0b",
          2118 => x"85",
          2119 => x"80",
          2120 => x"0b",
          2121 => x"a5",
          2122 => x"80",
          2123 => x"0b",
          2124 => x"c5",
          2125 => x"80",
          2126 => x"0b",
          2127 => x"e5",
          2128 => x"80",
          2129 => x"0b",
          2130 => x"85",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"c4",
          2177 => x"93",
          2178 => x"d5",
          2179 => x"93",
          2180 => x"80",
          2181 => x"93",
          2182 => x"df",
          2183 => x"93",
          2184 => x"80",
          2185 => x"93",
          2186 => x"e0",
          2187 => x"93",
          2188 => x"80",
          2189 => x"93",
          2190 => x"e0",
          2191 => x"93",
          2192 => x"80",
          2193 => x"93",
          2194 => x"e6",
          2195 => x"93",
          2196 => x"80",
          2197 => x"93",
          2198 => x"e8",
          2199 => x"93",
          2200 => x"80",
          2201 => x"93",
          2202 => x"e0",
          2203 => x"93",
          2204 => x"80",
          2205 => x"93",
          2206 => x"e8",
          2207 => x"93",
          2208 => x"80",
          2209 => x"93",
          2210 => x"ea",
          2211 => x"93",
          2212 => x"80",
          2213 => x"93",
          2214 => x"e6",
          2215 => x"93",
          2216 => x"80",
          2217 => x"93",
          2218 => x"e6",
          2219 => x"93",
          2220 => x"80",
          2221 => x"93",
          2222 => x"e6",
          2223 => x"93",
          2224 => x"80",
          2225 => x"93",
          2226 => x"d7",
          2227 => x"93",
          2228 => x"80",
          2229 => x"93",
          2230 => x"d7",
          2231 => x"93",
          2232 => x"80",
          2233 => x"93",
          2234 => x"cf",
          2235 => x"93",
          2236 => x"80",
          2237 => x"93",
          2238 => x"d1",
          2239 => x"93",
          2240 => x"80",
          2241 => x"93",
          2242 => x"d2",
          2243 => x"93",
          2244 => x"80",
          2245 => x"93",
          2246 => x"9e",
          2247 => x"93",
          2248 => x"80",
          2249 => x"93",
          2250 => x"ad",
          2251 => x"93",
          2252 => x"80",
          2253 => x"93",
          2254 => x"a3",
          2255 => x"93",
          2256 => x"80",
          2257 => x"93",
          2258 => x"a7",
          2259 => x"93",
          2260 => x"80",
          2261 => x"93",
          2262 => x"b3",
          2263 => x"93",
          2264 => x"80",
          2265 => x"93",
          2266 => x"bd",
          2267 => x"93",
          2268 => x"80",
          2269 => x"93",
          2270 => x"ac",
          2271 => x"93",
          2272 => x"80",
          2273 => x"93",
          2274 => x"b7",
          2275 => x"93",
          2276 => x"80",
          2277 => x"93",
          2278 => x"b8",
          2279 => x"93",
          2280 => x"80",
          2281 => x"93",
          2282 => x"b9",
          2283 => x"93",
          2284 => x"80",
          2285 => x"93",
          2286 => x"c2",
          2287 => x"93",
          2288 => x"80",
          2289 => x"93",
          2290 => x"bf",
          2291 => x"93",
          2292 => x"80",
          2293 => x"93",
          2294 => x"c4",
          2295 => x"93",
          2296 => x"80",
          2297 => x"93",
          2298 => x"ba",
          2299 => x"93",
          2300 => x"80",
          2301 => x"93",
          2302 => x"c7",
          2303 => x"93",
          2304 => x"80",
          2305 => x"93",
          2306 => x"c8",
          2307 => x"93",
          2308 => x"80",
          2309 => x"93",
          2310 => x"ae",
          2311 => x"93",
          2312 => x"80",
          2313 => x"93",
          2314 => x"ae",
          2315 => x"93",
          2316 => x"80",
          2317 => x"93",
          2318 => x"af",
          2319 => x"93",
          2320 => x"80",
          2321 => x"93",
          2322 => x"ba",
          2323 => x"93",
          2324 => x"80",
          2325 => x"93",
          2326 => x"c9",
          2327 => x"93",
          2328 => x"80",
          2329 => x"93",
          2330 => x"cc",
          2331 => x"93",
          2332 => x"80",
          2333 => x"93",
          2334 => x"cf",
          2335 => x"93",
          2336 => x"80",
          2337 => x"93",
          2338 => x"9e",
          2339 => x"93",
          2340 => x"80",
          2341 => x"93",
          2342 => x"d2",
          2343 => x"93",
          2344 => x"80",
          2345 => x"93",
          2346 => x"ed",
          2347 => x"93",
          2348 => x"80",
          2349 => x"93",
          2350 => x"ef",
          2351 => x"93",
          2352 => x"80",
          2353 => x"93",
          2354 => x"f1",
          2355 => x"93",
          2356 => x"80",
          2357 => x"93",
          2358 => x"d0",
          2359 => x"93",
          2360 => x"80",
          2361 => x"93",
          2362 => x"d0",
          2363 => x"93",
          2364 => x"80",
          2365 => x"93",
          2366 => x"d3",
          2367 => x"93",
          2368 => x"80",
          2369 => x"93",
          2370 => x"df",
          2371 => x"93",
          2372 => x"80",
          2373 => x"93",
          2374 => x"b6",
          2375 => x"38",
          2376 => x"84",
          2377 => x"0b",
          2378 => x"98",
          2379 => x"80",
          2380 => x"da",
          2381 => x"82",
          2382 => x"02",
          2383 => x"0c",
          2384 => x"80",
          2385 => x"d4",
          2386 => x"08",
          2387 => x"d4",
          2388 => x"08",
          2389 => x"3f",
          2390 => x"08",
          2391 => x"c8",
          2392 => x"3d",
          2393 => x"d4",
          2394 => x"93",
          2395 => x"82",
          2396 => x"fd",
          2397 => x"53",
          2398 => x"08",
          2399 => x"52",
          2400 => x"08",
          2401 => x"51",
          2402 => x"93",
          2403 => x"82",
          2404 => x"54",
          2405 => x"82",
          2406 => x"04",
          2407 => x"08",
          2408 => x"d4",
          2409 => x"0d",
          2410 => x"93",
          2411 => x"05",
          2412 => x"82",
          2413 => x"f8",
          2414 => x"93",
          2415 => x"05",
          2416 => x"d4",
          2417 => x"08",
          2418 => x"82",
          2419 => x"fc",
          2420 => x"2e",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"24",
          2424 => x"93",
          2425 => x"05",
          2426 => x"93",
          2427 => x"05",
          2428 => x"d4",
          2429 => x"08",
          2430 => x"d4",
          2431 => x"0c",
          2432 => x"82",
          2433 => x"fc",
          2434 => x"2e",
          2435 => x"82",
          2436 => x"8c",
          2437 => x"93",
          2438 => x"05",
          2439 => x"38",
          2440 => x"08",
          2441 => x"82",
          2442 => x"8c",
          2443 => x"82",
          2444 => x"88",
          2445 => x"93",
          2446 => x"05",
          2447 => x"d4",
          2448 => x"08",
          2449 => x"d4",
          2450 => x"0c",
          2451 => x"08",
          2452 => x"81",
          2453 => x"d4",
          2454 => x"0c",
          2455 => x"08",
          2456 => x"81",
          2457 => x"d4",
          2458 => x"0c",
          2459 => x"82",
          2460 => x"90",
          2461 => x"2e",
          2462 => x"93",
          2463 => x"05",
          2464 => x"93",
          2465 => x"05",
          2466 => x"39",
          2467 => x"08",
          2468 => x"70",
          2469 => x"08",
          2470 => x"51",
          2471 => x"08",
          2472 => x"82",
          2473 => x"85",
          2474 => x"93",
          2475 => x"fc",
          2476 => x"79",
          2477 => x"05",
          2478 => x"57",
          2479 => x"83",
          2480 => x"38",
          2481 => x"51",
          2482 => x"a4",
          2483 => x"52",
          2484 => x"93",
          2485 => x"70",
          2486 => x"34",
          2487 => x"71",
          2488 => x"81",
          2489 => x"74",
          2490 => x"0c",
          2491 => x"04",
          2492 => x"2b",
          2493 => x"71",
          2494 => x"51",
          2495 => x"72",
          2496 => x"72",
          2497 => x"05",
          2498 => x"71",
          2499 => x"53",
          2500 => x"70",
          2501 => x"0c",
          2502 => x"84",
          2503 => x"f0",
          2504 => x"8f",
          2505 => x"83",
          2506 => x"38",
          2507 => x"84",
          2508 => x"fc",
          2509 => x"83",
          2510 => x"70",
          2511 => x"39",
          2512 => x"77",
          2513 => x"07",
          2514 => x"54",
          2515 => x"38",
          2516 => x"08",
          2517 => x"71",
          2518 => x"80",
          2519 => x"75",
          2520 => x"33",
          2521 => x"06",
          2522 => x"80",
          2523 => x"72",
          2524 => x"75",
          2525 => x"06",
          2526 => x"12",
          2527 => x"33",
          2528 => x"06",
          2529 => x"52",
          2530 => x"72",
          2531 => x"81",
          2532 => x"81",
          2533 => x"71",
          2534 => x"c8",
          2535 => x"87",
          2536 => x"71",
          2537 => x"fb",
          2538 => x"06",
          2539 => x"82",
          2540 => x"51",
          2541 => x"97",
          2542 => x"84",
          2543 => x"54",
          2544 => x"75",
          2545 => x"38",
          2546 => x"52",
          2547 => x"80",
          2548 => x"c8",
          2549 => x"0d",
          2550 => x"0d",
          2551 => x"52",
          2552 => x"52",
          2553 => x"82",
          2554 => x"81",
          2555 => x"07",
          2556 => x"52",
          2557 => x"e8",
          2558 => x"93",
          2559 => x"3d",
          2560 => x"3d",
          2561 => x"08",
          2562 => x"55",
          2563 => x"80",
          2564 => x"33",
          2565 => x"2e",
          2566 => x"8c",
          2567 => x"70",
          2568 => x"70",
          2569 => x"38",
          2570 => x"39",
          2571 => x"80",
          2572 => x"53",
          2573 => x"83",
          2574 => x"70",
          2575 => x"2a",
          2576 => x"51",
          2577 => x"71",
          2578 => x"a0",
          2579 => x"06",
          2580 => x"72",
          2581 => x"54",
          2582 => x"0c",
          2583 => x"82",
          2584 => x"86",
          2585 => x"fc",
          2586 => x"53",
          2587 => x"2e",
          2588 => x"3d",
          2589 => x"72",
          2590 => x"3f",
          2591 => x"08",
          2592 => x"53",
          2593 => x"53",
          2594 => x"c8",
          2595 => x"0d",
          2596 => x"0d",
          2597 => x"33",
          2598 => x"5c",
          2599 => x"8b",
          2600 => x"38",
          2601 => x"ff",
          2602 => x"5b",
          2603 => x"81",
          2604 => x"1c",
          2605 => x"5b",
          2606 => x"81",
          2607 => x"1c",
          2608 => x"5b",
          2609 => x"81",
          2610 => x"1c",
          2611 => x"5b",
          2612 => x"81",
          2613 => x"1c",
          2614 => x"5b",
          2615 => x"26",
          2616 => x"8a",
          2617 => x"87",
          2618 => x"e7",
          2619 => x"38",
          2620 => x"59",
          2621 => x"58",
          2622 => x"57",
          2623 => x"56",
          2624 => x"55",
          2625 => x"54",
          2626 => x"53",
          2627 => x"81",
          2628 => x"94",
          2629 => x"c0",
          2630 => x"81",
          2631 => x"22",
          2632 => x"bc",
          2633 => x"33",
          2634 => x"b8",
          2635 => x"33",
          2636 => x"b4",
          2637 => x"33",
          2638 => x"b0",
          2639 => x"33",
          2640 => x"ac",
          2641 => x"33",
          2642 => x"a8",
          2643 => x"22",
          2644 => x"a4",
          2645 => x"22",
          2646 => x"a0",
          2647 => x"0c",
          2648 => x"82",
          2649 => x"8d",
          2650 => x"f5",
          2651 => x"5a",
          2652 => x"9c",
          2653 => x"0c",
          2654 => x"bc",
          2655 => x"7a",
          2656 => x"98",
          2657 => x"7a",
          2658 => x"87",
          2659 => x"08",
          2660 => x"1b",
          2661 => x"98",
          2662 => x"7a",
          2663 => x"87",
          2664 => x"08",
          2665 => x"1b",
          2666 => x"98",
          2667 => x"7a",
          2668 => x"87",
          2669 => x"08",
          2670 => x"1b",
          2671 => x"98",
          2672 => x"7a",
          2673 => x"80",
          2674 => x"1a",
          2675 => x"1a",
          2676 => x"1a",
          2677 => x"1a",
          2678 => x"1a",
          2679 => x"1a",
          2680 => x"1a",
          2681 => x"22",
          2682 => x"a8",
          2683 => x"3f",
          2684 => x"04",
          2685 => x"02",
          2686 => x"70",
          2687 => x"2a",
          2688 => x"70",
          2689 => x"8b",
          2690 => x"3d",
          2691 => x"3d",
          2692 => x"0b",
          2693 => x"33",
          2694 => x"c0",
          2695 => x"72",
          2696 => x"38",
          2697 => x"94",
          2698 => x"70",
          2699 => x"81",
          2700 => x"52",
          2701 => x"8c",
          2702 => x"2a",
          2703 => x"51",
          2704 => x"38",
          2705 => x"81",
          2706 => x"06",
          2707 => x"80",
          2708 => x"71",
          2709 => x"81",
          2710 => x"70",
          2711 => x"0b",
          2712 => x"c0",
          2713 => x"c0",
          2714 => x"70",
          2715 => x"38",
          2716 => x"90",
          2717 => x"0c",
          2718 => x"c8",
          2719 => x"0d",
          2720 => x"0d",
          2721 => x"33",
          2722 => x"8b",
          2723 => x"54",
          2724 => x"84",
          2725 => x"2e",
          2726 => x"c0",
          2727 => x"70",
          2728 => x"2a",
          2729 => x"51",
          2730 => x"80",
          2731 => x"71",
          2732 => x"81",
          2733 => x"70",
          2734 => x"96",
          2735 => x"70",
          2736 => x"51",
          2737 => x"8d",
          2738 => x"2a",
          2739 => x"51",
          2740 => x"bc",
          2741 => x"82",
          2742 => x"51",
          2743 => x"80",
          2744 => x"2e",
          2745 => x"c0",
          2746 => x"73",
          2747 => x"3d",
          2748 => x"3d",
          2749 => x"80",
          2750 => x"56",
          2751 => x"80",
          2752 => x"70",
          2753 => x"33",
          2754 => x"8b",
          2755 => x"55",
          2756 => x"84",
          2757 => x"2e",
          2758 => x"c0",
          2759 => x"70",
          2760 => x"2a",
          2761 => x"51",
          2762 => x"80",
          2763 => x"71",
          2764 => x"81",
          2765 => x"70",
          2766 => x"96",
          2767 => x"70",
          2768 => x"51",
          2769 => x"8d",
          2770 => x"2a",
          2771 => x"51",
          2772 => x"bc",
          2773 => x"82",
          2774 => x"51",
          2775 => x"80",
          2776 => x"2e",
          2777 => x"c0",
          2778 => x"74",
          2779 => x"16",
          2780 => x"56",
          2781 => x"38",
          2782 => x"c8",
          2783 => x"0d",
          2784 => x"0d",
          2785 => x"8b",
          2786 => x"87",
          2787 => x"51",
          2788 => x"86",
          2789 => x"94",
          2790 => x"08",
          2791 => x"70",
          2792 => x"51",
          2793 => x"2e",
          2794 => x"0b",
          2795 => x"33",
          2796 => x"94",
          2797 => x"80",
          2798 => x"87",
          2799 => x"52",
          2800 => x"81",
          2801 => x"93",
          2802 => x"83",
          2803 => x"ff",
          2804 => x"0b",
          2805 => x"33",
          2806 => x"94",
          2807 => x"80",
          2808 => x"87",
          2809 => x"52",
          2810 => x"82",
          2811 => x"06",
          2812 => x"ff",
          2813 => x"2e",
          2814 => x"0b",
          2815 => x"33",
          2816 => x"94",
          2817 => x"80",
          2818 => x"87",
          2819 => x"52",
          2820 => x"98",
          2821 => x"2c",
          2822 => x"71",
          2823 => x"0c",
          2824 => x"04",
          2825 => x"87",
          2826 => x"70",
          2827 => x"2a",
          2828 => x"52",
          2829 => x"2e",
          2830 => x"82",
          2831 => x"87",
          2832 => x"08",
          2833 => x"11",
          2834 => x"a0",
          2835 => x"52",
          2836 => x"c0",
          2837 => x"71",
          2838 => x"11",
          2839 => x"90",
          2840 => x"52",
          2841 => x"c0",
          2842 => x"71",
          2843 => x"11",
          2844 => x"98",
          2845 => x"52",
          2846 => x"c0",
          2847 => x"71",
          2848 => x"11",
          2849 => x"a8",
          2850 => x"52",
          2851 => x"c0",
          2852 => x"71",
          2853 => x"08",
          2854 => x"a4",
          2855 => x"12",
          2856 => x"84",
          2857 => x"51",
          2858 => x"13",
          2859 => x"52",
          2860 => x"c0",
          2861 => x"70",
          2862 => x"51",
          2863 => x"80",
          2864 => x"81",
          2865 => x"34",
          2866 => x"c0",
          2867 => x"70",
          2868 => x"06",
          2869 => x"70",
          2870 => x"38",
          2871 => x"82",
          2872 => x"80",
          2873 => x"9e",
          2874 => x"80",
          2875 => x"51",
          2876 => x"80",
          2877 => x"81",
          2878 => x"8b",
          2879 => x"0b",
          2880 => x"88",
          2881 => x"80",
          2882 => x"52",
          2883 => x"83",
          2884 => x"71",
          2885 => x"34",
          2886 => x"c0",
          2887 => x"70",
          2888 => x"51",
          2889 => x"80",
          2890 => x"81",
          2891 => x"8b",
          2892 => x"0b",
          2893 => x"88",
          2894 => x"80",
          2895 => x"52",
          2896 => x"83",
          2897 => x"71",
          2898 => x"34",
          2899 => x"c0",
          2900 => x"70",
          2901 => x"51",
          2902 => x"80",
          2903 => x"81",
          2904 => x"8b",
          2905 => x"0b",
          2906 => x"88",
          2907 => x"80",
          2908 => x"52",
          2909 => x"83",
          2910 => x"71",
          2911 => x"34",
          2912 => x"52",
          2913 => x"88",
          2914 => x"80",
          2915 => x"86",
          2916 => x"52",
          2917 => x"70",
          2918 => x"34",
          2919 => x"73",
          2920 => x"06",
          2921 => x"70",
          2922 => x"38",
          2923 => x"74",
          2924 => x"87",
          2925 => x"08",
          2926 => x"51",
          2927 => x"80",
          2928 => x"81",
          2929 => x"8b",
          2930 => x"c0",
          2931 => x"70",
          2932 => x"51",
          2933 => x"fc",
          2934 => x"0d",
          2935 => x"0d",
          2936 => x"51",
          2937 => x"82",
          2938 => x"54",
          2939 => x"88",
          2940 => x"d4",
          2941 => x"3f",
          2942 => x"51",
          2943 => x"82",
          2944 => x"33",
          2945 => x"80",
          2946 => x"d7",
          2947 => x"82",
          2948 => x"52",
          2949 => x"51",
          2950 => x"82",
          2951 => x"33",
          2952 => x"80",
          2953 => x"de",
          2954 => x"da",
          2955 => x"81",
          2956 => x"89",
          2957 => x"8b",
          2958 => x"55",
          2959 => x"38",
          2960 => x"54",
          2961 => x"93",
          2962 => x"d8",
          2963 => x"fc",
          2964 => x"54",
          2965 => x"51",
          2966 => x"82",
          2967 => x"54",
          2968 => x"88",
          2969 => x"f0",
          2970 => x"3f",
          2971 => x"33",
          2972 => x"2e",
          2973 => x"f7",
          2974 => x"a8",
          2975 => x"f7",
          2976 => x"80",
          2977 => x"81",
          2978 => x"83",
          2979 => x"8b",
          2980 => x"55",
          2981 => x"2e",
          2982 => x"15",
          2983 => x"f8",
          2984 => x"fa",
          2985 => x"fa",
          2986 => x"80",
          2987 => x"81",
          2988 => x"82",
          2989 => x"8b",
          2990 => x"55",
          2991 => x"2e",
          2992 => x"15",
          2993 => x"f8",
          2994 => x"d2",
          2995 => x"ec",
          2996 => x"3f",
          2997 => x"70",
          2998 => x"05",
          2999 => x"81",
          3000 => x"55",
          3001 => x"3f",
          3002 => x"81",
          3003 => x"88",
          3004 => x"15",
          3005 => x"f9",
          3006 => x"a2",
          3007 => x"22",
          3008 => x"f0",
          3009 => x"3f",
          3010 => x"52",
          3011 => x"51",
          3012 => x"86",
          3013 => x"ff",
          3014 => x"8e",
          3015 => x"71",
          3016 => x"38",
          3017 => x"0b",
          3018 => x"c4",
          3019 => x"08",
          3020 => x"c0",
          3021 => x"3f",
          3022 => x"fa",
          3023 => x"b2",
          3024 => x"81",
          3025 => x"f7",
          3026 => x"39",
          3027 => x"51",
          3028 => x"91",
          3029 => x"dc",
          3030 => x"3f",
          3031 => x"fa",
          3032 => x"8e",
          3033 => x"0d",
          3034 => x"80",
          3035 => x"0b",
          3036 => x"84",
          3037 => x"3d",
          3038 => x"96",
          3039 => x"52",
          3040 => x"0c",
          3041 => x"70",
          3042 => x"0c",
          3043 => x"3d",
          3044 => x"3d",
          3045 => x"96",
          3046 => x"82",
          3047 => x"52",
          3048 => x"73",
          3049 => x"8c",
          3050 => x"70",
          3051 => x"0c",
          3052 => x"83",
          3053 => x"82",
          3054 => x"87",
          3055 => x"0c",
          3056 => x"0d",
          3057 => x"33",
          3058 => x"2e",
          3059 => x"85",
          3060 => x"ed",
          3061 => x"e0",
          3062 => x"95",
          3063 => x"e0",
          3064 => x"72",
          3065 => x"e0",
          3066 => x"82",
          3067 => x"92",
          3068 => x"d8",
          3069 => x"8a",
          3070 => x"82",
          3071 => x"52",
          3072 => x"3d",
          3073 => x"3d",
          3074 => x"05",
          3075 => x"d8",
          3076 => x"93",
          3077 => x"51",
          3078 => x"72",
          3079 => x"0c",
          3080 => x"04",
          3081 => x"74",
          3082 => x"53",
          3083 => x"91",
          3084 => x"81",
          3085 => x"51",
          3086 => x"72",
          3087 => x"f1",
          3088 => x"0d",
          3089 => x"0d",
          3090 => x"d8",
          3091 => x"93",
          3092 => x"33",
          3093 => x"71",
          3094 => x"38",
          3095 => x"05",
          3096 => x"fe",
          3097 => x"33",
          3098 => x"38",
          3099 => x"d8",
          3100 => x"0d",
          3101 => x"0d",
          3102 => x"59",
          3103 => x"05",
          3104 => x"75",
          3105 => x"92",
          3106 => x"2e",
          3107 => x"51",
          3108 => x"e8",
          3109 => x"7a",
          3110 => x"5c",
          3111 => x"5a",
          3112 => x"09",
          3113 => x"38",
          3114 => x"81",
          3115 => x"57",
          3116 => x"75",
          3117 => x"81",
          3118 => x"82",
          3119 => x"05",
          3120 => x"5d",
          3121 => x"09",
          3122 => x"38",
          3123 => x"71",
          3124 => x"81",
          3125 => x"59",
          3126 => x"9f",
          3127 => x"53",
          3128 => x"97",
          3129 => x"29",
          3130 => x"79",
          3131 => x"5b",
          3132 => x"55",
          3133 => x"73",
          3134 => x"75",
          3135 => x"70",
          3136 => x"07",
          3137 => x"80",
          3138 => x"30",
          3139 => x"80",
          3140 => x"53",
          3141 => x"54",
          3142 => x"2e",
          3143 => x"84",
          3144 => x"81",
          3145 => x"57",
          3146 => x"2e",
          3147 => x"75",
          3148 => x"76",
          3149 => x"e0",
          3150 => x"ff",
          3151 => x"ff",
          3152 => x"72",
          3153 => x"98",
          3154 => x"10",
          3155 => x"05",
          3156 => x"04",
          3157 => x"71",
          3158 => x"53",
          3159 => x"54",
          3160 => x"2e",
          3161 => x"14",
          3162 => x"33",
          3163 => x"72",
          3164 => x"81",
          3165 => x"06",
          3166 => x"a3",
          3167 => x"15",
          3168 => x"7a",
          3169 => x"7c",
          3170 => x"06",
          3171 => x"fc",
          3172 => x"8b",
          3173 => x"15",
          3174 => x"73",
          3175 => x"74",
          3176 => x"3f",
          3177 => x"55",
          3178 => x"27",
          3179 => x"a0",
          3180 => x"3f",
          3181 => x"55",
          3182 => x"26",
          3183 => x"bc",
          3184 => x"1d",
          3185 => x"53",
          3186 => x"f5",
          3187 => x"39",
          3188 => x"39",
          3189 => x"39",
          3190 => x"39",
          3191 => x"39",
          3192 => x"dd",
          3193 => x"39",
          3194 => x"70",
          3195 => x"53",
          3196 => x"8b",
          3197 => x"1d",
          3198 => x"5d",
          3199 => x"74",
          3200 => x"09",
          3201 => x"38",
          3202 => x"71",
          3203 => x"53",
          3204 => x"84",
          3205 => x"59",
          3206 => x"80",
          3207 => x"30",
          3208 => x"80",
          3209 => x"7b",
          3210 => x"52",
          3211 => x"80",
          3212 => x"76",
          3213 => x"07",
          3214 => x"58",
          3215 => x"51",
          3216 => x"82",
          3217 => x"81",
          3218 => x"53",
          3219 => x"e5",
          3220 => x"93",
          3221 => x"89",
          3222 => x"38",
          3223 => x"70",
          3224 => x"57",
          3225 => x"80",
          3226 => x"38",
          3227 => x"81",
          3228 => x"53",
          3229 => x"05",
          3230 => x"16",
          3231 => x"74",
          3232 => x"77",
          3233 => x"07",
          3234 => x"9f",
          3235 => x"51",
          3236 => x"72",
          3237 => x"7c",
          3238 => x"81",
          3239 => x"72",
          3240 => x"38",
          3241 => x"05",
          3242 => x"ad",
          3243 => x"18",
          3244 => x"81",
          3245 => x"b0",
          3246 => x"38",
          3247 => x"81",
          3248 => x"06",
          3249 => x"a3",
          3250 => x"15",
          3251 => x"7a",
          3252 => x"7c",
          3253 => x"06",
          3254 => x"f9",
          3255 => x"8b",
          3256 => x"15",
          3257 => x"73",
          3258 => x"ff",
          3259 => x"e0",
          3260 => x"33",
          3261 => x"f9",
          3262 => x"ef",
          3263 => x"15",
          3264 => x"7a",
          3265 => x"38",
          3266 => x"b5",
          3267 => x"15",
          3268 => x"73",
          3269 => x"fa",
          3270 => x"3d",
          3271 => x"3d",
          3272 => x"70",
          3273 => x"52",
          3274 => x"73",
          3275 => x"3f",
          3276 => x"04",
          3277 => x"74",
          3278 => x"0c",
          3279 => x"05",
          3280 => x"fa",
          3281 => x"93",
          3282 => x"80",
          3283 => x"0b",
          3284 => x"0c",
          3285 => x"04",
          3286 => x"82",
          3287 => x"76",
          3288 => x"0c",
          3289 => x"05",
          3290 => x"53",
          3291 => x"72",
          3292 => x"0c",
          3293 => x"04",
          3294 => x"78",
          3295 => x"80",
          3296 => x"dc",
          3297 => x"80",
          3298 => x"39",
          3299 => x"f3",
          3300 => x"82",
          3301 => x"52",
          3302 => x"93",
          3303 => x"ff",
          3304 => x"80",
          3305 => x"73",
          3306 => x"ca",
          3307 => x"32",
          3308 => x"30",
          3309 => x"9f",
          3310 => x"25",
          3311 => x"51",
          3312 => x"2e",
          3313 => x"15",
          3314 => x"06",
          3315 => x"f1",
          3316 => x"9f",
          3317 => x"bb",
          3318 => x"52",
          3319 => x"ff",
          3320 => x"15",
          3321 => x"34",
          3322 => x"81",
          3323 => x"55",
          3324 => x"ff",
          3325 => x"17",
          3326 => x"34",
          3327 => x"c1",
          3328 => x"72",
          3329 => x"0c",
          3330 => x"04",
          3331 => x"82",
          3332 => x"75",
          3333 => x"0c",
          3334 => x"52",
          3335 => x"3f",
          3336 => x"dc",
          3337 => x"0d",
          3338 => x"0d",
          3339 => x"55",
          3340 => x"0c",
          3341 => x"33",
          3342 => x"73",
          3343 => x"81",
          3344 => x"74",
          3345 => x"75",
          3346 => x"70",
          3347 => x"73",
          3348 => x"38",
          3349 => x"09",
          3350 => x"38",
          3351 => x"11",
          3352 => x"08",
          3353 => x"54",
          3354 => x"2e",
          3355 => x"80",
          3356 => x"08",
          3357 => x"0c",
          3358 => x"33",
          3359 => x"80",
          3360 => x"38",
          3361 => x"2e",
          3362 => x"a1",
          3363 => x"81",
          3364 => x"75",
          3365 => x"56",
          3366 => x"c1",
          3367 => x"08",
          3368 => x"0c",
          3369 => x"33",
          3370 => x"b1",
          3371 => x"a0",
          3372 => x"82",
          3373 => x"53",
          3374 => x"57",
          3375 => x"9d",
          3376 => x"39",
          3377 => x"80",
          3378 => x"26",
          3379 => x"8b",
          3380 => x"80",
          3381 => x"56",
          3382 => x"8a",
          3383 => x"a0",
          3384 => x"c5",
          3385 => x"74",
          3386 => x"e0",
          3387 => x"ff",
          3388 => x"d0",
          3389 => x"ff",
          3390 => x"90",
          3391 => x"38",
          3392 => x"81",
          3393 => x"53",
          3394 => x"c5",
          3395 => x"27",
          3396 => x"76",
          3397 => x"08",
          3398 => x"0c",
          3399 => x"33",
          3400 => x"73",
          3401 => x"bd",
          3402 => x"2e",
          3403 => x"30",
          3404 => x"0c",
          3405 => x"82",
          3406 => x"8a",
          3407 => x"f8",
          3408 => x"7c",
          3409 => x"70",
          3410 => x"08",
          3411 => x"54",
          3412 => x"2e",
          3413 => x"92",
          3414 => x"81",
          3415 => x"74",
          3416 => x"55",
          3417 => x"2e",
          3418 => x"ad",
          3419 => x"06",
          3420 => x"75",
          3421 => x"0c",
          3422 => x"33",
          3423 => x"73",
          3424 => x"81",
          3425 => x"38",
          3426 => x"05",
          3427 => x"08",
          3428 => x"53",
          3429 => x"2e",
          3430 => x"80",
          3431 => x"81",
          3432 => x"90",
          3433 => x"76",
          3434 => x"70",
          3435 => x"57",
          3436 => x"82",
          3437 => x"05",
          3438 => x"08",
          3439 => x"54",
          3440 => x"81",
          3441 => x"27",
          3442 => x"d0",
          3443 => x"56",
          3444 => x"73",
          3445 => x"80",
          3446 => x"14",
          3447 => x"72",
          3448 => x"e8",
          3449 => x"80",
          3450 => x"39",
          3451 => x"dc",
          3452 => x"80",
          3453 => x"27",
          3454 => x"80",
          3455 => x"89",
          3456 => x"70",
          3457 => x"55",
          3458 => x"70",
          3459 => x"55",
          3460 => x"27",
          3461 => x"14",
          3462 => x"06",
          3463 => x"74",
          3464 => x"73",
          3465 => x"38",
          3466 => x"14",
          3467 => x"05",
          3468 => x"08",
          3469 => x"54",
          3470 => x"26",
          3471 => x"77",
          3472 => x"38",
          3473 => x"75",
          3474 => x"56",
          3475 => x"c8",
          3476 => x"0d",
          3477 => x"0d",
          3478 => x"33",
          3479 => x"70",
          3480 => x"38",
          3481 => x"11",
          3482 => x"82",
          3483 => x"83",
          3484 => x"fd",
          3485 => x"97",
          3486 => x"84",
          3487 => x"33",
          3488 => x"51",
          3489 => x"80",
          3490 => x"90",
          3491 => x"92",
          3492 => x"88",
          3493 => x"2e",
          3494 => x"88",
          3495 => x"0c",
          3496 => x"87",
          3497 => x"05",
          3498 => x"0c",
          3499 => x"c0",
          3500 => x"70",
          3501 => x"98",
          3502 => x"08",
          3503 => x"51",
          3504 => x"2e",
          3505 => x"08",
          3506 => x"38",
          3507 => x"87",
          3508 => x"05",
          3509 => x"80",
          3510 => x"51",
          3511 => x"87",
          3512 => x"08",
          3513 => x"2e",
          3514 => x"82",
          3515 => x"34",
          3516 => x"13",
          3517 => x"82",
          3518 => x"85",
          3519 => x"f2",
          3520 => x"63",
          3521 => x"05",
          3522 => x"33",
          3523 => x"58",
          3524 => x"5b",
          3525 => x"82",
          3526 => x"81",
          3527 => x"52",
          3528 => x"38",
          3529 => x"5d",
          3530 => x"8c",
          3531 => x"87",
          3532 => x"11",
          3533 => x"84",
          3534 => x"5c",
          3535 => x"85",
          3536 => x"c0",
          3537 => x"7c",
          3538 => x"84",
          3539 => x"08",
          3540 => x"70",
          3541 => x"53",
          3542 => x"2e",
          3543 => x"08",
          3544 => x"70",
          3545 => x"34",
          3546 => x"73",
          3547 => x"71",
          3548 => x"38",
          3549 => x"71",
          3550 => x"08",
          3551 => x"2e",
          3552 => x"84",
          3553 => x"38",
          3554 => x"87",
          3555 => x"1e",
          3556 => x"70",
          3557 => x"52",
          3558 => x"ff",
          3559 => x"39",
          3560 => x"81",
          3561 => x"ff",
          3562 => x"5c",
          3563 => x"90",
          3564 => x"80",
          3565 => x"71",
          3566 => x"7d",
          3567 => x"38",
          3568 => x"80",
          3569 => x"80",
          3570 => x"81",
          3571 => x"73",
          3572 => x"0c",
          3573 => x"04",
          3574 => x"60",
          3575 => x"8c",
          3576 => x"33",
          3577 => x"57",
          3578 => x"5a",
          3579 => x"82",
          3580 => x"81",
          3581 => x"52",
          3582 => x"38",
          3583 => x"c0",
          3584 => x"84",
          3585 => x"92",
          3586 => x"c0",
          3587 => x"72",
          3588 => x"5a",
          3589 => x"0c",
          3590 => x"80",
          3591 => x"0c",
          3592 => x"0c",
          3593 => x"08",
          3594 => x"70",
          3595 => x"53",
          3596 => x"2e",
          3597 => x"70",
          3598 => x"33",
          3599 => x"13",
          3600 => x"2a",
          3601 => x"51",
          3602 => x"2e",
          3603 => x"08",
          3604 => x"38",
          3605 => x"71",
          3606 => x"38",
          3607 => x"2e",
          3608 => x"75",
          3609 => x"92",
          3610 => x"72",
          3611 => x"06",
          3612 => x"f7",
          3613 => x"5a",
          3614 => x"1c",
          3615 => x"06",
          3616 => x"5d",
          3617 => x"80",
          3618 => x"73",
          3619 => x"06",
          3620 => x"38",
          3621 => x"fe",
          3622 => x"fc",
          3623 => x"52",
          3624 => x"83",
          3625 => x"71",
          3626 => x"93",
          3627 => x"3d",
          3628 => x"3d",
          3629 => x"84",
          3630 => x"33",
          3631 => x"b3",
          3632 => x"54",
          3633 => x"fb",
          3634 => x"93",
          3635 => x"06",
          3636 => x"71",
          3637 => x"54",
          3638 => x"a2",
          3639 => x"24",
          3640 => x"80",
          3641 => x"a7",
          3642 => x"2e",
          3643 => x"39",
          3644 => x"87",
          3645 => x"05",
          3646 => x"52",
          3647 => x"80",
          3648 => x"80",
          3649 => x"81",
          3650 => x"80",
          3651 => x"84",
          3652 => x"93",
          3653 => x"3d",
          3654 => x"3d",
          3655 => x"33",
          3656 => x"70",
          3657 => x"07",
          3658 => x"0c",
          3659 => x"83",
          3660 => x"fd",
          3661 => x"83",
          3662 => x"12",
          3663 => x"2b",
          3664 => x"07",
          3665 => x"71",
          3666 => x"71",
          3667 => x"82",
          3668 => x"51",
          3669 => x"52",
          3670 => x"04",
          3671 => x"73",
          3672 => x"92",
          3673 => x"52",
          3674 => x"81",
          3675 => x"70",
          3676 => x"70",
          3677 => x"3d",
          3678 => x"3d",
          3679 => x"52",
          3680 => x"70",
          3681 => x"34",
          3682 => x"51",
          3683 => x"81",
          3684 => x"70",
          3685 => x"70",
          3686 => x"05",
          3687 => x"88",
          3688 => x"72",
          3689 => x"0d",
          3690 => x"0d",
          3691 => x"54",
          3692 => x"80",
          3693 => x"71",
          3694 => x"53",
          3695 => x"81",
          3696 => x"ff",
          3697 => x"ef",
          3698 => x"0d",
          3699 => x"0d",
          3700 => x"54",
          3701 => x"72",
          3702 => x"54",
          3703 => x"51",
          3704 => x"84",
          3705 => x"fc",
          3706 => x"77",
          3707 => x"53",
          3708 => x"05",
          3709 => x"70",
          3710 => x"33",
          3711 => x"ff",
          3712 => x"52",
          3713 => x"2e",
          3714 => x"80",
          3715 => x"71",
          3716 => x"0c",
          3717 => x"04",
          3718 => x"74",
          3719 => x"53",
          3720 => x"80",
          3721 => x"70",
          3722 => x"38",
          3723 => x"33",
          3724 => x"80",
          3725 => x"70",
          3726 => x"81",
          3727 => x"71",
          3728 => x"c8",
          3729 => x"0d",
          3730 => x"82",
          3731 => x"04",
          3732 => x"93",
          3733 => x"f9",
          3734 => x"56",
          3735 => x"17",
          3736 => x"74",
          3737 => x"d7",
          3738 => x"b0",
          3739 => x"b4",
          3740 => x"81",
          3741 => x"57",
          3742 => x"82",
          3743 => x"78",
          3744 => x"06",
          3745 => x"93",
          3746 => x"17",
          3747 => x"08",
          3748 => x"31",
          3749 => x"17",
          3750 => x"38",
          3751 => x"55",
          3752 => x"09",
          3753 => x"38",
          3754 => x"16",
          3755 => x"08",
          3756 => x"52",
          3757 => x"51",
          3758 => x"83",
          3759 => x"77",
          3760 => x"0c",
          3761 => x"04",
          3762 => x"78",
          3763 => x"80",
          3764 => x"08",
          3765 => x"38",
          3766 => x"fb",
          3767 => x"c8",
          3768 => x"93",
          3769 => x"38",
          3770 => x"53",
          3771 => x"81",
          3772 => x"f8",
          3773 => x"93",
          3774 => x"2e",
          3775 => x"55",
          3776 => x"b0",
          3777 => x"82",
          3778 => x"88",
          3779 => x"f8",
          3780 => x"70",
          3781 => x"bf",
          3782 => x"c8",
          3783 => x"93",
          3784 => x"91",
          3785 => x"55",
          3786 => x"09",
          3787 => x"f0",
          3788 => x"33",
          3789 => x"2e",
          3790 => x"80",
          3791 => x"80",
          3792 => x"c8",
          3793 => x"17",
          3794 => x"fd",
          3795 => x"d4",
          3796 => x"b2",
          3797 => x"84",
          3798 => x"85",
          3799 => x"75",
          3800 => x"3f",
          3801 => x"e4",
          3802 => x"98",
          3803 => x"8a",
          3804 => x"08",
          3805 => x"17",
          3806 => x"3f",
          3807 => x"52",
          3808 => x"51",
          3809 => x"a0",
          3810 => x"05",
          3811 => x"0c",
          3812 => x"75",
          3813 => x"33",
          3814 => x"3f",
          3815 => x"34",
          3816 => x"52",
          3817 => x"51",
          3818 => x"82",
          3819 => x"80",
          3820 => x"81",
          3821 => x"93",
          3822 => x"3d",
          3823 => x"3d",
          3824 => x"1a",
          3825 => x"fe",
          3826 => x"54",
          3827 => x"73",
          3828 => x"8a",
          3829 => x"76",
          3830 => x"08",
          3831 => x"75",
          3832 => x"0c",
          3833 => x"04",
          3834 => x"7a",
          3835 => x"56",
          3836 => x"75",
          3837 => x"98",
          3838 => x"26",
          3839 => x"56",
          3840 => x"ff",
          3841 => x"56",
          3842 => x"80",
          3843 => x"82",
          3844 => x"72",
          3845 => x"38",
          3846 => x"72",
          3847 => x"8e",
          3848 => x"39",
          3849 => x"15",
          3850 => x"a4",
          3851 => x"53",
          3852 => x"fd",
          3853 => x"93",
          3854 => x"9f",
          3855 => x"ff",
          3856 => x"11",
          3857 => x"70",
          3858 => x"18",
          3859 => x"76",
          3860 => x"53",
          3861 => x"82",
          3862 => x"80",
          3863 => x"83",
          3864 => x"b4",
          3865 => x"88",
          3866 => x"77",
          3867 => x"84",
          3868 => x"5a",
          3869 => x"80",
          3870 => x"9f",
          3871 => x"80",
          3872 => x"88",
          3873 => x"08",
          3874 => x"51",
          3875 => x"82",
          3876 => x"80",
          3877 => x"15",
          3878 => x"74",
          3879 => x"51",
          3880 => x"82",
          3881 => x"83",
          3882 => x"56",
          3883 => x"87",
          3884 => x"08",
          3885 => x"51",
          3886 => x"82",
          3887 => x"9b",
          3888 => x"2b",
          3889 => x"74",
          3890 => x"51",
          3891 => x"82",
          3892 => x"f0",
          3893 => x"83",
          3894 => x"75",
          3895 => x"0c",
          3896 => x"04",
          3897 => x"7b",
          3898 => x"55",
          3899 => x"81",
          3900 => x"af",
          3901 => x"16",
          3902 => x"a7",
          3903 => x"53",
          3904 => x"81",
          3905 => x"77",
          3906 => x"72",
          3907 => x"38",
          3908 => x"72",
          3909 => x"c9",
          3910 => x"39",
          3911 => x"14",
          3912 => x"a4",
          3913 => x"53",
          3914 => x"fb",
          3915 => x"93",
          3916 => x"82",
          3917 => x"81",
          3918 => x"83",
          3919 => x"b4",
          3920 => x"76",
          3921 => x"5b",
          3922 => x"57",
          3923 => x"8f",
          3924 => x"2b",
          3925 => x"78",
          3926 => x"71",
          3927 => x"76",
          3928 => x"0b",
          3929 => x"78",
          3930 => x"16",
          3931 => x"74",
          3932 => x"3f",
          3933 => x"08",
          3934 => x"c8",
          3935 => x"38",
          3936 => x"06",
          3937 => x"75",
          3938 => x"84",
          3939 => x"51",
          3940 => x"38",
          3941 => x"78",
          3942 => x"06",
          3943 => x"06",
          3944 => x"78",
          3945 => x"83",
          3946 => x"f7",
          3947 => x"2a",
          3948 => x"05",
          3949 => x"fa",
          3950 => x"93",
          3951 => x"82",
          3952 => x"80",
          3953 => x"83",
          3954 => x"52",
          3955 => x"ff",
          3956 => x"b4",
          3957 => x"84",
          3958 => x"83",
          3959 => x"c3",
          3960 => x"2a",
          3961 => x"05",
          3962 => x"f9",
          3963 => x"93",
          3964 => x"82",
          3965 => x"ab",
          3966 => x"0a",
          3967 => x"2b",
          3968 => x"76",
          3969 => x"70",
          3970 => x"56",
          3971 => x"82",
          3972 => x"8f",
          3973 => x"07",
          3974 => x"f6",
          3975 => x"0b",
          3976 => x"76",
          3977 => x"0c",
          3978 => x"04",
          3979 => x"79",
          3980 => x"08",
          3981 => x"57",
          3982 => x"88",
          3983 => x"08",
          3984 => x"38",
          3985 => x"8e",
          3986 => x"2e",
          3987 => x"53",
          3988 => x"51",
          3989 => x"82",
          3990 => x"56",
          3991 => x"08",
          3992 => x"93",
          3993 => x"80",
          3994 => x"56",
          3995 => x"82",
          3996 => x"56",
          3997 => x"73",
          3998 => x"fa",
          3999 => x"93",
          4000 => x"82",
          4001 => x"80",
          4002 => x"38",
          4003 => x"08",
          4004 => x"38",
          4005 => x"08",
          4006 => x"38",
          4007 => x"52",
          4008 => x"c0",
          4009 => x"c8",
          4010 => x"98",
          4011 => x"05",
          4012 => x"08",
          4013 => x"38",
          4014 => x"81",
          4015 => x"0c",
          4016 => x"81",
          4017 => x"84",
          4018 => x"54",
          4019 => x"76",
          4020 => x"38",
          4021 => x"82",
          4022 => x"89",
          4023 => x"f5",
          4024 => x"7f",
          4025 => x"5c",
          4026 => x"38",
          4027 => x"58",
          4028 => x"88",
          4029 => x"08",
          4030 => x"38",
          4031 => x"39",
          4032 => x"51",
          4033 => x"81",
          4034 => x"93",
          4035 => x"82",
          4036 => x"93",
          4037 => x"82",
          4038 => x"ff",
          4039 => x"38",
          4040 => x"08",
          4041 => x"08",
          4042 => x"08",
          4043 => x"38",
          4044 => x"55",
          4045 => x"75",
          4046 => x"38",
          4047 => x"7b",
          4048 => x"06",
          4049 => x"81",
          4050 => x"19",
          4051 => x"83",
          4052 => x"76",
          4053 => x"f9",
          4054 => x"93",
          4055 => x"80",
          4056 => x"c8",
          4057 => x"09",
          4058 => x"38",
          4059 => x"08",
          4060 => x"32",
          4061 => x"72",
          4062 => x"70",
          4063 => x"53",
          4064 => x"54",
          4065 => x"38",
          4066 => x"95",
          4067 => x"08",
          4068 => x"27",
          4069 => x"98",
          4070 => x"83",
          4071 => x"80",
          4072 => x"de",
          4073 => x"81",
          4074 => x"19",
          4075 => x"89",
          4076 => x"76",
          4077 => x"b6",
          4078 => x"7b",
          4079 => x"3f",
          4080 => x"08",
          4081 => x"c8",
          4082 => x"b6",
          4083 => x"82",
          4084 => x"81",
          4085 => x"06",
          4086 => x"93",
          4087 => x"75",
          4088 => x"30",
          4089 => x"80",
          4090 => x"07",
          4091 => x"54",
          4092 => x"38",
          4093 => x"09",
          4094 => x"ab",
          4095 => x"80",
          4096 => x"53",
          4097 => x"51",
          4098 => x"82",
          4099 => x"82",
          4100 => x"30",
          4101 => x"c8",
          4102 => x"25",
          4103 => x"7f",
          4104 => x"72",
          4105 => x"51",
          4106 => x"80",
          4107 => x"76",
          4108 => x"78",
          4109 => x"3f",
          4110 => x"08",
          4111 => x"38",
          4112 => x"0c",
          4113 => x"fe",
          4114 => x"19",
          4115 => x"89",
          4116 => x"08",
          4117 => x"1a",
          4118 => x"33",
          4119 => x"73",
          4120 => x"94",
          4121 => x"75",
          4122 => x"38",
          4123 => x"55",
          4124 => x"55",
          4125 => x"57",
          4126 => x"82",
          4127 => x"8d",
          4128 => x"f7",
          4129 => x"70",
          4130 => x"cb",
          4131 => x"82",
          4132 => x"80",
          4133 => x"52",
          4134 => x"a2",
          4135 => x"c8",
          4136 => x"c8",
          4137 => x"0c",
          4138 => x"53",
          4139 => x"17",
          4140 => x"f2",
          4141 => x"59",
          4142 => x"56",
          4143 => x"16",
          4144 => x"22",
          4145 => x"27",
          4146 => x"54",
          4147 => x"78",
          4148 => x"33",
          4149 => x"3f",
          4150 => x"08",
          4151 => x"38",
          4152 => x"18",
          4153 => x"74",
          4154 => x"38",
          4155 => x"55",
          4156 => x"c8",
          4157 => x"0d",
          4158 => x"0d",
          4159 => x"08",
          4160 => x"74",
          4161 => x"26",
          4162 => x"9f",
          4163 => x"80",
          4164 => x"82",
          4165 => x"39",
          4166 => x"0c",
          4167 => x"54",
          4168 => x"75",
          4169 => x"73",
          4170 => x"a8",
          4171 => x"73",
          4172 => x"85",
          4173 => x"0b",
          4174 => x"5a",
          4175 => x"27",
          4176 => x"a8",
          4177 => x"18",
          4178 => x"39",
          4179 => x"70",
          4180 => x"58",
          4181 => x"b6",
          4182 => x"76",
          4183 => x"3f",
          4184 => x"08",
          4185 => x"c8",
          4186 => x"bf",
          4187 => x"82",
          4188 => x"27",
          4189 => x"16",
          4190 => x"c8",
          4191 => x"38",
          4192 => x"c1",
          4193 => x"31",
          4194 => x"27",
          4195 => x"52",
          4196 => x"aa",
          4197 => x"c8",
          4198 => x"0c",
          4199 => x"0c",
          4200 => x"17",
          4201 => x"9d",
          4202 => x"81",
          4203 => x"74",
          4204 => x"18",
          4205 => x"18",
          4206 => x"ff",
          4207 => x"05",
          4208 => x"80",
          4209 => x"93",
          4210 => x"3d",
          4211 => x"3d",
          4212 => x"71",
          4213 => x"08",
          4214 => x"59",
          4215 => x"80",
          4216 => x"86",
          4217 => x"98",
          4218 => x"53",
          4219 => x"80",
          4220 => x"38",
          4221 => x"06",
          4222 => x"c1",
          4223 => x"08",
          4224 => x"16",
          4225 => x"08",
          4226 => x"85",
          4227 => x"22",
          4228 => x"73",
          4229 => x"38",
          4230 => x"0c",
          4231 => x"ad",
          4232 => x"22",
          4233 => x"89",
          4234 => x"53",
          4235 => x"38",
          4236 => x"52",
          4237 => x"b0",
          4238 => x"c8",
          4239 => x"53",
          4240 => x"93",
          4241 => x"81",
          4242 => x"53",
          4243 => x"08",
          4244 => x"f9",
          4245 => x"08",
          4246 => x"08",
          4247 => x"38",
          4248 => x"77",
          4249 => x"84",
          4250 => x"39",
          4251 => x"52",
          4252 => x"eb",
          4253 => x"c8",
          4254 => x"53",
          4255 => x"08",
          4256 => x"c9",
          4257 => x"82",
          4258 => x"81",
          4259 => x"81",
          4260 => x"c8",
          4261 => x"b5",
          4262 => x"c8",
          4263 => x"51",
          4264 => x"81",
          4265 => x"c8",
          4266 => x"73",
          4267 => x"73",
          4268 => x"f2",
          4269 => x"93",
          4270 => x"16",
          4271 => x"16",
          4272 => x"ff",
          4273 => x"05",
          4274 => x"80",
          4275 => x"93",
          4276 => x"3d",
          4277 => x"3d",
          4278 => x"71",
          4279 => x"56",
          4280 => x"51",
          4281 => x"82",
          4282 => x"54",
          4283 => x"08",
          4284 => x"82",
          4285 => x"57",
          4286 => x"52",
          4287 => x"c8",
          4288 => x"c8",
          4289 => x"93",
          4290 => x"c7",
          4291 => x"c8",
          4292 => x"08",
          4293 => x"54",
          4294 => x"e5",
          4295 => x"06",
          4296 => x"55",
          4297 => x"80",
          4298 => x"51",
          4299 => x"2e",
          4300 => x"17",
          4301 => x"2e",
          4302 => x"39",
          4303 => x"52",
          4304 => x"8a",
          4305 => x"c8",
          4306 => x"93",
          4307 => x"2e",
          4308 => x"73",
          4309 => x"81",
          4310 => x"87",
          4311 => x"93",
          4312 => x"3d",
          4313 => x"3d",
          4314 => x"11",
          4315 => x"aa",
          4316 => x"c8",
          4317 => x"ff",
          4318 => x"33",
          4319 => x"71",
          4320 => x"81",
          4321 => x"94",
          4322 => x"8e",
          4323 => x"c8",
          4324 => x"73",
          4325 => x"82",
          4326 => x"85",
          4327 => x"fc",
          4328 => x"79",
          4329 => x"ff",
          4330 => x"12",
          4331 => x"eb",
          4332 => x"70",
          4333 => x"72",
          4334 => x"81",
          4335 => x"73",
          4336 => x"94",
          4337 => x"94",
          4338 => x"0d",
          4339 => x"0d",
          4340 => x"56",
          4341 => x"5a",
          4342 => x"08",
          4343 => x"86",
          4344 => x"08",
          4345 => x"ed",
          4346 => x"93",
          4347 => x"82",
          4348 => x"80",
          4349 => x"16",
          4350 => x"56",
          4351 => x"38",
          4352 => x"e2",
          4353 => x"08",
          4354 => x"70",
          4355 => x"81",
          4356 => x"51",
          4357 => x"86",
          4358 => x"81",
          4359 => x"30",
          4360 => x"70",
          4361 => x"06",
          4362 => x"51",
          4363 => x"73",
          4364 => x"38",
          4365 => x"96",
          4366 => x"df",
          4367 => x"72",
          4368 => x"81",
          4369 => x"81",
          4370 => x"2e",
          4371 => x"52",
          4372 => x"fa",
          4373 => x"c8",
          4374 => x"93",
          4375 => x"38",
          4376 => x"fe",
          4377 => x"80",
          4378 => x"80",
          4379 => x"0c",
          4380 => x"c8",
          4381 => x"0d",
          4382 => x"0d",
          4383 => x"59",
          4384 => x"75",
          4385 => x"3f",
          4386 => x"08",
          4387 => x"c8",
          4388 => x"38",
          4389 => x"57",
          4390 => x"98",
          4391 => x"77",
          4392 => x"3f",
          4393 => x"08",
          4394 => x"c8",
          4395 => x"38",
          4396 => x"70",
          4397 => x"73",
          4398 => x"38",
          4399 => x"8b",
          4400 => x"06",
          4401 => x"86",
          4402 => x"15",
          4403 => x"2a",
          4404 => x"51",
          4405 => x"93",
          4406 => x"a0",
          4407 => x"51",
          4408 => x"82",
          4409 => x"80",
          4410 => x"80",
          4411 => x"f9",
          4412 => x"93",
          4413 => x"82",
          4414 => x"80",
          4415 => x"38",
          4416 => x"82",
          4417 => x"8a",
          4418 => x"fb",
          4419 => x"70",
          4420 => x"81",
          4421 => x"fb",
          4422 => x"93",
          4423 => x"82",
          4424 => x"b4",
          4425 => x"08",
          4426 => x"eb",
          4427 => x"93",
          4428 => x"82",
          4429 => x"a0",
          4430 => x"82",
          4431 => x"52",
          4432 => x"51",
          4433 => x"8b",
          4434 => x"52",
          4435 => x"51",
          4436 => x"81",
          4437 => x"34",
          4438 => x"c8",
          4439 => x"0d",
          4440 => x"0d",
          4441 => x"98",
          4442 => x"70",
          4443 => x"ea",
          4444 => x"93",
          4445 => x"82",
          4446 => x"8d",
          4447 => x"08",
          4448 => x"34",
          4449 => x"16",
          4450 => x"93",
          4451 => x"3d",
          4452 => x"3d",
          4453 => x"57",
          4454 => x"89",
          4455 => x"17",
          4456 => x"81",
          4457 => x"70",
          4458 => x"17",
          4459 => x"33",
          4460 => x"54",
          4461 => x"2e",
          4462 => x"85",
          4463 => x"06",
          4464 => x"e5",
          4465 => x"2e",
          4466 => x"8e",
          4467 => x"88",
          4468 => x"0b",
          4469 => x"81",
          4470 => x"15",
          4471 => x"72",
          4472 => x"81",
          4473 => x"74",
          4474 => x"75",
          4475 => x"52",
          4476 => x"13",
          4477 => x"08",
          4478 => x"33",
          4479 => x"9c",
          4480 => x"05",
          4481 => x"3f",
          4482 => x"08",
          4483 => x"17",
          4484 => x"51",
          4485 => x"82",
          4486 => x"86",
          4487 => x"17",
          4488 => x"51",
          4489 => x"82",
          4490 => x"84",
          4491 => x"3d",
          4492 => x"3d",
          4493 => x"08",
          4494 => x"5d",
          4495 => x"53",
          4496 => x"51",
          4497 => x"80",
          4498 => x"88",
          4499 => x"5a",
          4500 => x"09",
          4501 => x"df",
          4502 => x"70",
          4503 => x"71",
          4504 => x"30",
          4505 => x"73",
          4506 => x"51",
          4507 => x"57",
          4508 => x"38",
          4509 => x"75",
          4510 => x"18",
          4511 => x"75",
          4512 => x"30",
          4513 => x"32",
          4514 => x"73",
          4515 => x"53",
          4516 => x"55",
          4517 => x"89",
          4518 => x"75",
          4519 => x"e4",
          4520 => x"7c",
          4521 => x"a0",
          4522 => x"38",
          4523 => x"8b",
          4524 => x"54",
          4525 => x"78",
          4526 => x"81",
          4527 => x"54",
          4528 => x"82",
          4529 => x"af",
          4530 => x"77",
          4531 => x"70",
          4532 => x"25",
          4533 => x"07",
          4534 => x"51",
          4535 => x"2e",
          4536 => x"39",
          4537 => x"80",
          4538 => x"33",
          4539 => x"73",
          4540 => x"81",
          4541 => x"81",
          4542 => x"1a",
          4543 => x"55",
          4544 => x"dc",
          4545 => x"06",
          4546 => x"55",
          4547 => x"54",
          4548 => x"81",
          4549 => x"ae",
          4550 => x"70",
          4551 => x"7d",
          4552 => x"51",
          4553 => x"2e",
          4554 => x"8b",
          4555 => x"77",
          4556 => x"30",
          4557 => x"71",
          4558 => x"53",
          4559 => x"55",
          4560 => x"38",
          4561 => x"5a",
          4562 => x"75",
          4563 => x"73",
          4564 => x"38",
          4565 => x"06",
          4566 => x"11",
          4567 => x"75",
          4568 => x"3f",
          4569 => x"08",
          4570 => x"38",
          4571 => x"33",
          4572 => x"54",
          4573 => x"e5",
          4574 => x"93",
          4575 => x"2e",
          4576 => x"1a",
          4577 => x"26",
          4578 => x"54",
          4579 => x"7a",
          4580 => x"74",
          4581 => x"7b",
          4582 => x"74",
          4583 => x"18",
          4584 => x"39",
          4585 => x"fa",
          4586 => x"ec",
          4587 => x"c8",
          4588 => x"38",
          4589 => x"54",
          4590 => x"89",
          4591 => x"70",
          4592 => x"57",
          4593 => x"54",
          4594 => x"81",
          4595 => x"e7",
          4596 => x"7c",
          4597 => x"77",
          4598 => x"38",
          4599 => x"73",
          4600 => x"09",
          4601 => x"38",
          4602 => x"84",
          4603 => x"27",
          4604 => x"39",
          4605 => x"39",
          4606 => x"39",
          4607 => x"8b",
          4608 => x"54",
          4609 => x"c8",
          4610 => x"0d",
          4611 => x"0d",
          4612 => x"58",
          4613 => x"70",
          4614 => x"55",
          4615 => x"83",
          4616 => x"80",
          4617 => x"51",
          4618 => x"80",
          4619 => x"38",
          4620 => x"74",
          4621 => x"80",
          4622 => x"94",
          4623 => x"17",
          4624 => x"81",
          4625 => x"7a",
          4626 => x"54",
          4627 => x"2e",
          4628 => x"83",
          4629 => x"80",
          4630 => x"51",
          4631 => x"80",
          4632 => x"81",
          4633 => x"81",
          4634 => x"07",
          4635 => x"38",
          4636 => x"17",
          4637 => x"33",
          4638 => x"9f",
          4639 => x"ff",
          4640 => x"17",
          4641 => x"75",
          4642 => x"3f",
          4643 => x"08",
          4644 => x"39",
          4645 => x"a5",
          4646 => x"84",
          4647 => x"51",
          4648 => x"82",
          4649 => x"55",
          4650 => x"08",
          4651 => x"75",
          4652 => x"3f",
          4653 => x"08",
          4654 => x"55",
          4655 => x"c8",
          4656 => x"80",
          4657 => x"93",
          4658 => x"2e",
          4659 => x"80",
          4660 => x"85",
          4661 => x"06",
          4662 => x"80",
          4663 => x"73",
          4664 => x"81",
          4665 => x"72",
          4666 => x"ad",
          4667 => x"0b",
          4668 => x"80",
          4669 => x"39",
          4670 => x"70",
          4671 => x"53",
          4672 => x"85",
          4673 => x"73",
          4674 => x"81",
          4675 => x"72",
          4676 => x"16",
          4677 => x"2a",
          4678 => x"51",
          4679 => x"80",
          4680 => x"38",
          4681 => x"83",
          4682 => x"b4",
          4683 => x"51",
          4684 => x"82",
          4685 => x"88",
          4686 => x"dd",
          4687 => x"93",
          4688 => x"3d",
          4689 => x"3d",
          4690 => x"ff",
          4691 => x"72",
          4692 => x"5a",
          4693 => x"81",
          4694 => x"70",
          4695 => x"33",
          4696 => x"70",
          4697 => x"26",
          4698 => x"06",
          4699 => x"53",
          4700 => x"72",
          4701 => x"81",
          4702 => x"38",
          4703 => x"11",
          4704 => x"89",
          4705 => x"82",
          4706 => x"ff",
          4707 => x"51",
          4708 => x"77",
          4709 => x"38",
          4710 => x"fb",
          4711 => x"77",
          4712 => x"70",
          4713 => x"57",
          4714 => x"70",
          4715 => x"33",
          4716 => x"05",
          4717 => x"9f",
          4718 => x"54",
          4719 => x"89",
          4720 => x"70",
          4721 => x"55",
          4722 => x"13",
          4723 => x"26",
          4724 => x"13",
          4725 => x"06",
          4726 => x"30",
          4727 => x"70",
          4728 => x"07",
          4729 => x"9f",
          4730 => x"55",
          4731 => x"ff",
          4732 => x"30",
          4733 => x"70",
          4734 => x"07",
          4735 => x"9f",
          4736 => x"55",
          4737 => x"80",
          4738 => x"81",
          4739 => x"78",
          4740 => x"38",
          4741 => x"83",
          4742 => x"77",
          4743 => x"5a",
          4744 => x"39",
          4745 => x"33",
          4746 => x"93",
          4747 => x"3d",
          4748 => x"3d",
          4749 => x"80",
          4750 => x"34",
          4751 => x"17",
          4752 => x"75",
          4753 => x"3f",
          4754 => x"93",
          4755 => x"84",
          4756 => x"16",
          4757 => x"3f",
          4758 => x"08",
          4759 => x"06",
          4760 => x"73",
          4761 => x"2e",
          4762 => x"80",
          4763 => x"0b",
          4764 => x"55",
          4765 => x"e9",
          4766 => x"06",
          4767 => x"55",
          4768 => x"32",
          4769 => x"80",
          4770 => x"51",
          4771 => x"8e",
          4772 => x"33",
          4773 => x"e8",
          4774 => x"06",
          4775 => x"53",
          4776 => x"52",
          4777 => x"51",
          4778 => x"82",
          4779 => x"55",
          4780 => x"08",
          4781 => x"38",
          4782 => x"fb",
          4783 => x"86",
          4784 => x"a3",
          4785 => x"c8",
          4786 => x"93",
          4787 => x"2e",
          4788 => x"55",
          4789 => x"c8",
          4790 => x"0d",
          4791 => x"0d",
          4792 => x"05",
          4793 => x"33",
          4794 => x"74",
          4795 => x"fc",
          4796 => x"93",
          4797 => x"8b",
          4798 => x"82",
          4799 => x"24",
          4800 => x"82",
          4801 => x"10",
          4802 => x"e4",
          4803 => x"56",
          4804 => x"74",
          4805 => x"88",
          4806 => x"0c",
          4807 => x"06",
          4808 => x"57",
          4809 => x"af",
          4810 => x"33",
          4811 => x"3f",
          4812 => x"08",
          4813 => x"70",
          4814 => x"54",
          4815 => x"76",
          4816 => x"38",
          4817 => x"70",
          4818 => x"53",
          4819 => x"86",
          4820 => x"56",
          4821 => x"80",
          4822 => x"81",
          4823 => x"52",
          4824 => x"51",
          4825 => x"82",
          4826 => x"81",
          4827 => x"81",
          4828 => x"83",
          4829 => x"a8",
          4830 => x"2e",
          4831 => x"82",
          4832 => x"06",
          4833 => x"56",
          4834 => x"38",
          4835 => x"75",
          4836 => x"9e",
          4837 => x"c8",
          4838 => x"06",
          4839 => x"2e",
          4840 => x"80",
          4841 => x"54",
          4842 => x"15",
          4843 => x"10",
          4844 => x"05",
          4845 => x"33",
          4846 => x"80",
          4847 => x"2e",
          4848 => x"fa",
          4849 => x"eb",
          4850 => x"c8",
          4851 => x"78",
          4852 => x"54",
          4853 => x"d0",
          4854 => x"8f",
          4855 => x"10",
          4856 => x"08",
          4857 => x"57",
          4858 => x"90",
          4859 => x"74",
          4860 => x"3f",
          4861 => x"08",
          4862 => x"57",
          4863 => x"89",
          4864 => x"54",
          4865 => x"d3",
          4866 => x"76",
          4867 => x"90",
          4868 => x"76",
          4869 => x"88",
          4870 => x"51",
          4871 => x"82",
          4872 => x"83",
          4873 => x"53",
          4874 => x"84",
          4875 => x"81",
          4876 => x"38",
          4877 => x"51",
          4878 => x"82",
          4879 => x"83",
          4880 => x"54",
          4881 => x"80",
          4882 => x"d9",
          4883 => x"93",
          4884 => x"73",
          4885 => x"80",
          4886 => x"82",
          4887 => x"c4",
          4888 => x"05",
          4889 => x"72",
          4890 => x"b4",
          4891 => x"33",
          4892 => x"80",
          4893 => x"52",
          4894 => x"8a",
          4895 => x"83",
          4896 => x"53",
          4897 => x"8b",
          4898 => x"73",
          4899 => x"80",
          4900 => x"8d",
          4901 => x"39",
          4902 => x"51",
          4903 => x"82",
          4904 => x"88",
          4905 => x"93",
          4906 => x"ff",
          4907 => x"06",
          4908 => x"72",
          4909 => x"80",
          4910 => x"d8",
          4911 => x"93",
          4912 => x"ff",
          4913 => x"72",
          4914 => x"d4",
          4915 => x"e3",
          4916 => x"c8",
          4917 => x"c2",
          4918 => x"be",
          4919 => x"c8",
          4920 => x"ff",
          4921 => x"56",
          4922 => x"83",
          4923 => x"15",
          4924 => x"71",
          4925 => x"59",
          4926 => x"77",
          4927 => x"a0",
          4928 => x"22",
          4929 => x"31",
          4930 => x"ab",
          4931 => x"c8",
          4932 => x"56",
          4933 => x"08",
          4934 => x"84",
          4935 => x"82",
          4936 => x"80",
          4937 => x"f5",
          4938 => x"83",
          4939 => x"ff",
          4940 => x"38",
          4941 => x"9f",
          4942 => x"38",
          4943 => x"56",
          4944 => x"82",
          4945 => x"13",
          4946 => x"79",
          4947 => x"79",
          4948 => x"0c",
          4949 => x"16",
          4950 => x"2e",
          4951 => x"b7",
          4952 => x"15",
          4953 => x"3f",
          4954 => x"08",
          4955 => x"06",
          4956 => x"72",
          4957 => x"88",
          4958 => x"8d",
          4959 => x"a0",
          4960 => x"15",
          4961 => x"3f",
          4962 => x"08",
          4963 => x"98",
          4964 => x"2b",
          4965 => x"88",
          4966 => x"8d",
          4967 => x"2e",
          4968 => x"a4",
          4969 => x"a8",
          4970 => x"82",
          4971 => x"06",
          4972 => x"15",
          4973 => x"94",
          4974 => x"08",
          4975 => x"08",
          4976 => x"2a",
          4977 => x"81",
          4978 => x"53",
          4979 => x"89",
          4980 => x"56",
          4981 => x"08",
          4982 => x"38",
          4983 => x"16",
          4984 => x"8c",
          4985 => x"80",
          4986 => x"34",
          4987 => x"09",
          4988 => x"92",
          4989 => x"15",
          4990 => x"3f",
          4991 => x"08",
          4992 => x"06",
          4993 => x"2e",
          4994 => x"80",
          4995 => x"1a",
          4996 => x"d9",
          4997 => x"93",
          4998 => x"ea",
          4999 => x"c8",
          5000 => x"34",
          5001 => x"51",
          5002 => x"82",
          5003 => x"83",
          5004 => x"53",
          5005 => x"d5",
          5006 => x"06",
          5007 => x"b4",
          5008 => x"ef",
          5009 => x"c8",
          5010 => x"85",
          5011 => x"09",
          5012 => x"38",
          5013 => x"51",
          5014 => x"82",
          5015 => x"86",
          5016 => x"f2",
          5017 => x"06",
          5018 => x"9c",
          5019 => x"c3",
          5020 => x"c8",
          5021 => x"0c",
          5022 => x"51",
          5023 => x"82",
          5024 => x"8c",
          5025 => x"75",
          5026 => x"f4",
          5027 => x"53",
          5028 => x"f4",
          5029 => x"16",
          5030 => x"94",
          5031 => x"56",
          5032 => x"c8",
          5033 => x"0d",
          5034 => x"0d",
          5035 => x"55",
          5036 => x"b5",
          5037 => x"80",
          5038 => x"73",
          5039 => x"53",
          5040 => x"2e",
          5041 => x"14",
          5042 => x"22",
          5043 => x"76",
          5044 => x"06",
          5045 => x"13",
          5046 => x"f9",
          5047 => x"c8",
          5048 => x"52",
          5049 => x"71",
          5050 => x"74",
          5051 => x"81",
          5052 => x"73",
          5053 => x"73",
          5054 => x"74",
          5055 => x"0c",
          5056 => x"04",
          5057 => x"02",
          5058 => x"7a",
          5059 => x"fc",
          5060 => x"f4",
          5061 => x"93",
          5062 => x"8b",
          5063 => x"82",
          5064 => x"24",
          5065 => x"82",
          5066 => x"10",
          5067 => x"e4",
          5068 => x"51",
          5069 => x"2e",
          5070 => x"74",
          5071 => x"2e",
          5072 => x"54",
          5073 => x"74",
          5074 => x"93",
          5075 => x"71",
          5076 => x"54",
          5077 => x"92",
          5078 => x"89",
          5079 => x"84",
          5080 => x"f9",
          5081 => x"c8",
          5082 => x"82",
          5083 => x"88",
          5084 => x"eb",
          5085 => x"02",
          5086 => x"e7",
          5087 => x"58",
          5088 => x"80",
          5089 => x"38",
          5090 => x"70",
          5091 => x"d0",
          5092 => x"3d",
          5093 => x"57",
          5094 => x"82",
          5095 => x"56",
          5096 => x"08",
          5097 => x"7a",
          5098 => x"97",
          5099 => x"51",
          5100 => x"82",
          5101 => x"56",
          5102 => x"08",
          5103 => x"80",
          5104 => x"70",
          5105 => x"59",
          5106 => x"83",
          5107 => x"76",
          5108 => x"74",
          5109 => x"c3",
          5110 => x"2e",
          5111 => x"84",
          5112 => x"06",
          5113 => x"3d",
          5114 => x"ea",
          5115 => x"93",
          5116 => x"76",
          5117 => x"a0",
          5118 => x"05",
          5119 => x"55",
          5120 => x"85",
          5121 => x"90",
          5122 => x"2a",
          5123 => x"51",
          5124 => x"2e",
          5125 => x"56",
          5126 => x"38",
          5127 => x"70",
          5128 => x"55",
          5129 => x"81",
          5130 => x"52",
          5131 => x"b6",
          5132 => x"c8",
          5133 => x"88",
          5134 => x"62",
          5135 => x"d2",
          5136 => x"55",
          5137 => x"16",
          5138 => x"62",
          5139 => x"e6",
          5140 => x"52",
          5141 => x"51",
          5142 => x"7a",
          5143 => x"83",
          5144 => x"80",
          5145 => x"38",
          5146 => x"08",
          5147 => x"54",
          5148 => x"05",
          5149 => x"db",
          5150 => x"93",
          5151 => x"82",
          5152 => x"82",
          5153 => x"52",
          5154 => x"bc",
          5155 => x"c8",
          5156 => x"1b",
          5157 => x"56",
          5158 => x"75",
          5159 => x"02",
          5160 => x"70",
          5161 => x"81",
          5162 => x"59",
          5163 => x"85",
          5164 => x"9c",
          5165 => x"2a",
          5166 => x"51",
          5167 => x"2e",
          5168 => x"b2",
          5169 => x"06",
          5170 => x"2e",
          5171 => x"56",
          5172 => x"38",
          5173 => x"70",
          5174 => x"55",
          5175 => x"86",
          5176 => x"c0",
          5177 => x"b0",
          5178 => x"1a",
          5179 => x"1a",
          5180 => x"81",
          5181 => x"52",
          5182 => x"ea",
          5183 => x"c8",
          5184 => x"0c",
          5185 => x"51",
          5186 => x"82",
          5187 => x"8c",
          5188 => x"78",
          5189 => x"22",
          5190 => x"76",
          5191 => x"75",
          5192 => x"75",
          5193 => x"75",
          5194 => x"84",
          5195 => x"52",
          5196 => x"d1",
          5197 => x"85",
          5198 => x"06",
          5199 => x"80",
          5200 => x"38",
          5201 => x"80",
          5202 => x"38",
          5203 => x"94",
          5204 => x"8a",
          5205 => x"89",
          5206 => x"08",
          5207 => x"5d",
          5208 => x"55",
          5209 => x"52",
          5210 => x"fc",
          5211 => x"c8",
          5212 => x"93",
          5213 => x"26",
          5214 => x"56",
          5215 => x"09",
          5216 => x"38",
          5217 => x"7a",
          5218 => x"30",
          5219 => x"80",
          5220 => x"7d",
          5221 => x"51",
          5222 => x"38",
          5223 => x"0c",
          5224 => x"38",
          5225 => x"06",
          5226 => x"2e",
          5227 => x"52",
          5228 => x"8a",
          5229 => x"c8",
          5230 => x"82",
          5231 => x"78",
          5232 => x"93",
          5233 => x"70",
          5234 => x"55",
          5235 => x"53",
          5236 => x"7a",
          5237 => x"52",
          5238 => x"3f",
          5239 => x"08",
          5240 => x"38",
          5241 => x"80",
          5242 => x"80",
          5243 => x"55",
          5244 => x"c8",
          5245 => x"0d",
          5246 => x"0d",
          5247 => x"63",
          5248 => x"57",
          5249 => x"8f",
          5250 => x"52",
          5251 => x"99",
          5252 => x"c8",
          5253 => x"93",
          5254 => x"38",
          5255 => x"55",
          5256 => x"86",
          5257 => x"83",
          5258 => x"17",
          5259 => x"55",
          5260 => x"80",
          5261 => x"38",
          5262 => x"0b",
          5263 => x"82",
          5264 => x"39",
          5265 => x"18",
          5266 => x"83",
          5267 => x"0b",
          5268 => x"82",
          5269 => x"39",
          5270 => x"18",
          5271 => x"82",
          5272 => x"0b",
          5273 => x"81",
          5274 => x"39",
          5275 => x"18",
          5276 => x"82",
          5277 => x"17",
          5278 => x"08",
          5279 => x"79",
          5280 => x"74",
          5281 => x"2e",
          5282 => x"94",
          5283 => x"83",
          5284 => x"56",
          5285 => x"38",
          5286 => x"22",
          5287 => x"89",
          5288 => x"55",
          5289 => x"75",
          5290 => x"17",
          5291 => x"39",
          5292 => x"52",
          5293 => x"b0",
          5294 => x"c8",
          5295 => x"75",
          5296 => x"38",
          5297 => x"fe",
          5298 => x"98",
          5299 => x"17",
          5300 => x"51",
          5301 => x"82",
          5302 => x"80",
          5303 => x"38",
          5304 => x"08",
          5305 => x"2a",
          5306 => x"80",
          5307 => x"38",
          5308 => x"8a",
          5309 => x"56",
          5310 => x"27",
          5311 => x"7b",
          5312 => x"54",
          5313 => x"52",
          5314 => x"33",
          5315 => x"ef",
          5316 => x"c8",
          5317 => x"38",
          5318 => x"70",
          5319 => x"56",
          5320 => x"9b",
          5321 => x"08",
          5322 => x"74",
          5323 => x"38",
          5324 => x"a8",
          5325 => x"84",
          5326 => x"51",
          5327 => x"79",
          5328 => x"80",
          5329 => x"17",
          5330 => x"80",
          5331 => x"17",
          5332 => x"2b",
          5333 => x"80",
          5334 => x"81",
          5335 => x"08",
          5336 => x"52",
          5337 => x"33",
          5338 => x"ec",
          5339 => x"c8",
          5340 => x"38",
          5341 => x"80",
          5342 => x"74",
          5343 => x"81",
          5344 => x"a8",
          5345 => x"81",
          5346 => x"55",
          5347 => x"82",
          5348 => x"fd",
          5349 => x"9c",
          5350 => x"17",
          5351 => x"06",
          5352 => x"31",
          5353 => x"76",
          5354 => x"78",
          5355 => x"94",
          5356 => x"ff",
          5357 => x"05",
          5358 => x"cb",
          5359 => x"76",
          5360 => x"17",
          5361 => x"1d",
          5362 => x"18",
          5363 => x"5d",
          5364 => x"b7",
          5365 => x"75",
          5366 => x"0c",
          5367 => x"04",
          5368 => x"7f",
          5369 => x"5f",
          5370 => x"80",
          5371 => x"3d",
          5372 => x"76",
          5373 => x"3f",
          5374 => x"08",
          5375 => x"c8",
          5376 => x"91",
          5377 => x"74",
          5378 => x"38",
          5379 => x"82",
          5380 => x"33",
          5381 => x"70",
          5382 => x"56",
          5383 => x"74",
          5384 => x"ee",
          5385 => x"82",
          5386 => x"34",
          5387 => x"e2",
          5388 => x"91",
          5389 => x"56",
          5390 => x"81",
          5391 => x"34",
          5392 => x"ce",
          5393 => x"91",
          5394 => x"56",
          5395 => x"81",
          5396 => x"34",
          5397 => x"ba",
          5398 => x"91",
          5399 => x"56",
          5400 => x"94",
          5401 => x"55",
          5402 => x"08",
          5403 => x"94",
          5404 => x"59",
          5405 => x"83",
          5406 => x"17",
          5407 => x"ff",
          5408 => x"74",
          5409 => x"7d",
          5410 => x"ff",
          5411 => x"2a",
          5412 => x"7a",
          5413 => x"75",
          5414 => x"17",
          5415 => x"a3",
          5416 => x"76",
          5417 => x"3f",
          5418 => x"08",
          5419 => x"98",
          5420 => x"76",
          5421 => x"3f",
          5422 => x"08",
          5423 => x"2e",
          5424 => x"74",
          5425 => x"df",
          5426 => x"2e",
          5427 => x"74",
          5428 => x"88",
          5429 => x"38",
          5430 => x"0c",
          5431 => x"70",
          5432 => x"58",
          5433 => x"a5",
          5434 => x"9c",
          5435 => x"a8",
          5436 => x"81",
          5437 => x"55",
          5438 => x"82",
          5439 => x"fe",
          5440 => x"17",
          5441 => x"06",
          5442 => x"18",
          5443 => x"08",
          5444 => x"cd",
          5445 => x"93",
          5446 => x"2e",
          5447 => x"82",
          5448 => x"1b",
          5449 => x"5b",
          5450 => x"2e",
          5451 => x"79",
          5452 => x"11",
          5453 => x"56",
          5454 => x"85",
          5455 => x"31",
          5456 => x"77",
          5457 => x"7d",
          5458 => x"52",
          5459 => x"3f",
          5460 => x"08",
          5461 => x"9c",
          5462 => x"31",
          5463 => x"27",
          5464 => x"80",
          5465 => x"80",
          5466 => x"a8",
          5467 => x"b9",
          5468 => x"33",
          5469 => x"55",
          5470 => x"34",
          5471 => x"56",
          5472 => x"9c",
          5473 => x"2e",
          5474 => x"17",
          5475 => x"08",
          5476 => x"81",
          5477 => x"a8",
          5478 => x"81",
          5479 => x"55",
          5480 => x"82",
          5481 => x"fd",
          5482 => x"9c",
          5483 => x"17",
          5484 => x"06",
          5485 => x"31",
          5486 => x"76",
          5487 => x"78",
          5488 => x"7b",
          5489 => x"08",
          5490 => x"17",
          5491 => x"c7",
          5492 => x"17",
          5493 => x"07",
          5494 => x"18",
          5495 => x"31",
          5496 => x"7e",
          5497 => x"94",
          5498 => x"70",
          5499 => x"8c",
          5500 => x"58",
          5501 => x"76",
          5502 => x"75",
          5503 => x"18",
          5504 => x"f6",
          5505 => x"33",
          5506 => x"55",
          5507 => x"34",
          5508 => x"82",
          5509 => x"8f",
          5510 => x"f7",
          5511 => x"8c",
          5512 => x"53",
          5513 => x"f1",
          5514 => x"93",
          5515 => x"82",
          5516 => x"81",
          5517 => x"18",
          5518 => x"2a",
          5519 => x"51",
          5520 => x"80",
          5521 => x"38",
          5522 => x"55",
          5523 => x"a7",
          5524 => x"9c",
          5525 => x"a8",
          5526 => x"81",
          5527 => x"55",
          5528 => x"81",
          5529 => x"c8",
          5530 => x"38",
          5531 => x"80",
          5532 => x"74",
          5533 => x"a0",
          5534 => x"79",
          5535 => x"3f",
          5536 => x"08",
          5537 => x"c8",
          5538 => x"38",
          5539 => x"8b",
          5540 => x"07",
          5541 => x"8b",
          5542 => x"18",
          5543 => x"52",
          5544 => x"d9",
          5545 => x"18",
          5546 => x"16",
          5547 => x"3f",
          5548 => x"0a",
          5549 => x"51",
          5550 => x"76",
          5551 => x"51",
          5552 => x"79",
          5553 => x"83",
          5554 => x"51",
          5555 => x"82",
          5556 => x"90",
          5557 => x"bf",
          5558 => x"74",
          5559 => x"76",
          5560 => x"93",
          5561 => x"3d",
          5562 => x"3d",
          5563 => x"52",
          5564 => x"3f",
          5565 => x"08",
          5566 => x"c8",
          5567 => x"86",
          5568 => x"52",
          5569 => x"a1",
          5570 => x"c8",
          5571 => x"93",
          5572 => x"38",
          5573 => x"08",
          5574 => x"82",
          5575 => x"86",
          5576 => x"fe",
          5577 => x"3d",
          5578 => x"3f",
          5579 => x"0b",
          5580 => x"08",
          5581 => x"82",
          5582 => x"82",
          5583 => x"80",
          5584 => x"93",
          5585 => x"3d",
          5586 => x"3d",
          5587 => x"93",
          5588 => x"52",
          5589 => x"e7",
          5590 => x"93",
          5591 => x"82",
          5592 => x"80",
          5593 => x"58",
          5594 => x"3d",
          5595 => x"e1",
          5596 => x"93",
          5597 => x"82",
          5598 => x"be",
          5599 => x"c7",
          5600 => x"98",
          5601 => x"73",
          5602 => x"38",
          5603 => x"12",
          5604 => x"39",
          5605 => x"33",
          5606 => x"70",
          5607 => x"55",
          5608 => x"2e",
          5609 => x"7f",
          5610 => x"54",
          5611 => x"82",
          5612 => x"94",
          5613 => x"39",
          5614 => x"84",
          5615 => x"06",
          5616 => x"55",
          5617 => x"c8",
          5618 => x"0d",
          5619 => x"0d",
          5620 => x"a3",
          5621 => x"5c",
          5622 => x"80",
          5623 => x"ff",
          5624 => x"a2",
          5625 => x"f5",
          5626 => x"c8",
          5627 => x"93",
          5628 => x"93",
          5629 => x"7b",
          5630 => x"08",
          5631 => x"56",
          5632 => x"2e",
          5633 => x"96",
          5634 => x"3d",
          5635 => x"a0",
          5636 => x"d1",
          5637 => x"93",
          5638 => x"82",
          5639 => x"81",
          5640 => x"52",
          5641 => x"a0",
          5642 => x"c8",
          5643 => x"93",
          5644 => x"cb",
          5645 => x"7e",
          5646 => x"3f",
          5647 => x"08",
          5648 => x"7a",
          5649 => x"3f",
          5650 => x"08",
          5651 => x"c8",
          5652 => x"38",
          5653 => x"52",
          5654 => x"f1",
          5655 => x"c8",
          5656 => x"93",
          5657 => x"38",
          5658 => x"51",
          5659 => x"82",
          5660 => x"75",
          5661 => x"76",
          5662 => x"d2",
          5663 => x"93",
          5664 => x"82",
          5665 => x"80",
          5666 => x"76",
          5667 => x"81",
          5668 => x"82",
          5669 => x"ef",
          5670 => x"ff",
          5671 => x"d4",
          5672 => x"ee",
          5673 => x"3d",
          5674 => x"81",
          5675 => x"52",
          5676 => x"73",
          5677 => x"38",
          5678 => x"16",
          5679 => x"51",
          5680 => x"f4",
          5681 => x"54",
          5682 => x"85",
          5683 => x"af",
          5684 => x"2e",
          5685 => x"58",
          5686 => x"3d",
          5687 => x"18",
          5688 => x"58",
          5689 => x"14",
          5690 => x"75",
          5691 => x"19",
          5692 => x"11",
          5693 => x"74",
          5694 => x"74",
          5695 => x"76",
          5696 => x"78",
          5697 => x"81",
          5698 => x"ff",
          5699 => x"08",
          5700 => x"af",
          5701 => x"70",
          5702 => x"33",
          5703 => x"81",
          5704 => x"70",
          5705 => x"52",
          5706 => x"57",
          5707 => x"2e",
          5708 => x"16",
          5709 => x"33",
          5710 => x"73",
          5711 => x"16",
          5712 => x"26",
          5713 => x"58",
          5714 => x"94",
          5715 => x"54",
          5716 => x"70",
          5717 => x"34",
          5718 => x"75",
          5719 => x"38",
          5720 => x"81",
          5721 => x"81",
          5722 => x"83",
          5723 => x"76",
          5724 => x"3d",
          5725 => x"1a",
          5726 => x"33",
          5727 => x"05",
          5728 => x"79",
          5729 => x"80",
          5730 => x"82",
          5731 => x"a1",
          5732 => x"f4",
          5733 => x"60",
          5734 => x"05",
          5735 => x"59",
          5736 => x"3f",
          5737 => x"08",
          5738 => x"c8",
          5739 => x"91",
          5740 => x"79",
          5741 => x"38",
          5742 => x"f9",
          5743 => x"08",
          5744 => x"38",
          5745 => x"70",
          5746 => x"81",
          5747 => x"56",
          5748 => x"8c",
          5749 => x"94",
          5750 => x"80",
          5751 => x"0c",
          5752 => x"2e",
          5753 => x"7c",
          5754 => x"70",
          5755 => x"51",
          5756 => x"2e",
          5757 => x"52",
          5758 => x"ff",
          5759 => x"82",
          5760 => x"ff",
          5761 => x"70",
          5762 => x"ff",
          5763 => x"82",
          5764 => x"75",
          5765 => x"78",
          5766 => x"94",
          5767 => x"94",
          5768 => x"98",
          5769 => x"58",
          5770 => x"88",
          5771 => x"75",
          5772 => x"52",
          5773 => x"a7",
          5774 => x"c8",
          5775 => x"93",
          5776 => x"2e",
          5777 => x"8b",
          5778 => x"91",
          5779 => x"55",
          5780 => x"82",
          5781 => x"ff",
          5782 => x"06",
          5783 => x"0b",
          5784 => x"81",
          5785 => x"39",
          5786 => x"08",
          5787 => x"75",
          5788 => x"75",
          5789 => x"a1",
          5790 => x"27",
          5791 => x"77",
          5792 => x"18",
          5793 => x"19",
          5794 => x"33",
          5795 => x"70",
          5796 => x"57",
          5797 => x"80",
          5798 => x"75",
          5799 => x"c8",
          5800 => x"93",
          5801 => x"82",
          5802 => x"94",
          5803 => x"c8",
          5804 => x"39",
          5805 => x"51",
          5806 => x"82",
          5807 => x"56",
          5808 => x"81",
          5809 => x"76",
          5810 => x"7c",
          5811 => x"08",
          5812 => x"38",
          5813 => x"18",
          5814 => x"81",
          5815 => x"98",
          5816 => x"79",
          5817 => x"38",
          5818 => x"18",
          5819 => x"77",
          5820 => x"55",
          5821 => x"a1",
          5822 => x"7c",
          5823 => x"3f",
          5824 => x"08",
          5825 => x"0b",
          5826 => x"82",
          5827 => x"39",
          5828 => x"82",
          5829 => x"05",
          5830 => x"08",
          5831 => x"27",
          5832 => x"17",
          5833 => x"0c",
          5834 => x"80",
          5835 => x"74",
          5836 => x"94",
          5837 => x"ff",
          5838 => x"80",
          5839 => x"38",
          5840 => x"7b",
          5841 => x"38",
          5842 => x"70",
          5843 => x"5c",
          5844 => x"b0",
          5845 => x"9c",
          5846 => x"a8",
          5847 => x"81",
          5848 => x"55",
          5849 => x"3f",
          5850 => x"08",
          5851 => x"38",
          5852 => x"18",
          5853 => x"bd",
          5854 => x"33",
          5855 => x"55",
          5856 => x"34",
          5857 => x"53",
          5858 => x"7c",
          5859 => x"52",
          5860 => x"eb",
          5861 => x"c8",
          5862 => x"93",
          5863 => x"91",
          5864 => x"55",
          5865 => x"0b",
          5866 => x"81",
          5867 => x"7a",
          5868 => x"79",
          5869 => x"93",
          5870 => x"3d",
          5871 => x"3d",
          5872 => x"89",
          5873 => x"2e",
          5874 => x"80",
          5875 => x"fc",
          5876 => x"3d",
          5877 => x"de",
          5878 => x"93",
          5879 => x"82",
          5880 => x"80",
          5881 => x"76",
          5882 => x"75",
          5883 => x"3f",
          5884 => x"08",
          5885 => x"c8",
          5886 => x"38",
          5887 => x"70",
          5888 => x"57",
          5889 => x"a6",
          5890 => x"33",
          5891 => x"70",
          5892 => x"55",
          5893 => x"2e",
          5894 => x"16",
          5895 => x"51",
          5896 => x"82",
          5897 => x"88",
          5898 => x"39",
          5899 => x"95",
          5900 => x"86",
          5901 => x"17",
          5902 => x"75",
          5903 => x"3f",
          5904 => x"08",
          5905 => x"2e",
          5906 => x"83",
          5907 => x"74",
          5908 => x"38",
          5909 => x"74",
          5910 => x"93",
          5911 => x"3d",
          5912 => x"3d",
          5913 => x"3d",
          5914 => x"70",
          5915 => x"b9",
          5916 => x"c8",
          5917 => x"93",
          5918 => x"38",
          5919 => x"08",
          5920 => x"82",
          5921 => x"86",
          5922 => x"fb",
          5923 => x"79",
          5924 => x"05",
          5925 => x"56",
          5926 => x"3f",
          5927 => x"08",
          5928 => x"c8",
          5929 => x"38",
          5930 => x"82",
          5931 => x"52",
          5932 => x"c5",
          5933 => x"c8",
          5934 => x"39",
          5935 => x"51",
          5936 => x"82",
          5937 => x"53",
          5938 => x"08",
          5939 => x"81",
          5940 => x"80",
          5941 => x"38",
          5942 => x"51",
          5943 => x"72",
          5944 => x"c9",
          5945 => x"93",
          5946 => x"82",
          5947 => x"84",
          5948 => x"06",
          5949 => x"53",
          5950 => x"c8",
          5951 => x"0d",
          5952 => x"0d",
          5953 => x"53",
          5954 => x"53",
          5955 => x"54",
          5956 => x"82",
          5957 => x"55",
          5958 => x"08",
          5959 => x"52",
          5960 => x"e9",
          5961 => x"c8",
          5962 => x"93",
          5963 => x"38",
          5964 => x"05",
          5965 => x"2b",
          5966 => x"80",
          5967 => x"86",
          5968 => x"75",
          5969 => x"38",
          5970 => x"3d",
          5971 => x"d0",
          5972 => x"82",
          5973 => x"93",
          5974 => x"f2",
          5975 => x"63",
          5976 => x"53",
          5977 => x"05",
          5978 => x"51",
          5979 => x"82",
          5980 => x"59",
          5981 => x"08",
          5982 => x"7a",
          5983 => x"08",
          5984 => x"fe",
          5985 => x"90",
          5986 => x"26",
          5987 => x"15",
          5988 => x"81",
          5989 => x"59",
          5990 => x"82",
          5991 => x"39",
          5992 => x"33",
          5993 => x"73",
          5994 => x"81",
          5995 => x"38",
          5996 => x"56",
          5997 => x"3d",
          5998 => x"ff",
          5999 => x"82",
          6000 => x"ff",
          6001 => x"82",
          6002 => x"81",
          6003 => x"82",
          6004 => x"30",
          6005 => x"c8",
          6006 => x"25",
          6007 => x"18",
          6008 => x"58",
          6009 => x"08",
          6010 => x"38",
          6011 => x"7a",
          6012 => x"a4",
          6013 => x"57",
          6014 => x"74",
          6015 => x"52",
          6016 => x"52",
          6017 => x"c0",
          6018 => x"c8",
          6019 => x"93",
          6020 => x"d5",
          6021 => x"33",
          6022 => x"82",
          6023 => x"06",
          6024 => x"15",
          6025 => x"ff",
          6026 => x"82",
          6027 => x"83",
          6028 => x"70",
          6029 => x"25",
          6030 => x"58",
          6031 => x"9d",
          6032 => x"b4",
          6033 => x"b5",
          6034 => x"93",
          6035 => x"0a",
          6036 => x"70",
          6037 => x"84",
          6038 => x"51",
          6039 => x"ff",
          6040 => x"57",
          6041 => x"93",
          6042 => x"0c",
          6043 => x"12",
          6044 => x"84",
          6045 => x"07",
          6046 => x"84",
          6047 => x"82",
          6048 => x"90",
          6049 => x"f8",
          6050 => x"8b",
          6051 => x"53",
          6052 => x"e0",
          6053 => x"93",
          6054 => x"82",
          6055 => x"8a",
          6056 => x"33",
          6057 => x"2e",
          6058 => x"56",
          6059 => x"90",
          6060 => x"81",
          6061 => x"06",
          6062 => x"87",
          6063 => x"2e",
          6064 => x"94",
          6065 => x"19",
          6066 => x"bc",
          6067 => x"08",
          6068 => x"53",
          6069 => x"52",
          6070 => x"be",
          6071 => x"93",
          6072 => x"80",
          6073 => x"0c",
          6074 => x"98",
          6075 => x"77",
          6076 => x"f4",
          6077 => x"c8",
          6078 => x"c8",
          6079 => x"70",
          6080 => x"07",
          6081 => x"57",
          6082 => x"93",
          6083 => x"2e",
          6084 => x"83",
          6085 => x"76",
          6086 => x"55",
          6087 => x"08",
          6088 => x"98",
          6089 => x"75",
          6090 => x"ff",
          6091 => x"82",
          6092 => x"57",
          6093 => x"8c",
          6094 => x"18",
          6095 => x"07",
          6096 => x"19",
          6097 => x"38",
          6098 => x"55",
          6099 => x"ab",
          6100 => x"9c",
          6101 => x"a8",
          6102 => x"81",
          6103 => x"55",
          6104 => x"3f",
          6105 => x"08",
          6106 => x"38",
          6107 => x"39",
          6108 => x"80",
          6109 => x"74",
          6110 => x"76",
          6111 => x"38",
          6112 => x"34",
          6113 => x"39",
          6114 => x"82",
          6115 => x"8a",
          6116 => x"e3",
          6117 => x"fb",
          6118 => x"96",
          6119 => x"53",
          6120 => x"a4",
          6121 => x"3d",
          6122 => x"3f",
          6123 => x"08",
          6124 => x"c8",
          6125 => x"38",
          6126 => x"51",
          6127 => x"3f",
          6128 => x"52",
          6129 => x"05",
          6130 => x"3f",
          6131 => x"08",
          6132 => x"52",
          6133 => x"9a",
          6134 => x"ae",
          6135 => x"f7",
          6136 => x"85",
          6137 => x"06",
          6138 => x"73",
          6139 => x"38",
          6140 => x"82",
          6141 => x"fb",
          6142 => x"95",
          6143 => x"80",
          6144 => x"70",
          6145 => x"55",
          6146 => x"85",
          6147 => x"90",
          6148 => x"d2",
          6149 => x"06",
          6150 => x"2e",
          6151 => x"56",
          6152 => x"38",
          6153 => x"51",
          6154 => x"82",
          6155 => x"02",
          6156 => x"d2",
          6157 => x"84",
          6158 => x"06",
          6159 => x"57",
          6160 => x"80",
          6161 => x"fb",
          6162 => x"95",
          6163 => x"78",
          6164 => x"14",
          6165 => x"80",
          6166 => x"fb",
          6167 => x"95",
          6168 => x"59",
          6169 => x"fb",
          6170 => x"95",
          6171 => x"52",
          6172 => x"52",
          6173 => x"3f",
          6174 => x"08",
          6175 => x"c8",
          6176 => x"38",
          6177 => x"08",
          6178 => x"c6",
          6179 => x"93",
          6180 => x"82",
          6181 => x"83",
          6182 => x"75",
          6183 => x"30",
          6184 => x"9f",
          6185 => x"58",
          6186 => x"80",
          6187 => x"fb",
          6188 => x"94",
          6189 => x"3d",
          6190 => x"c9",
          6191 => x"93",
          6192 => x"93",
          6193 => x"70",
          6194 => x"08",
          6195 => x"79",
          6196 => x"07",
          6197 => x"06",
          6198 => x"56",
          6199 => x"2e",
          6200 => x"fb",
          6201 => x"94",
          6202 => x"53",
          6203 => x"3d",
          6204 => x"ff",
          6205 => x"82",
          6206 => x"56",
          6207 => x"77",
          6208 => x"8b",
          6209 => x"c8",
          6210 => x"fb",
          6211 => x"93",
          6212 => x"82",
          6213 => x"9f",
          6214 => x"ea",
          6215 => x"53",
          6216 => x"05",
          6217 => x"51",
          6218 => x"82",
          6219 => x"55",
          6220 => x"08",
          6221 => x"77",
          6222 => x"98",
          6223 => x"51",
          6224 => x"82",
          6225 => x"55",
          6226 => x"08",
          6227 => x"55",
          6228 => x"09",
          6229 => x"93",
          6230 => x"db",
          6231 => x"85",
          6232 => x"06",
          6233 => x"73",
          6234 => x"38",
          6235 => x"84",
          6236 => x"06",
          6237 => x"77",
          6238 => x"98",
          6239 => x"51",
          6240 => x"3f",
          6241 => x"08",
          6242 => x"82",
          6243 => x"75",
          6244 => x"06",
          6245 => x"55",
          6246 => x"09",
          6247 => x"38",
          6248 => x"ff",
          6249 => x"06",
          6250 => x"55",
          6251 => x"0a",
          6252 => x"aa",
          6253 => x"77",
          6254 => x"c7",
          6255 => x"c8",
          6256 => x"93",
          6257 => x"96",
          6258 => x"a0",
          6259 => x"51",
          6260 => x"3f",
          6261 => x"0b",
          6262 => x"77",
          6263 => x"bf",
          6264 => x"52",
          6265 => x"51",
          6266 => x"3f",
          6267 => x"18",
          6268 => x"c3",
          6269 => x"53",
          6270 => x"80",
          6271 => x"ff",
          6272 => x"77",
          6273 => x"80",
          6274 => x"7e",
          6275 => x"18",
          6276 => x"c3",
          6277 => x"54",
          6278 => x"15",
          6279 => x"d4",
          6280 => x"e7",
          6281 => x"c8",
          6282 => x"93",
          6283 => x"38",
          6284 => x"96",
          6285 => x"ae",
          6286 => x"53",
          6287 => x"51",
          6288 => x"63",
          6289 => x"8b",
          6290 => x"54",
          6291 => x"15",
          6292 => x"ff",
          6293 => x"82",
          6294 => x"55",
          6295 => x"53",
          6296 => x"3d",
          6297 => x"ff",
          6298 => x"74",
          6299 => x"0c",
          6300 => x"04",
          6301 => x"a8",
          6302 => x"51",
          6303 => x"82",
          6304 => x"ff",
          6305 => x"a8",
          6306 => x"d1",
          6307 => x"c8",
          6308 => x"93",
          6309 => x"d7",
          6310 => x"a8",
          6311 => x"a7",
          6312 => x"51",
          6313 => x"82",
          6314 => x"55",
          6315 => x"08",
          6316 => x"02",
          6317 => x"33",
          6318 => x"54",
          6319 => x"83",
          6320 => x"74",
          6321 => x"a0",
          6322 => x"08",
          6323 => x"ff",
          6324 => x"ff",
          6325 => x"ac",
          6326 => x"d4",
          6327 => x"3d",
          6328 => x"ff",
          6329 => x"a9",
          6330 => x"73",
          6331 => x"3f",
          6332 => x"08",
          6333 => x"c8",
          6334 => x"62",
          6335 => x"81",
          6336 => x"84",
          6337 => x"3d",
          6338 => x"38",
          6339 => x"84",
          6340 => x"06",
          6341 => x"a7",
          6342 => x"05",
          6343 => x"3f",
          6344 => x"08",
          6345 => x"c8",
          6346 => x"38",
          6347 => x"53",
          6348 => x"95",
          6349 => x"16",
          6350 => x"ed",
          6351 => x"05",
          6352 => x"34",
          6353 => x"70",
          6354 => x"81",
          6355 => x"57",
          6356 => x"76",
          6357 => x"73",
          6358 => x"77",
          6359 => x"83",
          6360 => x"16",
          6361 => x"2a",
          6362 => x"51",
          6363 => x"80",
          6364 => x"38",
          6365 => x"80",
          6366 => x"52",
          6367 => x"bf",
          6368 => x"93",
          6369 => x"77",
          6370 => x"b2",
          6371 => x"82",
          6372 => x"80",
          6373 => x"82",
          6374 => x"52",
          6375 => x"ae",
          6376 => x"93",
          6377 => x"d4",
          6378 => x"82",
          6379 => x"bf",
          6380 => x"33",
          6381 => x"2e",
          6382 => x"92",
          6383 => x"75",
          6384 => x"ff",
          6385 => x"77",
          6386 => x"83",
          6387 => x"9f",
          6388 => x"d4",
          6389 => x"89",
          6390 => x"c8",
          6391 => x"93",
          6392 => x"38",
          6393 => x"ae",
          6394 => x"93",
          6395 => x"74",
          6396 => x"0c",
          6397 => x"04",
          6398 => x"02",
          6399 => x"33",
          6400 => x"80",
          6401 => x"57",
          6402 => x"95",
          6403 => x"52",
          6404 => x"cd",
          6405 => x"93",
          6406 => x"82",
          6407 => x"80",
          6408 => x"5a",
          6409 => x"3d",
          6410 => x"c7",
          6411 => x"93",
          6412 => x"82",
          6413 => x"bd",
          6414 => x"cf",
          6415 => x"a0",
          6416 => x"80",
          6417 => x"86",
          6418 => x"38",
          6419 => x"61",
          6420 => x"12",
          6421 => x"7a",
          6422 => x"51",
          6423 => x"74",
          6424 => x"78",
          6425 => x"83",
          6426 => x"51",
          6427 => x"3f",
          6428 => x"08",
          6429 => x"93",
          6430 => x"3d",
          6431 => x"3d",
          6432 => x"82",
          6433 => x"d0",
          6434 => x"3d",
          6435 => x"3f",
          6436 => x"08",
          6437 => x"c8",
          6438 => x"38",
          6439 => x"52",
          6440 => x"05",
          6441 => x"3f",
          6442 => x"08",
          6443 => x"c8",
          6444 => x"02",
          6445 => x"33",
          6446 => x"54",
          6447 => x"83",
          6448 => x"74",
          6449 => x"16",
          6450 => x"22",
          6451 => x"72",
          6452 => x"54",
          6453 => x"51",
          6454 => x"3f",
          6455 => x"0b",
          6456 => x"77",
          6457 => x"a7",
          6458 => x"c8",
          6459 => x"82",
          6460 => x"94",
          6461 => x"ea",
          6462 => x"6b",
          6463 => x"53",
          6464 => x"05",
          6465 => x"51",
          6466 => x"82",
          6467 => x"82",
          6468 => x"30",
          6469 => x"c8",
          6470 => x"25",
          6471 => x"7d",
          6472 => x"72",
          6473 => x"51",
          6474 => x"80",
          6475 => x"38",
          6476 => x"5f",
          6477 => x"3d",
          6478 => x"ff",
          6479 => x"82",
          6480 => x"56",
          6481 => x"08",
          6482 => x"81",
          6483 => x"ff",
          6484 => x"82",
          6485 => x"56",
          6486 => x"08",
          6487 => x"93",
          6488 => x"93",
          6489 => x"5c",
          6490 => x"17",
          6491 => x"1a",
          6492 => x"74",
          6493 => x"81",
          6494 => x"77",
          6495 => x"77",
          6496 => x"74",
          6497 => x"2e",
          6498 => x"18",
          6499 => x"33",
          6500 => x"73",
          6501 => x"38",
          6502 => x"09",
          6503 => x"38",
          6504 => x"80",
          6505 => x"70",
          6506 => x"25",
          6507 => x"7e",
          6508 => x"72",
          6509 => x"51",
          6510 => x"2e",
          6511 => x"a0",
          6512 => x"51",
          6513 => x"3f",
          6514 => x"08",
          6515 => x"c8",
          6516 => x"7b",
          6517 => x"54",
          6518 => x"73",
          6519 => x"38",
          6520 => x"73",
          6521 => x"38",
          6522 => x"18",
          6523 => x"ff",
          6524 => x"82",
          6525 => x"7b",
          6526 => x"93",
          6527 => x"3d",
          6528 => x"3d",
          6529 => x"9a",
          6530 => x"05",
          6531 => x"51",
          6532 => x"82",
          6533 => x"55",
          6534 => x"08",
          6535 => x"8b",
          6536 => x"9a",
          6537 => x"05",
          6538 => x"a1",
          6539 => x"70",
          6540 => x"57",
          6541 => x"74",
          6542 => x"38",
          6543 => x"81",
          6544 => x"81",
          6545 => x"56",
          6546 => x"3f",
          6547 => x"08",
          6548 => x"38",
          6549 => x"70",
          6550 => x"ff",
          6551 => x"82",
          6552 => x"80",
          6553 => x"75",
          6554 => x"07",
          6555 => x"4c",
          6556 => x"80",
          6557 => x"16",
          6558 => x"26",
          6559 => x"16",
          6560 => x"ff",
          6561 => x"80",
          6562 => x"87",
          6563 => x"f8",
          6564 => x"75",
          6565 => x"38",
          6566 => x"fc",
          6567 => x"a6",
          6568 => x"93",
          6569 => x"38",
          6570 => x"27",
          6571 => x"89",
          6572 => x"8b",
          6573 => x"27",
          6574 => x"55",
          6575 => x"81",
          6576 => x"93",
          6577 => x"77",
          6578 => x"05",
          6579 => x"55",
          6580 => x"34",
          6581 => x"9a",
          6582 => x"ff",
          6583 => x"75",
          6584 => x"17",
          6585 => x"56",
          6586 => x"9f",
          6587 => x"38",
          6588 => x"54",
          6589 => x"81",
          6590 => x"ea",
          6591 => x"2e",
          6592 => x"9f",
          6593 => x"12",
          6594 => x"52",
          6595 => x"a0",
          6596 => x"06",
          6597 => x"17",
          6598 => x"2e",
          6599 => x"15",
          6600 => x"54",
          6601 => x"ee",
          6602 => x"80",
          6603 => x"8f",
          6604 => x"55",
          6605 => x"3f",
          6606 => x"08",
          6607 => x"c8",
          6608 => x"38",
          6609 => x"51",
          6610 => x"3f",
          6611 => x"08",
          6612 => x"c8",
          6613 => x"76",
          6614 => x"38",
          6615 => x"3d",
          6616 => x"52",
          6617 => x"a4",
          6618 => x"39",
          6619 => x"74",
          6620 => x"81",
          6621 => x"34",
          6622 => x"a7",
          6623 => x"93",
          6624 => x"80",
          6625 => x"93",
          6626 => x"2e",
          6627 => x"80",
          6628 => x"54",
          6629 => x"80",
          6630 => x"52",
          6631 => x"05",
          6632 => x"b2",
          6633 => x"c8",
          6634 => x"93",
          6635 => x"38",
          6636 => x"93",
          6637 => x"65",
          6638 => x"91",
          6639 => x"88",
          6640 => x"34",
          6641 => x"3d",
          6642 => x"52",
          6643 => x"a3",
          6644 => x"54",
          6645 => x"15",
          6646 => x"ff",
          6647 => x"82",
          6648 => x"54",
          6649 => x"82",
          6650 => x"9a",
          6651 => x"f1",
          6652 => x"63",
          6653 => x"80",
          6654 => x"94",
          6655 => x"55",
          6656 => x"5c",
          6657 => x"3f",
          6658 => x"08",
          6659 => x"c8",
          6660 => x"91",
          6661 => x"76",
          6662 => x"38",
          6663 => x"b7",
          6664 => x"2e",
          6665 => x"18",
          6666 => x"90",
          6667 => x"81",
          6668 => x"06",
          6669 => x"73",
          6670 => x"54",
          6671 => x"82",
          6672 => x"39",
          6673 => x"84",
          6674 => x"11",
          6675 => x"2b",
          6676 => x"54",
          6677 => x"fe",
          6678 => x"ff",
          6679 => x"70",
          6680 => x"07",
          6681 => x"93",
          6682 => x"62",
          6683 => x"5d",
          6684 => x"55",
          6685 => x"79",
          6686 => x"98",
          6687 => x"26",
          6688 => x"59",
          6689 => x"5d",
          6690 => x"52",
          6691 => x"a6",
          6692 => x"93",
          6693 => x"16",
          6694 => x"56",
          6695 => x"75",
          6696 => x"82",
          6697 => x"2e",
          6698 => x"75",
          6699 => x"94",
          6700 => x"38",
          6701 => x"79",
          6702 => x"38",
          6703 => x"5d",
          6704 => x"79",
          6705 => x"06",
          6706 => x"57",
          6707 => x"38",
          6708 => x"b9",
          6709 => x"57",
          6710 => x"2e",
          6711 => x"15",
          6712 => x"2e",
          6713 => x"83",
          6714 => x"73",
          6715 => x"7f",
          6716 => x"f0",
          6717 => x"c8",
          6718 => x"93",
          6719 => x"38",
          6720 => x"ff",
          6721 => x"5f",
          6722 => x"84",
          6723 => x"5f",
          6724 => x"38",
          6725 => x"12",
          6726 => x"80",
          6727 => x"7c",
          6728 => x"7a",
          6729 => x"90",
          6730 => x"c0",
          6731 => x"90",
          6732 => x"98",
          6733 => x"05",
          6734 => x"15",
          6735 => x"95",
          6736 => x"08",
          6737 => x"16",
          6738 => x"11",
          6739 => x"55",
          6740 => x"16",
          6741 => x"73",
          6742 => x"0c",
          6743 => x"04",
          6744 => x"6a",
          6745 => x"80",
          6746 => x"9b",
          6747 => x"58",
          6748 => x"3f",
          6749 => x"08",
          6750 => x"80",
          6751 => x"c8",
          6752 => x"d1",
          6753 => x"c8",
          6754 => x"82",
          6755 => x"55",
          6756 => x"2e",
          6757 => x"08",
          6758 => x"34",
          6759 => x"06",
          6760 => x"79",
          6761 => x"cb",
          6762 => x"c8",
          6763 => x"06",
          6764 => x"56",
          6765 => x"74",
          6766 => x"75",
          6767 => x"81",
          6768 => x"8a",
          6769 => x"8d",
          6770 => x"fc",
          6771 => x"52",
          6772 => x"9d",
          6773 => x"93",
          6774 => x"38",
          6775 => x"93",
          6776 => x"80",
          6777 => x"38",
          6778 => x"67",
          6779 => x"80",
          6780 => x"81",
          6781 => x"5e",
          6782 => x"86",
          6783 => x"26",
          6784 => x"81",
          6785 => x"8b",
          6786 => x"78",
          6787 => x"80",
          6788 => x"93",
          6789 => x"39",
          6790 => x"51",
          6791 => x"3f",
          6792 => x"08",
          6793 => x"6e",
          6794 => x"fe",
          6795 => x"82",
          6796 => x"7e",
          6797 => x"08",
          6798 => x"70",
          6799 => x"25",
          6800 => x"08",
          6801 => x"93",
          6802 => x"80",
          6803 => x"52",
          6804 => x"46",
          6805 => x"75",
          6806 => x"98",
          6807 => x"53",
          6808 => x"51",
          6809 => x"3f",
          6810 => x"93",
          6811 => x"e5",
          6812 => x"2a",
          6813 => x"51",
          6814 => x"74",
          6815 => x"81",
          6816 => x"bf",
          6817 => x"63",
          6818 => x"c9",
          6819 => x"31",
          6820 => x"80",
          6821 => x"8a",
          6822 => x"57",
          6823 => x"26",
          6824 => x"7c",
          6825 => x"81",
          6826 => x"74",
          6827 => x"38",
          6828 => x"55",
          6829 => x"88",
          6830 => x"06",
          6831 => x"38",
          6832 => x"39",
          6833 => x"55",
          6834 => x"42",
          6835 => x"8a",
          6836 => x"59",
          6837 => x"09",
          6838 => x"f1",
          6839 => x"38",
          6840 => x"78",
          6841 => x"0b",
          6842 => x"70",
          6843 => x"58",
          6844 => x"80",
          6845 => x"74",
          6846 => x"38",
          6847 => x"10",
          6848 => x"70",
          6849 => x"5a",
          6850 => x"2e",
          6851 => x"75",
          6852 => x"78",
          6853 => x"fe",
          6854 => x"82",
          6855 => x"82",
          6856 => x"10",
          6857 => x"54",
          6858 => x"56",
          6859 => x"3f",
          6860 => x"08",
          6861 => x"80",
          6862 => x"8a",
          6863 => x"fd",
          6864 => x"75",
          6865 => x"38",
          6866 => x"89",
          6867 => x"38",
          6868 => x"78",
          6869 => x"0b",
          6870 => x"70",
          6871 => x"58",
          6872 => x"80",
          6873 => x"74",
          6874 => x"38",
          6875 => x"10",
          6876 => x"70",
          6877 => x"5a",
          6878 => x"2e",
          6879 => x"75",
          6880 => x"78",
          6881 => x"fe",
          6882 => x"82",
          6883 => x"10",
          6884 => x"82",
          6885 => x"9f",
          6886 => x"38",
          6887 => x"93",
          6888 => x"29",
          6889 => x"2a",
          6890 => x"58",
          6891 => x"76",
          6892 => x"51",
          6893 => x"3f",
          6894 => x"08",
          6895 => x"53",
          6896 => x"80",
          6897 => x"ef",
          6898 => x"c8",
          6899 => x"ff",
          6900 => x"1b",
          6901 => x"05",
          6902 => x"05",
          6903 => x"72",
          6904 => x"52",
          6905 => x"40",
          6906 => x"09",
          6907 => x"38",
          6908 => x"18",
          6909 => x"39",
          6910 => x"78",
          6911 => x"70",
          6912 => x"55",
          6913 => x"87",
          6914 => x"7b",
          6915 => x"79",
          6916 => x"31",
          6917 => x"f2",
          6918 => x"93",
          6919 => x"61",
          6920 => x"81",
          6921 => x"82",
          6922 => x"83",
          6923 => x"91",
          6924 => x"38",
          6925 => x"58",
          6926 => x"38",
          6927 => x"95",
          6928 => x"2e",
          6929 => x"80",
          6930 => x"ff",
          6931 => x"b4",
          6932 => x"38",
          6933 => x"74",
          6934 => x"86",
          6935 => x"fc",
          6936 => x"81",
          6937 => x"55",
          6938 => x"86",
          6939 => x"fc",
          6940 => x"8b",
          6941 => x"58",
          6942 => x"27",
          6943 => x"8e",
          6944 => x"39",
          6945 => x"26",
          6946 => x"8b",
          6947 => x"58",
          6948 => x"27",
          6949 => x"8e",
          6950 => x"39",
          6951 => x"81",
          6952 => x"06",
          6953 => x"55",
          6954 => x"26",
          6955 => x"8e",
          6956 => x"a1",
          6957 => x"80",
          6958 => x"ff",
          6959 => x"8b",
          6960 => x"b4",
          6961 => x"ff",
          6962 => x"7d",
          6963 => x"51",
          6964 => x"3f",
          6965 => x"05",
          6966 => x"ff",
          6967 => x"8e",
          6968 => x"98",
          6969 => x"7f",
          6970 => x"61",
          6971 => x"30",
          6972 => x"84",
          6973 => x"51",
          6974 => x"51",
          6975 => x"3f",
          6976 => x"ff",
          6977 => x"02",
          6978 => x"22",
          6979 => x"51",
          6980 => x"3f",
          6981 => x"52",
          6982 => x"ff",
          6983 => x"f8",
          6984 => x"34",
          6985 => x"1f",
          6986 => x"b0",
          6987 => x"52",
          6988 => x"ff",
          6989 => x"63",
          6990 => x"51",
          6991 => x"3f",
          6992 => x"09",
          6993 => x"cf",
          6994 => x"b2",
          6995 => x"c3",
          6996 => x"98",
          6997 => x"52",
          6998 => x"ff",
          6999 => x"82",
          7000 => x"51",
          7001 => x"3f",
          7002 => x"1f",
          7003 => x"ec",
          7004 => x"b2",
          7005 => x"97",
          7006 => x"80",
          7007 => x"05",
          7008 => x"80",
          7009 => x"93",
          7010 => x"c0",
          7011 => x"1f",
          7012 => x"95",
          7013 => x"82",
          7014 => x"52",
          7015 => x"ff",
          7016 => x"7b",
          7017 => x"06",
          7018 => x"51",
          7019 => x"3f",
          7020 => x"a4",
          7021 => x"7f",
          7022 => x"93",
          7023 => x"d4",
          7024 => x"51",
          7025 => x"3f",
          7026 => x"52",
          7027 => x"51",
          7028 => x"3f",
          7029 => x"53",
          7030 => x"51",
          7031 => x"3f",
          7032 => x"93",
          7033 => x"ed",
          7034 => x"2e",
          7035 => x"80",
          7036 => x"54",
          7037 => x"53",
          7038 => x"51",
          7039 => x"3f",
          7040 => x"52",
          7041 => x"97",
          7042 => x"8b",
          7043 => x"52",
          7044 => x"96",
          7045 => x"8a",
          7046 => x"52",
          7047 => x"51",
          7048 => x"3f",
          7049 => x"83",
          7050 => x"ff",
          7051 => x"82",
          7052 => x"1f",
          7053 => x"c2",
          7054 => x"d5",
          7055 => x"1f",
          7056 => x"98",
          7057 => x"63",
          7058 => x"7e",
          7059 => x"ff",
          7060 => x"81",
          7061 => x"05",
          7062 => x"79",
          7063 => x"f8",
          7064 => x"80",
          7065 => x"ff",
          7066 => x"7f",
          7067 => x"61",
          7068 => x"81",
          7069 => x"f8",
          7070 => x"ff",
          7071 => x"ff",
          7072 => x"51",
          7073 => x"3f",
          7074 => x"88",
          7075 => x"95",
          7076 => x"39",
          7077 => x"f8",
          7078 => x"2e",
          7079 => x"55",
          7080 => x"51",
          7081 => x"3f",
          7082 => x"57",
          7083 => x"83",
          7084 => x"76",
          7085 => x"7e",
          7086 => x"ff",
          7087 => x"82",
          7088 => x"82",
          7089 => x"53",
          7090 => x"51",
          7091 => x"3f",
          7092 => x"78",
          7093 => x"74",
          7094 => x"1b",
          7095 => x"2e",
          7096 => x"78",
          7097 => x"2e",
          7098 => x"55",
          7099 => x"61",
          7100 => x"74",
          7101 => x"75",
          7102 => x"79",
          7103 => x"d8",
          7104 => x"c8",
          7105 => x"38",
          7106 => x"78",
          7107 => x"74",
          7108 => x"57",
          7109 => x"93",
          7110 => x"65",
          7111 => x"26",
          7112 => x"57",
          7113 => x"83",
          7114 => x"7c",
          7115 => x"06",
          7116 => x"ff",
          7117 => x"77",
          7118 => x"ff",
          7119 => x"82",
          7120 => x"83",
          7121 => x"ff",
          7122 => x"83",
          7123 => x"77",
          7124 => x"0b",
          7125 => x"81",
          7126 => x"34",
          7127 => x"34",
          7128 => x"34",
          7129 => x"57",
          7130 => x"52",
          7131 => x"eb",
          7132 => x"0b",
          7133 => x"82",
          7134 => x"82",
          7135 => x"55",
          7136 => x"34",
          7137 => x"08",
          7138 => x"63",
          7139 => x"1f",
          7140 => x"e6",
          7141 => x"83",
          7142 => x"ff",
          7143 => x"81",
          7144 => x"7e",
          7145 => x"ff",
          7146 => x"81",
          7147 => x"c8",
          7148 => x"80",
          7149 => x"79",
          7150 => x"f6",
          7151 => x"82",
          7152 => x"91",
          7153 => x"8e",
          7154 => x"81",
          7155 => x"81",
          7156 => x"80",
          7157 => x"93",
          7158 => x"3d",
          7159 => x"3d",
          7160 => x"71",
          7161 => x"e2",
          7162 => x"10",
          7163 => x"05",
          7164 => x"04",
          7165 => x"51",
          7166 => x"3f",
          7167 => x"82",
          7168 => x"ff",
          7169 => x"81",
          7170 => x"82",
          7171 => x"80",
          7172 => x"be",
          7173 => x"ac",
          7174 => x"88",
          7175 => x"39",
          7176 => x"51",
          7177 => x"3f",
          7178 => x"82",
          7179 => x"fe",
          7180 => x"81",
          7181 => x"82",
          7182 => x"ff",
          7183 => x"92",
          7184 => x"f0",
          7185 => x"dc",
          7186 => x"39",
          7187 => x"51",
          7188 => x"3f",
          7189 => x"82",
          7190 => x"fe",
          7191 => x"80",
          7192 => x"83",
          7193 => x"ff",
          7194 => x"e6",
          7195 => x"d4",
          7196 => x"b0",
          7197 => x"39",
          7198 => x"51",
          7199 => x"3f",
          7200 => x"82",
          7201 => x"fe",
          7202 => x"80",
          7203 => x"84",
          7204 => x"ff",
          7205 => x"39",
          7206 => x"51",
          7207 => x"3f",
          7208 => x"84",
          7209 => x"fe",
          7210 => x"39",
          7211 => x"51",
          7212 => x"3f",
          7213 => x"85",
          7214 => x"fe",
          7215 => x"39",
          7216 => x"51",
          7217 => x"3f",
          7218 => x"85",
          7219 => x"fe",
          7220 => x"3d",
          7221 => x"3d",
          7222 => x"56",
          7223 => x"e7",
          7224 => x"74",
          7225 => x"e8",
          7226 => x"e8",
          7227 => x"93",
          7228 => x"9a",
          7229 => x"52",
          7230 => x"e8",
          7231 => x"93",
          7232 => x"75",
          7233 => x"af",
          7234 => x"c8",
          7235 => x"54",
          7236 => x"52",
          7237 => x"51",
          7238 => x"3f",
          7239 => x"04",
          7240 => x"0d",
          7241 => x"08",
          7242 => x"08",
          7243 => x"84",
          7244 => x"71",
          7245 => x"75",
          7246 => x"87",
          7247 => x"07",
          7248 => x"5c",
          7249 => x"55",
          7250 => x"38",
          7251 => x"52",
          7252 => x"fb",
          7253 => x"ff",
          7254 => x"82",
          7255 => x"58",
          7256 => x"08",
          7257 => x"93",
          7258 => x"c0",
          7259 => x"82",
          7260 => x"59",
          7261 => x"fb",
          7262 => x"55",
          7263 => x"76",
          7264 => x"15",
          7265 => x"3f",
          7266 => x"08",
          7267 => x"c8",
          7268 => x"7a",
          7269 => x"38",
          7270 => x"18",
          7271 => x"39",
          7272 => x"fb",
          7273 => x"ca",
          7274 => x"30",
          7275 => x"80",
          7276 => x"70",
          7277 => x"06",
          7278 => x"56",
          7279 => x"90",
          7280 => x"e4",
          7281 => x"98",
          7282 => x"78",
          7283 => x"3f",
          7284 => x"82",
          7285 => x"81",
          7286 => x"04",
          7287 => x"02",
          7288 => x"57",
          7289 => x"59",
          7290 => x"52",
          7291 => x"b0",
          7292 => x"c8",
          7293 => x"76",
          7294 => x"38",
          7295 => x"98",
          7296 => x"61",
          7297 => x"82",
          7298 => x"7f",
          7299 => x"75",
          7300 => x"c8",
          7301 => x"39",
          7302 => x"82",
          7303 => x"8a",
          7304 => x"fb",
          7305 => x"9f",
          7306 => x"85",
          7307 => x"85",
          7308 => x"ff",
          7309 => x"82",
          7310 => x"22",
          7311 => x"f9",
          7312 => x"86",
          7313 => x"86",
          7314 => x"15",
          7315 => x"86",
          7316 => x"81",
          7317 => x"80",
          7318 => x"fe",
          7319 => x"87",
          7320 => x"fe",
          7321 => x"c0",
          7322 => x"53",
          7323 => x"3f",
          7324 => x"ee",
          7325 => x"86",
          7326 => x"f0",
          7327 => x"51",
          7328 => x"3f",
          7329 => x"70",
          7330 => x"52",
          7331 => x"95",
          7332 => x"fe",
          7333 => x"82",
          7334 => x"fe",
          7335 => x"80",
          7336 => x"d0",
          7337 => x"2a",
          7338 => x"51",
          7339 => x"2e",
          7340 => x"51",
          7341 => x"3f",
          7342 => x"51",
          7343 => x"3f",
          7344 => x"ee",
          7345 => x"83",
          7346 => x"06",
          7347 => x"80",
          7348 => x"81",
          7349 => x"9c",
          7350 => x"f0",
          7351 => x"92",
          7352 => x"fe",
          7353 => x"72",
          7354 => x"81",
          7355 => x"71",
          7356 => x"38",
          7357 => x"ed",
          7358 => x"87",
          7359 => x"ef",
          7360 => x"51",
          7361 => x"3f",
          7362 => x"70",
          7363 => x"52",
          7364 => x"95",
          7365 => x"fe",
          7366 => x"82",
          7367 => x"fe",
          7368 => x"80",
          7369 => x"cc",
          7370 => x"2a",
          7371 => x"51",
          7372 => x"2e",
          7373 => x"51",
          7374 => x"3f",
          7375 => x"51",
          7376 => x"3f",
          7377 => x"ed",
          7378 => x"87",
          7379 => x"06",
          7380 => x"80",
          7381 => x"81",
          7382 => x"98",
          7383 => x"c0",
          7384 => x"8e",
          7385 => x"fe",
          7386 => x"72",
          7387 => x"81",
          7388 => x"71",
          7389 => x"38",
          7390 => x"ec",
          7391 => x"87",
          7392 => x"ee",
          7393 => x"51",
          7394 => x"3f",
          7395 => x"3f",
          7396 => x"04",
          7397 => x"78",
          7398 => x"55",
          7399 => x"80",
          7400 => x"38",
          7401 => x"77",
          7402 => x"33",
          7403 => x"39",
          7404 => x"80",
          7405 => x"54",
          7406 => x"83",
          7407 => x"72",
          7408 => x"2a",
          7409 => x"53",
          7410 => x"74",
          7411 => x"a0",
          7412 => x"06",
          7413 => x"75",
          7414 => x"57",
          7415 => x"75",
          7416 => x"8c",
          7417 => x"08",
          7418 => x"52",
          7419 => x"d0",
          7420 => x"c8",
          7421 => x"84",
          7422 => x"72",
          7423 => x"a6",
          7424 => x"70",
          7425 => x"57",
          7426 => x"27",
          7427 => x"53",
          7428 => x"c8",
          7429 => x"0d",
          7430 => x"0d",
          7431 => x"b6",
          7432 => x"0c",
          7433 => x"8c",
          7434 => x"7b",
          7435 => x"c3",
          7436 => x"c8",
          7437 => x"06",
          7438 => x"2e",
          7439 => x"9f",
          7440 => x"94",
          7441 => x"70",
          7442 => x"fd",
          7443 => x"53",
          7444 => x"b0",
          7445 => x"b5",
          7446 => x"93",
          7447 => x"79",
          7448 => x"38",
          7449 => x"51",
          7450 => x"3f",
          7451 => x"70",
          7452 => x"88",
          7453 => x"f7",
          7454 => x"3d",
          7455 => x"80",
          7456 => x"5a",
          7457 => x"51",
          7458 => x"3f",
          7459 => x"51",
          7460 => x"3f",
          7461 => x"f8",
          7462 => x"f8",
          7463 => x"c8",
          7464 => x"70",
          7465 => x"59",
          7466 => x"26",
          7467 => x"78",
          7468 => x"f2",
          7469 => x"78",
          7470 => x"3d",
          7471 => x"53",
          7472 => x"51",
          7473 => x"3f",
          7474 => x"08",
          7475 => x"88",
          7476 => x"fc",
          7477 => x"9a",
          7478 => x"fe",
          7479 => x"fe",
          7480 => x"fe",
          7481 => x"82",
          7482 => x"80",
          7483 => x"81",
          7484 => x"38",
          7485 => x"bf",
          7486 => x"02",
          7487 => x"33",
          7488 => x"ef",
          7489 => x"c8",
          7490 => x"06",
          7491 => x"38",
          7492 => x"51",
          7493 => x"3f",
          7494 => x"d6",
          7495 => x"f4",
          7496 => x"80",
          7497 => x"39",
          7498 => x"f4",
          7499 => x"f8",
          7500 => x"fd",
          7501 => x"93",
          7502 => x"2e",
          7503 => x"80",
          7504 => x"02",
          7505 => x"33",
          7506 => x"e6",
          7507 => x"c8",
          7508 => x"89",
          7509 => x"fb",
          7510 => x"96",
          7511 => x"fe",
          7512 => x"fe",
          7513 => x"fe",
          7514 => x"82",
          7515 => x"80",
          7516 => x"60",
          7517 => x"fa",
          7518 => x"fe",
          7519 => x"fe",
          7520 => x"fe",
          7521 => x"82",
          7522 => x"86",
          7523 => x"c8",
          7524 => x"53",
          7525 => x"52",
          7526 => x"52",
          7527 => x"94",
          7528 => x"05",
          7529 => x"52",
          7530 => x"29",
          7531 => x"05",
          7532 => x"d0",
          7533 => x"c8",
          7534 => x"8c",
          7535 => x"c8",
          7536 => x"9a",
          7537 => x"39",
          7538 => x"51",
          7539 => x"3f",
          7540 => x"9e",
          7541 => x"fe",
          7542 => x"fe",
          7543 => x"82",
          7544 => x"b5",
          7545 => x"05",
          7546 => x"e4",
          7547 => x"53",
          7548 => x"08",
          7549 => x"f6",
          7550 => x"93",
          7551 => x"2e",
          7552 => x"82",
          7553 => x"51",
          7554 => x"fc",
          7555 => x"3d",
          7556 => x"51",
          7557 => x"3f",
          7558 => x"08",
          7559 => x"f8",
          7560 => x"fe",
          7561 => x"82",
          7562 => x"b5",
          7563 => x"05",
          7564 => x"e4",
          7565 => x"93",
          7566 => x"3d",
          7567 => x"52",
          7568 => x"a3",
          7569 => x"c4",
          7570 => x"fc",
          7571 => x"80",
          7572 => x"c8",
          7573 => x"06",
          7574 => x"79",
          7575 => x"f6",
          7576 => x"93",
          7577 => x"2e",
          7578 => x"82",
          7579 => x"51",
          7580 => x"fb",
          7581 => x"89",
          7582 => x"f3",
          7583 => x"51",
          7584 => x"3f",
          7585 => x"82",
          7586 => x"fe",
          7587 => x"a2",
          7588 => x"e2",
          7589 => x"39",
          7590 => x"0b",
          7591 => x"84",
          7592 => x"81",
          7593 => x"94",
          7594 => x"89",
          7595 => x"f2",
          7596 => x"be",
          7597 => x"dc",
          7598 => x"e8",
          7599 => x"83",
          7600 => x"94",
          7601 => x"80",
          7602 => x"c0",
          7603 => x"fb",
          7604 => x"3d",
          7605 => x"53",
          7606 => x"51",
          7607 => x"3f",
          7608 => x"08",
          7609 => x"8a",
          7610 => x"82",
          7611 => x"fe",
          7612 => x"60",
          7613 => x"b4",
          7614 => x"11",
          7615 => x"05",
          7616 => x"a5",
          7617 => x"c8",
          7618 => x"fa",
          7619 => x"52",
          7620 => x"51",
          7621 => x"3f",
          7622 => x"2d",
          7623 => x"08",
          7624 => x"c8",
          7625 => x"fa",
          7626 => x"93",
          7627 => x"82",
          7628 => x"fe",
          7629 => x"fa",
          7630 => x"8a",
          7631 => x"f1",
          7632 => x"d1",
          7633 => x"aa",
          7634 => x"e0",
          7635 => x"d4",
          7636 => x"ff",
          7637 => x"ed",
          7638 => x"96",
          7639 => x"33",
          7640 => x"80",
          7641 => x"38",
          7642 => x"59",
          7643 => x"80",
          7644 => x"3d",
          7645 => x"51",
          7646 => x"3f",
          7647 => x"56",
          7648 => x"08",
          7649 => x"f8",
          7650 => x"82",
          7651 => x"a0",
          7652 => x"59",
          7653 => x"3f",
          7654 => x"58",
          7655 => x"57",
          7656 => x"81",
          7657 => x"55",
          7658 => x"80",
          7659 => x"80",
          7660 => x"51",
          7661 => x"82",
          7662 => x"5e",
          7663 => x"7c",
          7664 => x"59",
          7665 => x"7d",
          7666 => x"81",
          7667 => x"38",
          7668 => x"51",
          7669 => x"3f",
          7670 => x"80",
          7671 => x"0b",
          7672 => x"34",
          7673 => x"e4",
          7674 => x"94",
          7675 => x"90",
          7676 => x"87",
          7677 => x"0c",
          7678 => x"0b",
          7679 => x"84",
          7680 => x"83",
          7681 => x"94",
          7682 => x"d4",
          7683 => x"93",
          7684 => x"d7",
          7685 => x"93",
          7686 => x"e8",
          7687 => x"ee",
          7688 => x"8b",
          7689 => x"e5",
          7690 => x"8b",
          7691 => x"ef",
          7692 => x"e4",
          7693 => x"ee",
          7694 => x"51",
          7695 => x"f7",
          7696 => x"04",
          7697 => x"2f",
          7698 => x"2f",
          7699 => x"2f",
          7700 => x"2f",
          7701 => x"2f",
          7702 => x"2f",
          7703 => x"31",
          7704 => x"31",
          7705 => x"31",
          7706 => x"31",
          7707 => x"31",
          7708 => x"31",
          7709 => x"31",
          7710 => x"31",
          7711 => x"31",
          7712 => x"31",
          7713 => x"31",
          7714 => x"31",
          7715 => x"31",
          7716 => x"31",
          7717 => x"31",
          7718 => x"31",
          7719 => x"31",
          7720 => x"31",
          7721 => x"31",
          7722 => x"31",
          7723 => x"31",
          7724 => x"31",
          7725 => x"31",
          7726 => x"70",
          7727 => x"6f",
          7728 => x"6f",
          7729 => x"70",
          7730 => x"70",
          7731 => x"70",
          7732 => x"70",
          7733 => x"70",
          7734 => x"70",
          7735 => x"70",
          7736 => x"70",
          7737 => x"70",
          7738 => x"70",
          7739 => x"70",
          7740 => x"70",
          7741 => x"70",
          7742 => x"70",
          7743 => x"70",
          7744 => x"70",
          7745 => x"70",
          7746 => x"74",
          7747 => x"77",
          7748 => x"74",
          7749 => x"77",
          7750 => x"75",
          7751 => x"77",
          7752 => x"77",
          7753 => x"77",
          7754 => x"77",
          7755 => x"77",
          7756 => x"77",
          7757 => x"77",
          7758 => x"77",
          7759 => x"77",
          7760 => x"77",
          7761 => x"77",
          7762 => x"77",
          7763 => x"77",
          7764 => x"77",
          7765 => x"77",
          7766 => x"75",
          7767 => x"77",
          7768 => x"77",
          7769 => x"77",
          7770 => x"77",
          7771 => x"77",
          7772 => x"77",
          7773 => x"77",
          7774 => x"77",
          7775 => x"77",
          7776 => x"77",
          7777 => x"77",
          7778 => x"77",
          7779 => x"77",
          7780 => x"77",
          7781 => x"77",
          7782 => x"77",
          7783 => x"77",
          7784 => x"77",
          7785 => x"77",
          7786 => x"77",
          7787 => x"77",
          7788 => x"77",
          7789 => x"75",
          7790 => x"77",
          7791 => x"77",
          7792 => x"77",
          7793 => x"77",
          7794 => x"76",
          7795 => x"77",
          7796 => x"77",
          7797 => x"77",
          7798 => x"77",
          7799 => x"77",
          7800 => x"77",
          7801 => x"77",
          7802 => x"77",
          7803 => x"77",
          7804 => x"77",
          7805 => x"77",
          7806 => x"77",
          7807 => x"77",
          7808 => x"77",
          7809 => x"77",
          7810 => x"77",
          7811 => x"77",
          7812 => x"77",
          7813 => x"77",
          7814 => x"77",
          7815 => x"77",
          7816 => x"77",
          7817 => x"77",
          7818 => x"77",
          7819 => x"77",
          7820 => x"77",
          7821 => x"77",
          7822 => x"77",
          7823 => x"77",
          7824 => x"77",
          7825 => x"77",
          7826 => x"76",
          7827 => x"76",
          7828 => x"77",
          7829 => x"77",
          7830 => x"76",
          7831 => x"76",
          7832 => x"77",
          7833 => x"77",
          7834 => x"77",
          7835 => x"77",
          7836 => x"77",
          7837 => x"77",
          7838 => x"77",
          7839 => x"77",
          7840 => x"77",
          7841 => x"77",
          7842 => x"77",
          7843 => x"77",
          7844 => x"77",
          7845 => x"77",
          7846 => x"77",
          7847 => x"77",
          7848 => x"77",
          7849 => x"77",
          7850 => x"77",
          7851 => x"77",
          7852 => x"77",
          7853 => x"77",
          7854 => x"77",
          7855 => x"77",
          7856 => x"77",
          7857 => x"77",
          7858 => x"77",
          7859 => x"77",
          7860 => x"77",
          7861 => x"77",
          7862 => x"77",
          7863 => x"77",
          7864 => x"77",
          7865 => x"77",
          7866 => x"76",
          7867 => x"76",
          7868 => x"77",
          7869 => x"77",
          7870 => x"77",
          7871 => x"77",
          7872 => x"77",
          7873 => x"77",
          7874 => x"77",
          7875 => x"77",
          7876 => x"77",
          7877 => x"77",
          7878 => x"77",
          7879 => x"77",
          7880 => x"77",
          7881 => x"74",
          7882 => x"2f",
          7883 => x"25",
          7884 => x"64",
          7885 => x"3a",
          7886 => x"25",
          7887 => x"0a",
          7888 => x"43",
          7889 => x"6e",
          7890 => x"75",
          7891 => x"69",
          7892 => x"00",
          7893 => x"66",
          7894 => x"20",
          7895 => x"20",
          7896 => x"66",
          7897 => x"00",
          7898 => x"44",
          7899 => x"63",
          7900 => x"69",
          7901 => x"65",
          7902 => x"74",
          7903 => x"0a",
          7904 => x"20",
          7905 => x"53",
          7906 => x"52",
          7907 => x"28",
          7908 => x"72",
          7909 => x"30",
          7910 => x"20",
          7911 => x"65",
          7912 => x"38",
          7913 => x"0a",
          7914 => x"20",
          7915 => x"41",
          7916 => x"53",
          7917 => x"74",
          7918 => x"38",
          7919 => x"53",
          7920 => x"3d",
          7921 => x"58",
          7922 => x"00",
          7923 => x"20",
          7924 => x"4d",
          7925 => x"74",
          7926 => x"3d",
          7927 => x"58",
          7928 => x"69",
          7929 => x"25",
          7930 => x"29",
          7931 => x"00",
          7932 => x"20",
          7933 => x"43",
          7934 => x"00",
          7935 => x"20",
          7936 => x"32",
          7937 => x"00",
          7938 => x"20",
          7939 => x"49",
          7940 => x"00",
          7941 => x"20",
          7942 => x"20",
          7943 => x"64",
          7944 => x"65",
          7945 => x"65",
          7946 => x"30",
          7947 => x"2e",
          7948 => x"00",
          7949 => x"20",
          7950 => x"54",
          7951 => x"55",
          7952 => x"43",
          7953 => x"52",
          7954 => x"45",
          7955 => x"00",
          7956 => x"20",
          7957 => x"4d",
          7958 => x"20",
          7959 => x"6d",
          7960 => x"3d",
          7961 => x"58",
          7962 => x"00",
          7963 => x"64",
          7964 => x"73",
          7965 => x"0a",
          7966 => x"20",
          7967 => x"55",
          7968 => x"73",
          7969 => x"56",
          7970 => x"6f",
          7971 => x"64",
          7972 => x"73",
          7973 => x"20",
          7974 => x"58",
          7975 => x"00",
          7976 => x"20",
          7977 => x"55",
          7978 => x"6d",
          7979 => x"20",
          7980 => x"72",
          7981 => x"64",
          7982 => x"73",
          7983 => x"20",
          7984 => x"58",
          7985 => x"00",
          7986 => x"20",
          7987 => x"61",
          7988 => x"53",
          7989 => x"74",
          7990 => x"64",
          7991 => x"73",
          7992 => x"20",
          7993 => x"20",
          7994 => x"58",
          7995 => x"00",
          7996 => x"20",
          7997 => x"55",
          7998 => x"20",
          7999 => x"20",
          8000 => x"20",
          8001 => x"20",
          8002 => x"20",
          8003 => x"20",
          8004 => x"58",
          8005 => x"00",
          8006 => x"20",
          8007 => x"73",
          8008 => x"20",
          8009 => x"63",
          8010 => x"72",
          8011 => x"20",
          8012 => x"20",
          8013 => x"20",
          8014 => x"58",
          8015 => x"00",
          8016 => x"61",
          8017 => x"00",
          8018 => x"64",
          8019 => x"00",
          8020 => x"65",
          8021 => x"00",
          8022 => x"4f",
          8023 => x"4f",
          8024 => x"00",
          8025 => x"6b",
          8026 => x"6e",
          8027 => x"00",
          8028 => x"2b",
          8029 => x"3c",
          8030 => x"5b",
          8031 => x"00",
          8032 => x"54",
          8033 => x"54",
          8034 => x"00",
          8035 => x"00",
          8036 => x"00",
          8037 => x"00",
          8038 => x"00",
          8039 => x"00",
          8040 => x"00",
          8041 => x"00",
          8042 => x"00",
          8043 => x"00",
          8044 => x"0a",
          8045 => x"90",
          8046 => x"4f",
          8047 => x"30",
          8048 => x"20",
          8049 => x"45",
          8050 => x"20",
          8051 => x"33",
          8052 => x"20",
          8053 => x"20",
          8054 => x"45",
          8055 => x"20",
          8056 => x"20",
          8057 => x"20",
          8058 => x"7d",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"45",
          8063 => x"8f",
          8064 => x"45",
          8065 => x"8e",
          8066 => x"92",
          8067 => x"55",
          8068 => x"9a",
          8069 => x"9e",
          8070 => x"4f",
          8071 => x"a6",
          8072 => x"aa",
          8073 => x"ae",
          8074 => x"b2",
          8075 => x"b6",
          8076 => x"ba",
          8077 => x"be",
          8078 => x"c2",
          8079 => x"c6",
          8080 => x"ca",
          8081 => x"ce",
          8082 => x"d2",
          8083 => x"d6",
          8084 => x"da",
          8085 => x"de",
          8086 => x"e2",
          8087 => x"e6",
          8088 => x"ea",
          8089 => x"ee",
          8090 => x"f2",
          8091 => x"f6",
          8092 => x"fa",
          8093 => x"fe",
          8094 => x"2c",
          8095 => x"5d",
          8096 => x"2a",
          8097 => x"3f",
          8098 => x"00",
          8099 => x"00",
          8100 => x"00",
          8101 => x"02",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"54",
          8108 => x"00",
          8109 => x"54",
          8110 => x"00",
          8111 => x"46",
          8112 => x"00",
          8113 => x"53",
          8114 => x"4f",
          8115 => x"4e",
          8116 => x"4c",
          8117 => x"00",
          8118 => x"53",
          8119 => x"55",
          8120 => x"52",
          8121 => x"4e",
          8122 => x"4c",
          8123 => x"00",
          8124 => x"4c",
          8125 => x"53",
          8126 => x"20",
          8127 => x"54",
          8128 => x"53",
          8129 => x"4d",
          8130 => x"00",
          8131 => x"52",
          8132 => x"52",
          8133 => x"00",
          8134 => x"53",
          8135 => x"47",
          8136 => x"45",
          8137 => x"49",
          8138 => x"00",
          8139 => x"53",
          8140 => x"4f",
          8141 => x"4e",
          8142 => x"00",
          8143 => x"75",
          8144 => x"00",
          8145 => x"6e",
          8146 => x"00",
          8147 => x"74",
          8148 => x"00",
          8149 => x"6f",
          8150 => x"00",
          8151 => x"75",
          8152 => x"00",
          8153 => x"64",
          8154 => x"00",
          8155 => x"65",
          8156 => x"00",
          8157 => x"72",
          8158 => x"00",
          8159 => x"69",
          8160 => x"00",
          8161 => x"65",
          8162 => x"00",
          8163 => x"6e",
          8164 => x"00",
          8165 => x"70",
          8166 => x"00",
          8167 => x"6c",
          8168 => x"00",
          8169 => x"65",
          8170 => x"00",
          8171 => x"65",
          8172 => x"00",
          8173 => x"6e",
          8174 => x"63",
          8175 => x"00",
          8176 => x"72",
          8177 => x"00",
          8178 => x"72",
          8179 => x"00",
          8180 => x"6c",
          8181 => x"00",
          8182 => x"74",
          8183 => x"00",
          8184 => x"69",
          8185 => x"00",
          8186 => x"65",
          8187 => x"65",
          8188 => x"65",
          8189 => x"00",
          8190 => x"6b",
          8191 => x"00",
          8192 => x"74",
          8193 => x"00",
          8194 => x"69",
          8195 => x"00",
          8196 => x"61",
          8197 => x"00",
          8198 => x"70",
          8199 => x"6f",
          8200 => x"74",
          8201 => x"74",
          8202 => x"74",
          8203 => x"6f",
          8204 => x"00",
          8205 => x"78",
          8206 => x"00",
          8207 => x"61",
          8208 => x"00",
          8209 => x"75",
          8210 => x"00",
          8211 => x"64",
          8212 => x"72",
          8213 => x"00",
          8214 => x"68",
          8215 => x"69",
          8216 => x"00",
          8217 => x"61",
          8218 => x"00",
          8219 => x"6b",
          8220 => x"00",
          8221 => x"6c",
          8222 => x"00",
          8223 => x"75",
          8224 => x"00",
          8225 => x"62",
          8226 => x"68",
          8227 => x"77",
          8228 => x"64",
          8229 => x"65",
          8230 => x"00",
          8231 => x"00",
          8232 => x"64",
          8233 => x"65",
          8234 => x"72",
          8235 => x"00",
          8236 => x"72",
          8237 => x"72",
          8238 => x"00",
          8239 => x"6c",
          8240 => x"00",
          8241 => x"70",
          8242 => x"73",
          8243 => x"74",
          8244 => x"73",
          8245 => x"00",
          8246 => x"6c",
          8247 => x"00",
          8248 => x"66",
          8249 => x"00",
          8250 => x"6d",
          8251 => x"00",
          8252 => x"73",
          8253 => x"00",
          8254 => x"73",
          8255 => x"72",
          8256 => x"0a",
          8257 => x"74",
          8258 => x"61",
          8259 => x"72",
          8260 => x"2e",
          8261 => x"00",
          8262 => x"73",
          8263 => x"6f",
          8264 => x"65",
          8265 => x"2e",
          8266 => x"00",
          8267 => x"20",
          8268 => x"65",
          8269 => x"75",
          8270 => x"0a",
          8271 => x"20",
          8272 => x"68",
          8273 => x"75",
          8274 => x"0a",
          8275 => x"76",
          8276 => x"64",
          8277 => x"6c",
          8278 => x"6d",
          8279 => x"00",
          8280 => x"63",
          8281 => x"20",
          8282 => x"69",
          8283 => x"0a",
          8284 => x"6c",
          8285 => x"6c",
          8286 => x"64",
          8287 => x"78",
          8288 => x"73",
          8289 => x"00",
          8290 => x"6c",
          8291 => x"61",
          8292 => x"65",
          8293 => x"76",
          8294 => x"64",
          8295 => x"00",
          8296 => x"20",
          8297 => x"77",
          8298 => x"65",
          8299 => x"6f",
          8300 => x"74",
          8301 => x"0a",
          8302 => x"69",
          8303 => x"6e",
          8304 => x"65",
          8305 => x"73",
          8306 => x"76",
          8307 => x"64",
          8308 => x"00",
          8309 => x"73",
          8310 => x"6f",
          8311 => x"6e",
          8312 => x"65",
          8313 => x"00",
          8314 => x"20",
          8315 => x"70",
          8316 => x"62",
          8317 => x"66",
          8318 => x"73",
          8319 => x"65",
          8320 => x"6f",
          8321 => x"20",
          8322 => x"64",
          8323 => x"2e",
          8324 => x"00",
          8325 => x"72",
          8326 => x"20",
          8327 => x"72",
          8328 => x"2e",
          8329 => x"00",
          8330 => x"6d",
          8331 => x"74",
          8332 => x"70",
          8333 => x"74",
          8334 => x"20",
          8335 => x"63",
          8336 => x"65",
          8337 => x"00",
          8338 => x"6c",
          8339 => x"73",
          8340 => x"63",
          8341 => x"2e",
          8342 => x"00",
          8343 => x"73",
          8344 => x"69",
          8345 => x"6e",
          8346 => x"65",
          8347 => x"79",
          8348 => x"00",
          8349 => x"6f",
          8350 => x"6e",
          8351 => x"70",
          8352 => x"66",
          8353 => x"73",
          8354 => x"00",
          8355 => x"72",
          8356 => x"74",
          8357 => x"20",
          8358 => x"6f",
          8359 => x"63",
          8360 => x"00",
          8361 => x"63",
          8362 => x"73",
          8363 => x"00",
          8364 => x"6b",
          8365 => x"6e",
          8366 => x"72",
          8367 => x"0a",
          8368 => x"6c",
          8369 => x"79",
          8370 => x"20",
          8371 => x"61",
          8372 => x"6c",
          8373 => x"79",
          8374 => x"2f",
          8375 => x"2e",
          8376 => x"00",
          8377 => x"61",
          8378 => x"00",
          8379 => x"55",
          8380 => x"00",
          8381 => x"2a",
          8382 => x"20",
          8383 => x"00",
          8384 => x"2f",
          8385 => x"32",
          8386 => x"00",
          8387 => x"2e",
          8388 => x"00",
          8389 => x"50",
          8390 => x"72",
          8391 => x"25",
          8392 => x"29",
          8393 => x"20",
          8394 => x"2a",
          8395 => x"00",
          8396 => x"55",
          8397 => x"49",
          8398 => x"72",
          8399 => x"74",
          8400 => x"6e",
          8401 => x"72",
          8402 => x"00",
          8403 => x"6d",
          8404 => x"69",
          8405 => x"72",
          8406 => x"74",
          8407 => x"00",
          8408 => x"32",
          8409 => x"74",
          8410 => x"75",
          8411 => x"00",
          8412 => x"43",
          8413 => x"52",
          8414 => x"6e",
          8415 => x"72",
          8416 => x"0a",
          8417 => x"43",
          8418 => x"57",
          8419 => x"6e",
          8420 => x"72",
          8421 => x"0a",
          8422 => x"52",
          8423 => x"52",
          8424 => x"6e",
          8425 => x"72",
          8426 => x"0a",
          8427 => x"52",
          8428 => x"54",
          8429 => x"6e",
          8430 => x"72",
          8431 => x"0a",
          8432 => x"52",
          8433 => x"52",
          8434 => x"6e",
          8435 => x"72",
          8436 => x"0a",
          8437 => x"52",
          8438 => x"54",
          8439 => x"6e",
          8440 => x"72",
          8441 => x"0a",
          8442 => x"74",
          8443 => x"67",
          8444 => x"20",
          8445 => x"65",
          8446 => x"2e",
          8447 => x"00",
          8448 => x"61",
          8449 => x"6e",
          8450 => x"69",
          8451 => x"2e",
          8452 => x"00",
          8453 => x"00",
          8454 => x"69",
          8455 => x"20",
          8456 => x"69",
          8457 => x"69",
          8458 => x"73",
          8459 => x"64",
          8460 => x"72",
          8461 => x"2c",
          8462 => x"65",
          8463 => x"20",
          8464 => x"74",
          8465 => x"6e",
          8466 => x"6c",
          8467 => x"00",
          8468 => x"00",
          8469 => x"64",
          8470 => x"73",
          8471 => x"64",
          8472 => x"00",
          8473 => x"69",
          8474 => x"6c",
          8475 => x"64",
          8476 => x"00",
          8477 => x"69",
          8478 => x"20",
          8479 => x"69",
          8480 => x"69",
          8481 => x"73",
          8482 => x"00",
          8483 => x"3d",
          8484 => x"00",
          8485 => x"3a",
          8486 => x"73",
          8487 => x"69",
          8488 => x"69",
          8489 => x"72",
          8490 => x"74",
          8491 => x"00",
          8492 => x"61",
          8493 => x"6e",
          8494 => x"6e",
          8495 => x"72",
          8496 => x"73",
          8497 => x"00",
          8498 => x"73",
          8499 => x"65",
          8500 => x"61",
          8501 => x"66",
          8502 => x"0a",
          8503 => x"61",
          8504 => x"6e",
          8505 => x"61",
          8506 => x"66",
          8507 => x"0a",
          8508 => x"65",
          8509 => x"69",
          8510 => x"63",
          8511 => x"20",
          8512 => x"30",
          8513 => x"2e",
          8514 => x"00",
          8515 => x"6c",
          8516 => x"67",
          8517 => x"64",
          8518 => x"20",
          8519 => x"78",
          8520 => x"2e",
          8521 => x"00",
          8522 => x"6c",
          8523 => x"65",
          8524 => x"6e",
          8525 => x"63",
          8526 => x"20",
          8527 => x"29",
          8528 => x"00",
          8529 => x"73",
          8530 => x"74",
          8531 => x"20",
          8532 => x"6c",
          8533 => x"74",
          8534 => x"2e",
          8535 => x"00",
          8536 => x"6c",
          8537 => x"65",
          8538 => x"74",
          8539 => x"2e",
          8540 => x"00",
          8541 => x"55",
          8542 => x"6e",
          8543 => x"3a",
          8544 => x"5c",
          8545 => x"25",
          8546 => x"00",
          8547 => x"64",
          8548 => x"6d",
          8549 => x"64",
          8550 => x"00",
          8551 => x"6e",
          8552 => x"67",
          8553 => x"0a",
          8554 => x"61",
          8555 => x"6e",
          8556 => x"6e",
          8557 => x"72",
          8558 => x"73",
          8559 => x"0a",
          8560 => x"00",
          8561 => x"00",
          8562 => x"7f",
          8563 => x"00",
          8564 => x"7f",
          8565 => x"00",
          8566 => x"7f",
          8567 => x"00",
          8568 => x"00",
          8569 => x"78",
          8570 => x"00",
          8571 => x"e1",
          8572 => x"01",
          8573 => x"01",
          8574 => x"01",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"7f",
          8579 => x"01",
          8580 => x"00",
          8581 => x"00",
          8582 => x"7f",
          8583 => x"01",
          8584 => x"00",
          8585 => x"00",
          8586 => x"7f",
          8587 => x"01",
          8588 => x"00",
          8589 => x"00",
          8590 => x"7f",
          8591 => x"01",
          8592 => x"00",
          8593 => x"00",
          8594 => x"7f",
          8595 => x"02",
          8596 => x"00",
          8597 => x"00",
          8598 => x"7f",
          8599 => x"02",
          8600 => x"00",
          8601 => x"00",
          8602 => x"7f",
          8603 => x"02",
          8604 => x"00",
          8605 => x"00",
          8606 => x"7f",
          8607 => x"02",
          8608 => x"00",
          8609 => x"00",
          8610 => x"7f",
          8611 => x"02",
          8612 => x"00",
          8613 => x"00",
          8614 => x"7f",
          8615 => x"02",
          8616 => x"00",
          8617 => x"00",
          8618 => x"7f",
          8619 => x"03",
          8620 => x"00",
          8621 => x"00",
          8622 => x"7f",
          8623 => x"03",
          8624 => x"00",
          8625 => x"00",
          8626 => x"7f",
          8627 => x"03",
          8628 => x"00",
          8629 => x"00",
          8630 => x"7f",
          8631 => x"03",
          8632 => x"00",
          8633 => x"00",
          8634 => x"7f",
          8635 => x"03",
          8636 => x"00",
          8637 => x"00",
          8638 => x"7f",
          8639 => x"03",
          8640 => x"00",
          8641 => x"00",
          8642 => x"7f",
          8643 => x"03",
          8644 => x"00",
          8645 => x"00",
          8646 => x"7f",
          8647 => x"03",
          8648 => x"00",
          8649 => x"00",
          8650 => x"7f",
          8651 => x"03",
          8652 => x"00",
          8653 => x"00",
          8654 => x"7f",
          8655 => x"03",
          8656 => x"00",
          8657 => x"00",
          8658 => x"7f",
          8659 => x"03",
          8660 => x"00",
          8661 => x"00",
          8662 => x"7f",
          8663 => x"03",
          8664 => x"00",
          8665 => x"00",
          8666 => x"7f",
          8667 => x"03",
          8668 => x"00",
          8669 => x"00",
          8670 => x"7f",
          8671 => x"03",
          8672 => x"00",
          8673 => x"00",
          8674 => x"80",
          8675 => x"03",
          8676 => x"00",
          8677 => x"00",
          8678 => x"80",
          8679 => x"03",
          8680 => x"00",
          8681 => x"00",
          8682 => x"80",
          8683 => x"03",
          8684 => x"00",
          8685 => x"00",
          8686 => x"80",
          8687 => x"03",
          8688 => x"00",
          8689 => x"00",
          8690 => x"80",
          8691 => x"03",
          8692 => x"00",
          8693 => x"00",
          8694 => x"80",
          8695 => x"03",
          8696 => x"00",
          8697 => x"00",
          8698 => x"80",
          8699 => x"03",
          8700 => x"00",
          8701 => x"00",
          8702 => x"80",
          8703 => x"03",
          8704 => x"00",
          8705 => x"00",
          8706 => x"80",
          8707 => x"03",
          8708 => x"00",
          8709 => x"00",
          8710 => x"80",
          8711 => x"03",
          8712 => x"00",
          8713 => x"00",
          8714 => x"80",
          8715 => x"03",
          8716 => x"00",
          8717 => x"00",
          8718 => x"80",
          8719 => x"03",
          8720 => x"00",
          8721 => x"00",
          8722 => x"80",
          8723 => x"03",
          8724 => x"00",
          8725 => x"00",
          8726 => x"80",
          8727 => x"03",
          8728 => x"00",
          8729 => x"00",
          8730 => x"80",
          8731 => x"03",
          8732 => x"00",
          8733 => x"00",
          8734 => x"80",
          8735 => x"04",
          8736 => x"00",
          8737 => x"00",
          8738 => x"80",
          8739 => x"04",
          8740 => x"00",
          8741 => x"00",
          8742 => x"80",
          8743 => x"04",
          8744 => x"00",
          8745 => x"00",
          8746 => x"80",
          8747 => x"04",
          8748 => x"00",
          8749 => x"00",
          8750 => x"80",
          8751 => x"04",
          8752 => x"00",
          8753 => x"00",
          8754 => x"80",
          8755 => x"05",
          8756 => x"00",
          8757 => x"00",
          8758 => x"80",
          8759 => x"05",
          8760 => x"00",
          8761 => x"00",
          8762 => x"80",
          8763 => x"05",
          8764 => x"00",
          8765 => x"00",
          8766 => x"80",
          8767 => x"05",
          8768 => x"00",
          8769 => x"00",
          8770 => x"80",
          8771 => x"05",
          8772 => x"00",
          8773 => x"00",
          8774 => x"80",
          8775 => x"05",
          8776 => x"00",
          8777 => x"00",
          8778 => x"80",
          8779 => x"06",
          8780 => x"00",
          8781 => x"00",
          8782 => x"80",
          8783 => x"06",
          8784 => x"00",
          8785 => x"00",
          8786 => x"80",
          8787 => x"07",
          8788 => x"00",
          8789 => x"00",
          8790 => x"80",
          8791 => x"07",
          8792 => x"00",
          8793 => x"00",
          8794 => x"80",
          8795 => x"08",
          8796 => x"00",
          8797 => x"00",
          8798 => x"80",
          8799 => x"08",
          8800 => x"00",
          8801 => x"00",
          8802 => x"80",
          8803 => x"08",
          8804 => x"00",
          8805 => x"00",
          8806 => x"80",
          8807 => x"08",
          8808 => x"00",
          8809 => x"00",
          8810 => x"80",
          8811 => x"08",
          8812 => x"00",
          8813 => x"00",
          8814 => x"80",
          8815 => x"08",
          8816 => x"00",
          8817 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"04",
           281 => x"04",
           282 => x"9f",
           283 => x"dc",
           284 => x"80",
           285 => x"05",
           286 => x"eb",
           287 => x"51",
           288 => x"94",
           289 => x"0c",
           290 => x"80",
           291 => x"8c",
           292 => x"94",
           293 => x"08",
           294 => x"3f",
           295 => x"88",
           296 => x"3d",
           297 => x"04",
           298 => x"94",
           299 => x"0d",
           300 => x"08",
           301 => x"52",
           302 => x"05",
           303 => x"b9",
           304 => x"70",
           305 => x"85",
           306 => x"0c",
           307 => x"02",
           308 => x"3d",
           309 => x"94",
           310 => x"0c",
           311 => x"05",
           312 => x"ab",
           313 => x"88",
           314 => x"94",
           315 => x"0c",
           316 => x"08",
           317 => x"94",
           318 => x"08",
           319 => x"0b",
           320 => x"05",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"08",
           325 => x"38",
           326 => x"05",
           327 => x"08",
           328 => x"80",
           329 => x"f0",
           330 => x"08",
           331 => x"88",
           332 => x"94",
           333 => x"0c",
           334 => x"05",
           335 => x"fc",
           336 => x"53",
           337 => x"05",
           338 => x"08",
           339 => x"51",
           340 => x"88",
           341 => x"08",
           342 => x"54",
           343 => x"05",
           344 => x"8c",
           345 => x"f8",
           346 => x"94",
           347 => x"0c",
           348 => x"05",
           349 => x"0c",
           350 => x"0d",
           351 => x"94",
           352 => x"0c",
           353 => x"80",
           354 => x"fc",
           355 => x"08",
           356 => x"80",
           357 => x"94",
           358 => x"08",
           359 => x"88",
           360 => x"0b",
           361 => x"05",
           362 => x"8c",
           363 => x"25",
           364 => x"08",
           365 => x"30",
           366 => x"05",
           367 => x"94",
           368 => x"08",
           369 => x"88",
           370 => x"ad",
           371 => x"70",
           372 => x"05",
           373 => x"08",
           374 => x"80",
           375 => x"94",
           376 => x"08",
           377 => x"f8",
           378 => x"08",
           379 => x"70",
           380 => x"87",
           381 => x"0c",
           382 => x"02",
           383 => x"3d",
           384 => x"94",
           385 => x"0c",
           386 => x"08",
           387 => x"94",
           388 => x"08",
           389 => x"05",
           390 => x"38",
           391 => x"05",
           392 => x"a3",
           393 => x"94",
           394 => x"08",
           395 => x"94",
           396 => x"08",
           397 => x"8c",
           398 => x"08",
           399 => x"10",
           400 => x"05",
           401 => x"94",
           402 => x"08",
           403 => x"c9",
           404 => x"8c",
           405 => x"08",
           406 => x"26",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"88",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"f8",
           415 => x"08",
           416 => x"81",
           417 => x"fc",
           418 => x"08",
           419 => x"81",
           420 => x"8c",
           421 => x"af",
           422 => x"90",
           423 => x"2e",
           424 => x"08",
           425 => x"70",
           426 => x"05",
           427 => x"39",
           428 => x"05",
           429 => x"08",
           430 => x"51",
           431 => x"05",
           432 => x"85",
           433 => x"0c",
           434 => x"0d",
           435 => x"87",
           436 => x"0c",
           437 => x"c0",
           438 => x"85",
           439 => x"98",
           440 => x"c0",
           441 => x"70",
           442 => x"51",
           443 => x"8a",
           444 => x"98",
           445 => x"70",
           446 => x"c0",
           447 => x"fc",
           448 => x"52",
           449 => x"87",
           450 => x"08",
           451 => x"2e",
           452 => x"0b",
           453 => x"a8",
           454 => x"0b",
           455 => x"88",
           456 => x"0d",
           457 => x"0d",
           458 => x"56",
           459 => x"0b",
           460 => x"9f",
           461 => x"06",
           462 => x"52",
           463 => x"09",
           464 => x"9e",
           465 => x"87",
           466 => x"0c",
           467 => x"92",
           468 => x"0b",
           469 => x"8c",
           470 => x"92",
           471 => x"85",
           472 => x"06",
           473 => x"70",
           474 => x"38",
           475 => x"84",
           476 => x"ff",
           477 => x"27",
           478 => x"73",
           479 => x"38",
           480 => x"8b",
           481 => x"70",
           482 => x"34",
           483 => x"81",
           484 => x"a2",
           485 => x"80",
           486 => x"87",
           487 => x"08",
           488 => x"b5",
           489 => x"98",
           490 => x"70",
           491 => x"0b",
           492 => x"8c",
           493 => x"92",
           494 => x"82",
           495 => x"70",
           496 => x"73",
           497 => x"06",
           498 => x"72",
           499 => x"06",
           500 => x"c0",
           501 => x"51",
           502 => x"09",
           503 => x"38",
           504 => x"88",
           505 => x"0d",
           506 => x"0d",
           507 => x"33",
           508 => x"88",
           509 => x"0c",
           510 => x"3d",
           511 => x"3d",
           512 => x"11",
           513 => x"33",
           514 => x"71",
           515 => x"81",
           516 => x"72",
           517 => x"75",
           518 => x"88",
           519 => x"54",
           520 => x"85",
           521 => x"f9",
           522 => x"0b",
           523 => x"ac",
           524 => x"81",
           525 => x"ed",
           526 => x"17",
           527 => x"e5",
           528 => x"55",
           529 => x"89",
           530 => x"2e",
           531 => x"d5",
           532 => x"76",
           533 => x"06",
           534 => x"2a",
           535 => x"05",
           536 => x"70",
           537 => x"bd",
           538 => x"b9",
           539 => x"fe",
           540 => x"08",
           541 => x"06",
           542 => x"84",
           543 => x"2b",
           544 => x"53",
           545 => x"8c",
           546 => x"52",
           547 => x"52",
           548 => x"3f",
           549 => x"38",
           550 => x"e2",
           551 => x"f0",
           552 => x"83",
           553 => x"74",
           554 => x"3d",
           555 => x"3d",
           556 => x"0b",
           557 => x"fe",
           558 => x"08",
           559 => x"56",
           560 => x"74",
           561 => x"38",
           562 => x"75",
           563 => x"16",
           564 => x"53",
           565 => x"87",
           566 => x"fd",
           567 => x"54",
           568 => x"0b",
           569 => x"08",
           570 => x"53",
           571 => x"2e",
           572 => x"8c",
           573 => x"51",
           574 => x"88",
           575 => x"53",
           576 => x"fd",
           577 => x"08",
           578 => x"06",
           579 => x"0c",
           580 => x"04",
           581 => x"76",
           582 => x"9f",
           583 => x"55",
           584 => x"88",
           585 => x"72",
           586 => x"38",
           587 => x"73",
           588 => x"81",
           589 => x"72",
           590 => x"33",
           591 => x"2e",
           592 => x"85",
           593 => x"08",
           594 => x"16",
           595 => x"2e",
           596 => x"51",
           597 => x"88",
           598 => x"39",
           599 => x"52",
           600 => x"0c",
           601 => x"88",
           602 => x"0d",
           603 => x"0d",
           604 => x"0b",
           605 => x"71",
           606 => x"70",
           607 => x"06",
           608 => x"55",
           609 => x"88",
           610 => x"08",
           611 => x"38",
           612 => x"dc",
           613 => x"06",
           614 => x"cf",
           615 => x"90",
           616 => x"15",
           617 => x"8f",
           618 => x"84",
           619 => x"52",
           620 => x"bc",
           621 => x"82",
           622 => x"05",
           623 => x"06",
           624 => x"38",
           625 => x"df",
           626 => x"71",
           627 => x"a0",
           628 => x"88",
           629 => x"08",
           630 => x"88",
           631 => x"0c",
           632 => x"fd",
           633 => x"08",
           634 => x"73",
           635 => x"52",
           636 => x"88",
           637 => x"f2",
           638 => x"62",
           639 => x"5c",
           640 => x"74",
           641 => x"81",
           642 => x"81",
           643 => x"56",
           644 => x"70",
           645 => x"74",
           646 => x"81",
           647 => x"81",
           648 => x"0b",
           649 => x"62",
           650 => x"55",
           651 => x"8f",
           652 => x"fd",
           653 => x"08",
           654 => x"34",
           655 => x"93",
           656 => x"08",
           657 => x"5f",
           658 => x"76",
           659 => x"58",
           660 => x"55",
           661 => x"09",
           662 => x"38",
           663 => x"5b",
           664 => x"5f",
           665 => x"1c",
           666 => x"06",
           667 => x"33",
           668 => x"70",
           669 => x"27",
           670 => x"07",
           671 => x"5b",
           672 => x"55",
           673 => x"38",
           674 => x"09",
           675 => x"38",
           676 => x"7a",
           677 => x"55",
           678 => x"9f",
           679 => x"32",
           680 => x"ae",
           681 => x"70",
           682 => x"2a",
           683 => x"51",
           684 => x"38",
           685 => x"5a",
           686 => x"77",
           687 => x"81",
           688 => x"1c",
           689 => x"55",
           690 => x"ff",
           691 => x"1e",
           692 => x"55",
           693 => x"83",
           694 => x"74",
           695 => x"7b",
           696 => x"3f",
           697 => x"ef",
           698 => x"7b",
           699 => x"2b",
           700 => x"54",
           701 => x"08",
           702 => x"f8",
           703 => x"08",
           704 => x"80",
           705 => x"33",
           706 => x"2e",
           707 => x"8b",
           708 => x"83",
           709 => x"06",
           710 => x"74",
           711 => x"7d",
           712 => x"88",
           713 => x"5b",
           714 => x"58",
           715 => x"9a",
           716 => x"81",
           717 => x"79",
           718 => x"5b",
           719 => x"31",
           720 => x"75",
           721 => x"38",
           722 => x"80",
           723 => x"7b",
           724 => x"3f",
           725 => x"88",
           726 => x"08",
           727 => x"39",
           728 => x"1c",
           729 => x"33",
           730 => x"a5",
           731 => x"33",
           732 => x"70",
           733 => x"56",
           734 => x"38",
           735 => x"39",
           736 => x"39",
           737 => x"d3",
           738 => x"88",
           739 => x"af",
           740 => x"0c",
           741 => x"04",
           742 => x"79",
           743 => x"82",
           744 => x"53",
           745 => x"51",
           746 => x"83",
           747 => x"80",
           748 => x"51",
           749 => x"88",
           750 => x"ff",
           751 => x"56",
           752 => x"d5",
           753 => x"06",
           754 => x"75",
           755 => x"77",
           756 => x"f6",
           757 => x"08",
           758 => x"94",
           759 => x"f8",
           760 => x"08",
           761 => x"06",
           762 => x"82",
           763 => x"38",
           764 => x"d2",
           765 => x"76",
           766 => x"3f",
           767 => x"88",
           768 => x"76",
           769 => x"3f",
           770 => x"ff",
           771 => x"74",
           772 => x"2e",
           773 => x"56",
           774 => x"89",
           775 => x"ed",
           776 => x"59",
           777 => x"0b",
           778 => x"0c",
           779 => x"88",
           780 => x"55",
           781 => x"82",
           782 => x"75",
           783 => x"70",
           784 => x"fe",
           785 => x"08",
           786 => x"57",
           787 => x"09",
           788 => x"38",
           789 => x"be",
           790 => x"75",
           791 => x"3f",
           792 => x"38",
           793 => x"55",
           794 => x"ac",
           795 => x"e4",
           796 => x"8a",
           797 => x"88",
           798 => x"52",
           799 => x"3f",
           800 => x"ff",
           801 => x"83",
           802 => x"06",
           803 => x"56",
           804 => x"76",
           805 => x"38",
           806 => x"8f",
           807 => x"8d",
           808 => x"75",
           809 => x"3f",
           810 => x"08",
           811 => x"95",
           812 => x"51",
           813 => x"88",
           814 => x"ff",
           815 => x"8c",
           816 => x"f3",
           817 => x"b6",
           818 => x"58",
           819 => x"33",
           820 => x"02",
           821 => x"05",
           822 => x"59",
           823 => x"3f",
           824 => x"ff",
           825 => x"05",
           826 => x"8c",
           827 => x"1a",
           828 => x"e0",
           829 => x"f1",
           830 => x"84",
           831 => x"3d",
           832 => x"f5",
           833 => x"08",
           834 => x"06",
           835 => x"38",
           836 => x"05",
           837 => x"3f",
           838 => x"7a",
           839 => x"3f",
           840 => x"ff",
           841 => x"71",
           842 => x"84",
           843 => x"84",
           844 => x"33",
           845 => x"31",
           846 => x"51",
           847 => x"3f",
           848 => x"05",
           849 => x"0c",
           850 => x"8a",
           851 => x"74",
           852 => x"26",
           853 => x"57",
           854 => x"76",
           855 => x"83",
           856 => x"86",
           857 => x"2e",
           858 => x"76",
           859 => x"83",
           860 => x"06",
           861 => x"3d",
           862 => x"f5",
           863 => x"08",
           864 => x"88",
           865 => x"08",
           866 => x"0c",
           867 => x"ff",
           868 => x"08",
           869 => x"2a",
           870 => x"0c",
           871 => x"81",
           872 => x"0b",
           873 => x"ac",
           874 => x"75",
           875 => x"3d",
           876 => x"3d",
           877 => x"0b",
           878 => x"55",
           879 => x"80",
           880 => x"38",
           881 => x"16",
           882 => x"e0",
           883 => x"54",
           884 => x"54",
           885 => x"51",
           886 => x"88",
           887 => x"08",
           888 => x"88",
           889 => x"73",
           890 => x"38",
           891 => x"33",
           892 => x"70",
           893 => x"55",
           894 => x"2e",
           895 => x"54",
           896 => x"51",
           897 => x"88",
           898 => x"0c",
           899 => x"05",
           900 => x"3f",
           901 => x"16",
           902 => x"16",
           903 => x"81",
           904 => x"88",
           905 => x"0d",
           906 => x"0d",
           907 => x"0b",
           908 => x"ac",
           909 => x"5c",
           910 => x"0c",
           911 => x"80",
           912 => x"38",
           913 => x"81",
           914 => x"57",
           915 => x"81",
           916 => x"39",
           917 => x"34",
           918 => x"0b",
           919 => x"81",
           920 => x"39",
           921 => x"98",
           922 => x"55",
           923 => x"83",
           924 => x"77",
           925 => x"9a",
           926 => x"08",
           927 => x"06",
           928 => x"80",
           929 => x"16",
           930 => x"77",
           931 => x"70",
           932 => x"5b",
           933 => x"38",
           934 => x"a0",
           935 => x"8b",
           936 => x"08",
           937 => x"3f",
           938 => x"81",
           939 => x"aa",
           940 => x"17",
           941 => x"08",
           942 => x"3f",
           943 => x"88",
           944 => x"ff",
           945 => x"08",
           946 => x"0c",
           947 => x"83",
           948 => x"80",
           949 => x"55",
           950 => x"83",
           951 => x"74",
           952 => x"08",
           953 => x"53",
           954 => x"52",
           955 => x"b5",
           956 => x"fe",
           957 => x"16",
           958 => x"17",
           959 => x"31",
           960 => x"7c",
           961 => x"80",
           962 => x"38",
           963 => x"fe",
           964 => x"57",
           965 => x"8c",
           966 => x"fb",
           967 => x"90",
           968 => x"87",
           969 => x"0c",
           970 => x"e4",
           971 => x"94",
           972 => x"80",
           973 => x"c0",
           974 => x"8c",
           975 => x"87",
           976 => x"0c",
           977 => x"f9",
           978 => x"08",
           979 => x"98",
           980 => x"3f",
           981 => x"38",
           982 => x"88",
           983 => x"98",
           984 => x"87",
           985 => x"53",
           986 => x"74",
           987 => x"3f",
           988 => x"38",
           989 => x"80",
           990 => x"73",
           991 => x"39",
           992 => x"73",
           993 => x"fb",
           994 => x"ff",
           995 => x"00",
           996 => x"ff",
           997 => x"ff",
           998 => x"4f",
           999 => x"49",
          1000 => x"52",
          1001 => x"00",
          1002 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"ca",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"04",
          2058 => x"c4",
          2059 => x"0b",
          2060 => x"04",
          2061 => x"c4",
          2062 => x"0b",
          2063 => x"04",
          2064 => x"c4",
          2065 => x"0b",
          2066 => x"04",
          2067 => x"c4",
          2068 => x"0b",
          2069 => x"04",
          2070 => x"c5",
          2071 => x"0b",
          2072 => x"04",
          2073 => x"c5",
          2074 => x"0b",
          2075 => x"04",
          2076 => x"c5",
          2077 => x"0b",
          2078 => x"04",
          2079 => x"c5",
          2080 => x"0b",
          2081 => x"04",
          2082 => x"c6",
          2083 => x"0b",
          2084 => x"04",
          2085 => x"c6",
          2086 => x"0b",
          2087 => x"04",
          2088 => x"c6",
          2089 => x"0b",
          2090 => x"04",
          2091 => x"c6",
          2092 => x"0b",
          2093 => x"04",
          2094 => x"c7",
          2095 => x"0b",
          2096 => x"04",
          2097 => x"c7",
          2098 => x"0b",
          2099 => x"04",
          2100 => x"c7",
          2101 => x"0b",
          2102 => x"04",
          2103 => x"c7",
          2104 => x"0b",
          2105 => x"04",
          2106 => x"c8",
          2107 => x"0b",
          2108 => x"04",
          2109 => x"c8",
          2110 => x"0b",
          2111 => x"04",
          2112 => x"c8",
          2113 => x"0b",
          2114 => x"04",
          2115 => x"c8",
          2116 => x"0b",
          2117 => x"04",
          2118 => x"c9",
          2119 => x"0b",
          2120 => x"04",
          2121 => x"c9",
          2122 => x"0b",
          2123 => x"04",
          2124 => x"c9",
          2125 => x"0b",
          2126 => x"04",
          2127 => x"c9",
          2128 => x"0b",
          2129 => x"04",
          2130 => x"ca",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"82",
          2178 => x"80",
          2179 => x"82",
          2180 => x"83",
          2181 => x"82",
          2182 => x"80",
          2183 => x"82",
          2184 => x"83",
          2185 => x"82",
          2186 => x"80",
          2187 => x"82",
          2188 => x"83",
          2189 => x"82",
          2190 => x"80",
          2191 => x"82",
          2192 => x"83",
          2193 => x"82",
          2194 => x"80",
          2195 => x"82",
          2196 => x"83",
          2197 => x"82",
          2198 => x"80",
          2199 => x"82",
          2200 => x"83",
          2201 => x"82",
          2202 => x"80",
          2203 => x"82",
          2204 => x"83",
          2205 => x"82",
          2206 => x"80",
          2207 => x"82",
          2208 => x"83",
          2209 => x"82",
          2210 => x"80",
          2211 => x"82",
          2212 => x"83",
          2213 => x"82",
          2214 => x"80",
          2215 => x"82",
          2216 => x"83",
          2217 => x"82",
          2218 => x"80",
          2219 => x"82",
          2220 => x"83",
          2221 => x"82",
          2222 => x"80",
          2223 => x"82",
          2224 => x"83",
          2225 => x"82",
          2226 => x"80",
          2227 => x"82",
          2228 => x"83",
          2229 => x"82",
          2230 => x"80",
          2231 => x"82",
          2232 => x"83",
          2233 => x"82",
          2234 => x"80",
          2235 => x"82",
          2236 => x"83",
          2237 => x"82",
          2238 => x"80",
          2239 => x"82",
          2240 => x"83",
          2241 => x"82",
          2242 => x"80",
          2243 => x"82",
          2244 => x"83",
          2245 => x"82",
          2246 => x"81",
          2247 => x"82",
          2248 => x"83",
          2249 => x"82",
          2250 => x"81",
          2251 => x"82",
          2252 => x"83",
          2253 => x"82",
          2254 => x"81",
          2255 => x"82",
          2256 => x"83",
          2257 => x"82",
          2258 => x"81",
          2259 => x"82",
          2260 => x"83",
          2261 => x"82",
          2262 => x"81",
          2263 => x"82",
          2264 => x"83",
          2265 => x"82",
          2266 => x"81",
          2267 => x"82",
          2268 => x"83",
          2269 => x"82",
          2270 => x"81",
          2271 => x"82",
          2272 => x"83",
          2273 => x"82",
          2274 => x"81",
          2275 => x"82",
          2276 => x"83",
          2277 => x"82",
          2278 => x"81",
          2279 => x"82",
          2280 => x"83",
          2281 => x"82",
          2282 => x"81",
          2283 => x"82",
          2284 => x"83",
          2285 => x"82",
          2286 => x"81",
          2287 => x"82",
          2288 => x"83",
          2289 => x"82",
          2290 => x"81",
          2291 => x"82",
          2292 => x"83",
          2293 => x"82",
          2294 => x"81",
          2295 => x"82",
          2296 => x"83",
          2297 => x"82",
          2298 => x"81",
          2299 => x"82",
          2300 => x"83",
          2301 => x"82",
          2302 => x"81",
          2303 => x"82",
          2304 => x"83",
          2305 => x"82",
          2306 => x"81",
          2307 => x"82",
          2308 => x"83",
          2309 => x"82",
          2310 => x"81",
          2311 => x"82",
          2312 => x"83",
          2313 => x"82",
          2314 => x"81",
          2315 => x"82",
          2316 => x"83",
          2317 => x"82",
          2318 => x"81",
          2319 => x"82",
          2320 => x"83",
          2321 => x"82",
          2322 => x"81",
          2323 => x"82",
          2324 => x"83",
          2325 => x"82",
          2326 => x"81",
          2327 => x"82",
          2328 => x"83",
          2329 => x"82",
          2330 => x"81",
          2331 => x"82",
          2332 => x"83",
          2333 => x"82",
          2334 => x"81",
          2335 => x"82",
          2336 => x"83",
          2337 => x"82",
          2338 => x"81",
          2339 => x"82",
          2340 => x"83",
          2341 => x"82",
          2342 => x"81",
          2343 => x"82",
          2344 => x"83",
          2345 => x"82",
          2346 => x"80",
          2347 => x"82",
          2348 => x"83",
          2349 => x"82",
          2350 => x"80",
          2351 => x"82",
          2352 => x"83",
          2353 => x"82",
          2354 => x"80",
          2355 => x"82",
          2356 => x"83",
          2357 => x"82",
          2358 => x"80",
          2359 => x"82",
          2360 => x"83",
          2361 => x"82",
          2362 => x"80",
          2363 => x"82",
          2364 => x"83",
          2365 => x"82",
          2366 => x"80",
          2367 => x"82",
          2368 => x"83",
          2369 => x"82",
          2370 => x"81",
          2371 => x"82",
          2372 => x"83",
          2373 => x"82",
          2374 => x"82",
          2375 => x"8e",
          2376 => x"70",
          2377 => x"0c",
          2378 => x"ca",
          2379 => x"c4",
          2380 => x"ef",
          2381 => x"04",
          2382 => x"08",
          2383 => x"d4",
          2384 => x"0d",
          2385 => x"93",
          2386 => x"05",
          2387 => x"93",
          2388 => x"05",
          2389 => x"c5",
          2390 => x"c8",
          2391 => x"93",
          2392 => x"85",
          2393 => x"93",
          2394 => x"82",
          2395 => x"02",
          2396 => x"0c",
          2397 => x"81",
          2398 => x"d4",
          2399 => x"08",
          2400 => x"d4",
          2401 => x"08",
          2402 => x"82",
          2403 => x"70",
          2404 => x"0c",
          2405 => x"0d",
          2406 => x"0c",
          2407 => x"d4",
          2408 => x"93",
          2409 => x"3d",
          2410 => x"82",
          2411 => x"fc",
          2412 => x"0b",
          2413 => x"08",
          2414 => x"82",
          2415 => x"8c",
          2416 => x"93",
          2417 => x"05",
          2418 => x"38",
          2419 => x"08",
          2420 => x"80",
          2421 => x"80",
          2422 => x"d4",
          2423 => x"08",
          2424 => x"82",
          2425 => x"8c",
          2426 => x"82",
          2427 => x"8c",
          2428 => x"93",
          2429 => x"05",
          2430 => x"93",
          2431 => x"05",
          2432 => x"39",
          2433 => x"08",
          2434 => x"80",
          2435 => x"38",
          2436 => x"08",
          2437 => x"82",
          2438 => x"88",
          2439 => x"ad",
          2440 => x"d4",
          2441 => x"08",
          2442 => x"08",
          2443 => x"31",
          2444 => x"08",
          2445 => x"82",
          2446 => x"f8",
          2447 => x"93",
          2448 => x"05",
          2449 => x"93",
          2450 => x"05",
          2451 => x"d4",
          2452 => x"08",
          2453 => x"93",
          2454 => x"05",
          2455 => x"d4",
          2456 => x"08",
          2457 => x"93",
          2458 => x"05",
          2459 => x"39",
          2460 => x"08",
          2461 => x"80",
          2462 => x"82",
          2463 => x"88",
          2464 => x"82",
          2465 => x"f4",
          2466 => x"91",
          2467 => x"d4",
          2468 => x"08",
          2469 => x"d4",
          2470 => x"0c",
          2471 => x"d4",
          2472 => x"08",
          2473 => x"0c",
          2474 => x"82",
          2475 => x"04",
          2476 => x"76",
          2477 => x"8c",
          2478 => x"33",
          2479 => x"55",
          2480 => x"8a",
          2481 => x"06",
          2482 => x"2e",
          2483 => x"12",
          2484 => x"2e",
          2485 => x"73",
          2486 => x"55",
          2487 => x"52",
          2488 => x"09",
          2489 => x"38",
          2490 => x"c8",
          2491 => x"0d",
          2492 => x"88",
          2493 => x"70",
          2494 => x"07",
          2495 => x"8f",
          2496 => x"38",
          2497 => x"84",
          2498 => x"72",
          2499 => x"05",
          2500 => x"71",
          2501 => x"53",
          2502 => x"70",
          2503 => x"0c",
          2504 => x"71",
          2505 => x"38",
          2506 => x"90",
          2507 => x"70",
          2508 => x"0c",
          2509 => x"71",
          2510 => x"38",
          2511 => x"8e",
          2512 => x"0d",
          2513 => x"72",
          2514 => x"53",
          2515 => x"93",
          2516 => x"73",
          2517 => x"54",
          2518 => x"2e",
          2519 => x"73",
          2520 => x"71",
          2521 => x"ff",
          2522 => x"70",
          2523 => x"38",
          2524 => x"70",
          2525 => x"81",
          2526 => x"81",
          2527 => x"71",
          2528 => x"ff",
          2529 => x"54",
          2530 => x"38",
          2531 => x"73",
          2532 => x"75",
          2533 => x"71",
          2534 => x"93",
          2535 => x"52",
          2536 => x"04",
          2537 => x"f7",
          2538 => x"14",
          2539 => x"84",
          2540 => x"06",
          2541 => x"70",
          2542 => x"14",
          2543 => x"08",
          2544 => x"71",
          2545 => x"dc",
          2546 => x"54",
          2547 => x"39",
          2548 => x"93",
          2549 => x"3d",
          2550 => x"3d",
          2551 => x"54",
          2552 => x"2b",
          2553 => x"3f",
          2554 => x"08",
          2555 => x"72",
          2556 => x"54",
          2557 => x"25",
          2558 => x"82",
          2559 => x"84",
          2560 => x"fc",
          2561 => x"70",
          2562 => x"55",
          2563 => x"2e",
          2564 => x"73",
          2565 => x"a0",
          2566 => x"06",
          2567 => x"14",
          2568 => x"54",
          2569 => x"f6",
          2570 => x"84",
          2571 => x"52",
          2572 => x"52",
          2573 => x"2e",
          2574 => x"53",
          2575 => x"9f",
          2576 => x"51",
          2577 => x"38",
          2578 => x"70",
          2579 => x"81",
          2580 => x"80",
          2581 => x"05",
          2582 => x"75",
          2583 => x"70",
          2584 => x"0c",
          2585 => x"04",
          2586 => x"76",
          2587 => x"80",
          2588 => x"86",
          2589 => x"52",
          2590 => x"c4",
          2591 => x"c8",
          2592 => x"80",
          2593 => x"74",
          2594 => x"93",
          2595 => x"3d",
          2596 => x"3d",
          2597 => x"11",
          2598 => x"5b",
          2599 => x"79",
          2600 => x"bf",
          2601 => x"33",
          2602 => x"82",
          2603 => x"26",
          2604 => x"84",
          2605 => x"83",
          2606 => x"26",
          2607 => x"85",
          2608 => x"84",
          2609 => x"26",
          2610 => x"86",
          2611 => x"85",
          2612 => x"26",
          2613 => x"88",
          2614 => x"86",
          2615 => x"e7",
          2616 => x"38",
          2617 => x"5a",
          2618 => x"87",
          2619 => x"f3",
          2620 => x"22",
          2621 => x"22",
          2622 => x"33",
          2623 => x"33",
          2624 => x"33",
          2625 => x"33",
          2626 => x"33",
          2627 => x"52",
          2628 => x"51",
          2629 => x"87",
          2630 => x"5b",
          2631 => x"7b",
          2632 => x"98",
          2633 => x"1c",
          2634 => x"98",
          2635 => x"1c",
          2636 => x"98",
          2637 => x"1c",
          2638 => x"98",
          2639 => x"1c",
          2640 => x"98",
          2641 => x"1c",
          2642 => x"98",
          2643 => x"1c",
          2644 => x"98",
          2645 => x"1c",
          2646 => x"98",
          2647 => x"7b",
          2648 => x"7a",
          2649 => x"0c",
          2650 => x"04",
          2651 => x"7d",
          2652 => x"98",
          2653 => x"7c",
          2654 => x"98",
          2655 => x"7a",
          2656 => x"c0",
          2657 => x"5b",
          2658 => x"34",
          2659 => x"b4",
          2660 => x"83",
          2661 => x"c0",
          2662 => x"5b",
          2663 => x"34",
          2664 => x"ac",
          2665 => x"85",
          2666 => x"c0",
          2667 => x"5b",
          2668 => x"34",
          2669 => x"a4",
          2670 => x"88",
          2671 => x"c0",
          2672 => x"5b",
          2673 => x"23",
          2674 => x"8a",
          2675 => x"88",
          2676 => x"86",
          2677 => x"85",
          2678 => x"84",
          2679 => x"83",
          2680 => x"82",
          2681 => x"79",
          2682 => x"f6",
          2683 => x"af",
          2684 => x"0d",
          2685 => x"0d",
          2686 => x"33",
          2687 => x"9f",
          2688 => x"51",
          2689 => x"82",
          2690 => x"82",
          2691 => x"fd",
          2692 => x"0b",
          2693 => x"c0",
          2694 => x"87",
          2695 => x"51",
          2696 => x"86",
          2697 => x"94",
          2698 => x"08",
          2699 => x"70",
          2700 => x"52",
          2701 => x"2e",
          2702 => x"91",
          2703 => x"06",
          2704 => x"d7",
          2705 => x"2a",
          2706 => x"81",
          2707 => x"70",
          2708 => x"38",
          2709 => x"70",
          2710 => x"51",
          2711 => x"38",
          2712 => x"8b",
          2713 => x"87",
          2714 => x"52",
          2715 => x"86",
          2716 => x"94",
          2717 => x"72",
          2718 => x"93",
          2719 => x"3d",
          2720 => x"3d",
          2721 => x"05",
          2722 => x"82",
          2723 => x"54",
          2724 => x"94",
          2725 => x"80",
          2726 => x"87",
          2727 => x"51",
          2728 => x"96",
          2729 => x"06",
          2730 => x"70",
          2731 => x"38",
          2732 => x"70",
          2733 => x"51",
          2734 => x"71",
          2735 => x"32",
          2736 => x"51",
          2737 => x"2e",
          2738 => x"93",
          2739 => x"06",
          2740 => x"ff",
          2741 => x"0b",
          2742 => x"33",
          2743 => x"94",
          2744 => x"80",
          2745 => x"87",
          2746 => x"52",
          2747 => x"85",
          2748 => x"fb",
          2749 => x"54",
          2750 => x"52",
          2751 => x"2e",
          2752 => x"73",
          2753 => x"55",
          2754 => x"82",
          2755 => x"54",
          2756 => x"94",
          2757 => x"80",
          2758 => x"87",
          2759 => x"51",
          2760 => x"96",
          2761 => x"06",
          2762 => x"70",
          2763 => x"38",
          2764 => x"70",
          2765 => x"51",
          2766 => x"71",
          2767 => x"32",
          2768 => x"51",
          2769 => x"2e",
          2770 => x"93",
          2771 => x"06",
          2772 => x"ff",
          2773 => x"0b",
          2774 => x"33",
          2775 => x"94",
          2776 => x"80",
          2777 => x"87",
          2778 => x"52",
          2779 => x"81",
          2780 => x"52",
          2781 => x"8b",
          2782 => x"93",
          2783 => x"3d",
          2784 => x"3d",
          2785 => x"82",
          2786 => x"52",
          2787 => x"84",
          2788 => x"2e",
          2789 => x"c0",
          2790 => x"70",
          2791 => x"2a",
          2792 => x"51",
          2793 => x"80",
          2794 => x"0b",
          2795 => x"c0",
          2796 => x"c0",
          2797 => x"70",
          2798 => x"38",
          2799 => x"90",
          2800 => x"70",
          2801 => x"82",
          2802 => x"51",
          2803 => x"04",
          2804 => x"0b",
          2805 => x"c0",
          2806 => x"c0",
          2807 => x"70",
          2808 => x"38",
          2809 => x"94",
          2810 => x"70",
          2811 => x"81",
          2812 => x"51",
          2813 => x"80",
          2814 => x"0b",
          2815 => x"c0",
          2816 => x"c0",
          2817 => x"70",
          2818 => x"38",
          2819 => x"90",
          2820 => x"70",
          2821 => x"98",
          2822 => x"51",
          2823 => x"c8",
          2824 => x"0d",
          2825 => x"0d",
          2826 => x"80",
          2827 => x"9c",
          2828 => x"51",
          2829 => x"80",
          2830 => x"38",
          2831 => x"0b",
          2832 => x"9c",
          2833 => x"84",
          2834 => x"9e",
          2835 => x"0c",
          2836 => x"87",
          2837 => x"08",
          2838 => x"8c",
          2839 => x"9e",
          2840 => x"0c",
          2841 => x"87",
          2842 => x"08",
          2843 => x"94",
          2844 => x"9e",
          2845 => x"0c",
          2846 => x"87",
          2847 => x"08",
          2848 => x"9c",
          2849 => x"9e",
          2850 => x"0c",
          2851 => x"87",
          2852 => x"08",
          2853 => x"73",
          2854 => x"70",
          2855 => x"a8",
          2856 => x"9e",
          2857 => x"0c",
          2858 => x"ac",
          2859 => x"12",
          2860 => x"87",
          2861 => x"08",
          2862 => x"06",
          2863 => x"70",
          2864 => x"38",
          2865 => x"72",
          2866 => x"87",
          2867 => x"08",
          2868 => x"80",
          2869 => x"52",
          2870 => x"83",
          2871 => x"71",
          2872 => x"34",
          2873 => x"c0",
          2874 => x"70",
          2875 => x"06",
          2876 => x"70",
          2877 => x"38",
          2878 => x"82",
          2879 => x"80",
          2880 => x"9e",
          2881 => x"90",
          2882 => x"52",
          2883 => x"2e",
          2884 => x"52",
          2885 => x"f4",
          2886 => x"87",
          2887 => x"08",
          2888 => x"06",
          2889 => x"70",
          2890 => x"38",
          2891 => x"82",
          2892 => x"80",
          2893 => x"9e",
          2894 => x"84",
          2895 => x"52",
          2896 => x"2e",
          2897 => x"52",
          2898 => x"f6",
          2899 => x"87",
          2900 => x"08",
          2901 => x"06",
          2902 => x"70",
          2903 => x"38",
          2904 => x"82",
          2905 => x"80",
          2906 => x"9e",
          2907 => x"81",
          2908 => x"52",
          2909 => x"2e",
          2910 => x"52",
          2911 => x"f8",
          2912 => x"f9",
          2913 => x"9e",
          2914 => x"70",
          2915 => x"70",
          2916 => x"51",
          2917 => x"72",
          2918 => x"54",
          2919 => x"80",
          2920 => x"90",
          2921 => x"52",
          2922 => x"83",
          2923 => x"71",
          2924 => x"0b",
          2925 => x"88",
          2926 => x"06",
          2927 => x"70",
          2928 => x"38",
          2929 => x"82",
          2930 => x"87",
          2931 => x"08",
          2932 => x"51",
          2933 => x"8b",
          2934 => x"3d",
          2935 => x"3d",
          2936 => x"c0",
          2937 => x"3f",
          2938 => x"33",
          2939 => x"2e",
          2940 => x"f6",
          2941 => x"ad",
          2942 => x"e8",
          2943 => x"3f",
          2944 => x"70",
          2945 => x"73",
          2946 => x"38",
          2947 => x"53",
          2948 => x"08",
          2949 => x"80",
          2950 => x"3f",
          2951 => x"70",
          2952 => x"73",
          2953 => x"38",
          2954 => x"53",
          2955 => x"52",
          2956 => x"51",
          2957 => x"82",
          2958 => x"33",
          2959 => x"8a",
          2960 => x"33",
          2961 => x"2e",
          2962 => x"8b",
          2963 => x"54",
          2964 => x"53",
          2965 => x"cc",
          2966 => x"3f",
          2967 => x"33",
          2968 => x"2e",
          2969 => x"f7",
          2970 => x"b9",
          2971 => x"f6",
          2972 => x"80",
          2973 => x"81",
          2974 => x"83",
          2975 => x"8b",
          2976 => x"73",
          2977 => x"38",
          2978 => x"51",
          2979 => x"82",
          2980 => x"33",
          2981 => x"80",
          2982 => x"81",
          2983 => x"81",
          2984 => x"88",
          2985 => x"8b",
          2986 => x"73",
          2987 => x"38",
          2988 => x"51",
          2989 => x"82",
          2990 => x"33",
          2991 => x"80",
          2992 => x"81",
          2993 => x"81",
          2994 => x"88",
          2995 => x"f8",
          2996 => x"d1",
          2997 => x"dc",
          2998 => x"84",
          2999 => x"54",
          3000 => x"53",
          3001 => x"b7",
          3002 => x"52",
          3003 => x"51",
          3004 => x"88",
          3005 => x"81",
          3006 => x"88",
          3007 => x"15",
          3008 => x"f9",
          3009 => x"97",
          3010 => x"08",
          3011 => x"98",
          3012 => x"3f",
          3013 => x"04",
          3014 => x"02",
          3015 => x"52",
          3016 => x"bb",
          3017 => x"10",
          3018 => x"f0",
          3019 => x"71",
          3020 => x"fa",
          3021 => x"bb",
          3022 => x"81",
          3023 => x"f7",
          3024 => x"39",
          3025 => x"51",
          3026 => x"9a",
          3027 => x"d8",
          3028 => x"3f",
          3029 => x"fa",
          3030 => x"97",
          3031 => x"81",
          3032 => x"f7",
          3033 => x"3d",
          3034 => x"88",
          3035 => x"80",
          3036 => x"96",
          3037 => x"ff",
          3038 => x"c0",
          3039 => x"08",
          3040 => x"72",
          3041 => x"07",
          3042 => x"80",
          3043 => x"83",
          3044 => x"ff",
          3045 => x"c0",
          3046 => x"08",
          3047 => x"0c",
          3048 => x"0c",
          3049 => x"82",
          3050 => x"06",
          3051 => x"80",
          3052 => x"51",
          3053 => x"04",
          3054 => x"08",
          3055 => x"84",
          3056 => x"3d",
          3057 => x"05",
          3058 => x"8a",
          3059 => x"06",
          3060 => x"51",
          3061 => x"93",
          3062 => x"2e",
          3063 => x"93",
          3064 => x"72",
          3065 => x"93",
          3066 => x"05",
          3067 => x"0c",
          3068 => x"93",
          3069 => x"2e",
          3070 => x"51",
          3071 => x"08",
          3072 => x"84",
          3073 => x"fe",
          3074 => x"97",
          3075 => x"93",
          3076 => x"82",
          3077 => x"54",
          3078 => x"3f",
          3079 => x"d8",
          3080 => x"0d",
          3081 => x"0d",
          3082 => x"53",
          3083 => x"2e",
          3084 => x"70",
          3085 => x"33",
          3086 => x"3f",
          3087 => x"71",
          3088 => x"3d",
          3089 => x"3d",
          3090 => x"93",
          3091 => x"82",
          3092 => x"71",
          3093 => x"53",
          3094 => x"91",
          3095 => x"81",
          3096 => x"51",
          3097 => x"72",
          3098 => x"f1",
          3099 => x"93",
          3100 => x"3d",
          3101 => x"3d",
          3102 => x"5d",
          3103 => x"81",
          3104 => x"56",
          3105 => x"85",
          3106 => x"a5",
          3107 => x"75",
          3108 => x"3f",
          3109 => x"70",
          3110 => x"05",
          3111 => x"5e",
          3112 => x"2e",
          3113 => x"8c",
          3114 => x"70",
          3115 => x"33",
          3116 => x"39",
          3117 => x"09",
          3118 => x"38",
          3119 => x"81",
          3120 => x"57",
          3121 => x"2e",
          3122 => x"92",
          3123 => x"1d",
          3124 => x"70",
          3125 => x"33",
          3126 => x"53",
          3127 => x"16",
          3128 => x"26",
          3129 => x"8a",
          3130 => x"05",
          3131 => x"05",
          3132 => x"11",
          3133 => x"89",
          3134 => x"38",
          3135 => x"32",
          3136 => x"72",
          3137 => x"78",
          3138 => x"70",
          3139 => x"07",
          3140 => x"07",
          3141 => x"52",
          3142 => x"80",
          3143 => x"7c",
          3144 => x"70",
          3145 => x"33",
          3146 => x"80",
          3147 => x"38",
          3148 => x"e0",
          3149 => x"38",
          3150 => x"81",
          3151 => x"53",
          3152 => x"53",
          3153 => x"81",
          3154 => x"10",
          3155 => x"dc",
          3156 => x"08",
          3157 => x"1d",
          3158 => x"5d",
          3159 => x"33",
          3160 => x"74",
          3161 => x"81",
          3162 => x"70",
          3163 => x"54",
          3164 => x"7c",
          3165 => x"81",
          3166 => x"72",
          3167 => x"81",
          3168 => x"72",
          3169 => x"38",
          3170 => x"81",
          3171 => x"51",
          3172 => x"75",
          3173 => x"81",
          3174 => x"79",
          3175 => x"38",
          3176 => x"81",
          3177 => x"15",
          3178 => x"7a",
          3179 => x"38",
          3180 => x"8e",
          3181 => x"15",
          3182 => x"73",
          3183 => x"fd",
          3184 => x"84",
          3185 => x"33",
          3186 => x"fb",
          3187 => x"ad",
          3188 => x"95",
          3189 => x"91",
          3190 => x"8d",
          3191 => x"89",
          3192 => x"fb",
          3193 => x"95",
          3194 => x"2a",
          3195 => x"51",
          3196 => x"2e",
          3197 => x"84",
          3198 => x"59",
          3199 => x"39",
          3200 => x"2e",
          3201 => x"8b",
          3202 => x"1d",
          3203 => x"5d",
          3204 => x"7b",
          3205 => x"08",
          3206 => x"74",
          3207 => x"70",
          3208 => x"07",
          3209 => x"80",
          3210 => x"51",
          3211 => x"72",
          3212 => x"38",
          3213 => x"90",
          3214 => x"80",
          3215 => x"76",
          3216 => x"3f",
          3217 => x"08",
          3218 => x"7b",
          3219 => x"55",
          3220 => x"82",
          3221 => x"57",
          3222 => x"99",
          3223 => x"16",
          3224 => x"06",
          3225 => x"75",
          3226 => x"89",
          3227 => x"70",
          3228 => x"56",
          3229 => x"78",
          3230 => x"b0",
          3231 => x"72",
          3232 => x"18",
          3233 => x"79",
          3234 => x"70",
          3235 => x"06",
          3236 => x"58",
          3237 => x"38",
          3238 => x"70",
          3239 => x"53",
          3240 => x"8e",
          3241 => x"78",
          3242 => x"53",
          3243 => x"81",
          3244 => x"7d",
          3245 => x"54",
          3246 => x"83",
          3247 => x"7c",
          3248 => x"81",
          3249 => x"72",
          3250 => x"81",
          3251 => x"72",
          3252 => x"38",
          3253 => x"81",
          3254 => x"51",
          3255 => x"75",
          3256 => x"81",
          3257 => x"79",
          3258 => x"38",
          3259 => x"3d",
          3260 => x"70",
          3261 => x"58",
          3262 => x"77",
          3263 => x"81",
          3264 => x"72",
          3265 => x"f5",
          3266 => x"f9",
          3267 => x"81",
          3268 => x"79",
          3269 => x"38",
          3270 => x"96",
          3271 => x"fd",
          3272 => x"3d",
          3273 => x"05",
          3274 => x"52",
          3275 => x"c6",
          3276 => x"0d",
          3277 => x"0d",
          3278 => x"e0",
          3279 => x"88",
          3280 => x"51",
          3281 => x"82",
          3282 => x"53",
          3283 => x"80",
          3284 => x"e0",
          3285 => x"0d",
          3286 => x"0d",
          3287 => x"08",
          3288 => x"d8",
          3289 => x"88",
          3290 => x"52",
          3291 => x"3f",
          3292 => x"d8",
          3293 => x"0d",
          3294 => x"0d",
          3295 => x"57",
          3296 => x"93",
          3297 => x"2e",
          3298 => x"86",
          3299 => x"80",
          3300 => x"55",
          3301 => x"08",
          3302 => x"82",
          3303 => x"81",
          3304 => x"73",
          3305 => x"38",
          3306 => x"80",
          3307 => x"88",
          3308 => x"76",
          3309 => x"07",
          3310 => x"80",
          3311 => x"54",
          3312 => x"80",
          3313 => x"ff",
          3314 => x"ff",
          3315 => x"f7",
          3316 => x"39",
          3317 => x"ff",
          3318 => x"16",
          3319 => x"25",
          3320 => x"76",
          3321 => x"72",
          3322 => x"74",
          3323 => x"52",
          3324 => x"3f",
          3325 => x"74",
          3326 => x"72",
          3327 => x"f7",
          3328 => x"53",
          3329 => x"c8",
          3330 => x"0d",
          3331 => x"0d",
          3332 => x"08",
          3333 => x"dc",
          3334 => x"76",
          3335 => x"d9",
          3336 => x"93",
          3337 => x"3d",
          3338 => x"3d",
          3339 => x"5a",
          3340 => x"7a",
          3341 => x"70",
          3342 => x"58",
          3343 => x"09",
          3344 => x"38",
          3345 => x"05",
          3346 => x"08",
          3347 => x"53",
          3348 => x"f0",
          3349 => x"2e",
          3350 => x"8e",
          3351 => x"08",
          3352 => x"75",
          3353 => x"56",
          3354 => x"b0",
          3355 => x"06",
          3356 => x"74",
          3357 => x"75",
          3358 => x"70",
          3359 => x"73",
          3360 => x"9a",
          3361 => x"f8",
          3362 => x"06",
          3363 => x"0b",
          3364 => x"0c",
          3365 => x"33",
          3366 => x"80",
          3367 => x"75",
          3368 => x"76",
          3369 => x"70",
          3370 => x"57",
          3371 => x"56",
          3372 => x"81",
          3373 => x"14",
          3374 => x"88",
          3375 => x"27",
          3376 => x"f3",
          3377 => x"53",
          3378 => x"89",
          3379 => x"38",
          3380 => x"56",
          3381 => x"80",
          3382 => x"39",
          3383 => x"56",
          3384 => x"80",
          3385 => x"e0",
          3386 => x"38",
          3387 => x"81",
          3388 => x"53",
          3389 => x"81",
          3390 => x"53",
          3391 => x"8e",
          3392 => x"70",
          3393 => x"55",
          3394 => x"27",
          3395 => x"77",
          3396 => x"76",
          3397 => x"75",
          3398 => x"76",
          3399 => x"70",
          3400 => x"56",
          3401 => x"ff",
          3402 => x"80",
          3403 => x"75",
          3404 => x"79",
          3405 => x"75",
          3406 => x"0c",
          3407 => x"04",
          3408 => x"7a",
          3409 => x"80",
          3410 => x"75",
          3411 => x"56",
          3412 => x"a0",
          3413 => x"06",
          3414 => x"08",
          3415 => x"0c",
          3416 => x"33",
          3417 => x"a0",
          3418 => x"73",
          3419 => x"81",
          3420 => x"81",
          3421 => x"76",
          3422 => x"70",
          3423 => x"58",
          3424 => x"09",
          3425 => x"d3",
          3426 => x"81",
          3427 => x"74",
          3428 => x"55",
          3429 => x"e2",
          3430 => x"73",
          3431 => x"09",
          3432 => x"38",
          3433 => x"14",
          3434 => x"08",
          3435 => x"54",
          3436 => x"39",
          3437 => x"81",
          3438 => x"75",
          3439 => x"56",
          3440 => x"39",
          3441 => x"74",
          3442 => x"38",
          3443 => x"80",
          3444 => x"89",
          3445 => x"38",
          3446 => x"d0",
          3447 => x"56",
          3448 => x"80",
          3449 => x"39",
          3450 => x"e1",
          3451 => x"80",
          3452 => x"57",
          3453 => x"74",
          3454 => x"38",
          3455 => x"27",
          3456 => x"14",
          3457 => x"06",
          3458 => x"14",
          3459 => x"06",
          3460 => x"74",
          3461 => x"f9",
          3462 => x"ff",
          3463 => x"89",
          3464 => x"38",
          3465 => x"c5",
          3466 => x"29",
          3467 => x"81",
          3468 => x"75",
          3469 => x"56",
          3470 => x"a0",
          3471 => x"38",
          3472 => x"84",
          3473 => x"56",
          3474 => x"81",
          3475 => x"93",
          3476 => x"3d",
          3477 => x"3d",
          3478 => x"05",
          3479 => x"52",
          3480 => x"87",
          3481 => x"84",
          3482 => x"71",
          3483 => x"0c",
          3484 => x"04",
          3485 => x"02",
          3486 => x"02",
          3487 => x"05",
          3488 => x"83",
          3489 => x"26",
          3490 => x"72",
          3491 => x"c0",
          3492 => x"51",
          3493 => x"80",
          3494 => x"81",
          3495 => x"71",
          3496 => x"29",
          3497 => x"8c",
          3498 => x"71",
          3499 => x"87",
          3500 => x"0c",
          3501 => x"c0",
          3502 => x"71",
          3503 => x"06",
          3504 => x"80",
          3505 => x"73",
          3506 => x"ef",
          3507 => x"29",
          3508 => x"8c",
          3509 => x"fc",
          3510 => x"53",
          3511 => x"38",
          3512 => x"8c",
          3513 => x"80",
          3514 => x"71",
          3515 => x"14",
          3516 => x"84",
          3517 => x"70",
          3518 => x"0c",
          3519 => x"04",
          3520 => x"61",
          3521 => x"8c",
          3522 => x"05",
          3523 => x"5d",
          3524 => x"52",
          3525 => x"3f",
          3526 => x"08",
          3527 => x"55",
          3528 => x"ac",
          3529 => x"58",
          3530 => x"98",
          3531 => x"2b",
          3532 => x"8c",
          3533 => x"92",
          3534 => x"42",
          3535 => x"56",
          3536 => x"87",
          3537 => x"1a",
          3538 => x"52",
          3539 => x"74",
          3540 => x"2a",
          3541 => x"51",
          3542 => x"80",
          3543 => x"78",
          3544 => x"78",
          3545 => x"5a",
          3546 => x"57",
          3547 => x"52",
          3548 => x"87",
          3549 => x"52",
          3550 => x"75",
          3551 => x"80",
          3552 => x"76",
          3553 => x"99",
          3554 => x"0c",
          3555 => x"8c",
          3556 => x"08",
          3557 => x"51",
          3558 => x"38",
          3559 => x"8d",
          3560 => x"1c",
          3561 => x"81",
          3562 => x"53",
          3563 => x"2e",
          3564 => x"fc",
          3565 => x"52",
          3566 => x"7e",
          3567 => x"80",
          3568 => x"80",
          3569 => x"71",
          3570 => x"38",
          3571 => x"54",
          3572 => x"c8",
          3573 => x"0d",
          3574 => x"0d",
          3575 => x"02",
          3576 => x"05",
          3577 => x"5c",
          3578 => x"52",
          3579 => x"3f",
          3580 => x"08",
          3581 => x"55",
          3582 => x"ae",
          3583 => x"87",
          3584 => x"73",
          3585 => x"c0",
          3586 => x"87",
          3587 => x"12",
          3588 => x"57",
          3589 => x"76",
          3590 => x"92",
          3591 => x"71",
          3592 => x"75",
          3593 => x"74",
          3594 => x"2a",
          3595 => x"51",
          3596 => x"80",
          3597 => x"76",
          3598 => x"58",
          3599 => x"81",
          3600 => x"81",
          3601 => x"06",
          3602 => x"80",
          3603 => x"75",
          3604 => x"d3",
          3605 => x"52",
          3606 => x"87",
          3607 => x"80",
          3608 => x"81",
          3609 => x"c0",
          3610 => x"53",
          3611 => x"82",
          3612 => x"71",
          3613 => x"1a",
          3614 => x"81",
          3615 => x"ff",
          3616 => x"1d",
          3617 => x"79",
          3618 => x"38",
          3619 => x"80",
          3620 => x"87",
          3621 => x"26",
          3622 => x"73",
          3623 => x"06",
          3624 => x"2e",
          3625 => x"52",
          3626 => x"82",
          3627 => x"8f",
          3628 => x"f7",
          3629 => x"02",
          3630 => x"05",
          3631 => x"05",
          3632 => x"71",
          3633 => x"56",
          3634 => x"82",
          3635 => x"81",
          3636 => x"54",
          3637 => x"81",
          3638 => x"2e",
          3639 => x"74",
          3640 => x"72",
          3641 => x"38",
          3642 => x"83",
          3643 => x"a0",
          3644 => x"29",
          3645 => x"8c",
          3646 => x"51",
          3647 => x"88",
          3648 => x"0c",
          3649 => x"39",
          3650 => x"0c",
          3651 => x"39",
          3652 => x"82",
          3653 => x"8b",
          3654 => x"ff",
          3655 => x"70",
          3656 => x"33",
          3657 => x"72",
          3658 => x"c8",
          3659 => x"52",
          3660 => x"04",
          3661 => x"75",
          3662 => x"82",
          3663 => x"90",
          3664 => x"2b",
          3665 => x"33",
          3666 => x"33",
          3667 => x"07",
          3668 => x"0c",
          3669 => x"54",
          3670 => x"0d",
          3671 => x"0d",
          3672 => x"05",
          3673 => x"52",
          3674 => x"70",
          3675 => x"34",
          3676 => x"51",
          3677 => x"83",
          3678 => x"ff",
          3679 => x"75",
          3680 => x"72",
          3681 => x"54",
          3682 => x"2a",
          3683 => x"70",
          3684 => x"34",
          3685 => x"51",
          3686 => x"81",
          3687 => x"70",
          3688 => x"70",
          3689 => x"3d",
          3690 => x"3d",
          3691 => x"77",
          3692 => x"70",
          3693 => x"38",
          3694 => x"05",
          3695 => x"70",
          3696 => x"34",
          3697 => x"70",
          3698 => x"3d",
          3699 => x"3d",
          3700 => x"76",
          3701 => x"72",
          3702 => x"05",
          3703 => x"11",
          3704 => x"38",
          3705 => x"04",
          3706 => x"78",
          3707 => x"56",
          3708 => x"81",
          3709 => x"74",
          3710 => x"56",
          3711 => x"31",
          3712 => x"52",
          3713 => x"80",
          3714 => x"71",
          3715 => x"38",
          3716 => x"c8",
          3717 => x"0d",
          3718 => x"0d",
          3719 => x"33",
          3720 => x"70",
          3721 => x"38",
          3722 => x"94",
          3723 => x"70",
          3724 => x"70",
          3725 => x"38",
          3726 => x"09",
          3727 => x"38",
          3728 => x"93",
          3729 => x"3d",
          3730 => x"0b",
          3731 => x"0c",
          3732 => x"82",
          3733 => x"04",
          3734 => x"79",
          3735 => x"83",
          3736 => x"58",
          3737 => x"80",
          3738 => x"54",
          3739 => x"53",
          3740 => x"53",
          3741 => x"52",
          3742 => x"3f",
          3743 => x"08",
          3744 => x"81",
          3745 => x"82",
          3746 => x"83",
          3747 => x"16",
          3748 => x"08",
          3749 => x"9c",
          3750 => x"a4",
          3751 => x"33",
          3752 => x"2e",
          3753 => x"98",
          3754 => x"b0",
          3755 => x"17",
          3756 => x"76",
          3757 => x"33",
          3758 => x"3f",
          3759 => x"58",
          3760 => x"c8",
          3761 => x"0d",
          3762 => x"0d",
          3763 => x"57",
          3764 => x"17",
          3765 => x"af",
          3766 => x"fe",
          3767 => x"93",
          3768 => x"82",
          3769 => x"9f",
          3770 => x"74",
          3771 => x"52",
          3772 => x"51",
          3773 => x"82",
          3774 => x"80",
          3775 => x"ff",
          3776 => x"74",
          3777 => x"75",
          3778 => x"0c",
          3779 => x"04",
          3780 => x"7a",
          3781 => x"fe",
          3782 => x"93",
          3783 => x"82",
          3784 => x"81",
          3785 => x"33",
          3786 => x"2e",
          3787 => x"80",
          3788 => x"17",
          3789 => x"81",
          3790 => x"06",
          3791 => x"84",
          3792 => x"93",
          3793 => x"b4",
          3794 => x"56",
          3795 => x"82",
          3796 => x"84",
          3797 => x"fc",
          3798 => x"8b",
          3799 => x"52",
          3800 => x"97",
          3801 => x"85",
          3802 => x"84",
          3803 => x"fc",
          3804 => x"17",
          3805 => x"9c",
          3806 => x"ff",
          3807 => x"08",
          3808 => x"17",
          3809 => x"3f",
          3810 => x"81",
          3811 => x"19",
          3812 => x"53",
          3813 => x"17",
          3814 => x"bd",
          3815 => x"18",
          3816 => x"80",
          3817 => x"33",
          3818 => x"3f",
          3819 => x"08",
          3820 => x"38",
          3821 => x"82",
          3822 => x"8a",
          3823 => x"fb",
          3824 => x"fe",
          3825 => x"08",
          3826 => x"56",
          3827 => x"74",
          3828 => x"38",
          3829 => x"70",
          3830 => x"16",
          3831 => x"53",
          3832 => x"c8",
          3833 => x"0d",
          3834 => x"0d",
          3835 => x"08",
          3836 => x"81",
          3837 => x"38",
          3838 => x"75",
          3839 => x"81",
          3840 => x"39",
          3841 => x"54",
          3842 => x"2e",
          3843 => x"72",
          3844 => x"38",
          3845 => x"8d",
          3846 => x"39",
          3847 => x"81",
          3848 => x"b6",
          3849 => x"2a",
          3850 => x"2a",
          3851 => x"05",
          3852 => x"57",
          3853 => x"82",
          3854 => x"81",
          3855 => x"83",
          3856 => x"b4",
          3857 => x"19",
          3858 => x"a4",
          3859 => x"55",
          3860 => x"59",
          3861 => x"3f",
          3862 => x"08",
          3863 => x"76",
          3864 => x"14",
          3865 => x"70",
          3866 => x"07",
          3867 => x"71",
          3868 => x"52",
          3869 => x"72",
          3870 => x"77",
          3871 => x"56",
          3872 => x"74",
          3873 => x"15",
          3874 => x"73",
          3875 => x"3f",
          3876 => x"08",
          3877 => x"74",
          3878 => x"06",
          3879 => x"05",
          3880 => x"3f",
          3881 => x"08",
          3882 => x"06",
          3883 => x"74",
          3884 => x"15",
          3885 => x"73",
          3886 => x"3f",
          3887 => x"08",
          3888 => x"82",
          3889 => x"06",
          3890 => x"05",
          3891 => x"3f",
          3892 => x"08",
          3893 => x"56",
          3894 => x"56",
          3895 => x"c8",
          3896 => x"0d",
          3897 => x"0d",
          3898 => x"58",
          3899 => x"57",
          3900 => x"82",
          3901 => x"98",
          3902 => x"82",
          3903 => x"33",
          3904 => x"2e",
          3905 => x"72",
          3906 => x"38",
          3907 => x"8d",
          3908 => x"39",
          3909 => x"81",
          3910 => x"88",
          3911 => x"2a",
          3912 => x"2a",
          3913 => x"05",
          3914 => x"59",
          3915 => x"82",
          3916 => x"57",
          3917 => x"08",
          3918 => x"78",
          3919 => x"15",
          3920 => x"1b",
          3921 => x"56",
          3922 => x"75",
          3923 => x"2e",
          3924 => x"84",
          3925 => x"06",
          3926 => x"06",
          3927 => x"53",
          3928 => x"81",
          3929 => x"34",
          3930 => x"a4",
          3931 => x"52",
          3932 => x"d5",
          3933 => x"c8",
          3934 => x"93",
          3935 => x"a4",
          3936 => x"ff",
          3937 => x"11",
          3938 => x"78",
          3939 => x"55",
          3940 => x"8f",
          3941 => x"2a",
          3942 => x"8f",
          3943 => x"f0",
          3944 => x"73",
          3945 => x"0b",
          3946 => x"80",
          3947 => x"88",
          3948 => x"08",
          3949 => x"51",
          3950 => x"82",
          3951 => x"57",
          3952 => x"08",
          3953 => x"75",
          3954 => x"06",
          3955 => x"83",
          3956 => x"05",
          3957 => x"f7",
          3958 => x"0b",
          3959 => x"80",
          3960 => x"87",
          3961 => x"08",
          3962 => x"51",
          3963 => x"82",
          3964 => x"57",
          3965 => x"08",
          3966 => x"f0",
          3967 => x"82",
          3968 => x"06",
          3969 => x"05",
          3970 => x"54",
          3971 => x"3f",
          3972 => x"08",
          3973 => x"76",
          3974 => x"51",
          3975 => x"81",
          3976 => x"34",
          3977 => x"c8",
          3978 => x"0d",
          3979 => x"0d",
          3980 => x"72",
          3981 => x"55",
          3982 => x"27",
          3983 => x"15",
          3984 => x"86",
          3985 => x"81",
          3986 => x"80",
          3987 => x"ff",
          3988 => x"74",
          3989 => x"3f",
          3990 => x"08",
          3991 => x"c8",
          3992 => x"38",
          3993 => x"56",
          3994 => x"81",
          3995 => x"39",
          3996 => x"08",
          3997 => x"39",
          3998 => x"51",
          3999 => x"82",
          4000 => x"56",
          4001 => x"08",
          4002 => x"c9",
          4003 => x"c8",
          4004 => x"d2",
          4005 => x"c8",
          4006 => x"cf",
          4007 => x"73",
          4008 => x"fc",
          4009 => x"93",
          4010 => x"38",
          4011 => x"fe",
          4012 => x"15",
          4013 => x"93",
          4014 => x"08",
          4015 => x"16",
          4016 => x"33",
          4017 => x"73",
          4018 => x"75",
          4019 => x"08",
          4020 => x"a4",
          4021 => x"75",
          4022 => x"0c",
          4023 => x"04",
          4024 => x"7d",
          4025 => x"5b",
          4026 => x"95",
          4027 => x"08",
          4028 => x"2e",
          4029 => x"19",
          4030 => x"b7",
          4031 => x"b3",
          4032 => x"7b",
          4033 => x"3f",
          4034 => x"82",
          4035 => x"27",
          4036 => x"82",
          4037 => x"55",
          4038 => x"08",
          4039 => x"db",
          4040 => x"c8",
          4041 => x"19",
          4042 => x"c8",
          4043 => x"cb",
          4044 => x"80",
          4045 => x"08",
          4046 => x"bf",
          4047 => x"77",
          4048 => x"81",
          4049 => x"38",
          4050 => x"98",
          4051 => x"26",
          4052 => x"57",
          4053 => x"51",
          4054 => x"82",
          4055 => x"56",
          4056 => x"93",
          4057 => x"2e",
          4058 => x"86",
          4059 => x"c8",
          4060 => x"ff",
          4061 => x"70",
          4062 => x"25",
          4063 => x"79",
          4064 => x"56",
          4065 => x"f3",
          4066 => x"2e",
          4067 => x"19",
          4068 => x"76",
          4069 => x"75",
          4070 => x"27",
          4071 => x"58",
          4072 => x"80",
          4073 => x"57",
          4074 => x"98",
          4075 => x"26",
          4076 => x"57",
          4077 => x"81",
          4078 => x"52",
          4079 => x"a9",
          4080 => x"c8",
          4081 => x"93",
          4082 => x"2e",
          4083 => x"5a",
          4084 => x"08",
          4085 => x"81",
          4086 => x"82",
          4087 => x"5a",
          4088 => x"70",
          4089 => x"07",
          4090 => x"7d",
          4091 => x"56",
          4092 => x"ff",
          4093 => x"2e",
          4094 => x"ff",
          4095 => x"55",
          4096 => x"ff",
          4097 => x"78",
          4098 => x"3f",
          4099 => x"08",
          4100 => x"08",
          4101 => x"93",
          4102 => x"80",
          4103 => x"70",
          4104 => x"2a",
          4105 => x"57",
          4106 => x"74",
          4107 => x"38",
          4108 => x"52",
          4109 => x"ad",
          4110 => x"c8",
          4111 => x"a6",
          4112 => x"1a",
          4113 => x"08",
          4114 => x"90",
          4115 => x"26",
          4116 => x"19",
          4117 => x"90",
          4118 => x"19",
          4119 => x"54",
          4120 => x"34",
          4121 => x"57",
          4122 => x"8d",
          4123 => x"80",
          4124 => x"75",
          4125 => x"81",
          4126 => x"74",
          4127 => x"0c",
          4128 => x"04",
          4129 => x"7b",
          4130 => x"f3",
          4131 => x"55",
          4132 => x"08",
          4133 => x"7c",
          4134 => x"f6",
          4135 => x"93",
          4136 => x"93",
          4137 => x"19",
          4138 => x"80",
          4139 => x"b4",
          4140 => x"55",
          4141 => x"74",
          4142 => x"80",
          4143 => x"77",
          4144 => x"17",
          4145 => x"75",
          4146 => x"77",
          4147 => x"53",
          4148 => x"17",
          4149 => x"81",
          4150 => x"c8",
          4151 => x"df",
          4152 => x"8a",
          4153 => x"58",
          4154 => x"83",
          4155 => x"77",
          4156 => x"93",
          4157 => x"3d",
          4158 => x"3d",
          4159 => x"71",
          4160 => x"57",
          4161 => x"0a",
          4162 => x"74",
          4163 => x"72",
          4164 => x"38",
          4165 => x"ae",
          4166 => x"18",
          4167 => x"08",
          4168 => x"38",
          4169 => x"82",
          4170 => x"38",
          4171 => x"54",
          4172 => x"74",
          4173 => x"82",
          4174 => x"22",
          4175 => x"79",
          4176 => x"38",
          4177 => x"98",
          4178 => x"d1",
          4179 => x"22",
          4180 => x"54",
          4181 => x"26",
          4182 => x"52",
          4183 => x"89",
          4184 => x"c8",
          4185 => x"93",
          4186 => x"2e",
          4187 => x"0b",
          4188 => x"08",
          4189 => x"98",
          4190 => x"93",
          4191 => x"86",
          4192 => x"80",
          4193 => x"73",
          4194 => x"73",
          4195 => x"73",
          4196 => x"f4",
          4197 => x"93",
          4198 => x"18",
          4199 => x"18",
          4200 => x"98",
          4201 => x"2e",
          4202 => x"39",
          4203 => x"39",
          4204 => x"98",
          4205 => x"98",
          4206 => x"83",
          4207 => x"b4",
          4208 => x"0c",
          4209 => x"82",
          4210 => x"8a",
          4211 => x"f9",
          4212 => x"7b",
          4213 => x"13",
          4214 => x"59",
          4215 => x"f0",
          4216 => x"27",
          4217 => x"0b",
          4218 => x"84",
          4219 => x"08",
          4220 => x"da",
          4221 => x"ff",
          4222 => x"81",
          4223 => x"15",
          4224 => x"98",
          4225 => x"15",
          4226 => x"75",
          4227 => x"18",
          4228 => x"77",
          4229 => x"a6",
          4230 => x"16",
          4231 => x"81",
          4232 => x"17",
          4233 => x"77",
          4234 => x"51",
          4235 => x"8e",
          4236 => x"08",
          4237 => x"f3",
          4238 => x"93",
          4239 => x"82",
          4240 => x"82",
          4241 => x"27",
          4242 => x"81",
          4243 => x"c8",
          4244 => x"80",
          4245 => x"17",
          4246 => x"c8",
          4247 => x"cc",
          4248 => x"38",
          4249 => x"0c",
          4250 => x"e2",
          4251 => x"08",
          4252 => x"f8",
          4253 => x"93",
          4254 => x"87",
          4255 => x"c8",
          4256 => x"80",
          4257 => x"53",
          4258 => x"08",
          4259 => x"38",
          4260 => x"93",
          4261 => x"2e",
          4262 => x"93",
          4263 => x"76",
          4264 => x"3f",
          4265 => x"93",
          4266 => x"38",
          4267 => x"0c",
          4268 => x"51",
          4269 => x"82",
          4270 => x"98",
          4271 => x"90",
          4272 => x"83",
          4273 => x"b4",
          4274 => x"0c",
          4275 => x"82",
          4276 => x"89",
          4277 => x"f8",
          4278 => x"7c",
          4279 => x"5a",
          4280 => x"75",
          4281 => x"3f",
          4282 => x"08",
          4283 => x"c8",
          4284 => x"38",
          4285 => x"08",
          4286 => x"08",
          4287 => x"ef",
          4288 => x"93",
          4289 => x"82",
          4290 => x"80",
          4291 => x"93",
          4292 => x"17",
          4293 => x"51",
          4294 => x"81",
          4295 => x"81",
          4296 => x"81",
          4297 => x"70",
          4298 => x"07",
          4299 => x"80",
          4300 => x"81",
          4301 => x"79",
          4302 => x"83",
          4303 => x"81",
          4304 => x"fd",
          4305 => x"93",
          4306 => x"82",
          4307 => x"80",
          4308 => x"38",
          4309 => x"09",
          4310 => x"38",
          4311 => x"82",
          4312 => x"8a",
          4313 => x"fd",
          4314 => x"9a",
          4315 => x"eb",
          4316 => x"93",
          4317 => x"ff",
          4318 => x"70",
          4319 => x"53",
          4320 => x"09",
          4321 => x"38",
          4322 => x"eb",
          4323 => x"93",
          4324 => x"2b",
          4325 => x"72",
          4326 => x"0c",
          4327 => x"04",
          4328 => x"77",
          4329 => x"ff",
          4330 => x"9a",
          4331 => x"55",
          4332 => x"76",
          4333 => x"53",
          4334 => x"09",
          4335 => x"38",
          4336 => x"52",
          4337 => x"eb",
          4338 => x"3d",
          4339 => x"3d",
          4340 => x"5b",
          4341 => x"08",
          4342 => x"16",
          4343 => x"81",
          4344 => x"16",
          4345 => x"51",
          4346 => x"82",
          4347 => x"58",
          4348 => x"08",
          4349 => x"9c",
          4350 => x"33",
          4351 => x"86",
          4352 => x"80",
          4353 => x"16",
          4354 => x"33",
          4355 => x"70",
          4356 => x"5a",
          4357 => x"72",
          4358 => x"74",
          4359 => x"70",
          4360 => x"32",
          4361 => x"73",
          4362 => x"53",
          4363 => x"54",
          4364 => x"9b",
          4365 => x"2e",
          4366 => x"77",
          4367 => x"54",
          4368 => x"09",
          4369 => x"38",
          4370 => x"7a",
          4371 => x"80",
          4372 => x"fa",
          4373 => x"93",
          4374 => x"82",
          4375 => x"87",
          4376 => x"08",
          4377 => x"77",
          4378 => x"38",
          4379 => x"17",
          4380 => x"93",
          4381 => x"3d",
          4382 => x"3d",
          4383 => x"08",
          4384 => x"52",
          4385 => x"f2",
          4386 => x"c8",
          4387 => x"93",
          4388 => x"ef",
          4389 => x"84",
          4390 => x"39",
          4391 => x"52",
          4392 => x"a5",
          4393 => x"c8",
          4394 => x"93",
          4395 => x"d1",
          4396 => x"08",
          4397 => x"54",
          4398 => x"db",
          4399 => x"08",
          4400 => x"bf",
          4401 => x"73",
          4402 => x"8b",
          4403 => x"83",
          4404 => x"06",
          4405 => x"73",
          4406 => x"53",
          4407 => x"74",
          4408 => x"3f",
          4409 => x"08",
          4410 => x"38",
          4411 => x"51",
          4412 => x"82",
          4413 => x"57",
          4414 => x"08",
          4415 => x"9c",
          4416 => x"73",
          4417 => x"0c",
          4418 => x"04",
          4419 => x"77",
          4420 => x"54",
          4421 => x"51",
          4422 => x"82",
          4423 => x"55",
          4424 => x"08",
          4425 => x"14",
          4426 => x"51",
          4427 => x"82",
          4428 => x"55",
          4429 => x"08",
          4430 => x"53",
          4431 => x"08",
          4432 => x"08",
          4433 => x"3f",
          4434 => x"14",
          4435 => x"08",
          4436 => x"3f",
          4437 => x"17",
          4438 => x"93",
          4439 => x"3d",
          4440 => x"3d",
          4441 => x"08",
          4442 => x"54",
          4443 => x"53",
          4444 => x"82",
          4445 => x"54",
          4446 => x"08",
          4447 => x"13",
          4448 => x"73",
          4449 => x"83",
          4450 => x"82",
          4451 => x"86",
          4452 => x"fa",
          4453 => x"7a",
          4454 => x"0b",
          4455 => x"98",
          4456 => x"2e",
          4457 => x"80",
          4458 => x"9c",
          4459 => x"70",
          4460 => x"56",
          4461 => x"a0",
          4462 => x"72",
          4463 => x"81",
          4464 => x"81",
          4465 => x"89",
          4466 => x"06",
          4467 => x"15",
          4468 => x"ae",
          4469 => x"34",
          4470 => x"75",
          4471 => x"52",
          4472 => x"34",
          4473 => x"8a",
          4474 => x"38",
          4475 => x"05",
          4476 => x"81",
          4477 => x"17",
          4478 => x"12",
          4479 => x"34",
          4480 => x"9c",
          4481 => x"ac",
          4482 => x"c8",
          4483 => x"9c",
          4484 => x"05",
          4485 => x"3f",
          4486 => x"08",
          4487 => x"9c",
          4488 => x"05",
          4489 => x"3f",
          4490 => x"08",
          4491 => x"88",
          4492 => x"f5",
          4493 => x"70",
          4494 => x"05",
          4495 => x"8b",
          4496 => x"7a",
          4497 => x"3f",
          4498 => x"58",
          4499 => x"55",
          4500 => x"2e",
          4501 => x"80",
          4502 => x"17",
          4503 => x"19",
          4504 => x"70",
          4505 => x"2a",
          4506 => x"07",
          4507 => x"59",
          4508 => x"8c",
          4509 => x"54",
          4510 => x"81",
          4511 => x"39",
          4512 => x"70",
          4513 => x"dc",
          4514 => x"70",
          4515 => x"2a",
          4516 => x"51",
          4517 => x"2e",
          4518 => x"54",
          4519 => x"82",
          4520 => x"19",
          4521 => x"54",
          4522 => x"83",
          4523 => x"73",
          4524 => x"80",
          4525 => x"39",
          4526 => x"33",
          4527 => x"57",
          4528 => x"27",
          4529 => x"75",
          4530 => x"30",
          4531 => x"32",
          4532 => x"80",
          4533 => x"25",
          4534 => x"56",
          4535 => x"80",
          4536 => x"84",
          4537 => x"57",
          4538 => x"70",
          4539 => x"5a",
          4540 => x"09",
          4541 => x"38",
          4542 => x"77",
          4543 => x"51",
          4544 => x"80",
          4545 => x"81",
          4546 => x"81",
          4547 => x"07",
          4548 => x"38",
          4549 => x"75",
          4550 => x"30",
          4551 => x"7a",
          4552 => x"51",
          4553 => x"80",
          4554 => x"79",
          4555 => x"30",
          4556 => x"70",
          4557 => x"25",
          4558 => x"07",
          4559 => x"51",
          4560 => x"b1",
          4561 => x"8b",
          4562 => x"39",
          4563 => x"54",
          4564 => x"8c",
          4565 => x"ff",
          4566 => x"f8",
          4567 => x"54",
          4568 => x"e6",
          4569 => x"c8",
          4570 => x"b9",
          4571 => x"70",
          4572 => x"71",
          4573 => x"54",
          4574 => x"82",
          4575 => x"80",
          4576 => x"ff",
          4577 => x"78",
          4578 => x"86",
          4579 => x"39",
          4580 => x"75",
          4581 => x"18",
          4582 => x"58",
          4583 => x"81",
          4584 => x"94",
          4585 => x"81",
          4586 => x"e4",
          4587 => x"93",
          4588 => x"c5",
          4589 => x"16",
          4590 => x"26",
          4591 => x"16",
          4592 => x"06",
          4593 => x"18",
          4594 => x"34",
          4595 => x"fd",
          4596 => x"19",
          4597 => x"54",
          4598 => x"a9",
          4599 => x"54",
          4600 => x"2e",
          4601 => x"84",
          4602 => x"34",
          4603 => x"76",
          4604 => x"89",
          4605 => x"8d",
          4606 => x"89",
          4607 => x"73",
          4608 => x"80",
          4609 => x"93",
          4610 => x"3d",
          4611 => x"3d",
          4612 => x"08",
          4613 => x"7a",
          4614 => x"54",
          4615 => x"2e",
          4616 => x"55",
          4617 => x"33",
          4618 => x"72",
          4619 => x"83",
          4620 => x"74",
          4621 => x"72",
          4622 => x"38",
          4623 => x"88",
          4624 => x"39",
          4625 => x"80",
          4626 => x"51",
          4627 => x"af",
          4628 => x"06",
          4629 => x"55",
          4630 => x"33",
          4631 => x"72",
          4632 => x"09",
          4633 => x"38",
          4634 => x"74",
          4635 => x"d4",
          4636 => x"88",
          4637 => x"70",
          4638 => x"72",
          4639 => x"38",
          4640 => x"ab",
          4641 => x"52",
          4642 => x"ee",
          4643 => x"c8",
          4644 => x"aa",
          4645 => x"81",
          4646 => x"3d",
          4647 => x"75",
          4648 => x"3f",
          4649 => x"08",
          4650 => x"c8",
          4651 => x"38",
          4652 => x"c6",
          4653 => x"c8",
          4654 => x"33",
          4655 => x"93",
          4656 => x"2e",
          4657 => x"82",
          4658 => x"84",
          4659 => x"06",
          4660 => x"73",
          4661 => x"81",
          4662 => x"72",
          4663 => x"38",
          4664 => x"70",
          4665 => x"53",
          4666 => x"ff",
          4667 => x"80",
          4668 => x"34",
          4669 => x"c6",
          4670 => x"2a",
          4671 => x"51",
          4672 => x"38",
          4673 => x"39",
          4674 => x"70",
          4675 => x"53",
          4676 => x"86",
          4677 => x"84",
          4678 => x"06",
          4679 => x"72",
          4680 => x"f1",
          4681 => x"08",
          4682 => x"17",
          4683 => x"76",
          4684 => x"3f",
          4685 => x"08",
          4686 => x"fe",
          4687 => x"82",
          4688 => x"88",
          4689 => x"f6",
          4690 => x"59",
          4691 => x"70",
          4692 => x"56",
          4693 => x"2e",
          4694 => x"76",
          4695 => x"58",
          4696 => x"32",
          4697 => x"a0",
          4698 => x"2a",
          4699 => x"52",
          4700 => x"38",
          4701 => x"09",
          4702 => x"a9",
          4703 => x"d0",
          4704 => x"70",
          4705 => x"38",
          4706 => x"81",
          4707 => x"11",
          4708 => x"70",
          4709 => x"ff",
          4710 => x"81",
          4711 => x"58",
          4712 => x"1b",
          4713 => x"08",
          4714 => x"75",
          4715 => x"57",
          4716 => x"81",
          4717 => x"ff",
          4718 => x"54",
          4719 => x"26",
          4720 => x"14",
          4721 => x"06",
          4722 => x"9f",
          4723 => x"99",
          4724 => x"e0",
          4725 => x"ff",
          4726 => x"73",
          4727 => x"32",
          4728 => x"72",
          4729 => x"73",
          4730 => x"53",
          4731 => x"70",
          4732 => x"73",
          4733 => x"32",
          4734 => x"72",
          4735 => x"73",
          4736 => x"53",
          4737 => x"70",
          4738 => x"38",
          4739 => x"83",
          4740 => x"8c",
          4741 => x"77",
          4742 => x"38",
          4743 => x"0c",
          4744 => x"86",
          4745 => x"f8",
          4746 => x"82",
          4747 => x"8c",
          4748 => x"fb",
          4749 => x"56",
          4750 => x"17",
          4751 => x"b0",
          4752 => x"52",
          4753 => x"81",
          4754 => x"82",
          4755 => x"81",
          4756 => x"b2",
          4757 => x"c3",
          4758 => x"c8",
          4759 => x"ff",
          4760 => x"55",
          4761 => x"d5",
          4762 => x"06",
          4763 => x"80",
          4764 => x"33",
          4765 => x"81",
          4766 => x"81",
          4767 => x"81",
          4768 => x"eb",
          4769 => x"70",
          4770 => x"07",
          4771 => x"73",
          4772 => x"16",
          4773 => x"81",
          4774 => x"81",
          4775 => x"83",
          4776 => x"80",
          4777 => x"16",
          4778 => x"3f",
          4779 => x"08",
          4780 => x"c8",
          4781 => x"9d",
          4782 => x"81",
          4783 => x"81",
          4784 => x"de",
          4785 => x"93",
          4786 => x"82",
          4787 => x"80",
          4788 => x"82",
          4789 => x"93",
          4790 => x"3d",
          4791 => x"3d",
          4792 => x"84",
          4793 => x"05",
          4794 => x"80",
          4795 => x"51",
          4796 => x"82",
          4797 => x"58",
          4798 => x"0b",
          4799 => x"08",
          4800 => x"38",
          4801 => x"08",
          4802 => x"93",
          4803 => x"08",
          4804 => x"56",
          4805 => x"87",
          4806 => x"74",
          4807 => x"fe",
          4808 => x"54",
          4809 => x"2e",
          4810 => x"15",
          4811 => x"a6",
          4812 => x"c8",
          4813 => x"06",
          4814 => x"54",
          4815 => x"38",
          4816 => x"8f",
          4817 => x"2a",
          4818 => x"51",
          4819 => x"72",
          4820 => x"80",
          4821 => x"39",
          4822 => x"77",
          4823 => x"81",
          4824 => x"33",
          4825 => x"3f",
          4826 => x"08",
          4827 => x"70",
          4828 => x"54",
          4829 => x"86",
          4830 => x"80",
          4831 => x"73",
          4832 => x"81",
          4833 => x"8a",
          4834 => x"95",
          4835 => x"53",
          4836 => x"fd",
          4837 => x"93",
          4838 => x"ff",
          4839 => x"82",
          4840 => x"06",
          4841 => x"79",
          4842 => x"29",
          4843 => x"75",
          4844 => x"f0",
          4845 => x"12",
          4846 => x"56",
          4847 => x"77",
          4848 => x"83",
          4849 => x"da",
          4850 => x"93",
          4851 => x"76",
          4852 => x"14",
          4853 => x"27",
          4854 => x"54",
          4855 => x"10",
          4856 => x"11",
          4857 => x"83",
          4858 => x"2e",
          4859 => x"52",
          4860 => x"bf",
          4861 => x"c8",
          4862 => x"06",
          4863 => x"27",
          4864 => x"14",
          4865 => x"27",
          4866 => x"56",
          4867 => x"85",
          4868 => x"56",
          4869 => x"85",
          4870 => x"15",
          4871 => x"3f",
          4872 => x"08",
          4873 => x"06",
          4874 => x"72",
          4875 => x"09",
          4876 => x"ed",
          4877 => x"15",
          4878 => x"3f",
          4879 => x"08",
          4880 => x"06",
          4881 => x"38",
          4882 => x"51",
          4883 => x"82",
          4884 => x"54",
          4885 => x"0c",
          4886 => x"33",
          4887 => x"80",
          4888 => x"ff",
          4889 => x"56",
          4890 => x"84",
          4891 => x"15",
          4892 => x"29",
          4893 => x"33",
          4894 => x"72",
          4895 => x"72",
          4896 => x"06",
          4897 => x"2e",
          4898 => x"13",
          4899 => x"72",
          4900 => x"38",
          4901 => x"89",
          4902 => x"15",
          4903 => x"3f",
          4904 => x"08",
          4905 => x"82",
          4906 => x"83",
          4907 => x"8f",
          4908 => x"56",
          4909 => x"38",
          4910 => x"51",
          4911 => x"82",
          4912 => x"83",
          4913 => x"53",
          4914 => x"80",
          4915 => x"d8",
          4916 => x"93",
          4917 => x"80",
          4918 => x"d8",
          4919 => x"93",
          4920 => x"ff",
          4921 => x"8d",
          4922 => x"2e",
          4923 => x"88",
          4924 => x"1a",
          4925 => x"05",
          4926 => x"56",
          4927 => x"83",
          4928 => x"15",
          4929 => x"78",
          4930 => x"b0",
          4931 => x"93",
          4932 => x"8d",
          4933 => x"c8",
          4934 => x"83",
          4935 => x"57",
          4936 => x"08",
          4937 => x"ff",
          4938 => x"38",
          4939 => x"83",
          4940 => x"83",
          4941 => x"72",
          4942 => x"83",
          4943 => x"8d",
          4944 => x"2e",
          4945 => x"82",
          4946 => x"0c",
          4947 => x"0c",
          4948 => x"16",
          4949 => x"ac",
          4950 => x"83",
          4951 => x"06",
          4952 => x"de",
          4953 => x"b3",
          4954 => x"c8",
          4955 => x"ff",
          4956 => x"56",
          4957 => x"38",
          4958 => x"53",
          4959 => x"82",
          4960 => x"e0",
          4961 => x"ac",
          4962 => x"c8",
          4963 => x"0c",
          4964 => x"82",
          4965 => x"39",
          4966 => x"53",
          4967 => x"80",
          4968 => x"38",
          4969 => x"14",
          4970 => x"76",
          4971 => x"81",
          4972 => x"98",
          4973 => x"53",
          4974 => x"15",
          4975 => x"16",
          4976 => x"81",
          4977 => x"08",
          4978 => x"51",
          4979 => x"13",
          4980 => x"8d",
          4981 => x"16",
          4982 => x"c5",
          4983 => x"90",
          4984 => x"0b",
          4985 => x"ff",
          4986 => x"16",
          4987 => x"2e",
          4988 => x"81",
          4989 => x"e4",
          4990 => x"9f",
          4991 => x"c8",
          4992 => x"ff",
          4993 => x"81",
          4994 => x"06",
          4995 => x"81",
          4996 => x"51",
          4997 => x"82",
          4998 => x"80",
          4999 => x"93",
          5000 => x"16",
          5001 => x"15",
          5002 => x"3f",
          5003 => x"08",
          5004 => x"06",
          5005 => x"d4",
          5006 => x"81",
          5007 => x"38",
          5008 => x"d5",
          5009 => x"93",
          5010 => x"8b",
          5011 => x"2e",
          5012 => x"b3",
          5013 => x"15",
          5014 => x"3f",
          5015 => x"08",
          5016 => x"e4",
          5017 => x"81",
          5018 => x"84",
          5019 => x"d5",
          5020 => x"93",
          5021 => x"16",
          5022 => x"15",
          5023 => x"3f",
          5024 => x"08",
          5025 => x"76",
          5026 => x"93",
          5027 => x"05",
          5028 => x"93",
          5029 => x"86",
          5030 => x"0b",
          5031 => x"80",
          5032 => x"93",
          5033 => x"3d",
          5034 => x"3d",
          5035 => x"89",
          5036 => x"2e",
          5037 => x"08",
          5038 => x"38",
          5039 => x"33",
          5040 => x"80",
          5041 => x"84",
          5042 => x"14",
          5043 => x"71",
          5044 => x"81",
          5045 => x"81",
          5046 => x"ce",
          5047 => x"93",
          5048 => x"06",
          5049 => x"38",
          5050 => x"53",
          5051 => x"09",
          5052 => x"38",
          5053 => x"78",
          5054 => x"52",
          5055 => x"c8",
          5056 => x"0d",
          5057 => x"0d",
          5058 => x"33",
          5059 => x"3d",
          5060 => x"56",
          5061 => x"82",
          5062 => x"55",
          5063 => x"0b",
          5064 => x"08",
          5065 => x"38",
          5066 => x"08",
          5067 => x"93",
          5068 => x"08",
          5069 => x"80",
          5070 => x"80",
          5071 => x"80",
          5072 => x"78",
          5073 => x"34",
          5074 => x"82",
          5075 => x"79",
          5076 => x"75",
          5077 => x"2e",
          5078 => x"53",
          5079 => x"53",
          5080 => x"f6",
          5081 => x"93",
          5082 => x"73",
          5083 => x"0c",
          5084 => x"04",
          5085 => x"67",
          5086 => x"80",
          5087 => x"58",
          5088 => x"77",
          5089 => x"e9",
          5090 => x"06",
          5091 => x"3d",
          5092 => x"99",
          5093 => x"52",
          5094 => x"3f",
          5095 => x"08",
          5096 => x"c8",
          5097 => x"38",
          5098 => x"52",
          5099 => x"05",
          5100 => x"3f",
          5101 => x"08",
          5102 => x"c8",
          5103 => x"02",
          5104 => x"33",
          5105 => x"56",
          5106 => x"25",
          5107 => x"56",
          5108 => x"55",
          5109 => x"81",
          5110 => x"80",
          5111 => x"75",
          5112 => x"81",
          5113 => x"97",
          5114 => x"51",
          5115 => x"82",
          5116 => x"56",
          5117 => x"57",
          5118 => x"b2",
          5119 => x"06",
          5120 => x"2e",
          5121 => x"56",
          5122 => x"82",
          5123 => x"06",
          5124 => x"80",
          5125 => x"88",
          5126 => x"d0",
          5127 => x"2a",
          5128 => x"51",
          5129 => x"2e",
          5130 => x"62",
          5131 => x"e6",
          5132 => x"93",
          5133 => x"82",
          5134 => x"52",
          5135 => x"51",
          5136 => x"62",
          5137 => x"8b",
          5138 => x"53",
          5139 => x"51",
          5140 => x"75",
          5141 => x"05",
          5142 => x"3f",
          5143 => x"0b",
          5144 => x"78",
          5145 => x"e9",
          5146 => x"11",
          5147 => x"7a",
          5148 => x"d4",
          5149 => x"55",
          5150 => x"82",
          5151 => x"56",
          5152 => x"08",
          5153 => x"74",
          5154 => x"d4",
          5155 => x"93",
          5156 => x"ff",
          5157 => x"0c",
          5158 => x"39",
          5159 => x"38",
          5160 => x"33",
          5161 => x"70",
          5162 => x"56",
          5163 => x"2e",
          5164 => x"56",
          5165 => x"81",
          5166 => x"06",
          5167 => x"80",
          5168 => x"02",
          5169 => x"81",
          5170 => x"80",
          5171 => x"87",
          5172 => x"98",
          5173 => x"2a",
          5174 => x"51",
          5175 => x"2e",
          5176 => x"80",
          5177 => x"7a",
          5178 => x"a0",
          5179 => x"a4",
          5180 => x"75",
          5181 => x"62",
          5182 => x"e4",
          5183 => x"93",
          5184 => x"19",
          5185 => x"05",
          5186 => x"3f",
          5187 => x"08",
          5188 => x"74",
          5189 => x"15",
          5190 => x"23",
          5191 => x"34",
          5192 => x"34",
          5193 => x"0c",
          5194 => x"0c",
          5195 => x"75",
          5196 => x"51",
          5197 => x"76",
          5198 => x"81",
          5199 => x"74",
          5200 => x"a3",
          5201 => x"08",
          5202 => x"9b",
          5203 => x"08",
          5204 => x"7a",
          5205 => x"70",
          5206 => x"1b",
          5207 => x"08",
          5208 => x"51",
          5209 => x"76",
          5210 => x"d4",
          5211 => x"93",
          5212 => x"82",
          5213 => x"81",
          5214 => x"82",
          5215 => x"2e",
          5216 => x"83",
          5217 => x"78",
          5218 => x"75",
          5219 => x"07",
          5220 => x"7b",
          5221 => x"51",
          5222 => x"cb",
          5223 => x"19",
          5224 => x"c8",
          5225 => x"ff",
          5226 => x"80",
          5227 => x"76",
          5228 => x"d4",
          5229 => x"93",
          5230 => x"38",
          5231 => x"39",
          5232 => x"82",
          5233 => x"05",
          5234 => x"0c",
          5235 => x"74",
          5236 => x"52",
          5237 => x"33",
          5238 => x"a4",
          5239 => x"c8",
          5240 => x"83",
          5241 => x"75",
          5242 => x"38",
          5243 => x"75",
          5244 => x"93",
          5245 => x"3d",
          5246 => x"3d",
          5247 => x"64",
          5248 => x"5a",
          5249 => x"0c",
          5250 => x"05",
          5251 => x"f9",
          5252 => x"93",
          5253 => x"82",
          5254 => x"8a",
          5255 => x"33",
          5256 => x"2e",
          5257 => x"56",
          5258 => x"90",
          5259 => x"06",
          5260 => x"74",
          5261 => x"a0",
          5262 => x"82",
          5263 => x"34",
          5264 => x"94",
          5265 => x"91",
          5266 => x"56",
          5267 => x"82",
          5268 => x"34",
          5269 => x"80",
          5270 => x"91",
          5271 => x"56",
          5272 => x"81",
          5273 => x"34",
          5274 => x"ec",
          5275 => x"91",
          5276 => x"56",
          5277 => x"8c",
          5278 => x"18",
          5279 => x"74",
          5280 => x"38",
          5281 => x"80",
          5282 => x"38",
          5283 => x"70",
          5284 => x"56",
          5285 => x"83",
          5286 => x"11",
          5287 => x"77",
          5288 => x"5c",
          5289 => x"38",
          5290 => x"88",
          5291 => x"8f",
          5292 => x"08",
          5293 => x"d2",
          5294 => x"93",
          5295 => x"81",
          5296 => x"f7",
          5297 => x"2e",
          5298 => x"74",
          5299 => x"98",
          5300 => x"7d",
          5301 => x"3f",
          5302 => x"08",
          5303 => x"ef",
          5304 => x"c8",
          5305 => x"89",
          5306 => x"79",
          5307 => x"d7",
          5308 => x"7e",
          5309 => x"51",
          5310 => x"76",
          5311 => x"74",
          5312 => x"79",
          5313 => x"7b",
          5314 => x"11",
          5315 => x"c7",
          5316 => x"93",
          5317 => x"c1",
          5318 => x"33",
          5319 => x"56",
          5320 => x"25",
          5321 => x"17",
          5322 => x"55",
          5323 => x"90",
          5324 => x"53",
          5325 => x"74",
          5326 => x"1c",
          5327 => x"3f",
          5328 => x"56",
          5329 => x"9c",
          5330 => x"2e",
          5331 => x"90",
          5332 => x"98",
          5333 => x"74",
          5334 => x"38",
          5335 => x"17",
          5336 => x"17",
          5337 => x"11",
          5338 => x"c8",
          5339 => x"93",
          5340 => x"ef",
          5341 => x"33",
          5342 => x"55",
          5343 => x"34",
          5344 => x"53",
          5345 => x"7d",
          5346 => x"52",
          5347 => x"3f",
          5348 => x"08",
          5349 => x"77",
          5350 => x"94",
          5351 => x"ff",
          5352 => x"71",
          5353 => x"78",
          5354 => x"38",
          5355 => x"53",
          5356 => x"83",
          5357 => x"a8",
          5358 => x"51",
          5359 => x"78",
          5360 => x"08",
          5361 => x"76",
          5362 => x"08",
          5363 => x"0c",
          5364 => x"fd",
          5365 => x"56",
          5366 => x"c8",
          5367 => x"0d",
          5368 => x"0d",
          5369 => x"63",
          5370 => x"57",
          5371 => x"8f",
          5372 => x"52",
          5373 => x"b2",
          5374 => x"c8",
          5375 => x"93",
          5376 => x"38",
          5377 => x"55",
          5378 => x"86",
          5379 => x"84",
          5380 => x"17",
          5381 => x"2a",
          5382 => x"51",
          5383 => x"56",
          5384 => x"83",
          5385 => x"39",
          5386 => x"18",
          5387 => x"83",
          5388 => x"0b",
          5389 => x"81",
          5390 => x"39",
          5391 => x"18",
          5392 => x"83",
          5393 => x"0b",
          5394 => x"82",
          5395 => x"39",
          5396 => x"18",
          5397 => x"83",
          5398 => x"0b",
          5399 => x"81",
          5400 => x"39",
          5401 => x"19",
          5402 => x"18",
          5403 => x"38",
          5404 => x"09",
          5405 => x"2e",
          5406 => x"94",
          5407 => x"83",
          5408 => x"56",
          5409 => x"38",
          5410 => x"22",
          5411 => x"89",
          5412 => x"55",
          5413 => x"38",
          5414 => x"88",
          5415 => x"74",
          5416 => x"52",
          5417 => x"b8",
          5418 => x"c8",
          5419 => x"39",
          5420 => x"52",
          5421 => x"a8",
          5422 => x"c8",
          5423 => x"80",
          5424 => x"38",
          5425 => x"fe",
          5426 => x"ff",
          5427 => x"38",
          5428 => x"0c",
          5429 => x"85",
          5430 => x"18",
          5431 => x"33",
          5432 => x"56",
          5433 => x"25",
          5434 => x"54",
          5435 => x"53",
          5436 => x"7d",
          5437 => x"52",
          5438 => x"3f",
          5439 => x"08",
          5440 => x"90",
          5441 => x"ff",
          5442 => x"90",
          5443 => x"17",
          5444 => x"51",
          5445 => x"82",
          5446 => x"80",
          5447 => x"38",
          5448 => x"08",
          5449 => x"2a",
          5450 => x"80",
          5451 => x"38",
          5452 => x"8a",
          5453 => x"56",
          5454 => x"27",
          5455 => x"7b",
          5456 => x"54",
          5457 => x"52",
          5458 => x"33",
          5459 => x"89",
          5460 => x"c8",
          5461 => x"38",
          5462 => x"78",
          5463 => x"7a",
          5464 => x"84",
          5465 => x"84",
          5466 => x"52",
          5467 => x"c8",
          5468 => x"17",
          5469 => x"06",
          5470 => x"18",
          5471 => x"2b",
          5472 => x"39",
          5473 => x"78",
          5474 => x"94",
          5475 => x"18",
          5476 => x"38",
          5477 => x"53",
          5478 => x"7d",
          5479 => x"52",
          5480 => x"3f",
          5481 => x"08",
          5482 => x"77",
          5483 => x"94",
          5484 => x"ff",
          5485 => x"71",
          5486 => x"78",
          5487 => x"38",
          5488 => x"53",
          5489 => x"17",
          5490 => x"06",
          5491 => x"51",
          5492 => x"90",
          5493 => x"80",
          5494 => x"90",
          5495 => x"76",
          5496 => x"17",
          5497 => x"1d",
          5498 => x"18",
          5499 => x"0c",
          5500 => x"58",
          5501 => x"74",
          5502 => x"38",
          5503 => x"8c",
          5504 => x"fc",
          5505 => x"17",
          5506 => x"07",
          5507 => x"18",
          5508 => x"75",
          5509 => x"0c",
          5510 => x"04",
          5511 => x"7b",
          5512 => x"05",
          5513 => x"58",
          5514 => x"82",
          5515 => x"57",
          5516 => x"08",
          5517 => x"90",
          5518 => x"86",
          5519 => x"06",
          5520 => x"74",
          5521 => x"98",
          5522 => x"2b",
          5523 => x"25",
          5524 => x"54",
          5525 => x"53",
          5526 => x"79",
          5527 => x"52",
          5528 => x"3f",
          5529 => x"93",
          5530 => x"f6",
          5531 => x"33",
          5532 => x"55",
          5533 => x"34",
          5534 => x"52",
          5535 => x"c9",
          5536 => x"c8",
          5537 => x"93",
          5538 => x"d4",
          5539 => x"08",
          5540 => x"a0",
          5541 => x"74",
          5542 => x"88",
          5543 => x"75",
          5544 => x"51",
          5545 => x"8c",
          5546 => x"9c",
          5547 => x"cb",
          5548 => x"b2",
          5549 => x"16",
          5550 => x"3f",
          5551 => x"16",
          5552 => x"3f",
          5553 => x"0b",
          5554 => x"79",
          5555 => x"3f",
          5556 => x"08",
          5557 => x"81",
          5558 => x"57",
          5559 => x"34",
          5560 => x"82",
          5561 => x"8b",
          5562 => x"fc",
          5563 => x"70",
          5564 => x"a8",
          5565 => x"c8",
          5566 => x"93",
          5567 => x"38",
          5568 => x"05",
          5569 => x"ef",
          5570 => x"93",
          5571 => x"82",
          5572 => x"87",
          5573 => x"c8",
          5574 => x"72",
          5575 => x"0c",
          5576 => x"04",
          5577 => x"85",
          5578 => x"9b",
          5579 => x"80",
          5580 => x"c8",
          5581 => x"38",
          5582 => x"08",
          5583 => x"34",
          5584 => x"82",
          5585 => x"84",
          5586 => x"ef",
          5587 => x"53",
          5588 => x"05",
          5589 => x"51",
          5590 => x"82",
          5591 => x"55",
          5592 => x"08",
          5593 => x"76",
          5594 => x"93",
          5595 => x"51",
          5596 => x"82",
          5597 => x"55",
          5598 => x"08",
          5599 => x"80",
          5600 => x"70",
          5601 => x"56",
          5602 => x"89",
          5603 => x"94",
          5604 => x"a7",
          5605 => x"05",
          5606 => x"2a",
          5607 => x"51",
          5608 => x"80",
          5609 => x"76",
          5610 => x"52",
          5611 => x"3f",
          5612 => x"08",
          5613 => x"83",
          5614 => x"74",
          5615 => x"81",
          5616 => x"85",
          5617 => x"93",
          5618 => x"3d",
          5619 => x"3d",
          5620 => x"08",
          5621 => x"5b",
          5622 => x"34",
          5623 => x"3d",
          5624 => x"52",
          5625 => x"e5",
          5626 => x"93",
          5627 => x"82",
          5628 => x"83",
          5629 => x"46",
          5630 => x"11",
          5631 => x"68",
          5632 => x"80",
          5633 => x"38",
          5634 => x"94",
          5635 => x"5b",
          5636 => x"51",
          5637 => x"82",
          5638 => x"57",
          5639 => x"08",
          5640 => x"6b",
          5641 => x"c5",
          5642 => x"93",
          5643 => x"82",
          5644 => x"81",
          5645 => x"52",
          5646 => x"ab",
          5647 => x"c8",
          5648 => x"52",
          5649 => x"b2",
          5650 => x"c8",
          5651 => x"93",
          5652 => x"ac",
          5653 => x"80",
          5654 => x"d6",
          5655 => x"93",
          5656 => x"82",
          5657 => x"a4",
          5658 => x"7e",
          5659 => x"3f",
          5660 => x"08",
          5661 => x"38",
          5662 => x"51",
          5663 => x"82",
          5664 => x"57",
          5665 => x"08",
          5666 => x"38",
          5667 => x"09",
          5668 => x"38",
          5669 => x"81",
          5670 => x"3d",
          5671 => x"53",
          5672 => x"d9",
          5673 => x"93",
          5674 => x"12",
          5675 => x"51",
          5676 => x"56",
          5677 => x"8e",
          5678 => x"70",
          5679 => x"33",
          5680 => x"73",
          5681 => x"16",
          5682 => x"27",
          5683 => x"57",
          5684 => x"80",
          5685 => x"7d",
          5686 => x"a3",
          5687 => x"ff",
          5688 => x"57",
          5689 => x"81",
          5690 => x"34",
          5691 => x"ff",
          5692 => x"08",
          5693 => x"af",
          5694 => x"55",
          5695 => x"38",
          5696 => x"38",
          5697 => x"09",
          5698 => x"38",
          5699 => x"3d",
          5700 => x"59",
          5701 => x"80",
          5702 => x"f8",
          5703 => x"10",
          5704 => x"05",
          5705 => x"33",
          5706 => x"57",
          5707 => x"78",
          5708 => x"81",
          5709 => x"70",
          5710 => x"56",
          5711 => x"82",
          5712 => x"79",
          5713 => x"80",
          5714 => x"27",
          5715 => x"15",
          5716 => x"7a",
          5717 => x"5c",
          5718 => x"58",
          5719 => x"ee",
          5720 => x"70",
          5721 => x"34",
          5722 => x"77",
          5723 => x"57",
          5724 => x"a2",
          5725 => x"81",
          5726 => x"73",
          5727 => x"81",
          5728 => x"7b",
          5729 => x"38",
          5730 => x"76",
          5731 => x"0c",
          5732 => x"04",
          5733 => x"7e",
          5734 => x"fc",
          5735 => x"53",
          5736 => x"86",
          5737 => x"c8",
          5738 => x"93",
          5739 => x"38",
          5740 => x"5a",
          5741 => x"86",
          5742 => x"83",
          5743 => x"17",
          5744 => x"94",
          5745 => x"33",
          5746 => x"70",
          5747 => x"56",
          5748 => x"38",
          5749 => x"58",
          5750 => x"56",
          5751 => x"19",
          5752 => x"7b",
          5753 => x"38",
          5754 => x"22",
          5755 => x"5b",
          5756 => x"7b",
          5757 => x"78",
          5758 => x"51",
          5759 => x"3f",
          5760 => x"08",
          5761 => x"54",
          5762 => x"55",
          5763 => x"3f",
          5764 => x"08",
          5765 => x"38",
          5766 => x"06",
          5767 => x"77",
          5768 => x"31",
          5769 => x"57",
          5770 => x"39",
          5771 => x"56",
          5772 => x"75",
          5773 => x"c9",
          5774 => x"93",
          5775 => x"82",
          5776 => x"81",
          5777 => x"06",
          5778 => x"0b",
          5779 => x"82",
          5780 => x"39",
          5781 => x"08",
          5782 => x"81",
          5783 => x"81",
          5784 => x"34",
          5785 => x"ce",
          5786 => x"c8",
          5787 => x"0c",
          5788 => x"0c",
          5789 => x"81",
          5790 => x"78",
          5791 => x"38",
          5792 => x"94",
          5793 => x"94",
          5794 => x"18",
          5795 => x"2a",
          5796 => x"51",
          5797 => x"74",
          5798 => x"38",
          5799 => x"51",
          5800 => x"82",
          5801 => x"56",
          5802 => x"08",
          5803 => x"93",
          5804 => x"b5",
          5805 => x"76",
          5806 => x"3f",
          5807 => x"08",
          5808 => x"2e",
          5809 => x"81",
          5810 => x"38",
          5811 => x"15",
          5812 => x"8b",
          5813 => x"91",
          5814 => x"55",
          5815 => x"75",
          5816 => x"77",
          5817 => x"98",
          5818 => x"08",
          5819 => x"0c",
          5820 => x"06",
          5821 => x"2e",
          5822 => x"52",
          5823 => x"bf",
          5824 => x"c8",
          5825 => x"82",
          5826 => x"34",
          5827 => x"a6",
          5828 => x"2a",
          5829 => x"08",
          5830 => x"17",
          5831 => x"08",
          5832 => x"94",
          5833 => x"18",
          5834 => x"33",
          5835 => x"55",
          5836 => x"34",
          5837 => x"83",
          5838 => x"74",
          5839 => x"f4",
          5840 => x"08",
          5841 => x"ec",
          5842 => x"33",
          5843 => x"56",
          5844 => x"25",
          5845 => x"54",
          5846 => x"53",
          5847 => x"7c",
          5848 => x"52",
          5849 => x"f1",
          5850 => x"c8",
          5851 => x"8a",
          5852 => x"91",
          5853 => x"55",
          5854 => x"17",
          5855 => x"06",
          5856 => x"18",
          5857 => x"7a",
          5858 => x"52",
          5859 => x"33",
          5860 => x"b6",
          5861 => x"93",
          5862 => x"2e",
          5863 => x"0b",
          5864 => x"81",
          5865 => x"81",
          5866 => x"34",
          5867 => x"39",
          5868 => x"0c",
          5869 => x"82",
          5870 => x"8e",
          5871 => x"f9",
          5872 => x"56",
          5873 => x"80",
          5874 => x"38",
          5875 => x"3d",
          5876 => x"8a",
          5877 => x"51",
          5878 => x"82",
          5879 => x"55",
          5880 => x"08",
          5881 => x"77",
          5882 => x"52",
          5883 => x"9e",
          5884 => x"c8",
          5885 => x"93",
          5886 => x"ca",
          5887 => x"33",
          5888 => x"55",
          5889 => x"24",
          5890 => x"16",
          5891 => x"2a",
          5892 => x"51",
          5893 => x"80",
          5894 => x"9c",
          5895 => x"77",
          5896 => x"3f",
          5897 => x"08",
          5898 => x"83",
          5899 => x"74",
          5900 => x"54",
          5901 => x"84",
          5902 => x"52",
          5903 => x"ba",
          5904 => x"c8",
          5905 => x"84",
          5906 => x"06",
          5907 => x"55",
          5908 => x"84",
          5909 => x"0c",
          5910 => x"82",
          5911 => x"89",
          5912 => x"fc",
          5913 => x"87",
          5914 => x"53",
          5915 => x"e4",
          5916 => x"93",
          5917 => x"82",
          5918 => x"87",
          5919 => x"c8",
          5920 => x"72",
          5921 => x"0c",
          5922 => x"04",
          5923 => x"77",
          5924 => x"fc",
          5925 => x"53",
          5926 => x"8e",
          5927 => x"c8",
          5928 => x"93",
          5929 => x"d1",
          5930 => x"38",
          5931 => x"08",
          5932 => x"c8",
          5933 => x"93",
          5934 => x"bd",
          5935 => x"73",
          5936 => x"3f",
          5937 => x"08",
          5938 => x"c8",
          5939 => x"09",
          5940 => x"38",
          5941 => x"a1",
          5942 => x"73",
          5943 => x"3f",
          5944 => x"51",
          5945 => x"82",
          5946 => x"53",
          5947 => x"08",
          5948 => x"81",
          5949 => x"80",
          5950 => x"93",
          5951 => x"3d",
          5952 => x"3d",
          5953 => x"80",
          5954 => x"70",
          5955 => x"52",
          5956 => x"3f",
          5957 => x"08",
          5958 => x"c8",
          5959 => x"63",
          5960 => x"d5",
          5961 => x"93",
          5962 => x"82",
          5963 => x"a3",
          5964 => x"c7",
          5965 => x"98",
          5966 => x"73",
          5967 => x"38",
          5968 => x"39",
          5969 => x"8b",
          5970 => x"93",
          5971 => x"51",
          5972 => x"74",
          5973 => x"0c",
          5974 => x"04",
          5975 => x"61",
          5976 => x"80",
          5977 => x"ec",
          5978 => x"3d",
          5979 => x"3f",
          5980 => x"08",
          5981 => x"c8",
          5982 => x"38",
          5983 => x"73",
          5984 => x"08",
          5985 => x"55",
          5986 => x"74",
          5987 => x"90",
          5988 => x"0c",
          5989 => x"81",
          5990 => x"39",
          5991 => x"ca",
          5992 => x"70",
          5993 => x"57",
          5994 => x"09",
          5995 => x"c0",
          5996 => x"5d",
          5997 => x"90",
          5998 => x"51",
          5999 => x"3f",
          6000 => x"08",
          6001 => x"38",
          6002 => x"08",
          6003 => x"38",
          6004 => x"08",
          6005 => x"93",
          6006 => x"80",
          6007 => x"81",
          6008 => x"58",
          6009 => x"14",
          6010 => x"c9",
          6011 => x"39",
          6012 => x"08",
          6013 => x"5a",
          6014 => x"55",
          6015 => x"77",
          6016 => x"7b",
          6017 => x"b9",
          6018 => x"93",
          6019 => x"82",
          6020 => x"80",
          6021 => x"70",
          6022 => x"73",
          6023 => x"81",
          6024 => x"7a",
          6025 => x"51",
          6026 => x"3f",
          6027 => x"08",
          6028 => x"06",
          6029 => x"80",
          6030 => x"18",
          6031 => x"54",
          6032 => x"15",
          6033 => x"ff",
          6034 => x"82",
          6035 => x"f0",
          6036 => x"30",
          6037 => x"19",
          6038 => x"59",
          6039 => x"83",
          6040 => x"17",
          6041 => x"ff",
          6042 => x"7a",
          6043 => x"90",
          6044 => x"7a",
          6045 => x"81",
          6046 => x"73",
          6047 => x"78",
          6048 => x"0c",
          6049 => x"04",
          6050 => x"7a",
          6051 => x"05",
          6052 => x"58",
          6053 => x"82",
          6054 => x"57",
          6055 => x"08",
          6056 => x"18",
          6057 => x"80",
          6058 => x"76",
          6059 => x"39",
          6060 => x"70",
          6061 => x"81",
          6062 => x"56",
          6063 => x"80",
          6064 => x"38",
          6065 => x"8c",
          6066 => x"81",
          6067 => x"18",
          6068 => x"80",
          6069 => x"08",
          6070 => x"ff",
          6071 => x"82",
          6072 => x"57",
          6073 => x"19",
          6074 => x"39",
          6075 => x"52",
          6076 => x"b9",
          6077 => x"93",
          6078 => x"93",
          6079 => x"32",
          6080 => x"72",
          6081 => x"52",
          6082 => x"82",
          6083 => x"81",
          6084 => x"06",
          6085 => x"57",
          6086 => x"78",
          6087 => x"16",
          6088 => x"38",
          6089 => x"53",
          6090 => x"51",
          6091 => x"3f",
          6092 => x"08",
          6093 => x"08",
          6094 => x"90",
          6095 => x"c0",
          6096 => x"90",
          6097 => x"b9",
          6098 => x"2b",
          6099 => x"25",
          6100 => x"54",
          6101 => x"53",
          6102 => x"78",
          6103 => x"52",
          6104 => x"f5",
          6105 => x"c8",
          6106 => x"85",
          6107 => x"8c",
          6108 => x"33",
          6109 => x"55",
          6110 => x"34",
          6111 => x"89",
          6112 => x"19",
          6113 => x"83",
          6114 => x"75",
          6115 => x"0c",
          6116 => x"04",
          6117 => x"81",
          6118 => x"ff",
          6119 => x"82",
          6120 => x"ff",
          6121 => x"a0",
          6122 => x"b2",
          6123 => x"c8",
          6124 => x"93",
          6125 => x"d3",
          6126 => x"90",
          6127 => x"b3",
          6128 => x"6f",
          6129 => x"d4",
          6130 => x"c2",
          6131 => x"c8",
          6132 => x"94",
          6133 => x"96",
          6134 => x"82",
          6135 => x"80",
          6136 => x"70",
          6137 => x"81",
          6138 => x"55",
          6139 => x"83",
          6140 => x"75",
          6141 => x"81",
          6142 => x"ff",
          6143 => x"02",
          6144 => x"33",
          6145 => x"55",
          6146 => x"25",
          6147 => x"56",
          6148 => x"80",
          6149 => x"81",
          6150 => x"80",
          6151 => x"87",
          6152 => x"e7",
          6153 => x"77",
          6154 => x"3f",
          6155 => x"08",
          6156 => x"80",
          6157 => x"70",
          6158 => x"81",
          6159 => x"56",
          6160 => x"2e",
          6161 => x"81",
          6162 => x"ff",
          6163 => x"87",
          6164 => x"94",
          6165 => x"2e",
          6166 => x"81",
          6167 => x"ff",
          6168 => x"77",
          6169 => x"81",
          6170 => x"ff",
          6171 => x"80",
          6172 => x"70",
          6173 => x"82",
          6174 => x"c8",
          6175 => x"93",
          6176 => x"87",
          6177 => x"c8",
          6178 => x"51",
          6179 => x"82",
          6180 => x"56",
          6181 => x"08",
          6182 => x"56",
          6183 => x"70",
          6184 => x"07",
          6185 => x"06",
          6186 => x"75",
          6187 => x"81",
          6188 => x"ff",
          6189 => x"9f",
          6190 => x"51",
          6191 => x"82",
          6192 => x"82",
          6193 => x"30",
          6194 => x"c8",
          6195 => x"25",
          6196 => x"7b",
          6197 => x"72",
          6198 => x"51",
          6199 => x"80",
          6200 => x"81",
          6201 => x"ff",
          6202 => x"80",
          6203 => x"9f",
          6204 => x"51",
          6205 => x"3f",
          6206 => x"08",
          6207 => x"38",
          6208 => x"b4",
          6209 => x"93",
          6210 => x"81",
          6211 => x"ff",
          6212 => x"75",
          6213 => x"0c",
          6214 => x"04",
          6215 => x"82",
          6216 => x"c0",
          6217 => x"3d",
          6218 => x"3f",
          6219 => x"08",
          6220 => x"c8",
          6221 => x"38",
          6222 => x"52",
          6223 => x"05",
          6224 => x"3f",
          6225 => x"08",
          6226 => x"c8",
          6227 => x"88",
          6228 => x"2e",
          6229 => x"82",
          6230 => x"80",
          6231 => x"70",
          6232 => x"81",
          6233 => x"56",
          6234 => x"83",
          6235 => x"74",
          6236 => x"81",
          6237 => x"38",
          6238 => x"52",
          6239 => x"05",
          6240 => x"dc",
          6241 => x"c8",
          6242 => x"55",
          6243 => x"08",
          6244 => x"81",
          6245 => x"87",
          6246 => x"2e",
          6247 => x"83",
          6248 => x"75",
          6249 => x"81",
          6250 => x"81",
          6251 => x"b2",
          6252 => x"81",
          6253 => x"52",
          6254 => x"bd",
          6255 => x"93",
          6256 => x"82",
          6257 => x"81",
          6258 => x"53",
          6259 => x"18",
          6260 => x"fa",
          6261 => x"ae",
          6262 => x"34",
          6263 => x"0b",
          6264 => x"76",
          6265 => x"18",
          6266 => x"8f",
          6267 => x"b4",
          6268 => x"51",
          6269 => x"a0",
          6270 => x"52",
          6271 => x"51",
          6272 => x"3f",
          6273 => x"0b",
          6274 => x"34",
          6275 => x"d4",
          6276 => x"51",
          6277 => x"77",
          6278 => x"83",
          6279 => x"3d",
          6280 => x"c5",
          6281 => x"93",
          6282 => x"82",
          6283 => x"af",
          6284 => x"63",
          6285 => x"ff",
          6286 => x"75",
          6287 => x"77",
          6288 => x"3f",
          6289 => x"0b",
          6290 => x"77",
          6291 => x"83",
          6292 => x"51",
          6293 => x"3f",
          6294 => x"08",
          6295 => x"80",
          6296 => x"98",
          6297 => x"51",
          6298 => x"3f",
          6299 => x"c8",
          6300 => x"0d",
          6301 => x"0d",
          6302 => x"05",
          6303 => x"3f",
          6304 => x"3d",
          6305 => x"52",
          6306 => x"d0",
          6307 => x"93",
          6308 => x"82",
          6309 => x"82",
          6310 => x"4c",
          6311 => x"52",
          6312 => x"05",
          6313 => x"3f",
          6314 => x"08",
          6315 => x"c8",
          6316 => x"38",
          6317 => x"05",
          6318 => x"06",
          6319 => x"2e",
          6320 => x"55",
          6321 => x"38",
          6322 => x"3d",
          6323 => x"3d",
          6324 => x"51",
          6325 => x"3f",
          6326 => x"3d",
          6327 => x"91",
          6328 => x"54",
          6329 => x"3f",
          6330 => x"52",
          6331 => x"9e",
          6332 => x"c8",
          6333 => x"93",
          6334 => x"38",
          6335 => x"09",
          6336 => x"38",
          6337 => x"a1",
          6338 => x"83",
          6339 => x"74",
          6340 => x"81",
          6341 => x"38",
          6342 => x"a8",
          6343 => x"ec",
          6344 => x"c8",
          6345 => x"93",
          6346 => x"c4",
          6347 => x"93",
          6348 => x"ff",
          6349 => x"8d",
          6350 => x"ac",
          6351 => x"ab",
          6352 => x"17",
          6353 => x"33",
          6354 => x"70",
          6355 => x"55",
          6356 => x"38",
          6357 => x"54",
          6358 => x"34",
          6359 => x"0b",
          6360 => x"8b",
          6361 => x"84",
          6362 => x"06",
          6363 => x"73",
          6364 => x"db",
          6365 => x"2e",
          6366 => x"75",
          6367 => x"ff",
          6368 => x"82",
          6369 => x"52",
          6370 => x"b0",
          6371 => x"55",
          6372 => x"08",
          6373 => x"38",
          6374 => x"08",
          6375 => x"ff",
          6376 => x"82",
          6377 => x"80",
          6378 => x"55",
          6379 => x"08",
          6380 => x"16",
          6381 => x"ae",
          6382 => x"06",
          6383 => x"53",
          6384 => x"51",
          6385 => x"3f",
          6386 => x"0b",
          6387 => x"74",
          6388 => x"3d",
          6389 => x"c3",
          6390 => x"93",
          6391 => x"82",
          6392 => x"8c",
          6393 => x"ff",
          6394 => x"82",
          6395 => x"55",
          6396 => x"c8",
          6397 => x"0d",
          6398 => x"0d",
          6399 => x"05",
          6400 => x"05",
          6401 => x"33",
          6402 => x"53",
          6403 => x"05",
          6404 => x"51",
          6405 => x"82",
          6406 => x"55",
          6407 => x"08",
          6408 => x"78",
          6409 => x"95",
          6410 => x"51",
          6411 => x"82",
          6412 => x"55",
          6413 => x"08",
          6414 => x"80",
          6415 => x"81",
          6416 => x"73",
          6417 => x"38",
          6418 => x"aa",
          6419 => x"06",
          6420 => x"8b",
          6421 => x"06",
          6422 => x"07",
          6423 => x"56",
          6424 => x"34",
          6425 => x"0b",
          6426 => x"78",
          6427 => x"a0",
          6428 => x"c8",
          6429 => x"82",
          6430 => x"95",
          6431 => x"ee",
          6432 => x"56",
          6433 => x"3d",
          6434 => x"95",
          6435 => x"ce",
          6436 => x"c8",
          6437 => x"93",
          6438 => x"d3",
          6439 => x"64",
          6440 => x"d4",
          6441 => x"e6",
          6442 => x"c8",
          6443 => x"93",
          6444 => x"38",
          6445 => x"05",
          6446 => x"06",
          6447 => x"2e",
          6448 => x"55",
          6449 => x"86",
          6450 => x"17",
          6451 => x"2b",
          6452 => x"57",
          6453 => x"05",
          6454 => x"9f",
          6455 => x"81",
          6456 => x"34",
          6457 => x"ac",
          6458 => x"93",
          6459 => x"74",
          6460 => x"0c",
          6461 => x"04",
          6462 => x"69",
          6463 => x"80",
          6464 => x"d0",
          6465 => x"3d",
          6466 => x"3f",
          6467 => x"08",
          6468 => x"08",
          6469 => x"93",
          6470 => x"80",
          6471 => x"70",
          6472 => x"2a",
          6473 => x"57",
          6474 => x"74",
          6475 => x"f6",
          6476 => x"80",
          6477 => x"8d",
          6478 => x"54",
          6479 => x"3f",
          6480 => x"08",
          6481 => x"c8",
          6482 => x"38",
          6483 => x"51",
          6484 => x"3f",
          6485 => x"08",
          6486 => x"c8",
          6487 => x"82",
          6488 => x"82",
          6489 => x"65",
          6490 => x"79",
          6491 => x"7a",
          6492 => x"55",
          6493 => x"34",
          6494 => x"8a",
          6495 => x"38",
          6496 => x"80",
          6497 => x"80",
          6498 => x"ff",
          6499 => x"70",
          6500 => x"58",
          6501 => x"e8",
          6502 => x"2e",
          6503 => x"86",
          6504 => x"34",
          6505 => x"30",
          6506 => x"80",
          6507 => x"70",
          6508 => x"2a",
          6509 => x"56",
          6510 => x"80",
          6511 => x"7b",
          6512 => x"53",
          6513 => x"81",
          6514 => x"c8",
          6515 => x"93",
          6516 => x"38",
          6517 => x"51",
          6518 => x"58",
          6519 => x"8b",
          6520 => x"58",
          6521 => x"83",
          6522 => x"7b",
          6523 => x"51",
          6524 => x"3f",
          6525 => x"08",
          6526 => x"82",
          6527 => x"98",
          6528 => x"e8",
          6529 => x"53",
          6530 => x"b8",
          6531 => x"3d",
          6532 => x"3f",
          6533 => x"08",
          6534 => x"c8",
          6535 => x"38",
          6536 => x"52",
          6537 => x"bc",
          6538 => x"a7",
          6539 => x"6b",
          6540 => x"52",
          6541 => x"9f",
          6542 => x"b5",
          6543 => x"6b",
          6544 => x"70",
          6545 => x"52",
          6546 => x"fe",
          6547 => x"c8",
          6548 => x"a2",
          6549 => x"33",
          6550 => x"54",
          6551 => x"3f",
          6552 => x"08",
          6553 => x"38",
          6554 => x"74",
          6555 => x"05",
          6556 => x"39",
          6557 => x"9f",
          6558 => x"99",
          6559 => x"e0",
          6560 => x"ff",
          6561 => x"54",
          6562 => x"27",
          6563 => x"fa",
          6564 => x"56",
          6565 => x"a3",
          6566 => x"81",
          6567 => x"ff",
          6568 => x"82",
          6569 => x"93",
          6570 => x"76",
          6571 => x"76",
          6572 => x"38",
          6573 => x"77",
          6574 => x"86",
          6575 => x"39",
          6576 => x"27",
          6577 => x"3d",
          6578 => x"bc",
          6579 => x"2a",
          6580 => x"75",
          6581 => x"57",
          6582 => x"05",
          6583 => x"54",
          6584 => x"81",
          6585 => x"33",
          6586 => x"73",
          6587 => x"cd",
          6588 => x"33",
          6589 => x"73",
          6590 => x"81",
          6591 => x"80",
          6592 => x"02",
          6593 => x"78",
          6594 => x"51",
          6595 => x"73",
          6596 => x"81",
          6597 => x"ff",
          6598 => x"80",
          6599 => x"76",
          6600 => x"51",
          6601 => x"2e",
          6602 => x"5f",
          6603 => x"52",
          6604 => x"52",
          6605 => x"c2",
          6606 => x"c8",
          6607 => x"93",
          6608 => x"a1",
          6609 => x"74",
          6610 => x"82",
          6611 => x"c8",
          6612 => x"93",
          6613 => x"38",
          6614 => x"91",
          6615 => x"9a",
          6616 => x"05",
          6617 => x"ff",
          6618 => x"86",
          6619 => x"e5",
          6620 => x"54",
          6621 => x"15",
          6622 => x"ff",
          6623 => x"82",
          6624 => x"54",
          6625 => x"82",
          6626 => x"84",
          6627 => x"06",
          6628 => x"80",
          6629 => x"2e",
          6630 => x"81",
          6631 => x"d4",
          6632 => x"b6",
          6633 => x"93",
          6634 => x"82",
          6635 => x"b5",
          6636 => x"82",
          6637 => x"52",
          6638 => x"a4",
          6639 => x"54",
          6640 => x"15",
          6641 => x"9a",
          6642 => x"05",
          6643 => x"ff",
          6644 => x"77",
          6645 => x"83",
          6646 => x"51",
          6647 => x"3f",
          6648 => x"08",
          6649 => x"74",
          6650 => x"0c",
          6651 => x"04",
          6652 => x"61",
          6653 => x"05",
          6654 => x"33",
          6655 => x"05",
          6656 => x"5e",
          6657 => x"a2",
          6658 => x"c8",
          6659 => x"93",
          6660 => x"38",
          6661 => x"57",
          6662 => x"86",
          6663 => x"82",
          6664 => x"80",
          6665 => x"8c",
          6666 => x"38",
          6667 => x"70",
          6668 => x"81",
          6669 => x"55",
          6670 => x"87",
          6671 => x"39",
          6672 => x"89",
          6673 => x"81",
          6674 => x"8a",
          6675 => x"89",
          6676 => x"7d",
          6677 => x"54",
          6678 => x"3f",
          6679 => x"06",
          6680 => x"72",
          6681 => x"82",
          6682 => x"05",
          6683 => x"08",
          6684 => x"55",
          6685 => x"81",
          6686 => x"38",
          6687 => x"79",
          6688 => x"82",
          6689 => x"56",
          6690 => x"74",
          6691 => x"ff",
          6692 => x"82",
          6693 => x"81",
          6694 => x"56",
          6695 => x"08",
          6696 => x"38",
          6697 => x"81",
          6698 => x"38",
          6699 => x"ff",
          6700 => x"8b",
          6701 => x"5a",
          6702 => x"91",
          6703 => x"74",
          6704 => x"74",
          6705 => x"81",
          6706 => x"87",
          6707 => x"86",
          6708 => x"2e",
          6709 => x"7e",
          6710 => x"80",
          6711 => x"81",
          6712 => x"81",
          6713 => x"06",
          6714 => x"54",
          6715 => x"52",
          6716 => x"a7",
          6717 => x"93",
          6718 => x"82",
          6719 => x"91",
          6720 => x"16",
          6721 => x"56",
          6722 => x"38",
          6723 => x"1d",
          6724 => x"c2",
          6725 => x"8c",
          6726 => x"7b",
          6727 => x"38",
          6728 => x"0c",
          6729 => x"0c",
          6730 => x"80",
          6731 => x"73",
          6732 => x"7f",
          6733 => x"fe",
          6734 => x"90",
          6735 => x"26",
          6736 => x"15",
          6737 => x"90",
          6738 => x"84",
          6739 => x"07",
          6740 => x"84",
          6741 => x"54",
          6742 => x"c8",
          6743 => x"0d",
          6744 => x"0d",
          6745 => x"05",
          6746 => x"33",
          6747 => x"5e",
          6748 => x"d3",
          6749 => x"c8",
          6750 => x"57",
          6751 => x"93",
          6752 => x"8c",
          6753 => x"93",
          6754 => x"10",
          6755 => x"05",
          6756 => x"80",
          6757 => x"74",
          6758 => x"75",
          6759 => x"ff",
          6760 => x"52",
          6761 => x"99",
          6762 => x"93",
          6763 => x"ff",
          6764 => x"06",
          6765 => x"57",
          6766 => x"38",
          6767 => x"70",
          6768 => x"55",
          6769 => x"8c",
          6770 => x"3d",
          6771 => x"83",
          6772 => x"ff",
          6773 => x"82",
          6774 => x"98",
          6775 => x"2e",
          6776 => x"82",
          6777 => x"8c",
          6778 => x"05",
          6779 => x"74",
          6780 => x"38",
          6781 => x"80",
          6782 => x"2e",
          6783 => x"78",
          6784 => x"77",
          6785 => x"26",
          6786 => x"18",
          6787 => x"74",
          6788 => x"38",
          6789 => x"be",
          6790 => x"77",
          6791 => x"98",
          6792 => x"c8",
          6793 => x"54",
          6794 => x"58",
          6795 => x"3f",
          6796 => x"08",
          6797 => x"c8",
          6798 => x"30",
          6799 => x"80",
          6800 => x"c8",
          6801 => x"82",
          6802 => x"07",
          6803 => x"07",
          6804 => x"58",
          6805 => x"57",
          6806 => x"38",
          6807 => x"05",
          6808 => x"79",
          6809 => x"cb",
          6810 => x"82",
          6811 => x"8a",
          6812 => x"83",
          6813 => x"06",
          6814 => x"44",
          6815 => x"09",
          6816 => x"38",
          6817 => x"57",
          6818 => x"8a",
          6819 => x"64",
          6820 => x"57",
          6821 => x"27",
          6822 => x"93",
          6823 => x"80",
          6824 => x"38",
          6825 => x"70",
          6826 => x"55",
          6827 => x"95",
          6828 => x"06",
          6829 => x"2e",
          6830 => x"81",
          6831 => x"85",
          6832 => x"8f",
          6833 => x"06",
          6834 => x"82",
          6835 => x"2e",
          6836 => x"77",
          6837 => x"2e",
          6838 => x"80",
          6839 => x"b4",
          6840 => x"2a",
          6841 => x"81",
          6842 => x"9c",
          6843 => x"52",
          6844 => x"74",
          6845 => x"38",
          6846 => x"98",
          6847 => x"79",
          6848 => x"18",
          6849 => x"57",
          6850 => x"80",
          6851 => x"76",
          6852 => x"38",
          6853 => x"51",
          6854 => x"3f",
          6855 => x"08",
          6856 => x"08",
          6857 => x"7f",
          6858 => x"52",
          6859 => x"88",
          6860 => x"c8",
          6861 => x"5b",
          6862 => x"80",
          6863 => x"43",
          6864 => x"0a",
          6865 => x"8b",
          6866 => x"89",
          6867 => x"b4",
          6868 => x"2a",
          6869 => x"81",
          6870 => x"8c",
          6871 => x"52",
          6872 => x"74",
          6873 => x"38",
          6874 => x"98",
          6875 => x"79",
          6876 => x"18",
          6877 => x"57",
          6878 => x"80",
          6879 => x"76",
          6880 => x"38",
          6881 => x"51",
          6882 => x"3f",
          6883 => x"08",
          6884 => x"57",
          6885 => x"08",
          6886 => x"92",
          6887 => x"82",
          6888 => x"83",
          6889 => x"72",
          6890 => x"51",
          6891 => x"52",
          6892 => x"05",
          6893 => x"80",
          6894 => x"c8",
          6895 => x"7e",
          6896 => x"80",
          6897 => x"f2",
          6898 => x"93",
          6899 => x"ff",
          6900 => x"63",
          6901 => x"64",
          6902 => x"ff",
          6903 => x"70",
          6904 => x"31",
          6905 => x"57",
          6906 => x"2e",
          6907 => x"89",
          6908 => x"60",
          6909 => x"84",
          6910 => x"5c",
          6911 => x"16",
          6912 => x"51",
          6913 => x"26",
          6914 => x"65",
          6915 => x"31",
          6916 => x"64",
          6917 => x"fe",
          6918 => x"82",
          6919 => x"56",
          6920 => x"09",
          6921 => x"38",
          6922 => x"08",
          6923 => x"26",
          6924 => x"89",
          6925 => x"2a",
          6926 => x"97",
          6927 => x"87",
          6928 => x"82",
          6929 => x"06",
          6930 => x"83",
          6931 => x"27",
          6932 => x"8f",
          6933 => x"55",
          6934 => x"26",
          6935 => x"58",
          6936 => x"7c",
          6937 => x"06",
          6938 => x"2e",
          6939 => x"42",
          6940 => x"77",
          6941 => x"19",
          6942 => x"78",
          6943 => x"38",
          6944 => x"d2",
          6945 => x"f5",
          6946 => x"77",
          6947 => x"19",
          6948 => x"78",
          6949 => x"38",
          6950 => x"ba",
          6951 => x"61",
          6952 => x"81",
          6953 => x"61",
          6954 => x"f5",
          6955 => x"55",
          6956 => x"86",
          6957 => x"53",
          6958 => x"51",
          6959 => x"3f",
          6960 => x"fb",
          6961 => x"51",
          6962 => x"3f",
          6963 => x"1f",
          6964 => x"89",
          6965 => x"8d",
          6966 => x"83",
          6967 => x"52",
          6968 => x"ff",
          6969 => x"81",
          6970 => x"34",
          6971 => x"70",
          6972 => x"2a",
          6973 => x"54",
          6974 => x"1f",
          6975 => x"dd",
          6976 => x"ff",
          6977 => x"38",
          6978 => x"05",
          6979 => x"1f",
          6980 => x"c9",
          6981 => x"65",
          6982 => x"51",
          6983 => x"3f",
          6984 => x"05",
          6985 => x"98",
          6986 => x"98",
          6987 => x"ff",
          6988 => x"51",
          6989 => x"3f",
          6990 => x"1f",
          6991 => x"bb",
          6992 => x"2e",
          6993 => x"80",
          6994 => x"88",
          6995 => x"80",
          6996 => x"ff",
          6997 => x"7b",
          6998 => x"51",
          6999 => x"3f",
          7000 => x"1f",
          7001 => x"93",
          7002 => x"b0",
          7003 => x"97",
          7004 => x"52",
          7005 => x"ff",
          7006 => x"ff",
          7007 => x"c0",
          7008 => x"7f",
          7009 => x"34",
          7010 => x"fb",
          7011 => x"c7",
          7012 => x"98",
          7013 => x"39",
          7014 => x"0a",
          7015 => x"51",
          7016 => x"3f",
          7017 => x"ff",
          7018 => x"1f",
          7019 => x"ad",
          7020 => x"7f",
          7021 => x"a9",
          7022 => x"34",
          7023 => x"fb",
          7024 => x"1f",
          7025 => x"e2",
          7026 => x"d5",
          7027 => x"1f",
          7028 => x"89",
          7029 => x"63",
          7030 => x"79",
          7031 => x"f9",
          7032 => x"82",
          7033 => x"83",
          7034 => x"83",
          7035 => x"06",
          7036 => x"81",
          7037 => x"05",
          7038 => x"79",
          7039 => x"d9",
          7040 => x"80",
          7041 => x"ff",
          7042 => x"84",
          7043 => x"d2",
          7044 => x"ff",
          7045 => x"86",
          7046 => x"f2",
          7047 => x"1f",
          7048 => x"d7",
          7049 => x"52",
          7050 => x"51",
          7051 => x"3f",
          7052 => x"ec",
          7053 => x"96",
          7054 => x"d4",
          7055 => x"fe",
          7056 => x"96",
          7057 => x"54",
          7058 => x"53",
          7059 => x"51",
          7060 => x"3f",
          7061 => x"81",
          7062 => x"52",
          7063 => x"92",
          7064 => x"53",
          7065 => x"51",
          7066 => x"3f",
          7067 => x"5b",
          7068 => x"09",
          7069 => x"38",
          7070 => x"51",
          7071 => x"3f",
          7072 => x"1f",
          7073 => x"f3",
          7074 => x"52",
          7075 => x"ff",
          7076 => x"95",
          7077 => x"ff",
          7078 => x"81",
          7079 => x"f8",
          7080 => x"7e",
          7081 => x"d3",
          7082 => x"60",
          7083 => x"26",
          7084 => x"57",
          7085 => x"53",
          7086 => x"51",
          7087 => x"3f",
          7088 => x"08",
          7089 => x"7d",
          7090 => x"7e",
          7091 => x"fe",
          7092 => x"75",
          7093 => x"56",
          7094 => x"81",
          7095 => x"80",
          7096 => x"38",
          7097 => x"83",
          7098 => x"62",
          7099 => x"74",
          7100 => x"38",
          7101 => x"54",
          7102 => x"52",
          7103 => x"91",
          7104 => x"93",
          7105 => x"c8",
          7106 => x"75",
          7107 => x"56",
          7108 => x"8c",
          7109 => x"2e",
          7110 => x"57",
          7111 => x"ff",
          7112 => x"84",
          7113 => x"2e",
          7114 => x"57",
          7115 => x"81",
          7116 => x"80",
          7117 => x"53",
          7118 => x"51",
          7119 => x"3f",
          7120 => x"52",
          7121 => x"51",
          7122 => x"3f",
          7123 => x"56",
          7124 => x"81",
          7125 => x"34",
          7126 => x"17",
          7127 => x"17",
          7128 => x"17",
          7129 => x"05",
          7130 => x"c1",
          7131 => x"fe",
          7132 => x"fe",
          7133 => x"34",
          7134 => x"08",
          7135 => x"07",
          7136 => x"17",
          7137 => x"c8",
          7138 => x"34",
          7139 => x"c6",
          7140 => x"93",
          7141 => x"52",
          7142 => x"51",
          7143 => x"3f",
          7144 => x"53",
          7145 => x"51",
          7146 => x"3f",
          7147 => x"93",
          7148 => x"38",
          7149 => x"52",
          7150 => x"91",
          7151 => x"57",
          7152 => x"08",
          7153 => x"39",
          7154 => x"39",
          7155 => x"39",
          7156 => x"39",
          7157 => x"82",
          7158 => x"98",
          7159 => x"ff",
          7160 => x"52",
          7161 => x"81",
          7162 => x"10",
          7163 => x"b8",
          7164 => x"08",
          7165 => x"f8",
          7166 => x"a9",
          7167 => x"39",
          7168 => x"51",
          7169 => x"3f",
          7170 => x"82",
          7171 => x"ff",
          7172 => x"81",
          7173 => x"82",
          7174 => x"80",
          7175 => x"b3",
          7176 => x"bc",
          7177 => x"fd",
          7178 => x"39",
          7179 => x"51",
          7180 => x"3f",
          7181 => x"82",
          7182 => x"fe",
          7183 => x"81",
          7184 => x"82",
          7185 => x"ff",
          7186 => x"87",
          7187 => x"88",
          7188 => x"d1",
          7189 => x"39",
          7190 => x"51",
          7191 => x"3f",
          7192 => x"82",
          7193 => x"fe",
          7194 => x"80",
          7195 => x"83",
          7196 => x"ff",
          7197 => x"db",
          7198 => x"e8",
          7199 => x"a5",
          7200 => x"39",
          7201 => x"51",
          7202 => x"3f",
          7203 => x"82",
          7204 => x"fe",
          7205 => x"bb",
          7206 => x"c8",
          7207 => x"85",
          7208 => x"82",
          7209 => x"fe",
          7210 => x"a7",
          7211 => x"f4",
          7212 => x"f1",
          7213 => x"82",
          7214 => x"fe",
          7215 => x"93",
          7216 => x"a4",
          7217 => x"dd",
          7218 => x"82",
          7219 => x"fe",
          7220 => x"83",
          7221 => x"fb",
          7222 => x"79",
          7223 => x"87",
          7224 => x"38",
          7225 => x"87",
          7226 => x"fe",
          7227 => x"82",
          7228 => x"55",
          7229 => x"e8",
          7230 => x"fe",
          7231 => x"82",
          7232 => x"52",
          7233 => x"e8",
          7234 => x"93",
          7235 => x"74",
          7236 => x"75",
          7237 => x"c0",
          7238 => x"83",
          7239 => x"0d",
          7240 => x"3d",
          7241 => x"3d",
          7242 => x"3d",
          7243 => x"05",
          7244 => x"33",
          7245 => x"70",
          7246 => x"25",
          7247 => x"27",
          7248 => x"5a",
          7249 => x"93",
          7250 => x"87",
          7251 => x"77",
          7252 => x"3d",
          7253 => x"51",
          7254 => x"3f",
          7255 => x"08",
          7256 => x"c8",
          7257 => x"82",
          7258 => x"87",
          7259 => x"0c",
          7260 => x"08",
          7261 => x"3d",
          7262 => x"55",
          7263 => x"53",
          7264 => x"d8",
          7265 => x"f2",
          7266 => x"c8",
          7267 => x"93",
          7268 => x"38",
          7269 => x"89",
          7270 => x"7b",
          7271 => x"d5",
          7272 => x"3d",
          7273 => x"51",
          7274 => x"77",
          7275 => x"07",
          7276 => x"30",
          7277 => x"72",
          7278 => x"51",
          7279 => x"2e",
          7280 => x"85",
          7281 => x"c0",
          7282 => x"52",
          7283 => x"87",
          7284 => x"74",
          7285 => x"0c",
          7286 => x"0d",
          7287 => x"0d",
          7288 => x"33",
          7289 => x"57",
          7290 => x"7b",
          7291 => x"fe",
          7292 => x"93",
          7293 => x"38",
          7294 => x"88",
          7295 => x"2e",
          7296 => x"39",
          7297 => x"54",
          7298 => x"53",
          7299 => x"51",
          7300 => x"93",
          7301 => x"83",
          7302 => x"78",
          7303 => x"0c",
          7304 => x"04",
          7305 => x"02",
          7306 => x"82",
          7307 => x"82",
          7308 => x"56",
          7309 => x"3f",
          7310 => x"70",
          7311 => x"fe",
          7312 => x"82",
          7313 => x"82",
          7314 => x"81",
          7315 => x"82",
          7316 => x"ff",
          7317 => x"75",
          7318 => x"38",
          7319 => x"3f",
          7320 => x"04",
          7321 => x"87",
          7322 => x"08",
          7323 => x"ff",
          7324 => x"fe",
          7325 => x"82",
          7326 => x"fe",
          7327 => x"80",
          7328 => x"f1",
          7329 => x"2a",
          7330 => x"51",
          7331 => x"2e",
          7332 => x"51",
          7333 => x"3f",
          7334 => x"51",
          7335 => x"3f",
          7336 => x"ee",
          7337 => x"82",
          7338 => x"06",
          7339 => x"80",
          7340 => x"81",
          7341 => x"bd",
          7342 => x"e0",
          7343 => x"b3",
          7344 => x"fe",
          7345 => x"72",
          7346 => x"81",
          7347 => x"71",
          7348 => x"38",
          7349 => x"ee",
          7350 => x"86",
          7351 => x"f0",
          7352 => x"51",
          7353 => x"3f",
          7354 => x"70",
          7355 => x"52",
          7356 => x"95",
          7357 => x"fe",
          7358 => x"82",
          7359 => x"fe",
          7360 => x"80",
          7361 => x"ed",
          7362 => x"2a",
          7363 => x"51",
          7364 => x"2e",
          7365 => x"51",
          7366 => x"3f",
          7367 => x"51",
          7368 => x"3f",
          7369 => x"ed",
          7370 => x"86",
          7371 => x"06",
          7372 => x"80",
          7373 => x"81",
          7374 => x"b9",
          7375 => x"ac",
          7376 => x"af",
          7377 => x"fe",
          7378 => x"72",
          7379 => x"81",
          7380 => x"71",
          7381 => x"38",
          7382 => x"ed",
          7383 => x"87",
          7384 => x"ef",
          7385 => x"51",
          7386 => x"3f",
          7387 => x"70",
          7388 => x"52",
          7389 => x"95",
          7390 => x"fe",
          7391 => x"82",
          7392 => x"fe",
          7393 => x"80",
          7394 => x"e9",
          7395 => x"a8",
          7396 => x"0d",
          7397 => x"0d",
          7398 => x"70",
          7399 => x"74",
          7400 => x"ed",
          7401 => x"74",
          7402 => x"14",
          7403 => x"e1",
          7404 => x"55",
          7405 => x"54",
          7406 => x"2e",
          7407 => x"54",
          7408 => x"9f",
          7409 => x"51",
          7410 => x"38",
          7411 => x"72",
          7412 => x"81",
          7413 => x"80",
          7414 => x"05",
          7415 => x"56",
          7416 => x"82",
          7417 => x"77",
          7418 => x"08",
          7419 => x"e6",
          7420 => x"93",
          7421 => x"38",
          7422 => x"53",
          7423 => x"ff",
          7424 => x"16",
          7425 => x"06",
          7426 => x"76",
          7427 => x"ff",
          7428 => x"93",
          7429 => x"3d",
          7430 => x"3d",
          7431 => x"82",
          7432 => x"71",
          7433 => x"5c",
          7434 => x"52",
          7435 => x"84",
          7436 => x"93",
          7437 => x"ff",
          7438 => x"7c",
          7439 => x"06",
          7440 => x"88",
          7441 => x"3d",
          7442 => x"fe",
          7443 => x"7b",
          7444 => x"ea",
          7445 => x"ff",
          7446 => x"82",
          7447 => x"5a",
          7448 => x"8b",
          7449 => x"98",
          7450 => x"b3",
          7451 => x"81",
          7452 => x"82",
          7453 => x"fe",
          7454 => x"96",
          7455 => x"59",
          7456 => x"54",
          7457 => x"78",
          7458 => x"a4",
          7459 => x"61",
          7460 => x"e5",
          7461 => x"fe",
          7462 => x"fd",
          7463 => x"93",
          7464 => x"2b",
          7465 => x"51",
          7466 => x"87",
          7467 => x"38",
          7468 => x"81",
          7469 => x"59",
          7470 => x"b4",
          7471 => x"11",
          7472 => x"05",
          7473 => x"e2",
          7474 => x"c8",
          7475 => x"82",
          7476 => x"fe",
          7477 => x"ff",
          7478 => x"3d",
          7479 => x"53",
          7480 => x"51",
          7481 => x"3f",
          7482 => x"08",
          7483 => x"38",
          7484 => x"83",
          7485 => x"02",
          7486 => x"52",
          7487 => x"05",
          7488 => x"82",
          7489 => x"93",
          7490 => x"ff",
          7491 => x"8e",
          7492 => x"e4",
          7493 => x"8d",
          7494 => x"fe",
          7495 => x"88",
          7496 => x"f6",
          7497 => x"cb",
          7498 => x"fe",
          7499 => x"fe",
          7500 => x"fe",
          7501 => x"82",
          7502 => x"80",
          7503 => x"38",
          7504 => x"52",
          7505 => x"05",
          7506 => x"86",
          7507 => x"93",
          7508 => x"82",
          7509 => x"fe",
          7510 => x"fe",
          7511 => x"3d",
          7512 => x"53",
          7513 => x"51",
          7514 => x"3f",
          7515 => x"08",
          7516 => x"38",
          7517 => x"fd",
          7518 => x"3d",
          7519 => x"53",
          7520 => x"51",
          7521 => x"3f",
          7522 => x"08",
          7523 => x"93",
          7524 => x"60",
          7525 => x"94",
          7526 => x"70",
          7527 => x"fb",
          7528 => x"bf",
          7529 => x"78",
          7530 => x"b4",
          7531 => x"f8",
          7532 => x"b2",
          7533 => x"93",
          7534 => x"2e",
          7535 => x"93",
          7536 => x"f4",
          7537 => x"ab",
          7538 => x"e4",
          7539 => x"d5",
          7540 => x"fd",
          7541 => x"3d",
          7542 => x"51",
          7543 => x"3f",
          7544 => x"08",
          7545 => x"f8",
          7546 => x"fe",
          7547 => x"81",
          7548 => x"c8",
          7549 => x"51",
          7550 => x"82",
          7551 => x"80",
          7552 => x"38",
          7553 => x"08",
          7554 => x"3f",
          7555 => x"b4",
          7556 => x"05",
          7557 => x"eb",
          7558 => x"c8",
          7559 => x"fe",
          7560 => x"5b",
          7561 => x"3f",
          7562 => x"08",
          7563 => x"f8",
          7564 => x"fe",
          7565 => x"82",
          7566 => x"b5",
          7567 => x"05",
          7568 => x"e4",
          7569 => x"8b",
          7570 => x"93",
          7571 => x"56",
          7572 => x"93",
          7573 => x"ff",
          7574 => x"53",
          7575 => x"51",
          7576 => x"82",
          7577 => x"80",
          7578 => x"38",
          7579 => x"08",
          7580 => x"3f",
          7581 => x"82",
          7582 => x"fe",
          7583 => x"82",
          7584 => x"8f",
          7585 => x"39",
          7586 => x"51",
          7587 => x"3f",
          7588 => x"f1",
          7589 => x"db",
          7590 => x"81",
          7591 => x"94",
          7592 => x"80",
          7593 => x"c0",
          7594 => x"82",
          7595 => x"fe",
          7596 => x"fb",
          7597 => x"89",
          7598 => x"f2",
          7599 => x"80",
          7600 => x"c0",
          7601 => x"8c",
          7602 => x"87",
          7603 => x"0c",
          7604 => x"b4",
          7605 => x"11",
          7606 => x"05",
          7607 => x"ca",
          7608 => x"c8",
          7609 => x"fb",
          7610 => x"52",
          7611 => x"51",
          7612 => x"3f",
          7613 => x"04",
          7614 => x"f4",
          7615 => x"f8",
          7616 => x"fa",
          7617 => x"93",
          7618 => x"2e",
          7619 => x"60",
          7620 => x"8c",
          7621 => x"87",
          7622 => x"78",
          7623 => x"c8",
          7624 => x"93",
          7625 => x"2e",
          7626 => x"82",
          7627 => x"52",
          7628 => x"51",
          7629 => x"3f",
          7630 => x"82",
          7631 => x"fe",
          7632 => x"fe",
          7633 => x"fa",
          7634 => x"8a",
          7635 => x"f1",
          7636 => x"59",
          7637 => x"fe",
          7638 => x"fa",
          7639 => x"70",
          7640 => x"78",
          7641 => x"8b",
          7642 => x"06",
          7643 => x"2e",
          7644 => x"b4",
          7645 => x"05",
          7646 => x"87",
          7647 => x"f4",
          7648 => x"c8",
          7649 => x"8a",
          7650 => x"53",
          7651 => x"52",
          7652 => x"52",
          7653 => x"9d",
          7654 => x"c4",
          7655 => x"fc",
          7656 => x"61",
          7657 => x"61",
          7658 => x"83",
          7659 => x"83",
          7660 => x"78",
          7661 => x"3f",
          7662 => x"08",
          7663 => x"32",
          7664 => x"07",
          7665 => x"38",
          7666 => x"09",
          7667 => x"a3",
          7668 => x"8c",
          7669 => x"c7",
          7670 => x"39",
          7671 => x"80",
          7672 => x"fc",
          7673 => x"86",
          7674 => x"c0",
          7675 => x"9b",
          7676 => x"0b",
          7677 => x"9c",
          7678 => x"83",
          7679 => x"94",
          7680 => x"80",
          7681 => x"c0",
          7682 => x"80",
          7683 => x"82",
          7684 => x"80",
          7685 => x"82",
          7686 => x"fe",
          7687 => x"fe",
          7688 => x"82",
          7689 => x"fe",
          7690 => x"82",
          7691 => x"fe",
          7692 => x"81",
          7693 => x"fe",
          7694 => x"81",
          7695 => x"3f",
          7696 => x"80",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"00",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"00",
          7708 => x"00",
          7709 => x"00",
          7710 => x"00",
          7711 => x"00",
          7712 => x"00",
          7713 => x"00",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"00",
          7734 => x"00",
          7735 => x"00",
          7736 => x"00",
          7737 => x"00",
          7738 => x"00",
          7739 => x"00",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"00",
          7744 => x"00",
          7745 => x"00",
          7746 => x"00",
          7747 => x"00",
          7748 => x"00",
          7749 => x"00",
          7750 => x"00",
          7751 => x"00",
          7752 => x"00",
          7753 => x"00",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"00",
          7758 => x"00",
          7759 => x"00",
          7760 => x"00",
          7761 => x"00",
          7762 => x"00",
          7763 => x"00",
          7764 => x"00",
          7765 => x"00",
          7766 => x"00",
          7767 => x"00",
          7768 => x"00",
          7769 => x"00",
          7770 => x"00",
          7771 => x"00",
          7772 => x"00",
          7773 => x"00",
          7774 => x"00",
          7775 => x"00",
          7776 => x"00",
          7777 => x"00",
          7778 => x"00",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"00",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"00",
          7810 => x"00",
          7811 => x"00",
          7812 => x"00",
          7813 => x"00",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"00",
          7848 => x"00",
          7849 => x"00",
          7850 => x"00",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"00",
          7855 => x"00",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"00",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"00",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"00",
          7868 => x"00",
          7869 => x"00",
          7870 => x"00",
          7871 => x"00",
          7872 => x"00",
          7873 => x"00",
          7874 => x"00",
          7875 => x"00",
          7876 => x"00",
          7877 => x"00",
          7878 => x"00",
          7879 => x"00",
          7880 => x"00",
          7881 => x"00",
          7882 => x"64",
          7883 => x"2f",
          7884 => x"25",
          7885 => x"64",
          7886 => x"2e",
          7887 => x"64",
          7888 => x"6f",
          7889 => x"6f",
          7890 => x"67",
          7891 => x"74",
          7892 => x"00",
          7893 => x"28",
          7894 => x"6d",
          7895 => x"43",
          7896 => x"6e",
          7897 => x"29",
          7898 => x"0a",
          7899 => x"69",
          7900 => x"20",
          7901 => x"6c",
          7902 => x"6e",
          7903 => x"3a",
          7904 => x"20",
          7905 => x"4e",
          7906 => x"42",
          7907 => x"20",
          7908 => x"61",
          7909 => x"25",
          7910 => x"2c",
          7911 => x"7a",
          7912 => x"30",
          7913 => x"2e",
          7914 => x"20",
          7915 => x"52",
          7916 => x"28",
          7917 => x"72",
          7918 => x"30",
          7919 => x"20",
          7920 => x"65",
          7921 => x"38",
          7922 => x"0a",
          7923 => x"20",
          7924 => x"41",
          7925 => x"53",
          7926 => x"74",
          7927 => x"38",
          7928 => x"53",
          7929 => x"3d",
          7930 => x"58",
          7931 => x"00",
          7932 => x"20",
          7933 => x"4f",
          7934 => x"0a",
          7935 => x"20",
          7936 => x"53",
          7937 => x"00",
          7938 => x"20",
          7939 => x"50",
          7940 => x"00",
          7941 => x"20",
          7942 => x"44",
          7943 => x"72",
          7944 => x"44",
          7945 => x"63",
          7946 => x"25",
          7947 => x"29",
          7948 => x"00",
          7949 => x"20",
          7950 => x"4e",
          7951 => x"52",
          7952 => x"20",
          7953 => x"54",
          7954 => x"4c",
          7955 => x"00",
          7956 => x"20",
          7957 => x"49",
          7958 => x"31",
          7959 => x"69",
          7960 => x"73",
          7961 => x"31",
          7962 => x"0a",
          7963 => x"64",
          7964 => x"73",
          7965 => x"3a",
          7966 => x"20",
          7967 => x"50",
          7968 => x"65",
          7969 => x"20",
          7970 => x"74",
          7971 => x"41",
          7972 => x"65",
          7973 => x"3d",
          7974 => x"38",
          7975 => x"00",
          7976 => x"20",
          7977 => x"50",
          7978 => x"65",
          7979 => x"79",
          7980 => x"61",
          7981 => x"41",
          7982 => x"65",
          7983 => x"3d",
          7984 => x"38",
          7985 => x"00",
          7986 => x"20",
          7987 => x"74",
          7988 => x"20",
          7989 => x"72",
          7990 => x"64",
          7991 => x"73",
          7992 => x"20",
          7993 => x"3d",
          7994 => x"38",
          7995 => x"00",
          7996 => x"20",
          7997 => x"50",
          7998 => x"64",
          7999 => x"20",
          8000 => x"20",
          8001 => x"20",
          8002 => x"20",
          8003 => x"3d",
          8004 => x"38",
          8005 => x"00",
          8006 => x"20",
          8007 => x"79",
          8008 => x"6d",
          8009 => x"6f",
          8010 => x"46",
          8011 => x"20",
          8012 => x"20",
          8013 => x"3d",
          8014 => x"38",
          8015 => x"00",
          8016 => x"6d",
          8017 => x"00",
          8018 => x"65",
          8019 => x"6d",
          8020 => x"6c",
          8021 => x"00",
          8022 => x"56",
          8023 => x"56",
          8024 => x"6e",
          8025 => x"6e",
          8026 => x"77",
          8027 => x"44",
          8028 => x"2a",
          8029 => x"3b",
          8030 => x"3f",
          8031 => x"7f",
          8032 => x"41",
          8033 => x"41",
          8034 => x"00",
          8035 => x"0a",
          8036 => x"0a",
          8037 => x"0a",
          8038 => x"0a",
          8039 => x"0a",
          8040 => x"0a",
          8041 => x"0a",
          8042 => x"0a",
          8043 => x"0a",
          8044 => x"30",
          8045 => x"fe",
          8046 => x"44",
          8047 => x"2e",
          8048 => x"4f",
          8049 => x"4d",
          8050 => x"20",
          8051 => x"54",
          8052 => x"20",
          8053 => x"4f",
          8054 => x"4d",
          8055 => x"20",
          8056 => x"54",
          8057 => x"20",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"9a",
          8063 => x"41",
          8064 => x"45",
          8065 => x"49",
          8066 => x"92",
          8067 => x"4f",
          8068 => x"99",
          8069 => x"9d",
          8070 => x"49",
          8071 => x"a5",
          8072 => x"a9",
          8073 => x"ad",
          8074 => x"b1",
          8075 => x"b5",
          8076 => x"b9",
          8077 => x"bd",
          8078 => x"c1",
          8079 => x"c5",
          8080 => x"c9",
          8081 => x"cd",
          8082 => x"d1",
          8083 => x"d5",
          8084 => x"d9",
          8085 => x"dd",
          8086 => x"e1",
          8087 => x"e5",
          8088 => x"e9",
          8089 => x"ed",
          8090 => x"f1",
          8091 => x"f5",
          8092 => x"f9",
          8093 => x"fd",
          8094 => x"2e",
          8095 => x"5b",
          8096 => x"22",
          8097 => x"3e",
          8098 => x"00",
          8099 => x"01",
          8100 => x"10",
          8101 => x"00",
          8102 => x"00",
          8103 => x"01",
          8104 => x"04",
          8105 => x"10",
          8106 => x"00",
          8107 => x"41",
          8108 => x"00",
          8109 => x"41",
          8110 => x"00",
          8111 => x"78",
          8112 => x"00",
          8113 => x"49",
          8114 => x"49",
          8115 => x"4f",
          8116 => x"4f",
          8117 => x"00",
          8118 => x"49",
          8119 => x"42",
          8120 => x"45",
          8121 => x"4f",
          8122 => x"4f",
          8123 => x"00",
          8124 => x"49",
          8125 => x"59",
          8126 => x"4d",
          8127 => x"4e",
          8128 => x"4c",
          8129 => x"45",
          8130 => x"59",
          8131 => x"41",
          8132 => x"41",
          8133 => x"00",
          8134 => x"45",
          8135 => x"4e",
          8136 => x"58",
          8137 => x"54",
          8138 => x"00",
          8139 => x"49",
          8140 => x"43",
          8141 => x"41",
          8142 => x"00",
          8143 => x"64",
          8144 => x"00",
          8145 => x"69",
          8146 => x"00",
          8147 => x"73",
          8148 => x"00",
          8149 => x"69",
          8150 => x"6c",
          8151 => x"64",
          8152 => x"00",
          8153 => x"65",
          8154 => x"00",
          8155 => x"72",
          8156 => x"00",
          8157 => x"77",
          8158 => x"65",
          8159 => x"66",
          8160 => x"00",
          8161 => x"6c",
          8162 => x"00",
          8163 => x"69",
          8164 => x"00",
          8165 => x"6f",
          8166 => x"00",
          8167 => x"63",
          8168 => x"65",
          8169 => x"73",
          8170 => x"00",
          8171 => x"72",
          8172 => x"00",
          8173 => x"69",
          8174 => x"65",
          8175 => x"00",
          8176 => x"77",
          8177 => x"65",
          8178 => x"74",
          8179 => x"63",
          8180 => x"61",
          8181 => x"63",
          8182 => x"61",
          8183 => x"00",
          8184 => x"74",
          8185 => x"00",
          8186 => x"72",
          8187 => x"6d",
          8188 => x"64",
          8189 => x"00",
          8190 => x"6d",
          8191 => x"72",
          8192 => x"73",
          8193 => x"00",
          8194 => x"64",
          8195 => x"00",
          8196 => x"63",
          8197 => x"00",
          8198 => x"63",
          8199 => x"63",
          8200 => x"61",
          8201 => x"78",
          8202 => x"63",
          8203 => x"6c",
          8204 => x"00",
          8205 => x"65",
          8206 => x"00",
          8207 => x"73",
          8208 => x"00",
          8209 => x"64",
          8210 => x"00",
          8211 => x"63",
          8212 => x"64",
          8213 => x"65",
          8214 => x"73",
          8215 => x"64",
          8216 => x"00",
          8217 => x"6c",
          8218 => x"6c",
          8219 => x"6d",
          8220 => x"00",
          8221 => x"63",
          8222 => x"00",
          8223 => x"64",
          8224 => x"00",
          8225 => x"65",
          8226 => x"65",
          8227 => x"65",
          8228 => x"69",
          8229 => x"69",
          8230 => x"72",
          8231 => x"74",
          8232 => x"66",
          8233 => x"66",
          8234 => x"68",
          8235 => x"00",
          8236 => x"6f",
          8237 => x"61",
          8238 => x"00",
          8239 => x"61",
          8240 => x"00",
          8241 => x"6d",
          8242 => x"65",
          8243 => x"72",
          8244 => x"65",
          8245 => x"00",
          8246 => x"65",
          8247 => x"00",
          8248 => x"6e",
          8249 => x"00",
          8250 => x"69",
          8251 => x"00",
          8252 => x"65",
          8253 => x"00",
          8254 => x"69",
          8255 => x"45",
          8256 => x"72",
          8257 => x"6e",
          8258 => x"6e",
          8259 => x"65",
          8260 => x"72",
          8261 => x"00",
          8262 => x"69",
          8263 => x"6e",
          8264 => x"72",
          8265 => x"79",
          8266 => x"00",
          8267 => x"6f",
          8268 => x"6c",
          8269 => x"6f",
          8270 => x"2e",
          8271 => x"6f",
          8272 => x"74",
          8273 => x"6f",
          8274 => x"2e",
          8275 => x"6e",
          8276 => x"69",
          8277 => x"69",
          8278 => x"61",
          8279 => x"0a",
          8280 => x"63",
          8281 => x"73",
          8282 => x"6e",
          8283 => x"2e",
          8284 => x"69",
          8285 => x"61",
          8286 => x"61",
          8287 => x"65",
          8288 => x"74",
          8289 => x"00",
          8290 => x"69",
          8291 => x"68",
          8292 => x"6c",
          8293 => x"6e",
          8294 => x"69",
          8295 => x"00",
          8296 => x"44",
          8297 => x"20",
          8298 => x"74",
          8299 => x"72",
          8300 => x"63",
          8301 => x"2e",
          8302 => x"72",
          8303 => x"20",
          8304 => x"62",
          8305 => x"69",
          8306 => x"6e",
          8307 => x"69",
          8308 => x"00",
          8309 => x"69",
          8310 => x"6e",
          8311 => x"65",
          8312 => x"6c",
          8313 => x"0a",
          8314 => x"6f",
          8315 => x"6d",
          8316 => x"69",
          8317 => x"20",
          8318 => x"65",
          8319 => x"74",
          8320 => x"66",
          8321 => x"64",
          8322 => x"20",
          8323 => x"6b",
          8324 => x"00",
          8325 => x"6f",
          8326 => x"74",
          8327 => x"6f",
          8328 => x"64",
          8329 => x"00",
          8330 => x"69",
          8331 => x"75",
          8332 => x"6f",
          8333 => x"61",
          8334 => x"6e",
          8335 => x"6e",
          8336 => x"6c",
          8337 => x"0a",
          8338 => x"69",
          8339 => x"69",
          8340 => x"6f",
          8341 => x"64",
          8342 => x"00",
          8343 => x"6e",
          8344 => x"66",
          8345 => x"65",
          8346 => x"6d",
          8347 => x"72",
          8348 => x"00",
          8349 => x"6f",
          8350 => x"61",
          8351 => x"6f",
          8352 => x"20",
          8353 => x"65",
          8354 => x"00",
          8355 => x"61",
          8356 => x"65",
          8357 => x"73",
          8358 => x"63",
          8359 => x"65",
          8360 => x"0a",
          8361 => x"75",
          8362 => x"73",
          8363 => x"00",
          8364 => x"6e",
          8365 => x"77",
          8366 => x"72",
          8367 => x"2e",
          8368 => x"25",
          8369 => x"62",
          8370 => x"73",
          8371 => x"20",
          8372 => x"25",
          8373 => x"62",
          8374 => x"73",
          8375 => x"63",
          8376 => x"00",
          8377 => x"65",
          8378 => x"00",
          8379 => x"50",
          8380 => x"00",
          8381 => x"2a",
          8382 => x"73",
          8383 => x"00",
          8384 => x"38",
          8385 => x"2f",
          8386 => x"39",
          8387 => x"31",
          8388 => x"00",
          8389 => x"5a",
          8390 => x"20",
          8391 => x"20",
          8392 => x"78",
          8393 => x"73",
          8394 => x"20",
          8395 => x"0a",
          8396 => x"50",
          8397 => x"20",
          8398 => x"65",
          8399 => x"70",
          8400 => x"61",
          8401 => x"65",
          8402 => x"00",
          8403 => x"69",
          8404 => x"20",
          8405 => x"65",
          8406 => x"70",
          8407 => x"00",
          8408 => x"53",
          8409 => x"6e",
          8410 => x"72",
          8411 => x"0a",
          8412 => x"4f",
          8413 => x"20",
          8414 => x"69",
          8415 => x"72",
          8416 => x"74",
          8417 => x"4f",
          8418 => x"20",
          8419 => x"69",
          8420 => x"72",
          8421 => x"74",
          8422 => x"41",
          8423 => x"20",
          8424 => x"69",
          8425 => x"72",
          8426 => x"74",
          8427 => x"41",
          8428 => x"20",
          8429 => x"69",
          8430 => x"72",
          8431 => x"74",
          8432 => x"41",
          8433 => x"20",
          8434 => x"69",
          8435 => x"72",
          8436 => x"74",
          8437 => x"41",
          8438 => x"20",
          8439 => x"69",
          8440 => x"72",
          8441 => x"74",
          8442 => x"65",
          8443 => x"6e",
          8444 => x"70",
          8445 => x"6d",
          8446 => x"2e",
          8447 => x"00",
          8448 => x"6e",
          8449 => x"69",
          8450 => x"74",
          8451 => x"72",
          8452 => x"0a",
          8453 => x"3a",
          8454 => x"61",
          8455 => x"64",
          8456 => x"20",
          8457 => x"74",
          8458 => x"69",
          8459 => x"73",
          8460 => x"61",
          8461 => x"30",
          8462 => x"6c",
          8463 => x"65",
          8464 => x"69",
          8465 => x"61",
          8466 => x"6c",
          8467 => x"0a",
          8468 => x"20",
          8469 => x"61",
          8470 => x"69",
          8471 => x"69",
          8472 => x"00",
          8473 => x"6e",
          8474 => x"61",
          8475 => x"65",
          8476 => x"00",
          8477 => x"61",
          8478 => x"64",
          8479 => x"20",
          8480 => x"74",
          8481 => x"69",
          8482 => x"0a",
          8483 => x"63",
          8484 => x"0a",
          8485 => x"75",
          8486 => x"69",
          8487 => x"6c",
          8488 => x"20",
          8489 => x"65",
          8490 => x"70",
          8491 => x"00",
          8492 => x"6e",
          8493 => x"69",
          8494 => x"69",
          8495 => x"72",
          8496 => x"74",
          8497 => x"00",
          8498 => x"69",
          8499 => x"6c",
          8500 => x"75",
          8501 => x"20",
          8502 => x"6f",
          8503 => x"6e",
          8504 => x"69",
          8505 => x"75",
          8506 => x"20",
          8507 => x"6f",
          8508 => x"78",
          8509 => x"74",
          8510 => x"20",
          8511 => x"65",
          8512 => x"25",
          8513 => x"20",
          8514 => x"0a",
          8515 => x"61",
          8516 => x"6e",
          8517 => x"6f",
          8518 => x"40",
          8519 => x"38",
          8520 => x"2e",
          8521 => x"00",
          8522 => x"61",
          8523 => x"72",
          8524 => x"72",
          8525 => x"20",
          8526 => x"65",
          8527 => x"64",
          8528 => x"00",
          8529 => x"65",
          8530 => x"72",
          8531 => x"67",
          8532 => x"70",
          8533 => x"61",
          8534 => x"6e",
          8535 => x"0a",
          8536 => x"6f",
          8537 => x"72",
          8538 => x"6f",
          8539 => x"67",
          8540 => x"0a",
          8541 => x"50",
          8542 => x"69",
          8543 => x"64",
          8544 => x"73",
          8545 => x"2e",
          8546 => x"00",
          8547 => x"61",
          8548 => x"6f",
          8549 => x"6e",
          8550 => x"00",
          8551 => x"75",
          8552 => x"6e",
          8553 => x"2e",
          8554 => x"6e",
          8555 => x"69",
          8556 => x"69",
          8557 => x"72",
          8558 => x"74",
          8559 => x"2e",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"01",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"f5",
          8572 => x"01",
          8573 => x"01",
          8574 => x"01",
          8575 => x"00",
          8576 => x"00",
          8577 => x"00",
          8578 => x"00",
          8579 => x"01",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"02",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"03",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"04",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"0a",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"0b",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"0c",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"0d",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"0e",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"0f",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"14",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"17",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"18",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"19",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"1a",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"1c",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"1d",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"1e",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"22",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"23",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"24",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"1f",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"20",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"21",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"15",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"16",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"1b",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"25",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"2d",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"2e",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"2b",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"30",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"2f",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"2c",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"26",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"27",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"28",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"29",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"2a",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"3c",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"3d",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"3e",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"3f",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"40",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"50",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"51",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"52",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"53",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"54",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"55",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"64",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"65",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"79",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"78",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"82",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"83",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"84",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"85",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"86",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"87",
          8816 => x"00",
          8817 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"88",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cb",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"fd",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"80",
           281 => x"e2",
           282 => x"00",
           283 => x"9f",
           284 => x"38",
           285 => x"84",
           286 => x"88",
           287 => x"e2",
           288 => x"04",
           289 => x"94",
           290 => x"0d",
           291 => x"08",
           292 => x"52",
           293 => x"05",
           294 => x"de",
           295 => x"70",
           296 => x"85",
           297 => x"0c",
           298 => x"02",
           299 => x"3d",
           300 => x"94",
           301 => x"08",
           302 => x"88",
           303 => x"82",
           304 => x"08",
           305 => x"54",
           306 => x"94",
           307 => x"08",
           308 => x"f9",
           309 => x"0b",
           310 => x"05",
           311 => x"88",
           312 => x"25",
           313 => x"08",
           314 => x"30",
           315 => x"05",
           316 => x"94",
           317 => x"0c",
           318 => x"05",
           319 => x"81",
           320 => x"f4",
           321 => x"08",
           322 => x"94",
           323 => x"0c",
           324 => x"05",
           325 => x"ab",
           326 => x"8c",
           327 => x"94",
           328 => x"0c",
           329 => x"08",
           330 => x"94",
           331 => x"08",
           332 => x"0b",
           333 => x"05",
           334 => x"f0",
           335 => x"08",
           336 => x"80",
           337 => x"8c",
           338 => x"94",
           339 => x"08",
           340 => x"3f",
           341 => x"94",
           342 => x"0c",
           343 => x"fc",
           344 => x"2e",
           345 => x"08",
           346 => x"30",
           347 => x"05",
           348 => x"f8",
           349 => x"88",
           350 => x"3d",
           351 => x"04",
           352 => x"94",
           353 => x"0d",
           354 => x"08",
           355 => x"94",
           356 => x"08",
           357 => x"38",
           358 => x"05",
           359 => x"08",
           360 => x"81",
           361 => x"fc",
           362 => x"08",
           363 => x"80",
           364 => x"94",
           365 => x"08",
           366 => x"8c",
           367 => x"53",
           368 => x"05",
           369 => x"08",
           370 => x"51",
           371 => x"08",
           372 => x"f8",
           373 => x"94",
           374 => x"08",
           375 => x"38",
           376 => x"05",
           377 => x"08",
           378 => x"94",
           379 => x"08",
           380 => x"54",
           381 => x"94",
           382 => x"08",
           383 => x"fd",
           384 => x"0b",
           385 => x"05",
           386 => x"94",
           387 => x"0c",
           388 => x"05",
           389 => x"88",
           390 => x"ac",
           391 => x"fc",
           392 => x"2e",
           393 => x"0b",
           394 => x"05",
           395 => x"38",
           396 => x"05",
           397 => x"08",
           398 => x"94",
           399 => x"08",
           400 => x"fc",
           401 => x"39",
           402 => x"05",
           403 => x"80",
           404 => x"08",
           405 => x"94",
           406 => x"08",
           407 => x"94",
           408 => x"08",
           409 => x"05",
           410 => x"08",
           411 => x"94",
           412 => x"08",
           413 => x"05",
           414 => x"08",
           415 => x"94",
           416 => x"08",
           417 => x"08",
           418 => x"94",
           419 => x"08",
           420 => x"08",
           421 => x"ff",
           422 => x"08",
           423 => x"80",
           424 => x"94",
           425 => x"08",
           426 => x"f4",
           427 => x"8d",
           428 => x"f8",
           429 => x"94",
           430 => x"0c",
           431 => x"f4",
           432 => x"0c",
           433 => x"94",
           434 => x"3d",
           435 => x"0b",
           436 => x"8c",
           437 => x"87",
           438 => x"0c",
           439 => x"c0",
           440 => x"87",
           441 => x"08",
           442 => x"51",
           443 => x"2e",
           444 => x"c0",
           445 => x"51",
           446 => x"87",
           447 => x"08",
           448 => x"06",
           449 => x"38",
           450 => x"8c",
           451 => x"80",
           452 => x"71",
           453 => x"9f",
           454 => x"0b",
           455 => x"33",
           456 => x"3d",
           457 => x"3d",
           458 => x"7d",
           459 => x"80",
           460 => x"0b",
           461 => x"81",
           462 => x"82",
           463 => x"2e",
           464 => x"81",
           465 => x"0b",
           466 => x"8c",
           467 => x"c0",
           468 => x"84",
           469 => x"92",
           470 => x"c0",
           471 => x"70",
           472 => x"81",
           473 => x"53",
           474 => x"a7",
           475 => x"92",
           476 => x"81",
           477 => x"79",
           478 => x"51",
           479 => x"90",
           480 => x"2e",
           481 => x"76",
           482 => x"58",
           483 => x"54",
           484 => x"72",
           485 => x"70",
           486 => x"38",
           487 => x"8c",
           488 => x"ff",
           489 => x"c0",
           490 => x"51",
           491 => x"81",
           492 => x"92",
           493 => x"c0",
           494 => x"70",
           495 => x"51",
           496 => x"80",
           497 => x"80",
           498 => x"70",
           499 => x"81",
           500 => x"87",
           501 => x"08",
           502 => x"2e",
           503 => x"83",
           504 => x"71",
           505 => x"3d",
           506 => x"3d",
           507 => x"11",
           508 => x"71",
           509 => x"88",
           510 => x"84",
           511 => x"fd",
           512 => x"83",
           513 => x"12",
           514 => x"2b",
           515 => x"07",
           516 => x"70",
           517 => x"2b",
           518 => x"07",
           519 => x"53",
           520 => x"52",
           521 => x"04",
           522 => x"79",
           523 => x"9f",
           524 => x"57",
           525 => x"80",
           526 => x"88",
           527 => x"80",
           528 => x"33",
           529 => x"2e",
           530 => x"83",
           531 => x"80",
           532 => x"54",
           533 => x"fe",
           534 => x"88",
           535 => x"08",
           536 => x"3d",
           537 => x"fd",
           538 => x"08",
           539 => x"51",
           540 => x"88",
           541 => x"ff",
           542 => x"39",
           543 => x"82",
           544 => x"06",
           545 => x"2a",
           546 => x"05",
           547 => x"70",
           548 => x"92",
           549 => x"8e",
           550 => x"fe",
           551 => x"08",
           552 => x"55",
           553 => x"55",
           554 => x"89",
           555 => x"fb",
           556 => x"0b",
           557 => x"08",
           558 => x"12",
           559 => x"55",
           560 => x"56",
           561 => x"8d",
           562 => x"33",
           563 => x"94",
           564 => x"57",
           565 => x"0c",
           566 => x"04",
           567 => x"75",
           568 => x"0b",
           569 => x"ac",
           570 => x"51",
           571 => x"83",
           572 => x"06",
           573 => x"14",
           574 => x"3f",
           575 => x"2b",
           576 => x"51",
           577 => x"88",
           578 => x"ff",
           579 => x"88",
           580 => x"0d",
           581 => x"0d",
           582 => x"0b",
           583 => x"55",
           584 => x"23",
           585 => x"53",
           586 => x"88",
           587 => x"08",
           588 => x"38",
           589 => x"39",
           590 => x"73",
           591 => x"83",
           592 => x"06",
           593 => x"14",
           594 => x"8c",
           595 => x"80",
           596 => x"72",
           597 => x"3f",
           598 => x"85",
           599 => x"08",
           600 => x"16",
           601 => x"71",
           602 => x"3d",
           603 => x"3d",
           604 => x"0b",
           605 => x"08",
           606 => x"05",
           607 => x"ff",
           608 => x"57",
           609 => x"2e",
           610 => x"15",
           611 => x"86",
           612 => x"80",
           613 => x"8f",
           614 => x"80",
           615 => x"13",
           616 => x"8c",
           617 => x"72",
           618 => x"0b",
           619 => x"57",
           620 => x"27",
           621 => x"39",
           622 => x"ff",
           623 => x"2a",
           624 => x"a8",
           625 => x"fc",
           626 => x"52",
           627 => x"27",
           628 => x"52",
           629 => x"17",
           630 => x"38",
           631 => x"16",
           632 => x"51",
           633 => x"88",
           634 => x"0c",
           635 => x"80",
           636 => x"0c",
           637 => x"04",
           638 => x"60",
           639 => x"5e",
           640 => x"55",
           641 => x"09",
           642 => x"38",
           643 => x"44",
           644 => x"62",
           645 => x"56",
           646 => x"09",
           647 => x"38",
           648 => x"80",
           649 => x"0c",
           650 => x"51",
           651 => x"26",
           652 => x"51",
           653 => x"88",
           654 => x"7d",
           655 => x"39",
           656 => x"1d",
           657 => x"5a",
           658 => x"a0",
           659 => x"05",
           660 => x"15",
           661 => x"2e",
           662 => x"ef",
           663 => x"59",
           664 => x"08",
           665 => x"81",
           666 => x"ff",
           667 => x"70",
           668 => x"32",
           669 => x"73",
           670 => x"25",
           671 => x"52",
           672 => x"57",
           673 => x"c7",
           674 => x"2e",
           675 => x"83",
           676 => x"77",
           677 => x"07",
           678 => x"2e",
           679 => x"88",
           680 => x"78",
           681 => x"30",
           682 => x"9f",
           683 => x"57",
           684 => x"9b",
           685 => x"8b",
           686 => x"39",
           687 => x"70",
           688 => x"72",
           689 => x"57",
           690 => x"34",
           691 => x"7a",
           692 => x"80",
           693 => x"26",
           694 => x"55",
           695 => x"34",
           696 => x"b1",
           697 => x"80",
           698 => x"54",
           699 => x"85",
           700 => x"06",
           701 => x"1c",
           702 => x"51",
           703 => x"88",
           704 => x"08",
           705 => x"7c",
           706 => x"80",
           707 => x"38",
           708 => x"70",
           709 => x"81",
           710 => x"56",
           711 => x"8b",
           712 => x"08",
           713 => x"5b",
           714 => x"18",
           715 => x"2e",
           716 => x"70",
           717 => x"33",
           718 => x"05",
           719 => x"71",
           720 => x"56",
           721 => x"e2",
           722 => x"75",
           723 => x"38",
           724 => x"9a",
           725 => x"39",
           726 => x"88",
           727 => x"83",
           728 => x"84",
           729 => x"11",
           730 => x"74",
           731 => x"1d",
           732 => x"2a",
           733 => x"51",
           734 => x"89",
           735 => x"92",
           736 => x"8e",
           737 => x"fa",
           738 => x"08",
           739 => x"fd",
           740 => x"88",
           741 => x"0d",
           742 => x"0d",
           743 => x"57",
           744 => x"fe",
           745 => x"76",
           746 => x"3f",
           747 => x"08",
           748 => x"76",
           749 => x"3f",
           750 => x"ff",
           751 => x"82",
           752 => x"d4",
           753 => x"81",
           754 => x"38",
           755 => x"53",
           756 => x"51",
           757 => x"88",
           758 => x"08",
           759 => x"51",
           760 => x"88",
           761 => x"ff",
           762 => x"81",
           763 => x"a9",
           764 => x"80",
           765 => x"52",
           766 => x"aa",
           767 => x"56",
           768 => x"38",
           769 => x"e2",
           770 => x"83",
           771 => x"55",
           772 => x"c6",
           773 => x"81",
           774 => x"0c",
           775 => x"04",
           776 => x"65",
           777 => x"0b",
           778 => x"ac",
           779 => x"3f",
           780 => x"06",
           781 => x"74",
           782 => x"74",
           783 => x"3d",
           784 => x"5a",
           785 => x"88",
           786 => x"06",
           787 => x"2e",
           788 => x"b3",
           789 => x"83",
           790 => x"52",
           791 => x"c6",
           792 => x"ab",
           793 => x"33",
           794 => x"2e",
           795 => x"3d",
           796 => x"f7",
           797 => x"08",
           798 => x"76",
           799 => x"99",
           800 => x"81",
           801 => x"76",
           802 => x"81",
           803 => x"81",
           804 => x"39",
           805 => x"86",
           806 => x"82",
           807 => x"54",
           808 => x"52",
           809 => x"fe",
           810 => x"88",
           811 => x"38",
           812 => x"05",
           813 => x"3f",
           814 => x"ff",
           815 => x"77",
           816 => x"3d",
           817 => x"f6",
           818 => x"08",
           819 => x"05",
           820 => x"29",
           821 => x"ad",
           822 => x"52",
           823 => x"8a",
           824 => x"83",
           825 => x"7a",
           826 => x"0c",
           827 => x"82",
           828 => x"3d",
           829 => x"f5",
           830 => x"08",
           831 => x"95",
           832 => x"51",
           833 => x"88",
           834 => x"ff",
           835 => x"8c",
           836 => x"ef",
           837 => x"e7",
           838 => x"56",
           839 => x"ca",
           840 => x"83",
           841 => x"76",
           842 => x"31",
           843 => x"70",
           844 => x"1d",
           845 => x"71",
           846 => x"5c",
           847 => x"c4",
           848 => x"82",
           849 => x"1b",
           850 => x"e0",
           851 => x"56",
           852 => x"fe",
           853 => x"82",
           854 => x"f6",
           855 => x"38",
           856 => x"39",
           857 => x"80",
           858 => x"38",
           859 => x"76",
           860 => x"81",
           861 => x"95",
           862 => x"51",
           863 => x"88",
           864 => x"0c",
           865 => x"19",
           866 => x"1a",
           867 => x"ff",
           868 => x"1a",
           869 => x"84",
           870 => x"1b",
           871 => x"0b",
           872 => x"78",
           873 => x"9f",
           874 => x"56",
           875 => x"95",
           876 => x"ea",
           877 => x"0b",
           878 => x"08",
           879 => x"74",
           880 => x"df",
           881 => x"81",
           882 => x"3d",
           883 => x"69",
           884 => x"70",
           885 => x"05",
           886 => x"3f",
           887 => x"88",
           888 => x"38",
           889 => x"54",
           890 => x"93",
           891 => x"05",
           892 => x"2a",
           893 => x"51",
           894 => x"80",
           895 => x"83",
           896 => x"75",
           897 => x"3f",
           898 => x"16",
           899 => x"dc",
           900 => x"eb",
           901 => x"9c",
           902 => x"98",
           903 => x"0b",
           904 => x"73",
           905 => x"3d",
           906 => x"3d",
           907 => x"7e",
           908 => x"9f",
           909 => x"5b",
           910 => x"7b",
           911 => x"75",
           912 => x"d1",
           913 => x"33",
           914 => x"84",
           915 => x"2e",
           916 => x"91",
           917 => x"17",
           918 => x"80",
           919 => x"34",
           920 => x"b1",
           921 => x"08",
           922 => x"31",
           923 => x"27",
           924 => x"58",
           925 => x"81",
           926 => x"16",
           927 => x"ff",
           928 => x"74",
           929 => x"82",
           930 => x"05",
           931 => x"06",
           932 => x"06",
           933 => x"9e",
           934 => x"38",
           935 => x"55",
           936 => x"16",
           937 => x"80",
           938 => x"55",
           939 => x"ff",
           940 => x"a4",
           941 => x"16",
           942 => x"f3",
           943 => x"55",
           944 => x"2e",
           945 => x"88",
           946 => x"17",
           947 => x"08",
           948 => x"84",
           949 => x"51",
           950 => x"27",
           951 => x"55",
           952 => x"16",
           953 => x"06",
           954 => x"08",
           955 => x"f0",
           956 => x"08",
           957 => x"98",
           958 => x"98",
           959 => x"75",
           960 => x"16",
           961 => x"78",
           962 => x"e8",
           963 => x"59",
           964 => x"80",
           965 => x"0c",
           966 => x"04",
           967 => x"9b",
           968 => x"0b",
           969 => x"8c",
           970 => x"86",
           971 => x"c0",
           972 => x"8c",
           973 => x"87",
           974 => x"0c",
           975 => x"0b",
           976 => x"94",
           977 => x"51",
           978 => x"88",
           979 => x"9f",
           980 => x"df",
           981 => x"ae",
           982 => x"0b",
           983 => x"c0",
           984 => x"55",
           985 => x"05",
           986 => x"52",
           987 => x"ba",
           988 => x"8d",
           989 => x"73",
           990 => x"38",
           991 => x"e4",
           992 => x"54",
           993 => x"54",
           994 => x"00",
           995 => x"ff",
           996 => x"ff",
           997 => x"ff",
           998 => x"42",
           999 => x"54",
          1000 => x"2e",
          1001 => x"00",
          1002 => x"01",
          2048 => x"0b",
          2049 => x"80",
          2050 => x"80",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"80",
          2058 => x"80",
          2059 => x"0b",
          2060 => x"95",
          2061 => x"80",
          2062 => x"0b",
          2063 => x"b5",
          2064 => x"80",
          2065 => x"0b",
          2066 => x"d5",
          2067 => x"80",
          2068 => x"0b",
          2069 => x"f5",
          2070 => x"80",
          2071 => x"0b",
          2072 => x"95",
          2073 => x"80",
          2074 => x"0b",
          2075 => x"b5",
          2076 => x"80",
          2077 => x"0b",
          2078 => x"d5",
          2079 => x"80",
          2080 => x"0b",
          2081 => x"f5",
          2082 => x"80",
          2083 => x"0b",
          2084 => x"95",
          2085 => x"80",
          2086 => x"0b",
          2087 => x"b5",
          2088 => x"80",
          2089 => x"0b",
          2090 => x"d5",
          2091 => x"80",
          2092 => x"0b",
          2093 => x"f5",
          2094 => x"80",
          2095 => x"0b",
          2096 => x"95",
          2097 => x"80",
          2098 => x"0b",
          2099 => x"b5",
          2100 => x"80",
          2101 => x"0b",
          2102 => x"d5",
          2103 => x"80",
          2104 => x"0b",
          2105 => x"f5",
          2106 => x"80",
          2107 => x"0b",
          2108 => x"95",
          2109 => x"80",
          2110 => x"0b",
          2111 => x"b5",
          2112 => x"80",
          2113 => x"0b",
          2114 => x"d5",
          2115 => x"80",
          2116 => x"0b",
          2117 => x"f5",
          2118 => x"80",
          2119 => x"0b",
          2120 => x"95",
          2121 => x"80",
          2122 => x"0b",
          2123 => x"b5",
          2124 => x"80",
          2125 => x"0b",
          2126 => x"d5",
          2127 => x"80",
          2128 => x"0b",
          2129 => x"f5",
          2130 => x"80",
          2131 => x"00",
          2132 => x"00",
          2133 => x"00",
          2134 => x"00",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"00",
          2177 => x"04",
          2178 => x"0c",
          2179 => x"2d",
          2180 => x"08",
          2181 => x"04",
          2182 => x"0c",
          2183 => x"2d",
          2184 => x"08",
          2185 => x"04",
          2186 => x"0c",
          2187 => x"2d",
          2188 => x"08",
          2189 => x"04",
          2190 => x"0c",
          2191 => x"2d",
          2192 => x"08",
          2193 => x"04",
          2194 => x"0c",
          2195 => x"2d",
          2196 => x"08",
          2197 => x"04",
          2198 => x"0c",
          2199 => x"2d",
          2200 => x"08",
          2201 => x"04",
          2202 => x"0c",
          2203 => x"2d",
          2204 => x"08",
          2205 => x"04",
          2206 => x"0c",
          2207 => x"2d",
          2208 => x"08",
          2209 => x"04",
          2210 => x"0c",
          2211 => x"2d",
          2212 => x"08",
          2213 => x"04",
          2214 => x"0c",
          2215 => x"2d",
          2216 => x"08",
          2217 => x"04",
          2218 => x"0c",
          2219 => x"2d",
          2220 => x"08",
          2221 => x"04",
          2222 => x"0c",
          2223 => x"2d",
          2224 => x"08",
          2225 => x"04",
          2226 => x"0c",
          2227 => x"2d",
          2228 => x"08",
          2229 => x"04",
          2230 => x"0c",
          2231 => x"2d",
          2232 => x"08",
          2233 => x"04",
          2234 => x"0c",
          2235 => x"2d",
          2236 => x"08",
          2237 => x"04",
          2238 => x"0c",
          2239 => x"2d",
          2240 => x"08",
          2241 => x"04",
          2242 => x"0c",
          2243 => x"2d",
          2244 => x"08",
          2245 => x"04",
          2246 => x"0c",
          2247 => x"2d",
          2248 => x"08",
          2249 => x"04",
          2250 => x"0c",
          2251 => x"2d",
          2252 => x"08",
          2253 => x"04",
          2254 => x"0c",
          2255 => x"2d",
          2256 => x"08",
          2257 => x"04",
          2258 => x"0c",
          2259 => x"2d",
          2260 => x"08",
          2261 => x"04",
          2262 => x"0c",
          2263 => x"2d",
          2264 => x"08",
          2265 => x"04",
          2266 => x"0c",
          2267 => x"2d",
          2268 => x"08",
          2269 => x"04",
          2270 => x"0c",
          2271 => x"2d",
          2272 => x"08",
          2273 => x"04",
          2274 => x"0c",
          2275 => x"2d",
          2276 => x"08",
          2277 => x"04",
          2278 => x"0c",
          2279 => x"2d",
          2280 => x"08",
          2281 => x"04",
          2282 => x"0c",
          2283 => x"2d",
          2284 => x"08",
          2285 => x"04",
          2286 => x"0c",
          2287 => x"2d",
          2288 => x"08",
          2289 => x"04",
          2290 => x"0c",
          2291 => x"2d",
          2292 => x"08",
          2293 => x"04",
          2294 => x"0c",
          2295 => x"2d",
          2296 => x"08",
          2297 => x"04",
          2298 => x"0c",
          2299 => x"2d",
          2300 => x"08",
          2301 => x"04",
          2302 => x"0c",
          2303 => x"2d",
          2304 => x"08",
          2305 => x"04",
          2306 => x"0c",
          2307 => x"2d",
          2308 => x"08",
          2309 => x"04",
          2310 => x"0c",
          2311 => x"2d",
          2312 => x"08",
          2313 => x"04",
          2314 => x"0c",
          2315 => x"2d",
          2316 => x"08",
          2317 => x"04",
          2318 => x"0c",
          2319 => x"2d",
          2320 => x"08",
          2321 => x"04",
          2322 => x"0c",
          2323 => x"2d",
          2324 => x"08",
          2325 => x"04",
          2326 => x"0c",
          2327 => x"2d",
          2328 => x"08",
          2329 => x"04",
          2330 => x"0c",
          2331 => x"2d",
          2332 => x"08",
          2333 => x"04",
          2334 => x"0c",
          2335 => x"2d",
          2336 => x"08",
          2337 => x"04",
          2338 => x"0c",
          2339 => x"2d",
          2340 => x"08",
          2341 => x"04",
          2342 => x"0c",
          2343 => x"2d",
          2344 => x"08",
          2345 => x"04",
          2346 => x"0c",
          2347 => x"2d",
          2348 => x"08",
          2349 => x"04",
          2350 => x"0c",
          2351 => x"2d",
          2352 => x"08",
          2353 => x"04",
          2354 => x"0c",
          2355 => x"2d",
          2356 => x"08",
          2357 => x"04",
          2358 => x"0c",
          2359 => x"2d",
          2360 => x"08",
          2361 => x"04",
          2362 => x"0c",
          2363 => x"2d",
          2364 => x"08",
          2365 => x"04",
          2366 => x"0c",
          2367 => x"2d",
          2368 => x"08",
          2369 => x"04",
          2370 => x"0c",
          2371 => x"2d",
          2372 => x"08",
          2373 => x"04",
          2374 => x"70",
          2375 => x"27",
          2376 => x"71",
          2377 => x"53",
          2378 => x"80",
          2379 => x"80",
          2380 => x"81",
          2381 => x"3c",
          2382 => x"d4",
          2383 => x"93",
          2384 => x"3d",
          2385 => x"82",
          2386 => x"8c",
          2387 => x"82",
          2388 => x"88",
          2389 => x"80",
          2390 => x"93",
          2391 => x"82",
          2392 => x"54",
          2393 => x"82",
          2394 => x"04",
          2395 => x"08",
          2396 => x"d4",
          2397 => x"0d",
          2398 => x"93",
          2399 => x"05",
          2400 => x"93",
          2401 => x"05",
          2402 => x"3f",
          2403 => x"08",
          2404 => x"c8",
          2405 => x"3d",
          2406 => x"d4",
          2407 => x"93",
          2408 => x"82",
          2409 => x"fd",
          2410 => x"0b",
          2411 => x"08",
          2412 => x"80",
          2413 => x"d4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"82",
          2417 => x"88",
          2418 => x"b9",
          2419 => x"d4",
          2420 => x"08",
          2421 => x"38",
          2422 => x"93",
          2423 => x"05",
          2424 => x"38",
          2425 => x"08",
          2426 => x"10",
          2427 => x"08",
          2428 => x"82",
          2429 => x"fc",
          2430 => x"82",
          2431 => x"fc",
          2432 => x"b8",
          2433 => x"d4",
          2434 => x"08",
          2435 => x"e1",
          2436 => x"d4",
          2437 => x"08",
          2438 => x"08",
          2439 => x"26",
          2440 => x"93",
          2441 => x"05",
          2442 => x"d4",
          2443 => x"08",
          2444 => x"d4",
          2445 => x"0c",
          2446 => x"08",
          2447 => x"82",
          2448 => x"fc",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"93",
          2452 => x"05",
          2453 => x"82",
          2454 => x"fc",
          2455 => x"93",
          2456 => x"05",
          2457 => x"82",
          2458 => x"8c",
          2459 => x"95",
          2460 => x"d4",
          2461 => x"08",
          2462 => x"38",
          2463 => x"08",
          2464 => x"70",
          2465 => x"08",
          2466 => x"51",
          2467 => x"93",
          2468 => x"05",
          2469 => x"93",
          2470 => x"05",
          2471 => x"93",
          2472 => x"05",
          2473 => x"c8",
          2474 => x"0d",
          2475 => x"0c",
          2476 => x"0d",
          2477 => x"02",
          2478 => x"05",
          2479 => x"53",
          2480 => x"27",
          2481 => x"83",
          2482 => x"80",
          2483 => x"ff",
          2484 => x"ff",
          2485 => x"73",
          2486 => x"05",
          2487 => x"12",
          2488 => x"2e",
          2489 => x"ef",
          2490 => x"93",
          2491 => x"3d",
          2492 => x"74",
          2493 => x"07",
          2494 => x"2b",
          2495 => x"51",
          2496 => x"a5",
          2497 => x"70",
          2498 => x"0c",
          2499 => x"84",
          2500 => x"72",
          2501 => x"05",
          2502 => x"71",
          2503 => x"53",
          2504 => x"52",
          2505 => x"dd",
          2506 => x"27",
          2507 => x"71",
          2508 => x"53",
          2509 => x"52",
          2510 => x"f2",
          2511 => x"ff",
          2512 => x"3d",
          2513 => x"70",
          2514 => x"06",
          2515 => x"70",
          2516 => x"73",
          2517 => x"56",
          2518 => x"08",
          2519 => x"38",
          2520 => x"52",
          2521 => x"81",
          2522 => x"54",
          2523 => x"9d",
          2524 => x"55",
          2525 => x"09",
          2526 => x"38",
          2527 => x"14",
          2528 => x"81",
          2529 => x"56",
          2530 => x"e5",
          2531 => x"55",
          2532 => x"06",
          2533 => x"06",
          2534 => x"82",
          2535 => x"52",
          2536 => x"0d",
          2537 => x"70",
          2538 => x"ff",
          2539 => x"f8",
          2540 => x"80",
          2541 => x"51",
          2542 => x"84",
          2543 => x"71",
          2544 => x"54",
          2545 => x"2e",
          2546 => x"75",
          2547 => x"94",
          2548 => x"82",
          2549 => x"87",
          2550 => x"fe",
          2551 => x"70",
          2552 => x"88",
          2553 => x"9b",
          2554 => x"c8",
          2555 => x"06",
          2556 => x"14",
          2557 => x"73",
          2558 => x"71",
          2559 => x"0c",
          2560 => x"04",
          2561 => x"76",
          2562 => x"53",
          2563 => x"80",
          2564 => x"38",
          2565 => x"70",
          2566 => x"81",
          2567 => x"81",
          2568 => x"52",
          2569 => x"2e",
          2570 => x"52",
          2571 => x"12",
          2572 => x"33",
          2573 => x"a0",
          2574 => x"81",
          2575 => x"70",
          2576 => x"06",
          2577 => x"e6",
          2578 => x"51",
          2579 => x"09",
          2580 => x"38",
          2581 => x"81",
          2582 => x"71",
          2583 => x"51",
          2584 => x"c8",
          2585 => x"0d",
          2586 => x"0d",
          2587 => x"08",
          2588 => x"38",
          2589 => x"05",
          2590 => x"99",
          2591 => x"93",
          2592 => x"38",
          2593 => x"39",
          2594 => x"82",
          2595 => x"86",
          2596 => x"f5",
          2597 => x"82",
          2598 => x"05",
          2599 => x"5b",
          2600 => x"81",
          2601 => x"1c",
          2602 => x"5a",
          2603 => x"9e",
          2604 => x"38",
          2605 => x"5a",
          2606 => x"97",
          2607 => x"38",
          2608 => x"5a",
          2609 => x"bb",
          2610 => x"38",
          2611 => x"5a",
          2612 => x"bb",
          2613 => x"38",
          2614 => x"5a",
          2615 => x"87",
          2616 => x"80",
          2617 => x"22",
          2618 => x"79",
          2619 => x"80",
          2620 => x"1c",
          2621 => x"1c",
          2622 => x"1c",
          2623 => x"1c",
          2624 => x"1c",
          2625 => x"1c",
          2626 => x"1c",
          2627 => x"22",
          2628 => x"a8",
          2629 => x"3f",
          2630 => x"9c",
          2631 => x"0c",
          2632 => x"c0",
          2633 => x"82",
          2634 => x"c0",
          2635 => x"83",
          2636 => x"c0",
          2637 => x"84",
          2638 => x"c0",
          2639 => x"85",
          2640 => x"c0",
          2641 => x"86",
          2642 => x"c0",
          2643 => x"88",
          2644 => x"c0",
          2645 => x"8a",
          2646 => x"c0",
          2647 => x"80",
          2648 => x"5b",
          2649 => x"c8",
          2650 => x"0d",
          2651 => x"0d",
          2652 => x"c0",
          2653 => x"81",
          2654 => x"c0",
          2655 => x"5b",
          2656 => x"87",
          2657 => x"08",
          2658 => x"1b",
          2659 => x"98",
          2660 => x"7a",
          2661 => x"87",
          2662 => x"08",
          2663 => x"1b",
          2664 => x"98",
          2665 => x"7a",
          2666 => x"87",
          2667 => x"08",
          2668 => x"1b",
          2669 => x"98",
          2670 => x"7a",
          2671 => x"87",
          2672 => x"08",
          2673 => x"1b",
          2674 => x"0c",
          2675 => x"59",
          2676 => x"58",
          2677 => x"57",
          2678 => x"56",
          2679 => x"55",
          2680 => x"54",
          2681 => x"53",
          2682 => x"81",
          2683 => x"92",
          2684 => x"3d",
          2685 => x"3d",
          2686 => x"05",
          2687 => x"70",
          2688 => x"51",
          2689 => x"0b",
          2690 => x"34",
          2691 => x"04",
          2692 => x"75",
          2693 => x"8b",
          2694 => x"54",
          2695 => x"84",
          2696 => x"2e",
          2697 => x"c0",
          2698 => x"70",
          2699 => x"2a",
          2700 => x"51",
          2701 => x"80",
          2702 => x"71",
          2703 => x"81",
          2704 => x"70",
          2705 => x"96",
          2706 => x"70",
          2707 => x"51",
          2708 => x"8d",
          2709 => x"2a",
          2710 => x"51",
          2711 => x"bc",
          2712 => x"82",
          2713 => x"51",
          2714 => x"80",
          2715 => x"2e",
          2716 => x"c0",
          2717 => x"73",
          2718 => x"82",
          2719 => x"85",
          2720 => x"fd",
          2721 => x"97",
          2722 => x"0b",
          2723 => x"33",
          2724 => x"c0",
          2725 => x"72",
          2726 => x"38",
          2727 => x"94",
          2728 => x"70",
          2729 => x"81",
          2730 => x"52",
          2731 => x"8c",
          2732 => x"2a",
          2733 => x"51",
          2734 => x"38",
          2735 => x"81",
          2736 => x"06",
          2737 => x"80",
          2738 => x"71",
          2739 => x"81",
          2740 => x"70",
          2741 => x"0b",
          2742 => x"c0",
          2743 => x"c0",
          2744 => x"70",
          2745 => x"38",
          2746 => x"90",
          2747 => x"0c",
          2748 => x"04",
          2749 => x"77",
          2750 => x"33",
          2751 => x"76",
          2752 => x"38",
          2753 => x"05",
          2754 => x"0b",
          2755 => x"33",
          2756 => x"c0",
          2757 => x"72",
          2758 => x"38",
          2759 => x"94",
          2760 => x"70",
          2761 => x"81",
          2762 => x"52",
          2763 => x"8c",
          2764 => x"2a",
          2765 => x"51",
          2766 => x"38",
          2767 => x"81",
          2768 => x"06",
          2769 => x"80",
          2770 => x"71",
          2771 => x"81",
          2772 => x"70",
          2773 => x"0b",
          2774 => x"c0",
          2775 => x"c0",
          2776 => x"70",
          2777 => x"38",
          2778 => x"90",
          2779 => x"0c",
          2780 => x"33",
          2781 => x"ff",
          2782 => x"82",
          2783 => x"87",
          2784 => x"ff",
          2785 => x"0b",
          2786 => x"33",
          2787 => x"94",
          2788 => x"80",
          2789 => x"87",
          2790 => x"51",
          2791 => x"82",
          2792 => x"06",
          2793 => x"70",
          2794 => x"38",
          2795 => x"8b",
          2796 => x"87",
          2797 => x"52",
          2798 => x"86",
          2799 => x"94",
          2800 => x"08",
          2801 => x"06",
          2802 => x"0c",
          2803 => x"0d",
          2804 => x"0d",
          2805 => x"8b",
          2806 => x"87",
          2807 => x"52",
          2808 => x"86",
          2809 => x"94",
          2810 => x"08",
          2811 => x"70",
          2812 => x"51",
          2813 => x"70",
          2814 => x"38",
          2815 => x"8b",
          2816 => x"87",
          2817 => x"52",
          2818 => x"86",
          2819 => x"94",
          2820 => x"08",
          2821 => x"70",
          2822 => x"53",
          2823 => x"93",
          2824 => x"3d",
          2825 => x"3d",
          2826 => x"9e",
          2827 => x"70",
          2828 => x"06",
          2829 => x"70",
          2830 => x"9f",
          2831 => x"c4",
          2832 => x"9e",
          2833 => x"0c",
          2834 => x"c0",
          2835 => x"71",
          2836 => x"11",
          2837 => x"8c",
          2838 => x"52",
          2839 => x"c0",
          2840 => x"71",
          2841 => x"11",
          2842 => x"94",
          2843 => x"52",
          2844 => x"c0",
          2845 => x"71",
          2846 => x"11",
          2847 => x"a4",
          2848 => x"52",
          2849 => x"c0",
          2850 => x"71",
          2851 => x"11",
          2852 => x"ac",
          2853 => x"52",
          2854 => x"52",
          2855 => x"23",
          2856 => x"c0",
          2857 => x"71",
          2858 => x"0b",
          2859 => x"ad",
          2860 => x"0b",
          2861 => x"88",
          2862 => x"80",
          2863 => x"53",
          2864 => x"83",
          2865 => x"72",
          2866 => x"0b",
          2867 => x"88",
          2868 => x"80",
          2869 => x"52",
          2870 => x"2e",
          2871 => x"52",
          2872 => x"f2",
          2873 => x"87",
          2874 => x"08",
          2875 => x"80",
          2876 => x"52",
          2877 => x"83",
          2878 => x"71",
          2879 => x"34",
          2880 => x"c0",
          2881 => x"70",
          2882 => x"51",
          2883 => x"80",
          2884 => x"81",
          2885 => x"8b",
          2886 => x"0b",
          2887 => x"88",
          2888 => x"80",
          2889 => x"52",
          2890 => x"83",
          2891 => x"71",
          2892 => x"34",
          2893 => x"c0",
          2894 => x"70",
          2895 => x"51",
          2896 => x"80",
          2897 => x"81",
          2898 => x"8b",
          2899 => x"0b",
          2900 => x"88",
          2901 => x"80",
          2902 => x"52",
          2903 => x"83",
          2904 => x"71",
          2905 => x"34",
          2906 => x"c0",
          2907 => x"70",
          2908 => x"51",
          2909 => x"80",
          2910 => x"81",
          2911 => x"8b",
          2912 => x"8b",
          2913 => x"c0",
          2914 => x"08",
          2915 => x"06",
          2916 => x"51",
          2917 => x"70",
          2918 => x"05",
          2919 => x"54",
          2920 => x"70",
          2921 => x"52",
          2922 => x"2e",
          2923 => x"52",
          2924 => x"80",
          2925 => x"9e",
          2926 => x"88",
          2927 => x"52",
          2928 => x"83",
          2929 => x"71",
          2930 => x"34",
          2931 => x"88",
          2932 => x"06",
          2933 => x"82",
          2934 => x"85",
          2935 => x"fc",
          2936 => x"f6",
          2937 => x"be",
          2938 => x"f0",
          2939 => x"80",
          2940 => x"81",
          2941 => x"84",
          2942 => x"f6",
          2943 => x"a6",
          2944 => x"f1",
          2945 => x"55",
          2946 => x"91",
          2947 => x"08",
          2948 => x"c4",
          2949 => x"f7",
          2950 => x"84",
          2951 => x"f2",
          2952 => x"55",
          2953 => x"90",
          2954 => x"08",
          2955 => x"08",
          2956 => x"a8",
          2957 => x"3f",
          2958 => x"70",
          2959 => x"73",
          2960 => x"15",
          2961 => x"80",
          2962 => x"82",
          2963 => x"08",
          2964 => x"08",
          2965 => x"f7",
          2966 => x"c4",
          2967 => x"f5",
          2968 => x"80",
          2969 => x"81",
          2970 => x"83",
          2971 => x"8b",
          2972 => x"73",
          2973 => x"38",
          2974 => x"51",
          2975 => x"82",
          2976 => x"54",
          2977 => x"88",
          2978 => x"88",
          2979 => x"3f",
          2980 => x"70",
          2981 => x"73",
          2982 => x"38",
          2983 => x"52",
          2984 => x"51",
          2985 => x"82",
          2986 => x"54",
          2987 => x"88",
          2988 => x"b4",
          2989 => x"3f",
          2990 => x"70",
          2991 => x"73",
          2992 => x"38",
          2993 => x"52",
          2994 => x"51",
          2995 => x"81",
          2996 => x"82",
          2997 => x"8b",
          2998 => x"70",
          2999 => x"08",
          3000 => x"f8",
          3001 => x"88",
          3002 => x"08",
          3003 => x"a0",
          3004 => x"3f",
          3005 => x"52",
          3006 => x"51",
          3007 => x"8c",
          3008 => x"81",
          3009 => x"88",
          3010 => x"15",
          3011 => x"fa",
          3012 => x"8c",
          3013 => x"0d",
          3014 => x"0d",
          3015 => x"33",
          3016 => x"26",
          3017 => x"10",
          3018 => x"81",
          3019 => x"52",
          3020 => x"81",
          3021 => x"f7",
          3022 => x"39",
          3023 => x"51",
          3024 => x"a3",
          3025 => x"d0",
          3026 => x"3f",
          3027 => x"fa",
          3028 => x"a0",
          3029 => x"81",
          3030 => x"f7",
          3031 => x"39",
          3032 => x"51",
          3033 => x"83",
          3034 => x"71",
          3035 => x"04",
          3036 => x"c0",
          3037 => x"04",
          3038 => x"87",
          3039 => x"70",
          3040 => x"80",
          3041 => x"74",
          3042 => x"8c",
          3043 => x"0c",
          3044 => x"04",
          3045 => x"87",
          3046 => x"70",
          3047 => x"80",
          3048 => x"72",
          3049 => x"70",
          3050 => x"08",
          3051 => x"8c",
          3052 => x"0c",
          3053 => x"0d",
          3054 => x"80",
          3055 => x"96",
          3056 => x"fe",
          3057 => x"93",
          3058 => x"72",
          3059 => x"81",
          3060 => x"8d",
          3061 => x"82",
          3062 => x"80",
          3063 => x"82",
          3064 => x"52",
          3065 => x"82",
          3066 => x"81",
          3067 => x"e0",
          3068 => x"82",
          3069 => x"80",
          3070 => x"72",
          3071 => x"d8",
          3072 => x"2d",
          3073 => x"04",
          3074 => x"02",
          3075 => x"82",
          3076 => x"76",
          3077 => x"0c",
          3078 => x"a7",
          3079 => x"93",
          3080 => x"3d",
          3081 => x"3d",
          3082 => x"33",
          3083 => x"80",
          3084 => x"72",
          3085 => x"54",
          3086 => x"87",
          3087 => x"52",
          3088 => x"84",
          3089 => x"fd",
          3090 => x"82",
          3091 => x"77",
          3092 => x"0c",
          3093 => x"55",
          3094 => x"2e",
          3095 => x"70",
          3096 => x"33",
          3097 => x"3f",
          3098 => x"71",
          3099 => x"82",
          3100 => x"85",
          3101 => x"ec",
          3102 => x"68",
          3103 => x"70",
          3104 => x"33",
          3105 => x"2e",
          3106 => x"75",
          3107 => x"38",
          3108 => x"af",
          3109 => x"80",
          3110 => x"81",
          3111 => x"58",
          3112 => x"b0",
          3113 => x"06",
          3114 => x"79",
          3115 => x"5b",
          3116 => x"92",
          3117 => x"2e",
          3118 => x"8a",
          3119 => x"70",
          3120 => x"33",
          3121 => x"aa",
          3122 => x"06",
          3123 => x"84",
          3124 => x"7b",
          3125 => x"5d",
          3126 => x"5d",
          3127 => x"d0",
          3128 => x"89",
          3129 => x"79",
          3130 => x"d0",
          3131 => x"81",
          3132 => x"d0",
          3133 => x"5a",
          3134 => x"eb",
          3135 => x"ec",
          3136 => x"70",
          3137 => x"25",
          3138 => x"32",
          3139 => x"72",
          3140 => x"73",
          3141 => x"52",
          3142 => x"73",
          3143 => x"38",
          3144 => x"79",
          3145 => x"5b",
          3146 => x"75",
          3147 => x"ec",
          3148 => x"80",
          3149 => x"89",
          3150 => x"70",
          3151 => x"56",
          3152 => x"15",
          3153 => x"26",
          3154 => x"72",
          3155 => x"f0",
          3156 => x"72",
          3157 => x"84",
          3158 => x"57",
          3159 => x"75",
          3160 => x"72",
          3161 => x"38",
          3162 => x"16",
          3163 => x"54",
          3164 => x"38",
          3165 => x"70",
          3166 => x"53",
          3167 => x"73",
          3168 => x"53",
          3169 => x"99",
          3170 => x"2a",
          3171 => x"a0",
          3172 => x"3f",
          3173 => x"73",
          3174 => x"53",
          3175 => x"ef",
          3176 => x"fd",
          3177 => x"81",
          3178 => x"72",
          3179 => x"ce",
          3180 => x"fc",
          3181 => x"81",
          3182 => x"79",
          3183 => x"38",
          3184 => x"7b",
          3185 => x"12",
          3186 => x"53",
          3187 => x"fd",
          3188 => x"5b",
          3189 => x"5b",
          3190 => x"5b",
          3191 => x"5b",
          3192 => x"51",
          3193 => x"fd",
          3194 => x"82",
          3195 => x"06",
          3196 => x"80",
          3197 => x"7b",
          3198 => x"08",
          3199 => x"9c",
          3200 => x"c4",
          3201 => x"06",
          3202 => x"84",
          3203 => x"59",
          3204 => x"39",
          3205 => x"71",
          3206 => x"53",
          3207 => x"32",
          3208 => x"72",
          3209 => x"70",
          3210 => x"06",
          3211 => x"53",
          3212 => x"88",
          3213 => x"7d",
          3214 => x"57",
          3215 => x"52",
          3216 => x"a8",
          3217 => x"c8",
          3218 => x"06",
          3219 => x"52",
          3220 => x"3f",
          3221 => x"08",
          3222 => x"27",
          3223 => x"a7",
          3224 => x"ff",
          3225 => x"54",
          3226 => x"2e",
          3227 => x"14",
          3228 => x"06",
          3229 => x"3d",
          3230 => x"05",
          3231 => x"54",
          3232 => x"81",
          3233 => x"70",
          3234 => x"2a",
          3235 => x"27",
          3236 => x"54",
          3237 => x"a6",
          3238 => x"2a",
          3239 => x"51",
          3240 => x"2e",
          3241 => x"3d",
          3242 => x"05",
          3243 => x"34",
          3244 => x"77",
          3245 => x"54",
          3246 => x"72",
          3247 => x"55",
          3248 => x"70",
          3249 => x"53",
          3250 => x"73",
          3251 => x"53",
          3252 => x"99",
          3253 => x"2a",
          3254 => x"74",
          3255 => x"3f",
          3256 => x"73",
          3257 => x"53",
          3258 => x"ef",
          3259 => x"97",
          3260 => x"11",
          3261 => x"54",
          3262 => x"3f",
          3263 => x"73",
          3264 => x"53",
          3265 => x"fa",
          3266 => x"51",
          3267 => x"73",
          3268 => x"53",
          3269 => x"f2",
          3270 => x"39",
          3271 => x"04",
          3272 => x"86",
          3273 => x"84",
          3274 => x"55",
          3275 => x"fa",
          3276 => x"3d",
          3277 => x"3d",
          3278 => x"93",
          3279 => x"3d",
          3280 => x"75",
          3281 => x"3f",
          3282 => x"08",
          3283 => x"34",
          3284 => x"93",
          3285 => x"3d",
          3286 => x"3d",
          3287 => x"d8",
          3288 => x"93",
          3289 => x"3d",
          3290 => x"77",
          3291 => x"87",
          3292 => x"93",
          3293 => x"3d",
          3294 => x"3d",
          3295 => x"57",
          3296 => x"82",
          3297 => x"73",
          3298 => x"38",
          3299 => x"53",
          3300 => x"80",
          3301 => x"dc",
          3302 => x"2d",
          3303 => x"08",
          3304 => x"54",
          3305 => x"e6",
          3306 => x"2e",
          3307 => x"73",
          3308 => x"30",
          3309 => x"78",
          3310 => x"72",
          3311 => x"52",
          3312 => x"72",
          3313 => x"38",
          3314 => x"81",
          3315 => x"55",
          3316 => x"c1",
          3317 => x"25",
          3318 => x"ff",
          3319 => x"72",
          3320 => x"38",
          3321 => x"73",
          3322 => x"15",
          3323 => x"06",
          3324 => x"cf",
          3325 => x"39",
          3326 => x"80",
          3327 => x"51",
          3328 => x"81",
          3329 => x"93",
          3330 => x"3d",
          3331 => x"3d",
          3332 => x"dc",
          3333 => x"93",
          3334 => x"53",
          3335 => x"fe",
          3336 => x"82",
          3337 => x"84",
          3338 => x"f8",
          3339 => x"7c",
          3340 => x"70",
          3341 => x"08",
          3342 => x"54",
          3343 => x"2e",
          3344 => x"92",
          3345 => x"81",
          3346 => x"74",
          3347 => x"55",
          3348 => x"2e",
          3349 => x"ad",
          3350 => x"06",
          3351 => x"75",
          3352 => x"0c",
          3353 => x"33",
          3354 => x"73",
          3355 => x"81",
          3356 => x"38",
          3357 => x"05",
          3358 => x"08",
          3359 => x"53",
          3360 => x"2e",
          3361 => x"80",
          3362 => x"81",
          3363 => x"90",
          3364 => x"76",
          3365 => x"70",
          3366 => x"57",
          3367 => x"82",
          3368 => x"05",
          3369 => x"08",
          3370 => x"54",
          3371 => x"81",
          3372 => x"27",
          3373 => x"d0",
          3374 => x"56",
          3375 => x"73",
          3376 => x"80",
          3377 => x"14",
          3378 => x"72",
          3379 => x"e8",
          3380 => x"80",
          3381 => x"39",
          3382 => x"dc",
          3383 => x"80",
          3384 => x"27",
          3385 => x"80",
          3386 => x"89",
          3387 => x"70",
          3388 => x"55",
          3389 => x"70",
          3390 => x"55",
          3391 => x"27",
          3392 => x"14",
          3393 => x"06",
          3394 => x"74",
          3395 => x"73",
          3396 => x"38",
          3397 => x"14",
          3398 => x"05",
          3399 => x"08",
          3400 => x"54",
          3401 => x"26",
          3402 => x"77",
          3403 => x"38",
          3404 => x"75",
          3405 => x"56",
          3406 => x"c8",
          3407 => x"0d",
          3408 => x"0d",
          3409 => x"55",
          3410 => x"0c",
          3411 => x"33",
          3412 => x"73",
          3413 => x"81",
          3414 => x"74",
          3415 => x"75",
          3416 => x"70",
          3417 => x"73",
          3418 => x"38",
          3419 => x"09",
          3420 => x"38",
          3421 => x"11",
          3422 => x"08",
          3423 => x"54",
          3424 => x"2e",
          3425 => x"80",
          3426 => x"08",
          3427 => x"0c",
          3428 => x"33",
          3429 => x"80",
          3430 => x"38",
          3431 => x"2e",
          3432 => x"a1",
          3433 => x"81",
          3434 => x"75",
          3435 => x"56",
          3436 => x"c1",
          3437 => x"08",
          3438 => x"0c",
          3439 => x"33",
          3440 => x"b1",
          3441 => x"a0",
          3442 => x"82",
          3443 => x"53",
          3444 => x"57",
          3445 => x"9d",
          3446 => x"39",
          3447 => x"80",
          3448 => x"26",
          3449 => x"8b",
          3450 => x"80",
          3451 => x"56",
          3452 => x"8a",
          3453 => x"a0",
          3454 => x"c5",
          3455 => x"74",
          3456 => x"e0",
          3457 => x"ff",
          3458 => x"d0",
          3459 => x"ff",
          3460 => x"90",
          3461 => x"38",
          3462 => x"81",
          3463 => x"53",
          3464 => x"c5",
          3465 => x"27",
          3466 => x"76",
          3467 => x"08",
          3468 => x"0c",
          3469 => x"33",
          3470 => x"73",
          3471 => x"bd",
          3472 => x"2e",
          3473 => x"30",
          3474 => x"0c",
          3475 => x"82",
          3476 => x"8a",
          3477 => x"ff",
          3478 => x"8f",
          3479 => x"81",
          3480 => x"26",
          3481 => x"8c",
          3482 => x"52",
          3483 => x"c8",
          3484 => x"0d",
          3485 => x"0d",
          3486 => x"33",
          3487 => x"9b",
          3488 => x"53",
          3489 => x"81",
          3490 => x"38",
          3491 => x"87",
          3492 => x"05",
          3493 => x"73",
          3494 => x"38",
          3495 => x"71",
          3496 => x"90",
          3497 => x"92",
          3498 => x"81",
          3499 => x"0b",
          3500 => x"8c",
          3501 => x"87",
          3502 => x"54",
          3503 => x"82",
          3504 => x"70",
          3505 => x"38",
          3506 => x"70",
          3507 => x"90",
          3508 => x"92",
          3509 => x"08",
          3510 => x"06",
          3511 => x"92",
          3512 => x"98",
          3513 => x"70",
          3514 => x"38",
          3515 => x"84",
          3516 => x"8c",
          3517 => x"51",
          3518 => x"c8",
          3519 => x"0d",
          3520 => x"0d",
          3521 => x"02",
          3522 => x"c3",
          3523 => x"41",
          3524 => x"73",
          3525 => x"bf",
          3526 => x"c8",
          3527 => x"7b",
          3528 => x"81",
          3529 => x"70",
          3530 => x"c0",
          3531 => x"84",
          3532 => x"92",
          3533 => x"c0",
          3534 => x"72",
          3535 => x"5b",
          3536 => x"0c",
          3537 => x"80",
          3538 => x"0c",
          3539 => x"0c",
          3540 => x"85",
          3541 => x"06",
          3542 => x"71",
          3543 => x"38",
          3544 => x"71",
          3545 => x"05",
          3546 => x"17",
          3547 => x"06",
          3548 => x"2e",
          3549 => x"08",
          3550 => x"38",
          3551 => x"71",
          3552 => x"38",
          3553 => x"2e",
          3554 => x"75",
          3555 => x"92",
          3556 => x"72",
          3557 => x"06",
          3558 => x"f7",
          3559 => x"5b",
          3560 => x"80",
          3561 => x"70",
          3562 => x"5f",
          3563 => x"80",
          3564 => x"73",
          3565 => x"06",
          3566 => x"38",
          3567 => x"ff",
          3568 => x"fc",
          3569 => x"52",
          3570 => x"83",
          3571 => x"71",
          3572 => x"93",
          3573 => x"3d",
          3574 => x"3d",
          3575 => x"64",
          3576 => x"bf",
          3577 => x"40",
          3578 => x"73",
          3579 => x"e7",
          3580 => x"c8",
          3581 => x"7a",
          3582 => x"81",
          3583 => x"5c",
          3584 => x"8c",
          3585 => x"87",
          3586 => x"11",
          3587 => x"84",
          3588 => x"5b",
          3589 => x"85",
          3590 => x"c0",
          3591 => x"7b",
          3592 => x"82",
          3593 => x"53",
          3594 => x"84",
          3595 => x"06",
          3596 => x"71",
          3597 => x"38",
          3598 => x"05",
          3599 => x"0c",
          3600 => x"73",
          3601 => x"81",
          3602 => x"71",
          3603 => x"38",
          3604 => x"71",
          3605 => x"08",
          3606 => x"2e",
          3607 => x"84",
          3608 => x"38",
          3609 => x"87",
          3610 => x"1d",
          3611 => x"70",
          3612 => x"52",
          3613 => x"ff",
          3614 => x"39",
          3615 => x"81",
          3616 => x"80",
          3617 => x"52",
          3618 => x"90",
          3619 => x"80",
          3620 => x"71",
          3621 => x"7c",
          3622 => x"38",
          3623 => x"80",
          3624 => x"80",
          3625 => x"81",
          3626 => x"73",
          3627 => x"0c",
          3628 => x"04",
          3629 => x"7d",
          3630 => x"af",
          3631 => x"88",
          3632 => x"33",
          3633 => x"56",
          3634 => x"3f",
          3635 => x"08",
          3636 => x"83",
          3637 => x"38",
          3638 => x"74",
          3639 => x"72",
          3640 => x"38",
          3641 => x"8a",
          3642 => x"72",
          3643 => x"38",
          3644 => x"90",
          3645 => x"92",
          3646 => x"08",
          3647 => x"39",
          3648 => x"76",
          3649 => x"8b",
          3650 => x"76",
          3651 => x"83",
          3652 => x"73",
          3653 => x"0c",
          3654 => x"04",
          3655 => x"73",
          3656 => x"12",
          3657 => x"2b",
          3658 => x"93",
          3659 => x"52",
          3660 => x"0d",
          3661 => x"0d",
          3662 => x"33",
          3663 => x"71",
          3664 => x"88",
          3665 => x"14",
          3666 => x"74",
          3667 => x"2b",
          3668 => x"c8",
          3669 => x"56",
          3670 => x"3d",
          3671 => x"3d",
          3672 => x"84",
          3673 => x"22",
          3674 => x"72",
          3675 => x"54",
          3676 => x"2a",
          3677 => x"34",
          3678 => x"04",
          3679 => x"73",
          3680 => x"70",
          3681 => x"05",
          3682 => x"88",
          3683 => x"72",
          3684 => x"54",
          3685 => x"2a",
          3686 => x"70",
          3687 => x"34",
          3688 => x"51",
          3689 => x"83",
          3690 => x"fe",
          3691 => x"75",
          3692 => x"51",
          3693 => x"93",
          3694 => x"81",
          3695 => x"73",
          3696 => x"55",
          3697 => x"51",
          3698 => x"84",
          3699 => x"fe",
          3700 => x"77",
          3701 => x"53",
          3702 => x"81",
          3703 => x"ff",
          3704 => x"f4",
          3705 => x"0d",
          3706 => x"0d",
          3707 => x"56",
          3708 => x"70",
          3709 => x"33",
          3710 => x"05",
          3711 => x"71",
          3712 => x"56",
          3713 => x"72",
          3714 => x"38",
          3715 => x"e2",
          3716 => x"93",
          3717 => x"3d",
          3718 => x"3d",
          3719 => x"71",
          3720 => x"52",
          3721 => x"99",
          3722 => x"2e",
          3723 => x"12",
          3724 => x"52",
          3725 => x"89",
          3726 => x"2e",
          3727 => x"ee",
          3728 => x"82",
          3729 => x"84",
          3730 => x"80",
          3731 => x"c8",
          3732 => x"0b",
          3733 => x"0c",
          3734 => x"0d",
          3735 => x"0b",
          3736 => x"56",
          3737 => x"2e",
          3738 => x"81",
          3739 => x"08",
          3740 => x"70",
          3741 => x"33",
          3742 => x"de",
          3743 => x"c8",
          3744 => x"09",
          3745 => x"38",
          3746 => x"08",
          3747 => x"b0",
          3748 => x"17",
          3749 => x"74",
          3750 => x"27",
          3751 => x"16",
          3752 => x"82",
          3753 => x"06",
          3754 => x"54",
          3755 => x"9c",
          3756 => x"53",
          3757 => x"16",
          3758 => x"9e",
          3759 => x"81",
          3760 => x"93",
          3761 => x"3d",
          3762 => x"3d",
          3763 => x"56",
          3764 => x"b0",
          3765 => x"2e",
          3766 => x"51",
          3767 => x"82",
          3768 => x"56",
          3769 => x"08",
          3770 => x"54",
          3771 => x"17",
          3772 => x"33",
          3773 => x"3f",
          3774 => x"08",
          3775 => x"38",
          3776 => x"56",
          3777 => x"0c",
          3778 => x"c8",
          3779 => x"0d",
          3780 => x"0d",
          3781 => x"57",
          3782 => x"82",
          3783 => x"58",
          3784 => x"08",
          3785 => x"76",
          3786 => x"83",
          3787 => x"06",
          3788 => x"84",
          3789 => x"78",
          3790 => x"81",
          3791 => x"38",
          3792 => x"82",
          3793 => x"52",
          3794 => x"52",
          3795 => x"3f",
          3796 => x"52",
          3797 => x"51",
          3798 => x"84",
          3799 => x"d2",
          3800 => x"fc",
          3801 => x"8a",
          3802 => x"52",
          3803 => x"51",
          3804 => x"90",
          3805 => x"84",
          3806 => x"fb",
          3807 => x"17",
          3808 => x"a0",
          3809 => x"f4",
          3810 => x"08",
          3811 => x"b0",
          3812 => x"55",
          3813 => x"81",
          3814 => x"f8",
          3815 => x"84",
          3816 => x"53",
          3817 => x"17",
          3818 => x"88",
          3819 => x"c8",
          3820 => x"83",
          3821 => x"77",
          3822 => x"0c",
          3823 => x"04",
          3824 => x"77",
          3825 => x"12",
          3826 => x"55",
          3827 => x"56",
          3828 => x"8d",
          3829 => x"22",
          3830 => x"ac",
          3831 => x"57",
          3832 => x"93",
          3833 => x"3d",
          3834 => x"3d",
          3835 => x"70",
          3836 => x"55",
          3837 => x"88",
          3838 => x"08",
          3839 => x"38",
          3840 => x"d9",
          3841 => x"33",
          3842 => x"82",
          3843 => x"38",
          3844 => x"89",
          3845 => x"2e",
          3846 => x"bf",
          3847 => x"2e",
          3848 => x"81",
          3849 => x"81",
          3850 => x"89",
          3851 => x"08",
          3852 => x"52",
          3853 => x"3f",
          3854 => x"08",
          3855 => x"76",
          3856 => x"14",
          3857 => x"81",
          3858 => x"2a",
          3859 => x"05",
          3860 => x"59",
          3861 => x"f2",
          3862 => x"c8",
          3863 => x"38",
          3864 => x"06",
          3865 => x"33",
          3866 => x"7a",
          3867 => x"06",
          3868 => x"5a",
          3869 => x"53",
          3870 => x"38",
          3871 => x"06",
          3872 => x"39",
          3873 => x"a4",
          3874 => x"52",
          3875 => x"ba",
          3876 => x"c8",
          3877 => x"38",
          3878 => x"ff",
          3879 => x"b4",
          3880 => x"f8",
          3881 => x"c8",
          3882 => x"ff",
          3883 => x"39",
          3884 => x"a4",
          3885 => x"52",
          3886 => x"8e",
          3887 => x"c8",
          3888 => x"74",
          3889 => x"fc",
          3890 => x"b4",
          3891 => x"e5",
          3892 => x"c8",
          3893 => x"06",
          3894 => x"81",
          3895 => x"93",
          3896 => x"3d",
          3897 => x"3d",
          3898 => x"7f",
          3899 => x"82",
          3900 => x"27",
          3901 => x"73",
          3902 => x"27",
          3903 => x"74",
          3904 => x"77",
          3905 => x"38",
          3906 => x"89",
          3907 => x"2e",
          3908 => x"91",
          3909 => x"2e",
          3910 => x"82",
          3911 => x"81",
          3912 => x"89",
          3913 => x"08",
          3914 => x"52",
          3915 => x"3f",
          3916 => x"08",
          3917 => x"c8",
          3918 => x"38",
          3919 => x"06",
          3920 => x"81",
          3921 => x"06",
          3922 => x"58",
          3923 => x"80",
          3924 => x"75",
          3925 => x"f0",
          3926 => x"8f",
          3927 => x"58",
          3928 => x"34",
          3929 => x"16",
          3930 => x"2a",
          3931 => x"05",
          3932 => x"fa",
          3933 => x"93",
          3934 => x"82",
          3935 => x"81",
          3936 => x"83",
          3937 => x"b4",
          3938 => x"06",
          3939 => x"57",
          3940 => x"72",
          3941 => x"88",
          3942 => x"57",
          3943 => x"81",
          3944 => x"54",
          3945 => x"81",
          3946 => x"34",
          3947 => x"73",
          3948 => x"16",
          3949 => x"74",
          3950 => x"3f",
          3951 => x"08",
          3952 => x"c8",
          3953 => x"38",
          3954 => x"ff",
          3955 => x"14",
          3956 => x"75",
          3957 => x"51",
          3958 => x"81",
          3959 => x"34",
          3960 => x"73",
          3961 => x"16",
          3962 => x"74",
          3963 => x"3f",
          3964 => x"08",
          3965 => x"c8",
          3966 => x"75",
          3967 => x"74",
          3968 => x"fc",
          3969 => x"b4",
          3970 => x"51",
          3971 => x"a5",
          3972 => x"c8",
          3973 => x"06",
          3974 => x"72",
          3975 => x"3f",
          3976 => x"16",
          3977 => x"93",
          3978 => x"3d",
          3979 => x"3d",
          3980 => x"7d",
          3981 => x"58",
          3982 => x"74",
          3983 => x"98",
          3984 => x"26",
          3985 => x"56",
          3986 => x"75",
          3987 => x"38",
          3988 => x"52",
          3989 => x"8e",
          3990 => x"c8",
          3991 => x"93",
          3992 => x"f4",
          3993 => x"82",
          3994 => x"39",
          3995 => x"e8",
          3996 => x"c8",
          3997 => x"e0",
          3998 => x"76",
          3999 => x"3f",
          4000 => x"08",
          4001 => x"c8",
          4002 => x"80",
          4003 => x"93",
          4004 => x"2e",
          4005 => x"93",
          4006 => x"2e",
          4007 => x"53",
          4008 => x"51",
          4009 => x"82",
          4010 => x"c5",
          4011 => x"08",
          4012 => x"90",
          4013 => x"27",
          4014 => x"15",
          4015 => x"90",
          4016 => x"15",
          4017 => x"54",
          4018 => x"34",
          4019 => x"15",
          4020 => x"ff",
          4021 => x"56",
          4022 => x"c8",
          4023 => x"0d",
          4024 => x"0d",
          4025 => x"08",
          4026 => x"7a",
          4027 => x"19",
          4028 => x"80",
          4029 => x"98",
          4030 => x"26",
          4031 => x"58",
          4032 => x"52",
          4033 => x"e2",
          4034 => x"74",
          4035 => x"08",
          4036 => x"38",
          4037 => x"08",
          4038 => x"c8",
          4039 => x"82",
          4040 => x"93",
          4041 => x"98",
          4042 => x"93",
          4043 => x"82",
          4044 => x"58",
          4045 => x"19",
          4046 => x"82",
          4047 => x"57",
          4048 => x"09",
          4049 => x"db",
          4050 => x"57",
          4051 => x"77",
          4052 => x"82",
          4053 => x"7b",
          4054 => x"3f",
          4055 => x"08",
          4056 => x"82",
          4057 => x"81",
          4058 => x"06",
          4059 => x"93",
          4060 => x"75",
          4061 => x"30",
          4062 => x"80",
          4063 => x"07",
          4064 => x"52",
          4065 => x"81",
          4066 => x"80",
          4067 => x"8c",
          4068 => x"81",
          4069 => x"38",
          4070 => x"08",
          4071 => x"75",
          4072 => x"76",
          4073 => x"77",
          4074 => x"57",
          4075 => x"77",
          4076 => x"82",
          4077 => x"26",
          4078 => x"76",
          4079 => x"f8",
          4080 => x"93",
          4081 => x"82",
          4082 => x"80",
          4083 => x"80",
          4084 => x"c8",
          4085 => x"09",
          4086 => x"38",
          4087 => x"08",
          4088 => x"32",
          4089 => x"72",
          4090 => x"70",
          4091 => x"52",
          4092 => x"80",
          4093 => x"78",
          4094 => x"06",
          4095 => x"80",
          4096 => x"39",
          4097 => x"52",
          4098 => x"da",
          4099 => x"c8",
          4100 => x"c8",
          4101 => x"82",
          4102 => x"07",
          4103 => x"30",
          4104 => x"9f",
          4105 => x"52",
          4106 => x"56",
          4107 => x"8f",
          4108 => x"7a",
          4109 => x"f9",
          4110 => x"93",
          4111 => x"75",
          4112 => x"8c",
          4113 => x"19",
          4114 => x"54",
          4115 => x"74",
          4116 => x"90",
          4117 => x"05",
          4118 => x"84",
          4119 => x"07",
          4120 => x"1a",
          4121 => x"ff",
          4122 => x"2e",
          4123 => x"39",
          4124 => x"39",
          4125 => x"39",
          4126 => x"55",
          4127 => x"c8",
          4128 => x"0d",
          4129 => x"0d",
          4130 => x"57",
          4131 => x"81",
          4132 => x"c8",
          4133 => x"38",
          4134 => x"51",
          4135 => x"82",
          4136 => x"82",
          4137 => x"b0",
          4138 => x"84",
          4139 => x"52",
          4140 => x"52",
          4141 => x"3f",
          4142 => x"58",
          4143 => x"39",
          4144 => x"8a",
          4145 => x"75",
          4146 => x"38",
          4147 => x"1a",
          4148 => x"81",
          4149 => x"ee",
          4150 => x"93",
          4151 => x"2e",
          4152 => x"0b",
          4153 => x"56",
          4154 => x"2e",
          4155 => x"58",
          4156 => x"82",
          4157 => x"8b",
          4158 => x"f8",
          4159 => x"7c",
          4160 => x"56",
          4161 => x"80",
          4162 => x"38",
          4163 => x"53",
          4164 => x"86",
          4165 => x"81",
          4166 => x"90",
          4167 => x"17",
          4168 => x"aa",
          4169 => x"53",
          4170 => x"85",
          4171 => x"08",
          4172 => x"38",
          4173 => x"53",
          4174 => x"17",
          4175 => x"72",
          4176 => x"83",
          4177 => x"08",
          4178 => x"80",
          4179 => x"16",
          4180 => x"2b",
          4181 => x"75",
          4182 => x"73",
          4183 => x"f5",
          4184 => x"93",
          4185 => x"82",
          4186 => x"ff",
          4187 => x"81",
          4188 => x"c8",
          4189 => x"38",
          4190 => x"82",
          4191 => x"26",
          4192 => x"58",
          4193 => x"74",
          4194 => x"74",
          4195 => x"38",
          4196 => x"51",
          4197 => x"82",
          4198 => x"98",
          4199 => x"94",
          4200 => x"58",
          4201 => x"80",
          4202 => x"85",
          4203 => x"97",
          4204 => x"2a",
          4205 => x"05",
          4206 => x"74",
          4207 => x"16",
          4208 => x"18",
          4209 => x"77",
          4210 => x"0c",
          4211 => x"04",
          4212 => x"79",
          4213 => x"90",
          4214 => x"05",
          4215 => x"55",
          4216 => x"76",
          4217 => x"80",
          4218 => x"0c",
          4219 => x"15",
          4220 => x"81",
          4221 => x"83",
          4222 => x"73",
          4223 => x"98",
          4224 => x"05",
          4225 => x"94",
          4226 => x"38",
          4227 => x"88",
          4228 => x"53",
          4229 => x"81",
          4230 => x"98",
          4231 => x"53",
          4232 => x"8a",
          4233 => x"11",
          4234 => x"06",
          4235 => x"81",
          4236 => x"15",
          4237 => x"51",
          4238 => x"82",
          4239 => x"54",
          4240 => x"0b",
          4241 => x"08",
          4242 => x"38",
          4243 => x"93",
          4244 => x"2e",
          4245 => x"98",
          4246 => x"93",
          4247 => x"80",
          4248 => x"8a",
          4249 => x"16",
          4250 => x"80",
          4251 => x"15",
          4252 => x"51",
          4253 => x"82",
          4254 => x"54",
          4255 => x"93",
          4256 => x"2e",
          4257 => x"82",
          4258 => x"c8",
          4259 => x"bf",
          4260 => x"82",
          4261 => x"ff",
          4262 => x"82",
          4263 => x"52",
          4264 => x"e1",
          4265 => x"82",
          4266 => x"a3",
          4267 => x"16",
          4268 => x"76",
          4269 => x"3f",
          4270 => x"08",
          4271 => x"75",
          4272 => x"75",
          4273 => x"17",
          4274 => x"16",
          4275 => x"72",
          4276 => x"0c",
          4277 => x"04",
          4278 => x"7a",
          4279 => x"5a",
          4280 => x"52",
          4281 => x"93",
          4282 => x"c8",
          4283 => x"93",
          4284 => x"e1",
          4285 => x"c8",
          4286 => x"16",
          4287 => x"51",
          4288 => x"82",
          4289 => x"54",
          4290 => x"08",
          4291 => x"82",
          4292 => x"9c",
          4293 => x"33",
          4294 => x"72",
          4295 => x"09",
          4296 => x"38",
          4297 => x"30",
          4298 => x"76",
          4299 => x"72",
          4300 => x"38",
          4301 => x"76",
          4302 => x"38",
          4303 => x"57",
          4304 => x"51",
          4305 => x"82",
          4306 => x"54",
          4307 => x"08",
          4308 => x"a6",
          4309 => x"2e",
          4310 => x"83",
          4311 => x"73",
          4312 => x"0c",
          4313 => x"04",
          4314 => x"76",
          4315 => x"54",
          4316 => x"82",
          4317 => x"83",
          4318 => x"76",
          4319 => x"53",
          4320 => x"2e",
          4321 => x"90",
          4322 => x"51",
          4323 => x"82",
          4324 => x"90",
          4325 => x"53",
          4326 => x"c8",
          4327 => x"0d",
          4328 => x"0d",
          4329 => x"83",
          4330 => x"54",
          4331 => x"55",
          4332 => x"3f",
          4333 => x"51",
          4334 => x"2e",
          4335 => x"8b",
          4336 => x"2a",
          4337 => x"51",
          4338 => x"86",
          4339 => x"f7",
          4340 => x"7d",
          4341 => x"76",
          4342 => x"98",
          4343 => x"2e",
          4344 => x"98",
          4345 => x"78",
          4346 => x"3f",
          4347 => x"08",
          4348 => x"c8",
          4349 => x"38",
          4350 => x"70",
          4351 => x"74",
          4352 => x"58",
          4353 => x"9c",
          4354 => x"11",
          4355 => x"06",
          4356 => x"06",
          4357 => x"53",
          4358 => x"34",
          4359 => x"32",
          4360 => x"ae",
          4361 => x"70",
          4362 => x"2a",
          4363 => x"51",
          4364 => x"2e",
          4365 => x"8f",
          4366 => x"80",
          4367 => x"54",
          4368 => x"2e",
          4369 => x"83",
          4370 => x"73",
          4371 => x"38",
          4372 => x"51",
          4373 => x"82",
          4374 => x"58",
          4375 => x"08",
          4376 => x"16",
          4377 => x"38",
          4378 => x"86",
          4379 => x"98",
          4380 => x"82",
          4381 => x"8b",
          4382 => x"f8",
          4383 => x"70",
          4384 => x"80",
          4385 => x"f8",
          4386 => x"93",
          4387 => x"82",
          4388 => x"80",
          4389 => x"39",
          4390 => x"e6",
          4391 => x"08",
          4392 => x"ec",
          4393 => x"93",
          4394 => x"82",
          4395 => x"80",
          4396 => x"16",
          4397 => x"51",
          4398 => x"2e",
          4399 => x"16",
          4400 => x"33",
          4401 => x"55",
          4402 => x"34",
          4403 => x"70",
          4404 => x"81",
          4405 => x"59",
          4406 => x"8b",
          4407 => x"52",
          4408 => x"85",
          4409 => x"c8",
          4410 => x"96",
          4411 => x"75",
          4412 => x"3f",
          4413 => x"08",
          4414 => x"c8",
          4415 => x"ff",
          4416 => x"54",
          4417 => x"c8",
          4418 => x"0d",
          4419 => x"0d",
          4420 => x"57",
          4421 => x"73",
          4422 => x"3f",
          4423 => x"08",
          4424 => x"c8",
          4425 => x"98",
          4426 => x"75",
          4427 => x"3f",
          4428 => x"08",
          4429 => x"c8",
          4430 => x"a0",
          4431 => x"c8",
          4432 => x"14",
          4433 => x"87",
          4434 => x"a0",
          4435 => x"14",
          4436 => x"d7",
          4437 => x"83",
          4438 => x"82",
          4439 => x"87",
          4440 => x"fc",
          4441 => x"70",
          4442 => x"08",
          4443 => x"56",
          4444 => x"3f",
          4445 => x"08",
          4446 => x"c8",
          4447 => x"9c",
          4448 => x"e5",
          4449 => x"0b",
          4450 => x"73",
          4451 => x"0c",
          4452 => x"04",
          4453 => x"78",
          4454 => x"80",
          4455 => x"34",
          4456 => x"80",
          4457 => x"38",
          4458 => x"55",
          4459 => x"14",
          4460 => x"16",
          4461 => x"72",
          4462 => x"38",
          4463 => x"09",
          4464 => x"38",
          4465 => x"73",
          4466 => x"81",
          4467 => x"75",
          4468 => x"52",
          4469 => x"13",
          4470 => x"55",
          4471 => x"05",
          4472 => x"13",
          4473 => x"55",
          4474 => x"c0",
          4475 => x"88",
          4476 => x"0b",
          4477 => x"9c",
          4478 => x"8b",
          4479 => x"17",
          4480 => x"08",
          4481 => x"e6",
          4482 => x"93",
          4483 => x"0c",
          4484 => x"96",
          4485 => x"84",
          4486 => x"c8",
          4487 => x"23",
          4488 => x"98",
          4489 => x"f4",
          4490 => x"c8",
          4491 => x"23",
          4492 => x"04",
          4493 => x"7e",
          4494 => x"a0",
          4495 => x"5c",
          4496 => x"52",
          4497 => x"87",
          4498 => x"58",
          4499 => x"33",
          4500 => x"ae",
          4501 => x"06",
          4502 => x"78",
          4503 => x"81",
          4504 => x"32",
          4505 => x"9f",
          4506 => x"26",
          4507 => x"53",
          4508 => x"73",
          4509 => x"18",
          4510 => x"34",
          4511 => x"db",
          4512 => x"32",
          4513 => x"80",
          4514 => x"30",
          4515 => x"9f",
          4516 => x"56",
          4517 => x"80",
          4518 => x"86",
          4519 => x"26",
          4520 => x"76",
          4521 => x"a4",
          4522 => x"27",
          4523 => x"54",
          4524 => x"34",
          4525 => x"ce",
          4526 => x"70",
          4527 => x"59",
          4528 => x"76",
          4529 => x"38",
          4530 => x"70",
          4531 => x"dc",
          4532 => x"72",
          4533 => x"80",
          4534 => x"51",
          4535 => x"74",
          4536 => x"38",
          4537 => x"17",
          4538 => x"1a",
          4539 => x"55",
          4540 => x"2e",
          4541 => x"83",
          4542 => x"80",
          4543 => x"33",
          4544 => x"73",
          4545 => x"09",
          4546 => x"38",
          4547 => x"75",
          4548 => x"d2",
          4549 => x"39",
          4550 => x"70",
          4551 => x"25",
          4552 => x"07",
          4553 => x"73",
          4554 => x"38",
          4555 => x"70",
          4556 => x"32",
          4557 => x"80",
          4558 => x"2a",
          4559 => x"56",
          4560 => x"81",
          4561 => x"58",
          4562 => x"ed",
          4563 => x"2b",
          4564 => x"25",
          4565 => x"80",
          4566 => x"fb",
          4567 => x"57",
          4568 => x"e5",
          4569 => x"93",
          4570 => x"2e",
          4571 => x"17",
          4572 => x"19",
          4573 => x"56",
          4574 => x"3f",
          4575 => x"08",
          4576 => x"38",
          4577 => x"73",
          4578 => x"38",
          4579 => x"f6",
          4580 => x"54",
          4581 => x"81",
          4582 => x"55",
          4583 => x"34",
          4584 => x"fe",
          4585 => x"52",
          4586 => x"51",
          4587 => x"82",
          4588 => x"80",
          4589 => x"9f",
          4590 => x"99",
          4591 => x"e0",
          4592 => x"ff",
          4593 => x"7a",
          4594 => x"74",
          4595 => x"58",
          4596 => x"76",
          4597 => x"86",
          4598 => x"2e",
          4599 => x"33",
          4600 => x"e5",
          4601 => x"06",
          4602 => x"7b",
          4603 => x"a0",
          4604 => x"38",
          4605 => x"54",
          4606 => x"54",
          4607 => x"54",
          4608 => x"34",
          4609 => x"82",
          4610 => x"8d",
          4611 => x"fa",
          4612 => x"70",
          4613 => x"80",
          4614 => x"51",
          4615 => x"af",
          4616 => x"81",
          4617 => x"70",
          4618 => x"54",
          4619 => x"2e",
          4620 => x"54",
          4621 => x"53",
          4622 => x"8c",
          4623 => x"08",
          4624 => x"b3",
          4625 => x"5a",
          4626 => x"33",
          4627 => x"72",
          4628 => x"81",
          4629 => x"81",
          4630 => x"70",
          4631 => x"54",
          4632 => x"2e",
          4633 => x"83",
          4634 => x"74",
          4635 => x"72",
          4636 => x"0b",
          4637 => x"79",
          4638 => x"53",
          4639 => x"9b",
          4640 => x"0b",
          4641 => x"80",
          4642 => x"f0",
          4643 => x"93",
          4644 => x"81",
          4645 => x"55",
          4646 => x"89",
          4647 => x"52",
          4648 => x"90",
          4649 => x"c8",
          4650 => x"93",
          4651 => x"8f",
          4652 => x"f7",
          4653 => x"93",
          4654 => x"17",
          4655 => x"82",
          4656 => x"80",
          4657 => x"38",
          4658 => x"08",
          4659 => x"81",
          4660 => x"38",
          4661 => x"70",
          4662 => x"53",
          4663 => x"9a",
          4664 => x"2a",
          4665 => x"51",
          4666 => x"2e",
          4667 => x"ff",
          4668 => x"17",
          4669 => x"80",
          4670 => x"82",
          4671 => x"06",
          4672 => x"bb",
          4673 => x"b7",
          4674 => x"2a",
          4675 => x"51",
          4676 => x"38",
          4677 => x"70",
          4678 => x"81",
          4679 => x"54",
          4680 => x"fe",
          4681 => x"16",
          4682 => x"06",
          4683 => x"52",
          4684 => x"b4",
          4685 => x"c8",
          4686 => x"0c",
          4687 => x"74",
          4688 => x"0c",
          4689 => x"04",
          4690 => x"7c",
          4691 => x"08",
          4692 => x"59",
          4693 => x"80",
          4694 => x"38",
          4695 => x"05",
          4696 => x"ba",
          4697 => x"72",
          4698 => x"9f",
          4699 => x"51",
          4700 => x"e8",
          4701 => x"2e",
          4702 => x"81",
          4703 => x"33",
          4704 => x"52",
          4705 => x"92",
          4706 => x"72",
          4707 => x"d0",
          4708 => x"51",
          4709 => x"80",
          4710 => x"0b",
          4711 => x"5c",
          4712 => x"10",
          4713 => x"7a",
          4714 => x"51",
          4715 => x"05",
          4716 => x"70",
          4717 => x"33",
          4718 => x"53",
          4719 => x"99",
          4720 => x"e0",
          4721 => x"ff",
          4722 => x"ff",
          4723 => x"70",
          4724 => x"38",
          4725 => x"81",
          4726 => x"51",
          4727 => x"74",
          4728 => x"70",
          4729 => x"25",
          4730 => x"06",
          4731 => x"51",
          4732 => x"38",
          4733 => x"78",
          4734 => x"70",
          4735 => x"2a",
          4736 => x"07",
          4737 => x"51",
          4738 => x"8c",
          4739 => x"58",
          4740 => x"ff",
          4741 => x"39",
          4742 => x"86",
          4743 => x"7a",
          4744 => x"51",
          4745 => x"93",
          4746 => x"70",
          4747 => x"0c",
          4748 => x"04",
          4749 => x"77",
          4750 => x"83",
          4751 => x"0b",
          4752 => x"78",
          4753 => x"e1",
          4754 => x"55",
          4755 => x"08",
          4756 => x"84",
          4757 => x"dd",
          4758 => x"93",
          4759 => x"ff",
          4760 => x"83",
          4761 => x"d4",
          4762 => x"81",
          4763 => x"38",
          4764 => x"17",
          4765 => x"73",
          4766 => x"09",
          4767 => x"38",
          4768 => x"81",
          4769 => x"30",
          4770 => x"77",
          4771 => x"54",
          4772 => x"b4",
          4773 => x"73",
          4774 => x"09",
          4775 => x"38",
          4776 => x"fb",
          4777 => x"ea",
          4778 => x"bd",
          4779 => x"c8",
          4780 => x"93",
          4781 => x"2e",
          4782 => x"53",
          4783 => x"52",
          4784 => x"51",
          4785 => x"82",
          4786 => x"55",
          4787 => x"08",
          4788 => x"38",
          4789 => x"82",
          4790 => x"87",
          4791 => x"f3",
          4792 => x"02",
          4793 => x"c7",
          4794 => x"54",
          4795 => x"7f",
          4796 => x"3f",
          4797 => x"08",
          4798 => x"80",
          4799 => x"c8",
          4800 => x"9e",
          4801 => x"c8",
          4802 => x"82",
          4803 => x"70",
          4804 => x"8c",
          4805 => x"2e",
          4806 => x"74",
          4807 => x"81",
          4808 => x"33",
          4809 => x"80",
          4810 => x"81",
          4811 => x"d6",
          4812 => x"93",
          4813 => x"ff",
          4814 => x"06",
          4815 => x"99",
          4816 => x"2e",
          4817 => x"82",
          4818 => x"06",
          4819 => x"56",
          4820 => x"38",
          4821 => x"ca",
          4822 => x"34",
          4823 => x"34",
          4824 => x"15",
          4825 => x"8d",
          4826 => x"c8",
          4827 => x"06",
          4828 => x"54",
          4829 => x"72",
          4830 => x"76",
          4831 => x"38",
          4832 => x"70",
          4833 => x"53",
          4834 => x"86",
          4835 => x"70",
          4836 => x"5a",
          4837 => x"82",
          4838 => x"81",
          4839 => x"76",
          4840 => x"81",
          4841 => x"38",
          4842 => x"90",
          4843 => x"3d",
          4844 => x"05",
          4845 => x"f6",
          4846 => x"59",
          4847 => x"72",
          4848 => x"38",
          4849 => x"51",
          4850 => x"82",
          4851 => x"57",
          4852 => x"81",
          4853 => x"74",
          4854 => x"80",
          4855 => x"74",
          4856 => x"f0",
          4857 => x"53",
          4858 => x"80",
          4859 => x"79",
          4860 => x"fc",
          4861 => x"93",
          4862 => x"ff",
          4863 => x"77",
          4864 => x"81",
          4865 => x"74",
          4866 => x"81",
          4867 => x"2e",
          4868 => x"8d",
          4869 => x"26",
          4870 => x"bf",
          4871 => x"fc",
          4872 => x"c8",
          4873 => x"ff",
          4874 => x"56",
          4875 => x"2e",
          4876 => x"84",
          4877 => x"ca",
          4878 => x"e0",
          4879 => x"c8",
          4880 => x"ff",
          4881 => x"8d",
          4882 => x"15",
          4883 => x"3f",
          4884 => x"08",
          4885 => x"16",
          4886 => x"15",
          4887 => x"34",
          4888 => x"33",
          4889 => x"8d",
          4890 => x"26",
          4891 => x"82",
          4892 => x"71",
          4893 => x"17",
          4894 => x"53",
          4895 => x"23",
          4896 => x"ff",
          4897 => x"80",
          4898 => x"ff",
          4899 => x"53",
          4900 => x"86",
          4901 => x"84",
          4902 => x"c5",
          4903 => x"fc",
          4904 => x"c8",
          4905 => x"23",
          4906 => x"08",
          4907 => x"06",
          4908 => x"8d",
          4909 => x"ea",
          4910 => x"15",
          4911 => x"3f",
          4912 => x"08",
          4913 => x"06",
          4914 => x"38",
          4915 => x"51",
          4916 => x"82",
          4917 => x"53",
          4918 => x"51",
          4919 => x"82",
          4920 => x"83",
          4921 => x"59",
          4922 => x"80",
          4923 => x"38",
          4924 => x"74",
          4925 => x"2a",
          4926 => x"8d",
          4927 => x"26",
          4928 => x"8a",
          4929 => x"72",
          4930 => x"ff",
          4931 => x"82",
          4932 => x"53",
          4933 => x"93",
          4934 => x"2e",
          4935 => x"80",
          4936 => x"c8",
          4937 => x"ff",
          4938 => x"83",
          4939 => x"72",
          4940 => x"26",
          4941 => x"57",
          4942 => x"26",
          4943 => x"57",
          4944 => x"80",
          4945 => x"38",
          4946 => x"16",
          4947 => x"16",
          4948 => x"a4",
          4949 => x"1a",
          4950 => x"76",
          4951 => x"81",
          4952 => x"80",
          4953 => x"d7",
          4954 => x"93",
          4955 => x"ff",
          4956 => x"8d",
          4957 => x"aa",
          4958 => x"22",
          4959 => x"72",
          4960 => x"80",
          4961 => x"d7",
          4962 => x"93",
          4963 => x"16",
          4964 => x"08",
          4965 => x"b6",
          4966 => x"22",
          4967 => x"72",
          4968 => x"fe",
          4969 => x"08",
          4970 => x"0c",
          4971 => x"09",
          4972 => x"38",
          4973 => x"10",
          4974 => x"98",
          4975 => x"98",
          4976 => x"70",
          4977 => x"17",
          4978 => x"05",
          4979 => x"ff",
          4980 => x"53",
          4981 => x"9c",
          4982 => x"81",
          4983 => x"0b",
          4984 => x"ff",
          4985 => x"0c",
          4986 => x"84",
          4987 => x"83",
          4988 => x"06",
          4989 => x"80",
          4990 => x"d6",
          4991 => x"93",
          4992 => x"ff",
          4993 => x"72",
          4994 => x"81",
          4995 => x"38",
          4996 => x"74",
          4997 => x"3f",
          4998 => x"08",
          4999 => x"82",
          5000 => x"84",
          5001 => x"b2",
          5002 => x"f0",
          5003 => x"c8",
          5004 => x"ff",
          5005 => x"82",
          5006 => x"09",
          5007 => x"c8",
          5008 => x"51",
          5009 => x"82",
          5010 => x"84",
          5011 => x"d2",
          5012 => x"06",
          5013 => x"98",
          5014 => x"d9",
          5015 => x"c8",
          5016 => x"85",
          5017 => x"09",
          5018 => x"38",
          5019 => x"51",
          5020 => x"82",
          5021 => x"90",
          5022 => x"a0",
          5023 => x"b5",
          5024 => x"c8",
          5025 => x"0c",
          5026 => x"82",
          5027 => x"81",
          5028 => x"82",
          5029 => x"72",
          5030 => x"80",
          5031 => x"0c",
          5032 => x"82",
          5033 => x"8f",
          5034 => x"fb",
          5035 => x"54",
          5036 => x"80",
          5037 => x"73",
          5038 => x"af",
          5039 => x"70",
          5040 => x"71",
          5041 => x"38",
          5042 => x"86",
          5043 => x"52",
          5044 => x"09",
          5045 => x"38",
          5046 => x"51",
          5047 => x"82",
          5048 => x"81",
          5049 => x"83",
          5050 => x"80",
          5051 => x"2e",
          5052 => x"84",
          5053 => x"53",
          5054 => x"0c",
          5055 => x"93",
          5056 => x"3d",
          5057 => x"3d",
          5058 => x"05",
          5059 => x"89",
          5060 => x"52",
          5061 => x"3f",
          5062 => x"08",
          5063 => x"80",
          5064 => x"c8",
          5065 => x"c4",
          5066 => x"c8",
          5067 => x"82",
          5068 => x"70",
          5069 => x"73",
          5070 => x"38",
          5071 => x"78",
          5072 => x"38",
          5073 => x"74",
          5074 => x"10",
          5075 => x"05",
          5076 => x"54",
          5077 => x"80",
          5078 => x"80",
          5079 => x"70",
          5080 => x"51",
          5081 => x"82",
          5082 => x"54",
          5083 => x"c8",
          5084 => x"0d",
          5085 => x"0d",
          5086 => x"05",
          5087 => x"33",
          5088 => x"55",
          5089 => x"84",
          5090 => x"bf",
          5091 => x"98",
          5092 => x"53",
          5093 => x"05",
          5094 => x"c3",
          5095 => x"c8",
          5096 => x"93",
          5097 => x"c5",
          5098 => x"68",
          5099 => x"d4",
          5100 => x"db",
          5101 => x"c8",
          5102 => x"93",
          5103 => x"38",
          5104 => x"05",
          5105 => x"2b",
          5106 => x"80",
          5107 => x"86",
          5108 => x"06",
          5109 => x"2e",
          5110 => x"75",
          5111 => x"38",
          5112 => x"09",
          5113 => x"38",
          5114 => x"05",
          5115 => x"3f",
          5116 => x"08",
          5117 => x"07",
          5118 => x"02",
          5119 => x"91",
          5120 => x"80",
          5121 => x"87",
          5122 => x"76",
          5123 => x"81",
          5124 => x"74",
          5125 => x"38",
          5126 => x"83",
          5127 => x"83",
          5128 => x"06",
          5129 => x"80",
          5130 => x"38",
          5131 => x"51",
          5132 => x"82",
          5133 => x"59",
          5134 => x"0a",
          5135 => x"05",
          5136 => x"3f",
          5137 => x"0b",
          5138 => x"75",
          5139 => x"7a",
          5140 => x"3f",
          5141 => x"9c",
          5142 => x"a0",
          5143 => x"81",
          5144 => x"34",
          5145 => x"80",
          5146 => x"b0",
          5147 => x"55",
          5148 => x"3d",
          5149 => x"51",
          5150 => x"3f",
          5151 => x"08",
          5152 => x"c8",
          5153 => x"38",
          5154 => x"51",
          5155 => x"82",
          5156 => x"7b",
          5157 => x"12",
          5158 => x"b6",
          5159 => x"cd",
          5160 => x"05",
          5161 => x"2a",
          5162 => x"51",
          5163 => x"80",
          5164 => x"84",
          5165 => x"76",
          5166 => x"81",
          5167 => x"74",
          5168 => x"38",
          5169 => x"33",
          5170 => x"74",
          5171 => x"38",
          5172 => x"82",
          5173 => x"83",
          5174 => x"06",
          5175 => x"80",
          5176 => x"76",
          5177 => x"57",
          5178 => x"08",
          5179 => x"63",
          5180 => x"55",
          5181 => x"38",
          5182 => x"51",
          5183 => x"82",
          5184 => x"88",
          5185 => x"9c",
          5186 => x"a9",
          5187 => x"c8",
          5188 => x"0c",
          5189 => x"86",
          5190 => x"19",
          5191 => x"19",
          5192 => x"19",
          5193 => x"19",
          5194 => x"19",
          5195 => x"53",
          5196 => x"18",
          5197 => x"3f",
          5198 => x"70",
          5199 => x"55",
          5200 => x"81",
          5201 => x"18",
          5202 => x"81",
          5203 => x"18",
          5204 => x"0c",
          5205 => x"22",
          5206 => x"88",
          5207 => x"1c",
          5208 => x"5c",
          5209 => x"39",
          5210 => x"51",
          5211 => x"82",
          5212 => x"57",
          5213 => x"08",
          5214 => x"38",
          5215 => x"ff",
          5216 => x"06",
          5217 => x"56",
          5218 => x"59",
          5219 => x"77",
          5220 => x"70",
          5221 => x"06",
          5222 => x"74",
          5223 => x"98",
          5224 => x"80",
          5225 => x"83",
          5226 => x"74",
          5227 => x"38",
          5228 => x"51",
          5229 => x"82",
          5230 => x"85",
          5231 => x"a8",
          5232 => x"2a",
          5233 => x"08",
          5234 => x"1a",
          5235 => x"54",
          5236 => x"18",
          5237 => x"11",
          5238 => x"ca",
          5239 => x"93",
          5240 => x"2e",
          5241 => x"56",
          5242 => x"84",
          5243 => x"0c",
          5244 => x"82",
          5245 => x"97",
          5246 => x"f3",
          5247 => x"62",
          5248 => x"5f",
          5249 => x"7d",
          5250 => x"fc",
          5251 => x"51",
          5252 => x"82",
          5253 => x"55",
          5254 => x"08",
          5255 => x"17",
          5256 => x"80",
          5257 => x"74",
          5258 => x"39",
          5259 => x"81",
          5260 => x"56",
          5261 => x"83",
          5262 => x"39",
          5263 => x"18",
          5264 => x"83",
          5265 => x"0b",
          5266 => x"81",
          5267 => x"39",
          5268 => x"18",
          5269 => x"83",
          5270 => x"0b",
          5271 => x"81",
          5272 => x"39",
          5273 => x"18",
          5274 => x"82",
          5275 => x"0b",
          5276 => x"81",
          5277 => x"39",
          5278 => x"94",
          5279 => x"55",
          5280 => x"83",
          5281 => x"78",
          5282 => x"cb",
          5283 => x"08",
          5284 => x"06",
          5285 => x"82",
          5286 => x"8a",
          5287 => x"05",
          5288 => x"06",
          5289 => x"a8",
          5290 => x"38",
          5291 => x"55",
          5292 => x"17",
          5293 => x"51",
          5294 => x"82",
          5295 => x"55",
          5296 => x"fe",
          5297 => x"ff",
          5298 => x"38",
          5299 => x"0c",
          5300 => x"52",
          5301 => x"e8",
          5302 => x"c8",
          5303 => x"fe",
          5304 => x"93",
          5305 => x"79",
          5306 => x"58",
          5307 => x"80",
          5308 => x"1b",
          5309 => x"22",
          5310 => x"74",
          5311 => x"38",
          5312 => x"5a",
          5313 => x"53",
          5314 => x"81",
          5315 => x"55",
          5316 => x"82",
          5317 => x"fe",
          5318 => x"17",
          5319 => x"2b",
          5320 => x"80",
          5321 => x"9c",
          5322 => x"31",
          5323 => x"27",
          5324 => x"80",
          5325 => x"52",
          5326 => x"29",
          5327 => x"eb",
          5328 => x"2b",
          5329 => x"39",
          5330 => x"78",
          5331 => x"38",
          5332 => x"70",
          5333 => x"56",
          5334 => x"a5",
          5335 => x"9c",
          5336 => x"a8",
          5337 => x"81",
          5338 => x"55",
          5339 => x"82",
          5340 => x"fd",
          5341 => x"17",
          5342 => x"06",
          5343 => x"18",
          5344 => x"77",
          5345 => x"52",
          5346 => x"33",
          5347 => x"f1",
          5348 => x"c8",
          5349 => x"38",
          5350 => x"0c",
          5351 => x"83",
          5352 => x"80",
          5353 => x"55",
          5354 => x"83",
          5355 => x"75",
          5356 => x"08",
          5357 => x"17",
          5358 => x"7b",
          5359 => x"3f",
          5360 => x"7d",
          5361 => x"0c",
          5362 => x"19",
          5363 => x"1a",
          5364 => x"78",
          5365 => x"80",
          5366 => x"93",
          5367 => x"3d",
          5368 => x"3d",
          5369 => x"64",
          5370 => x"5a",
          5371 => x"0c",
          5372 => x"05",
          5373 => x"f5",
          5374 => x"93",
          5375 => x"82",
          5376 => x"8a",
          5377 => x"33",
          5378 => x"2e",
          5379 => x"56",
          5380 => x"90",
          5381 => x"81",
          5382 => x"06",
          5383 => x"87",
          5384 => x"2e",
          5385 => x"bd",
          5386 => x"91",
          5387 => x"56",
          5388 => x"81",
          5389 => x"34",
          5390 => x"d8",
          5391 => x"91",
          5392 => x"56",
          5393 => x"82",
          5394 => x"34",
          5395 => x"c4",
          5396 => x"91",
          5397 => x"56",
          5398 => x"81",
          5399 => x"34",
          5400 => x"b0",
          5401 => x"08",
          5402 => x"94",
          5403 => x"86",
          5404 => x"08",
          5405 => x"80",
          5406 => x"38",
          5407 => x"70",
          5408 => x"56",
          5409 => x"a8",
          5410 => x"11",
          5411 => x"77",
          5412 => x"5c",
          5413 => x"c6",
          5414 => x"38",
          5415 => x"55",
          5416 => x"7a",
          5417 => x"d4",
          5418 => x"93",
          5419 => x"8f",
          5420 => x"08",
          5421 => x"d4",
          5422 => x"93",
          5423 => x"74",
          5424 => x"c3",
          5425 => x"2e",
          5426 => x"74",
          5427 => x"e3",
          5428 => x"18",
          5429 => x"08",
          5430 => x"88",
          5431 => x"17",
          5432 => x"2b",
          5433 => x"80",
          5434 => x"81",
          5435 => x"08",
          5436 => x"52",
          5437 => x"33",
          5438 => x"de",
          5439 => x"c8",
          5440 => x"38",
          5441 => x"80",
          5442 => x"74",
          5443 => x"98",
          5444 => x"7d",
          5445 => x"3f",
          5446 => x"08",
          5447 => x"a7",
          5448 => x"c8",
          5449 => x"89",
          5450 => x"79",
          5451 => x"d5",
          5452 => x"7e",
          5453 => x"51",
          5454 => x"76",
          5455 => x"74",
          5456 => x"79",
          5457 => x"7b",
          5458 => x"11",
          5459 => x"c5",
          5460 => x"93",
          5461 => x"f9",
          5462 => x"08",
          5463 => x"74",
          5464 => x"38",
          5465 => x"74",
          5466 => x"1c",
          5467 => x"51",
          5468 => x"90",
          5469 => x"ff",
          5470 => x"90",
          5471 => x"89",
          5472 => x"db",
          5473 => x"08",
          5474 => x"38",
          5475 => x"8c",
          5476 => x"98",
          5477 => x"77",
          5478 => x"52",
          5479 => x"33",
          5480 => x"dd",
          5481 => x"c8",
          5482 => x"38",
          5483 => x"0c",
          5484 => x"83",
          5485 => x"80",
          5486 => x"55",
          5487 => x"83",
          5488 => x"75",
          5489 => x"94",
          5490 => x"ff",
          5491 => x"05",
          5492 => x"3f",
          5493 => x"ff",
          5494 => x"74",
          5495 => x"78",
          5496 => x"08",
          5497 => x"76",
          5498 => x"08",
          5499 => x"1b",
          5500 => x"08",
          5501 => x"59",
          5502 => x"83",
          5503 => x"74",
          5504 => x"78",
          5505 => x"90",
          5506 => x"c0",
          5507 => x"90",
          5508 => x"56",
          5509 => x"c8",
          5510 => x"0d",
          5511 => x"0d",
          5512 => x"fc",
          5513 => x"52",
          5514 => x"3f",
          5515 => x"08",
          5516 => x"c8",
          5517 => x"38",
          5518 => x"70",
          5519 => x"81",
          5520 => x"56",
          5521 => x"81",
          5522 => x"98",
          5523 => x"80",
          5524 => x"81",
          5525 => x"08",
          5526 => x"52",
          5527 => x"33",
          5528 => x"f6",
          5529 => x"82",
          5530 => x"80",
          5531 => x"18",
          5532 => x"06",
          5533 => x"19",
          5534 => x"08",
          5535 => x"c8",
          5536 => x"93",
          5537 => x"82",
          5538 => x"80",
          5539 => x"18",
          5540 => x"33",
          5541 => x"56",
          5542 => x"34",
          5543 => x"53",
          5544 => x"08",
          5545 => x"3f",
          5546 => x"52",
          5547 => x"c5",
          5548 => x"88",
          5549 => x"96",
          5550 => x"c0",
          5551 => x"92",
          5552 => x"9a",
          5553 => x"81",
          5554 => x"34",
          5555 => x"c1",
          5556 => x"c8",
          5557 => x"33",
          5558 => x"56",
          5559 => x"19",
          5560 => x"74",
          5561 => x"0c",
          5562 => x"04",
          5563 => x"76",
          5564 => x"fe",
          5565 => x"93",
          5566 => x"82",
          5567 => x"9c",
          5568 => x"fc",
          5569 => x"51",
          5570 => x"82",
          5571 => x"53",
          5572 => x"08",
          5573 => x"93",
          5574 => x"0c",
          5575 => x"c8",
          5576 => x"0d",
          5577 => x"0d",
          5578 => x"e4",
          5579 => x"53",
          5580 => x"93",
          5581 => x"8b",
          5582 => x"c8",
          5583 => x"f8",
          5584 => x"72",
          5585 => x"0c",
          5586 => x"04",
          5587 => x"80",
          5588 => x"d0",
          5589 => x"3d",
          5590 => x"3f",
          5591 => x"08",
          5592 => x"c8",
          5593 => x"38",
          5594 => x"52",
          5595 => x"05",
          5596 => x"3f",
          5597 => x"08",
          5598 => x"c8",
          5599 => x"02",
          5600 => x"33",
          5601 => x"55",
          5602 => x"25",
          5603 => x"7a",
          5604 => x"54",
          5605 => x"a2",
          5606 => x"84",
          5607 => x"06",
          5608 => x"73",
          5609 => x"38",
          5610 => x"70",
          5611 => x"b8",
          5612 => x"c8",
          5613 => x"0c",
          5614 => x"55",
          5615 => x"09",
          5616 => x"38",
          5617 => x"82",
          5618 => x"93",
          5619 => x"e1",
          5620 => x"3d",
          5621 => x"08",
          5622 => x"7a",
          5623 => x"a1",
          5624 => x"05",
          5625 => x"51",
          5626 => x"82",
          5627 => x"57",
          5628 => x"08",
          5629 => x"7e",
          5630 => x"94",
          5631 => x"55",
          5632 => x"74",
          5633 => x"f9",
          5634 => x"70",
          5635 => x"5e",
          5636 => x"7a",
          5637 => x"3f",
          5638 => x"08",
          5639 => x"c8",
          5640 => x"38",
          5641 => x"51",
          5642 => x"82",
          5643 => x"57",
          5644 => x"08",
          5645 => x"6c",
          5646 => x"d6",
          5647 => x"93",
          5648 => x"76",
          5649 => x"d1",
          5650 => x"93",
          5651 => x"82",
          5652 => x"81",
          5653 => x"54",
          5654 => x"51",
          5655 => x"82",
          5656 => x"57",
          5657 => x"08",
          5658 => x"52",
          5659 => x"f8",
          5660 => x"c8",
          5661 => x"95",
          5662 => x"73",
          5663 => x"3f",
          5664 => x"08",
          5665 => x"c8",
          5666 => x"cc",
          5667 => x"2e",
          5668 => x"83",
          5669 => x"76",
          5670 => x"a1",
          5671 => x"11",
          5672 => x"51",
          5673 => x"76",
          5674 => x"79",
          5675 => x"33",
          5676 => x"55",
          5677 => x"2e",
          5678 => x"16",
          5679 => x"11",
          5680 => x"56",
          5681 => x"81",
          5682 => x"74",
          5683 => x"91",
          5684 => x"75",
          5685 => x"38",
          5686 => x"19",
          5687 => x"11",
          5688 => x"1b",
          5689 => x"59",
          5690 => x"75",
          5691 => x"38",
          5692 => x"3d",
          5693 => x"59",
          5694 => x"67",
          5695 => x"91",
          5696 => x"85",
          5697 => x"2e",
          5698 => x"8c",
          5699 => x"a3",
          5700 => x"55",
          5701 => x"34",
          5702 => x"93",
          5703 => x"10",
          5704 => x"e8",
          5705 => x"70",
          5706 => x"57",
          5707 => x"73",
          5708 => x"38",
          5709 => x"16",
          5710 => x"55",
          5711 => x"38",
          5712 => x"73",
          5713 => x"38",
          5714 => x"76",
          5715 => x"77",
          5716 => x"33",
          5717 => x"05",
          5718 => x"18",
          5719 => x"26",
          5720 => x"7a",
          5721 => x"5c",
          5722 => x"58",
          5723 => x"91",
          5724 => x"38",
          5725 => x"19",
          5726 => x"54",
          5727 => x"70",
          5728 => x"34",
          5729 => x"ec",
          5730 => x"34",
          5731 => x"c8",
          5732 => x"0d",
          5733 => x"0d",
          5734 => x"3d",
          5735 => x"71",
          5736 => x"ea",
          5737 => x"93",
          5738 => x"82",
          5739 => x"8a",
          5740 => x"33",
          5741 => x"2e",
          5742 => x"55",
          5743 => x"8c",
          5744 => x"27",
          5745 => x"17",
          5746 => x"2a",
          5747 => x"51",
          5748 => x"85",
          5749 => x"08",
          5750 => x"08",
          5751 => x"94",
          5752 => x"77",
          5753 => x"b3",
          5754 => x"11",
          5755 => x"2b",
          5756 => x"75",
          5757 => x"38",
          5758 => x"18",
          5759 => x"b9",
          5760 => x"c8",
          5761 => x"7a",
          5762 => x"57",
          5763 => x"a9",
          5764 => x"c8",
          5765 => x"95",
          5766 => x"76",
          5767 => x"0c",
          5768 => x"08",
          5769 => x"08",
          5770 => x"c9",
          5771 => x"08",
          5772 => x"38",
          5773 => x"51",
          5774 => x"82",
          5775 => x"56",
          5776 => x"08",
          5777 => x"81",
          5778 => x"82",
          5779 => x"34",
          5780 => x"e3",
          5781 => x"c8",
          5782 => x"09",
          5783 => x"38",
          5784 => x"18",
          5785 => x"82",
          5786 => x"93",
          5787 => x"18",
          5788 => x"18",
          5789 => x"2e",
          5790 => x"78",
          5791 => x"ea",
          5792 => x"31",
          5793 => x"1a",
          5794 => x"90",
          5795 => x"81",
          5796 => x"06",
          5797 => x"58",
          5798 => x"9a",
          5799 => x"76",
          5800 => x"3f",
          5801 => x"08",
          5802 => x"c8",
          5803 => x"82",
          5804 => x"58",
          5805 => x"52",
          5806 => x"ae",
          5807 => x"c8",
          5808 => x"ff",
          5809 => x"38",
          5810 => x"8a",
          5811 => x"98",
          5812 => x"26",
          5813 => x"0b",
          5814 => x"82",
          5815 => x"39",
          5816 => x"0c",
          5817 => x"ff",
          5818 => x"17",
          5819 => x"18",
          5820 => x"ff",
          5821 => x"80",
          5822 => x"75",
          5823 => x"c1",
          5824 => x"93",
          5825 => x"38",
          5826 => x"18",
          5827 => x"81",
          5828 => x"89",
          5829 => x"c8",
          5830 => x"8c",
          5831 => x"18",
          5832 => x"38",
          5833 => x"8c",
          5834 => x"17",
          5835 => x"07",
          5836 => x"18",
          5837 => x"08",
          5838 => x"55",
          5839 => x"80",
          5840 => x"17",
          5841 => x"80",
          5842 => x"17",
          5843 => x"2b",
          5844 => x"80",
          5845 => x"81",
          5846 => x"08",
          5847 => x"52",
          5848 => x"33",
          5849 => x"b8",
          5850 => x"93",
          5851 => x"2e",
          5852 => x"0b",
          5853 => x"81",
          5854 => x"90",
          5855 => x"ff",
          5856 => x"90",
          5857 => x"54",
          5858 => x"17",
          5859 => x"11",
          5860 => x"ff",
          5861 => x"82",
          5862 => x"80",
          5863 => x"81",
          5864 => x"34",
          5865 => x"39",
          5866 => x"18",
          5867 => x"87",
          5868 => x"18",
          5869 => x"74",
          5870 => x"0c",
          5871 => x"04",
          5872 => x"79",
          5873 => x"75",
          5874 => x"8f",
          5875 => x"89",
          5876 => x"52",
          5877 => x"05",
          5878 => x"3f",
          5879 => x"08",
          5880 => x"c8",
          5881 => x"38",
          5882 => x"7a",
          5883 => x"d8",
          5884 => x"93",
          5885 => x"82",
          5886 => x"80",
          5887 => x"16",
          5888 => x"2b",
          5889 => x"74",
          5890 => x"86",
          5891 => x"84",
          5892 => x"06",
          5893 => x"73",
          5894 => x"38",
          5895 => x"52",
          5896 => x"c4",
          5897 => x"c8",
          5898 => x"0c",
          5899 => x"55",
          5900 => x"77",
          5901 => x"22",
          5902 => x"74",
          5903 => x"c9",
          5904 => x"93",
          5905 => x"74",
          5906 => x"81",
          5907 => x"85",
          5908 => x"2e",
          5909 => x"76",
          5910 => x"73",
          5911 => x"0c",
          5912 => x"04",
          5913 => x"76",
          5914 => x"05",
          5915 => x"54",
          5916 => x"82",
          5917 => x"53",
          5918 => x"08",
          5919 => x"93",
          5920 => x"0c",
          5921 => x"c8",
          5922 => x"0d",
          5923 => x"0d",
          5924 => x"3d",
          5925 => x"71",
          5926 => x"e4",
          5927 => x"93",
          5928 => x"82",
          5929 => x"80",
          5930 => x"92",
          5931 => x"c8",
          5932 => x"51",
          5933 => x"82",
          5934 => x"53",
          5935 => x"52",
          5936 => x"8b",
          5937 => x"c8",
          5938 => x"93",
          5939 => x"2e",
          5940 => x"83",
          5941 => x"72",
          5942 => x"52",
          5943 => x"b4",
          5944 => x"73",
          5945 => x"3f",
          5946 => x"08",
          5947 => x"c8",
          5948 => x"09",
          5949 => x"38",
          5950 => x"82",
          5951 => x"87",
          5952 => x"ef",
          5953 => x"56",
          5954 => x"3d",
          5955 => x"3d",
          5956 => x"cb",
          5957 => x"c8",
          5958 => x"93",
          5959 => x"38",
          5960 => x"51",
          5961 => x"82",
          5962 => x"55",
          5963 => x"08",
          5964 => x"80",
          5965 => x"70",
          5966 => x"57",
          5967 => x"85",
          5968 => x"90",
          5969 => x"2e",
          5970 => x"52",
          5971 => x"05",
          5972 => x"3f",
          5973 => x"c8",
          5974 => x"0d",
          5975 => x"0d",
          5976 => x"5a",
          5977 => x"3d",
          5978 => x"91",
          5979 => x"ef",
          5980 => x"c8",
          5981 => x"93",
          5982 => x"84",
          5983 => x"0c",
          5984 => x"11",
          5985 => x"55",
          5986 => x"08",
          5987 => x"38",
          5988 => x"7a",
          5989 => x"39",
          5990 => x"cf",
          5991 => x"81",
          5992 => x"7b",
          5993 => x"56",
          5994 => x"2e",
          5995 => x"80",
          5996 => x"75",
          5997 => x"52",
          5998 => x"05",
          5999 => x"aa",
          6000 => x"c8",
          6001 => x"d0",
          6002 => x"c8",
          6003 => x"cd",
          6004 => x"c8",
          6005 => x"82",
          6006 => x"07",
          6007 => x"05",
          6008 => x"53",
          6009 => x"98",
          6010 => x"26",
          6011 => x"fb",
          6012 => x"11",
          6013 => x"08",
          6014 => x"80",
          6015 => x"38",
          6016 => x"18",
          6017 => x"ff",
          6018 => x"82",
          6019 => x"59",
          6020 => x"08",
          6021 => x"7a",
          6022 => x"54",
          6023 => x"09",
          6024 => x"38",
          6025 => x"05",
          6026 => x"f0",
          6027 => x"c8",
          6028 => x"ff",
          6029 => x"70",
          6030 => x"82",
          6031 => x"51",
          6032 => x"7a",
          6033 => x"51",
          6034 => x"3f",
          6035 => x"08",
          6036 => x"70",
          6037 => x"25",
          6038 => x"58",
          6039 => x"74",
          6040 => x"ff",
          6041 => x"75",
          6042 => x"76",
          6043 => x"77",
          6044 => x"54",
          6045 => x"33",
          6046 => x"55",
          6047 => x"34",
          6048 => x"c8",
          6049 => x"0d",
          6050 => x"0d",
          6051 => x"fc",
          6052 => x"52",
          6053 => x"3f",
          6054 => x"08",
          6055 => x"c8",
          6056 => x"91",
          6057 => x"76",
          6058 => x"38",
          6059 => x"dc",
          6060 => x"33",
          6061 => x"70",
          6062 => x"56",
          6063 => x"74",
          6064 => x"c8",
          6065 => x"08",
          6066 => x"27",
          6067 => x"94",
          6068 => x"38",
          6069 => x"18",
          6070 => x"51",
          6071 => x"3f",
          6072 => x"08",
          6073 => x"88",
          6074 => x"ca",
          6075 => x"08",
          6076 => x"ff",
          6077 => x"82",
          6078 => x"82",
          6079 => x"ff",
          6080 => x"70",
          6081 => x"25",
          6082 => x"56",
          6083 => x"08",
          6084 => x"81",
          6085 => x"82",
          6086 => x"38",
          6087 => x"98",
          6088 => x"92",
          6089 => x"08",
          6090 => x"77",
          6091 => x"fe",
          6092 => x"c8",
          6093 => x"18",
          6094 => x"0c",
          6095 => x"80",
          6096 => x"74",
          6097 => x"76",
          6098 => x"98",
          6099 => x"80",
          6100 => x"81",
          6101 => x"08",
          6102 => x"52",
          6103 => x"33",
          6104 => x"b0",
          6105 => x"93",
          6106 => x"2e",
          6107 => x"57",
          6108 => x"18",
          6109 => x"06",
          6110 => x"19",
          6111 => x"2e",
          6112 => x"91",
          6113 => x"56",
          6114 => x"56",
          6115 => x"c8",
          6116 => x"0d",
          6117 => x"0d",
          6118 => x"51",
          6119 => x"3f",
          6120 => x"3d",
          6121 => x"52",
          6122 => x"d6",
          6123 => x"93",
          6124 => x"82",
          6125 => x"82",
          6126 => x"fb",
          6127 => x"96",
          6128 => x"44",
          6129 => x"3d",
          6130 => x"d0",
          6131 => x"93",
          6132 => x"fb",
          6133 => x"ff",
          6134 => x"75",
          6135 => x"02",
          6136 => x"33",
          6137 => x"70",
          6138 => x"55",
          6139 => x"2e",
          6140 => x"56",
          6141 => x"38",
          6142 => x"51",
          6143 => x"3f",
          6144 => x"05",
          6145 => x"2b",
          6146 => x"80",
          6147 => x"86",
          6148 => x"02",
          6149 => x"33",
          6150 => x"73",
          6151 => x"38",
          6152 => x"81",
          6153 => x"52",
          6154 => x"bc",
          6155 => x"c8",
          6156 => x"05",
          6157 => x"33",
          6158 => x"70",
          6159 => x"56",
          6160 => x"80",
          6161 => x"38",
          6162 => x"51",
          6163 => x"3f",
          6164 => x"56",
          6165 => x"77",
          6166 => x"38",
          6167 => x"51",
          6168 => x"3f",
          6169 => x"5b",
          6170 => x"51",
          6171 => x"3f",
          6172 => x"3d",
          6173 => x"c1",
          6174 => x"93",
          6175 => x"82",
          6176 => x"81",
          6177 => x"93",
          6178 => x"73",
          6179 => x"3f",
          6180 => x"08",
          6181 => x"c8",
          6182 => x"87",
          6183 => x"32",
          6184 => x"72",
          6185 => x"78",
          6186 => x"54",
          6187 => x"38",
          6188 => x"51",
          6189 => x"3f",
          6190 => x"05",
          6191 => x"3f",
          6192 => x"08",
          6193 => x"08",
          6194 => x"93",
          6195 => x"80",
          6196 => x"70",
          6197 => x"2a",
          6198 => x"57",
          6199 => x"74",
          6200 => x"38",
          6201 => x"51",
          6202 => x"3f",
          6203 => x"52",
          6204 => x"05",
          6205 => x"b6",
          6206 => x"c8",
          6207 => x"8c",
          6208 => x"ff",
          6209 => x"82",
          6210 => x"56",
          6211 => x"51",
          6212 => x"3f",
          6213 => x"c8",
          6214 => x"0d",
          6215 => x"0d",
          6216 => x"3d",
          6217 => x"99",
          6218 => x"b3",
          6219 => x"c8",
          6220 => x"93",
          6221 => x"b5",
          6222 => x"68",
          6223 => x"d4",
          6224 => x"cb",
          6225 => x"c8",
          6226 => x"93",
          6227 => x"38",
          6228 => x"84",
          6229 => x"06",
          6230 => x"02",
          6231 => x"33",
          6232 => x"70",
          6233 => x"55",
          6234 => x"2e",
          6235 => x"55",
          6236 => x"09",
          6237 => x"f5",
          6238 => x"80",
          6239 => x"c4",
          6240 => x"ba",
          6241 => x"93",
          6242 => x"80",
          6243 => x"c8",
          6244 => x"09",
          6245 => x"38",
          6246 => x"81",
          6247 => x"06",
          6248 => x"55",
          6249 => x"09",
          6250 => x"38",
          6251 => x"88",
          6252 => x"74",
          6253 => x"75",
          6254 => x"ff",
          6255 => x"82",
          6256 => x"55",
          6257 => x"08",
          6258 => x"8b",
          6259 => x"b4",
          6260 => x"af",
          6261 => x"54",
          6262 => x"15",
          6263 => x"90",
          6264 => x"34",
          6265 => x"ca",
          6266 => x"af",
          6267 => x"53",
          6268 => x"77",
          6269 => x"3f",
          6270 => x"18",
          6271 => x"18",
          6272 => x"a7",
          6273 => x"ae",
          6274 => x"15",
          6275 => x"80",
          6276 => x"77",
          6277 => x"3f",
          6278 => x"0b",
          6279 => x"98",
          6280 => x"51",
          6281 => x"82",
          6282 => x"55",
          6283 => x"08",
          6284 => x"52",
          6285 => x"51",
          6286 => x"3f",
          6287 => x"52",
          6288 => x"dd",
          6289 => x"90",
          6290 => x"34",
          6291 => x"0b",
          6292 => x"77",
          6293 => x"b9",
          6294 => x"c8",
          6295 => x"39",
          6296 => x"52",
          6297 => x"05",
          6298 => x"c2",
          6299 => x"93",
          6300 => x"3d",
          6301 => x"3d",
          6302 => x"84",
          6303 => x"c8",
          6304 => x"a7",
          6305 => x"05",
          6306 => x"51",
          6307 => x"82",
          6308 => x"55",
          6309 => x"08",
          6310 => x"77",
          6311 => x"08",
          6312 => x"d4",
          6313 => x"e7",
          6314 => x"c8",
          6315 => x"93",
          6316 => x"bd",
          6317 => x"97",
          6318 => x"a0",
          6319 => x"80",
          6320 => x"86",
          6321 => x"a9",
          6322 => x"a3",
          6323 => x"a7",
          6324 => x"05",
          6325 => x"d3",
          6326 => x"a7",
          6327 => x"52",
          6328 => x"52",
          6329 => x"c3",
          6330 => x"08",
          6331 => x"ca",
          6332 => x"93",
          6333 => x"82",
          6334 => x"94",
          6335 => x"2e",
          6336 => x"8a",
          6337 => x"64",
          6338 => x"2e",
          6339 => x"55",
          6340 => x"09",
          6341 => x"b8",
          6342 => x"ff",
          6343 => x"c3",
          6344 => x"93",
          6345 => x"82",
          6346 => x"81",
          6347 => x"56",
          6348 => x"3d",
          6349 => x"52",
          6350 => x"ff",
          6351 => x"02",
          6352 => x"8b",
          6353 => x"16",
          6354 => x"2a",
          6355 => x"51",
          6356 => x"89",
          6357 => x"07",
          6358 => x"17",
          6359 => x"81",
          6360 => x"34",
          6361 => x"70",
          6362 => x"81",
          6363 => x"57",
          6364 => x"80",
          6365 => x"63",
          6366 => x"38",
          6367 => x"51",
          6368 => x"3f",
          6369 => x"08",
          6370 => x"ff",
          6371 => x"82",
          6372 => x"c8",
          6373 => x"b8",
          6374 => x"c8",
          6375 => x"51",
          6376 => x"3f",
          6377 => x"08",
          6378 => x"57",
          6379 => x"c8",
          6380 => x"81",
          6381 => x"73",
          6382 => x"81",
          6383 => x"62",
          6384 => x"77",
          6385 => x"d9",
          6386 => x"81",
          6387 => x"34",
          6388 => x"a7",
          6389 => x"51",
          6390 => x"82",
          6391 => x"55",
          6392 => x"08",
          6393 => x"51",
          6394 => x"3f",
          6395 => x"08",
          6396 => x"93",
          6397 => x"3d",
          6398 => x"3d",
          6399 => x"db",
          6400 => x"84",
          6401 => x"05",
          6402 => x"82",
          6403 => x"d0",
          6404 => x"3d",
          6405 => x"3f",
          6406 => x"08",
          6407 => x"c8",
          6408 => x"38",
          6409 => x"52",
          6410 => x"05",
          6411 => x"3f",
          6412 => x"08",
          6413 => x"c8",
          6414 => x"02",
          6415 => x"33",
          6416 => x"54",
          6417 => x"83",
          6418 => x"74",
          6419 => x"a7",
          6420 => x"09",
          6421 => x"71",
          6422 => x"06",
          6423 => x"55",
          6424 => x"15",
          6425 => x"81",
          6426 => x"34",
          6427 => x"ad",
          6428 => x"93",
          6429 => x"74",
          6430 => x"0c",
          6431 => x"04",
          6432 => x"65",
          6433 => x"94",
          6434 => x"52",
          6435 => x"cc",
          6436 => x"93",
          6437 => x"82",
          6438 => x"80",
          6439 => x"59",
          6440 => x"3d",
          6441 => x"c6",
          6442 => x"93",
          6443 => x"82",
          6444 => x"bc",
          6445 => x"cb",
          6446 => x"a0",
          6447 => x"80",
          6448 => x"86",
          6449 => x"38",
          6450 => x"84",
          6451 => x"90",
          6452 => x"54",
          6453 => x"96",
          6454 => x"a9",
          6455 => x"54",
          6456 => x"15",
          6457 => x"ff",
          6458 => x"82",
          6459 => x"55",
          6460 => x"c8",
          6461 => x"0d",
          6462 => x"0d",
          6463 => x"59",
          6464 => x"3d",
          6465 => x"99",
          6466 => x"d3",
          6467 => x"c8",
          6468 => x"c8",
          6469 => x"82",
          6470 => x"07",
          6471 => x"30",
          6472 => x"9f",
          6473 => x"52",
          6474 => x"56",
          6475 => x"80",
          6476 => x"5d",
          6477 => x"52",
          6478 => x"52",
          6479 => x"bb",
          6480 => x"c8",
          6481 => x"93",
          6482 => x"ce",
          6483 => x"73",
          6484 => x"fb",
          6485 => x"c8",
          6486 => x"93",
          6487 => x"38",
          6488 => x"08",
          6489 => x"08",
          6490 => x"58",
          6491 => x"18",
          6492 => x"58",
          6493 => x"74",
          6494 => x"58",
          6495 => x"ec",
          6496 => x"54",
          6497 => x"77",
          6498 => x"38",
          6499 => x"11",
          6500 => x"55",
          6501 => x"2e",
          6502 => x"84",
          6503 => x"06",
          6504 => x"79",
          6505 => x"75",
          6506 => x"07",
          6507 => x"30",
          6508 => x"9f",
          6509 => x"52",
          6510 => x"74",
          6511 => x"38",
          6512 => x"08",
          6513 => x"aa",
          6514 => x"93",
          6515 => x"82",
          6516 => x"a7",
          6517 => x"33",
          6518 => x"c3",
          6519 => x"2e",
          6520 => x"e4",
          6521 => x"2e",
          6522 => x"58",
          6523 => x"05",
          6524 => x"c1",
          6525 => x"c8",
          6526 => x"75",
          6527 => x"0c",
          6528 => x"04",
          6529 => x"82",
          6530 => x"ff",
          6531 => x"9b",
          6532 => x"cb",
          6533 => x"c8",
          6534 => x"93",
          6535 => x"c8",
          6536 => x"a0",
          6537 => x"ff",
          6538 => x"ff",
          6539 => x"80",
          6540 => x"33",
          6541 => x"57",
          6542 => x"81",
          6543 => x"33",
          6544 => x"4c",
          6545 => x"06",
          6546 => x"a7",
          6547 => x"93",
          6548 => x"2e",
          6549 => x"70",
          6550 => x"51",
          6551 => x"f2",
          6552 => x"c8",
          6553 => x"8d",
          6554 => x"2b",
          6555 => x"81",
          6556 => x"83",
          6557 => x"ff",
          6558 => x"73",
          6559 => x"38",
          6560 => x"83",
          6561 => x"57",
          6562 => x"76",
          6563 => x"81",
          6564 => x"33",
          6565 => x"2e",
          6566 => x"52",
          6567 => x"51",
          6568 => x"3f",
          6569 => x"08",
          6570 => x"ff",
          6571 => x"38",
          6572 => x"88",
          6573 => x"8a",
          6574 => x"38",
          6575 => x"a8",
          6576 => x"76",
          6577 => x"9a",
          6578 => x"ff",
          6579 => x"88",
          6580 => x"73",
          6581 => x"17",
          6582 => x"77",
          6583 => x"05",
          6584 => x"34",
          6585 => x"70",
          6586 => x"57",
          6587 => x"fe",
          6588 => x"3d",
          6589 => x"55",
          6590 => x"2e",
          6591 => x"76",
          6592 => x"38",
          6593 => x"70",
          6594 => x"33",
          6595 => x"54",
          6596 => x"09",
          6597 => x"38",
          6598 => x"76",
          6599 => x"38",
          6600 => x"33",
          6601 => x"a0",
          6602 => x"77",
          6603 => x"80",
          6604 => x"70",
          6605 => x"b3",
          6606 => x"93",
          6607 => x"82",
          6608 => x"81",
          6609 => x"52",
          6610 => x"b9",
          6611 => x"93",
          6612 => x"82",
          6613 => x"b0",
          6614 => x"2e",
          6615 => x"53",
          6616 => x"bc",
          6617 => x"51",
          6618 => x"3f",
          6619 => x"54",
          6620 => x"77",
          6621 => x"83",
          6622 => x"51",
          6623 => x"3f",
          6624 => x"08",
          6625 => x"39",
          6626 => x"08",
          6627 => x"81",
          6628 => x"38",
          6629 => x"74",
          6630 => x"38",
          6631 => x"3d",
          6632 => x"ff",
          6633 => x"82",
          6634 => x"54",
          6635 => x"08",
          6636 => x"53",
          6637 => x"08",
          6638 => x"ff",
          6639 => x"65",
          6640 => x"8b",
          6641 => x"53",
          6642 => x"bc",
          6643 => x"51",
          6644 => x"3f",
          6645 => x"0b",
          6646 => x"77",
          6647 => x"b1",
          6648 => x"c8",
          6649 => x"55",
          6650 => x"c8",
          6651 => x"0d",
          6652 => x"0d",
          6653 => x"88",
          6654 => x"05",
          6655 => x"fc",
          6656 => x"54",
          6657 => x"cd",
          6658 => x"93",
          6659 => x"82",
          6660 => x"8a",
          6661 => x"33",
          6662 => x"2e",
          6663 => x"54",
          6664 => x"7a",
          6665 => x"38",
          6666 => x"90",
          6667 => x"33",
          6668 => x"70",
          6669 => x"55",
          6670 => x"38",
          6671 => x"99",
          6672 => x"81",
          6673 => x"57",
          6674 => x"7f",
          6675 => x"70",
          6676 => x"55",
          6677 => x"51",
          6678 => x"dd",
          6679 => x"7b",
          6680 => x"70",
          6681 => x"2a",
          6682 => x"08",
          6683 => x"11",
          6684 => x"40",
          6685 => x"5f",
          6686 => x"88",
          6687 => x"08",
          6688 => x"38",
          6689 => x"79",
          6690 => x"5a",
          6691 => x"51",
          6692 => x"3f",
          6693 => x"08",
          6694 => x"56",
          6695 => x"14",
          6696 => x"83",
          6697 => x"75",
          6698 => x"95",
          6699 => x"2e",
          6700 => x"75",
          6701 => x"1a",
          6702 => x"2e",
          6703 => x"39",
          6704 => x"5a",
          6705 => x"09",
          6706 => x"38",
          6707 => x"81",
          6708 => x"80",
          6709 => x"7c",
          6710 => x"7d",
          6711 => x"38",
          6712 => x"75",
          6713 => x"81",
          6714 => x"ff",
          6715 => x"74",
          6716 => x"ff",
          6717 => x"82",
          6718 => x"57",
          6719 => x"08",
          6720 => x"81",
          6721 => x"58",
          6722 => x"d4",
          6723 => x"ff",
          6724 => x"80",
          6725 => x"7f",
          6726 => x"54",
          6727 => x"b7",
          6728 => x"19",
          6729 => x"19",
          6730 => x"33",
          6731 => x"54",
          6732 => x"34",
          6733 => x"08",
          6734 => x"55",
          6735 => x"74",
          6736 => x"90",
          6737 => x"31",
          6738 => x"7f",
          6739 => x"81",
          6740 => x"73",
          6741 => x"76",
          6742 => x"93",
          6743 => x"3d",
          6744 => x"3d",
          6745 => x"84",
          6746 => x"05",
          6747 => x"53",
          6748 => x"bf",
          6749 => x"93",
          6750 => x"8b",
          6751 => x"82",
          6752 => x"24",
          6753 => x"82",
          6754 => x"10",
          6755 => x"e4",
          6756 => x"08",
          6757 => x"38",
          6758 => x"80",
          6759 => x"81",
          6760 => x"81",
          6761 => x"ff",
          6762 => x"82",
          6763 => x"81",
          6764 => x"81",
          6765 => x"83",
          6766 => x"9b",
          6767 => x"2a",
          6768 => x"51",
          6769 => x"74",
          6770 => x"98",
          6771 => x"53",
          6772 => x"51",
          6773 => x"3f",
          6774 => x"08",
          6775 => x"80",
          6776 => x"66",
          6777 => x"26",
          6778 => x"ff",
          6779 => x"55",
          6780 => x"83",
          6781 => x"84",
          6782 => x"80",
          6783 => x"7d",
          6784 => x"38",
          6785 => x"0a",
          6786 => x"ff",
          6787 => x"55",
          6788 => x"86",
          6789 => x"8b",
          6790 => x"52",
          6791 => x"f6",
          6792 => x"93",
          6793 => x"7f",
          6794 => x"40",
          6795 => x"89",
          6796 => x"c8",
          6797 => x"93",
          6798 => x"60",
          6799 => x"07",
          6800 => x"93",
          6801 => x"70",
          6802 => x"08",
          6803 => x"72",
          6804 => x"51",
          6805 => x"91",
          6806 => x"fb",
          6807 => x"f8",
          6808 => x"52",
          6809 => x"9c",
          6810 => x"57",
          6811 => x"08",
          6812 => x"7c",
          6813 => x"81",
          6814 => x"80",
          6815 => x"2e",
          6816 => x"83",
          6817 => x"8e",
          6818 => x"26",
          6819 => x"65",
          6820 => x"8e",
          6821 => x"66",
          6822 => x"38",
          6823 => x"81",
          6824 => x"b3",
          6825 => x"2a",
          6826 => x"51",
          6827 => x"2e",
          6828 => x"87",
          6829 => x"82",
          6830 => x"7c",
          6831 => x"74",
          6832 => x"42",
          6833 => x"81",
          6834 => x"57",
          6835 => x"80",
          6836 => x"38",
          6837 => x"83",
          6838 => x"06",
          6839 => x"77",
          6840 => x"91",
          6841 => x"57",
          6842 => x"fd",
          6843 => x"22",
          6844 => x"59",
          6845 => x"9d",
          6846 => x"26",
          6847 => x"1b",
          6848 => x"10",
          6849 => x"51",
          6850 => x"74",
          6851 => x"38",
          6852 => x"ea",
          6853 => x"65",
          6854 => x"9d",
          6855 => x"c8",
          6856 => x"c8",
          6857 => x"1f",
          6858 => x"05",
          6859 => x"f4",
          6860 => x"93",
          6861 => x"a0",
          6862 => x"fc",
          6863 => x"56",
          6864 => x"f0",
          6865 => x"81",
          6866 => x"57",
          6867 => x"77",
          6868 => x"8c",
          6869 => x"57",
          6870 => x"fd",
          6871 => x"22",
          6872 => x"59",
          6873 => x"9d",
          6874 => x"26",
          6875 => x"1b",
          6876 => x"10",
          6877 => x"51",
          6878 => x"74",
          6879 => x"38",
          6880 => x"ea",
          6881 => x"65",
          6882 => x"ad",
          6883 => x"c8",
          6884 => x"05",
          6885 => x"c8",
          6886 => x"26",
          6887 => x"0b",
          6888 => x"08",
          6889 => x"70",
          6890 => x"05",
          6891 => x"7d",
          6892 => x"ff",
          6893 => x"f3",
          6894 => x"93",
          6895 => x"81",
          6896 => x"81",
          6897 => x"fe",
          6898 => x"82",
          6899 => x"83",
          6900 => x"43",
          6901 => x"11",
          6902 => x"11",
          6903 => x"30",
          6904 => x"73",
          6905 => x"59",
          6906 => x"83",
          6907 => x"06",
          6908 => x"1b",
          6909 => x"5b",
          6910 => x"1c",
          6911 => x"29",
          6912 => x"31",
          6913 => x"66",
          6914 => x"38",
          6915 => x"7c",
          6916 => x"70",
          6917 => x"56",
          6918 => x"3f",
          6919 => x"08",
          6920 => x"2e",
          6921 => x"9b",
          6922 => x"c8",
          6923 => x"f5",
          6924 => x"77",
          6925 => x"81",
          6926 => x"fd",
          6927 => x"57",
          6928 => x"61",
          6929 => x"81",
          6930 => x"38",
          6931 => x"76",
          6932 => x"77",
          6933 => x"19",
          6934 => x"c0",
          6935 => x"74",
          6936 => x"39",
          6937 => x"81",
          6938 => x"80",
          6939 => x"83",
          6940 => x"39",
          6941 => x"78",
          6942 => x"80",
          6943 => x"d4",
          6944 => x"86",
          6945 => x"9f",
          6946 => x"38",
          6947 => x"78",
          6948 => x"80",
          6949 => x"bc",
          6950 => x"86",
          6951 => x"55",
          6952 => x"09",
          6953 => x"38",
          6954 => x"9f",
          6955 => x"06",
          6956 => x"74",
          6957 => x"7d",
          6958 => x"7e",
          6959 => x"8f",
          6960 => x"81",
          6961 => x"7e",
          6962 => x"df",
          6963 => x"8b",
          6964 => x"99",
          6965 => x"7f",
          6966 => x"7a",
          6967 => x"06",
          6968 => x"51",
          6969 => x"3f",
          6970 => x"05",
          6971 => x"32",
          6972 => x"96",
          6973 => x"06",
          6974 => x"91",
          6975 => x"98",
          6976 => x"83",
          6977 => x"90",
          6978 => x"d6",
          6979 => x"93",
          6980 => x"98",
          6981 => x"39",
          6982 => x"1f",
          6983 => x"dc",
          6984 => x"95",
          6985 => x"52",
          6986 => x"ff",
          6987 => x"81",
          6988 => x"1f",
          6989 => x"a6",
          6990 => x"9c",
          6991 => x"98",
          6992 => x"83",
          6993 => x"06",
          6994 => x"82",
          6995 => x"52",
          6996 => x"51",
          6997 => x"3f",
          6998 => x"1f",
          6999 => x"9c",
          7000 => x"ac",
          7001 => x"98",
          7002 => x"52",
          7003 => x"ff",
          7004 => x"86",
          7005 => x"51",
          7006 => x"3f",
          7007 => x"80",
          7008 => x"a9",
          7009 => x"05",
          7010 => x"81",
          7011 => x"80",
          7012 => x"ff",
          7013 => x"b2",
          7014 => x"b2",
          7015 => x"1f",
          7016 => x"d8",
          7017 => x"ff",
          7018 => x"96",
          7019 => x"97",
          7020 => x"80",
          7021 => x"34",
          7022 => x"05",
          7023 => x"81",
          7024 => x"ab",
          7025 => x"97",
          7026 => x"d4",
          7027 => x"fe",
          7028 => x"97",
          7029 => x"54",
          7030 => x"52",
          7031 => x"93",
          7032 => x"57",
          7033 => x"08",
          7034 => x"61",
          7035 => x"81",
          7036 => x"38",
          7037 => x"86",
          7038 => x"52",
          7039 => x"93",
          7040 => x"53",
          7041 => x"51",
          7042 => x"3f",
          7043 => x"a4",
          7044 => x"51",
          7045 => x"3f",
          7046 => x"e4",
          7047 => x"e4",
          7048 => x"96",
          7049 => x"16",
          7050 => x"1f",
          7051 => x"cc",
          7052 => x"83",
          7053 => x"ff",
          7054 => x"82",
          7055 => x"83",
          7056 => x"ff",
          7057 => x"81",
          7058 => x"05",
          7059 => x"79",
          7060 => x"86",
          7061 => x"63",
          7062 => x"7e",
          7063 => x"ff",
          7064 => x"64",
          7065 => x"7e",
          7066 => x"e3",
          7067 => x"80",
          7068 => x"2e",
          7069 => x"9e",
          7070 => x"7e",
          7071 => x"fc",
          7072 => x"84",
          7073 => x"95",
          7074 => x"0a",
          7075 => x"51",
          7076 => x"3f",
          7077 => x"ff",
          7078 => x"61",
          7079 => x"38",
          7080 => x"52",
          7081 => x"95",
          7082 => x"55",
          7083 => x"61",
          7084 => x"74",
          7085 => x"75",
          7086 => x"79",
          7087 => x"9a",
          7088 => x"c8",
          7089 => x"38",
          7090 => x"52",
          7091 => x"95",
          7092 => x"16",
          7093 => x"56",
          7094 => x"38",
          7095 => x"7a",
          7096 => x"8d",
          7097 => x"61",
          7098 => x"38",
          7099 => x"57",
          7100 => x"83",
          7101 => x"76",
          7102 => x"7e",
          7103 => x"ff",
          7104 => x"82",
          7105 => x"81",
          7106 => x"16",
          7107 => x"56",
          7108 => x"38",
          7109 => x"83",
          7110 => x"86",
          7111 => x"ff",
          7112 => x"38",
          7113 => x"82",
          7114 => x"81",
          7115 => x"2a",
          7116 => x"77",
          7117 => x"7d",
          7118 => x"7e",
          7119 => x"8f",
          7120 => x"d5",
          7121 => x"1f",
          7122 => x"92",
          7123 => x"1f",
          7124 => x"34",
          7125 => x"17",
          7126 => x"82",
          7127 => x"83",
          7128 => x"84",
          7129 => x"66",
          7130 => x"fd",
          7131 => x"51",
          7132 => x"3f",
          7133 => x"17",
          7134 => x"c8",
          7135 => x"bf",
          7136 => x"86",
          7137 => x"93",
          7138 => x"17",
          7139 => x"83",
          7140 => x"ff",
          7141 => x"65",
          7142 => x"1f",
          7143 => x"dc",
          7144 => x"77",
          7145 => x"79",
          7146 => x"ae",
          7147 => x"82",
          7148 => x"a3",
          7149 => x"80",
          7150 => x"ff",
          7151 => x"81",
          7152 => x"c8",
          7153 => x"8d",
          7154 => x"8b",
          7155 => x"87",
          7156 => x"83",
          7157 => x"76",
          7158 => x"0c",
          7159 => x"04",
          7160 => x"73",
          7161 => x"26",
          7162 => x"71",
          7163 => x"f1",
          7164 => x"71",
          7165 => x"81",
          7166 => x"80",
          7167 => x"d4",
          7168 => x"84",
          7169 => x"9e",
          7170 => x"39",
          7171 => x"51",
          7172 => x"3f",
          7173 => x"82",
          7174 => x"ff",
          7175 => x"81",
          7176 => x"82",
          7177 => x"ff",
          7178 => x"a8",
          7179 => x"cc",
          7180 => x"f2",
          7181 => x"39",
          7182 => x"51",
          7183 => x"3f",
          7184 => x"82",
          7185 => x"fe",
          7186 => x"81",
          7187 => x"83",
          7188 => x"ff",
          7189 => x"fc",
          7190 => x"a0",
          7191 => x"c6",
          7192 => x"39",
          7193 => x"51",
          7194 => x"3f",
          7195 => x"82",
          7196 => x"fe",
          7197 => x"80",
          7198 => x"83",
          7199 => x"ff",
          7200 => x"d0",
          7201 => x"94",
          7202 => x"9a",
          7203 => x"39",
          7204 => x"51",
          7205 => x"3f",
          7206 => x"84",
          7207 => x"ff",
          7208 => x"39",
          7209 => x"51",
          7210 => x"3f",
          7211 => x"84",
          7212 => x"fe",
          7213 => x"39",
          7214 => x"51",
          7215 => x"3f",
          7216 => x"85",
          7217 => x"fe",
          7218 => x"39",
          7219 => x"51",
          7220 => x"3f",
          7221 => x"04",
          7222 => x"77",
          7223 => x"74",
          7224 => x"93",
          7225 => x"75",
          7226 => x"51",
          7227 => x"3f",
          7228 => x"08",
          7229 => x"87",
          7230 => x"51",
          7231 => x"3f",
          7232 => x"08",
          7233 => x"fe",
          7234 => x"82",
          7235 => x"55",
          7236 => x"53",
          7237 => x"85",
          7238 => x"84",
          7239 => x"3d",
          7240 => x"ec",
          7241 => x"97",
          7242 => x"99",
          7243 => x"88",
          7244 => x"05",
          7245 => x"30",
          7246 => x"80",
          7247 => x"75",
          7248 => x"59",
          7249 => x"58",
          7250 => x"81",
          7251 => x"53",
          7252 => x"96",
          7253 => x"05",
          7254 => x"99",
          7255 => x"c8",
          7256 => x"93",
          7257 => x"38",
          7258 => x"08",
          7259 => x"88",
          7260 => x"c8",
          7261 => x"96",
          7262 => x"11",
          7263 => x"80",
          7264 => x"fb",
          7265 => x"c0",
          7266 => x"93",
          7267 => x"82",
          7268 => x"8e",
          7269 => x"2e",
          7270 => x"19",
          7271 => x"59",
          7272 => x"96",
          7273 => x"05",
          7274 => x"3f",
          7275 => x"79",
          7276 => x"7b",
          7277 => x"2a",
          7278 => x"57",
          7279 => x"80",
          7280 => x"82",
          7281 => x"87",
          7282 => x"08",
          7283 => x"fe",
          7284 => x"55",
          7285 => x"c8",
          7286 => x"3d",
          7287 => x"3d",
          7288 => x"05",
          7289 => x"7d",
          7290 => x"53",
          7291 => x"51",
          7292 => x"82",
          7293 => x"a4",
          7294 => x"2e",
          7295 => x"81",
          7296 => x"98",
          7297 => x"60",
          7298 => x"c8",
          7299 => x"7e",
          7300 => x"82",
          7301 => x"59",
          7302 => x"04",
          7303 => x"c8",
          7304 => x"0d",
          7305 => x"0d",
          7306 => x"33",
          7307 => x"53",
          7308 => x"52",
          7309 => x"e8",
          7310 => x"e8",
          7311 => x"55",
          7312 => x"3f",
          7313 => x"54",
          7314 => x"53",
          7315 => x"52",
          7316 => x"51",
          7317 => x"3f",
          7318 => x"85",
          7319 => x"ff",
          7320 => x"0d",
          7321 => x"0d",
          7322 => x"80",
          7323 => x"f9",
          7324 => x"51",
          7325 => x"3f",
          7326 => x"51",
          7327 => x"3f",
          7328 => x"ee",
          7329 => x"81",
          7330 => x"06",
          7331 => x"80",
          7332 => x"81",
          7333 => x"de",
          7334 => x"cc",
          7335 => x"d4",
          7336 => x"fe",
          7337 => x"72",
          7338 => x"81",
          7339 => x"71",
          7340 => x"38",
          7341 => x"ee",
          7342 => x"86",
          7343 => x"f0",
          7344 => x"51",
          7345 => x"3f",
          7346 => x"70",
          7347 => x"52",
          7348 => x"95",
          7349 => x"fe",
          7350 => x"82",
          7351 => x"fe",
          7352 => x"80",
          7353 => x"8e",
          7354 => x"2a",
          7355 => x"51",
          7356 => x"2e",
          7357 => x"51",
          7358 => x"3f",
          7359 => x"51",
          7360 => x"3f",
          7361 => x"ed",
          7362 => x"85",
          7363 => x"06",
          7364 => x"80",
          7365 => x"81",
          7366 => x"da",
          7367 => x"98",
          7368 => x"d0",
          7369 => x"fe",
          7370 => x"72",
          7371 => x"81",
          7372 => x"71",
          7373 => x"38",
          7374 => x"ed",
          7375 => x"87",
          7376 => x"ef",
          7377 => x"51",
          7378 => x"3f",
          7379 => x"70",
          7380 => x"52",
          7381 => x"95",
          7382 => x"fe",
          7383 => x"82",
          7384 => x"fe",
          7385 => x"80",
          7386 => x"8a",
          7387 => x"2a",
          7388 => x"51",
          7389 => x"2e",
          7390 => x"51",
          7391 => x"3f",
          7392 => x"51",
          7393 => x"3f",
          7394 => x"ec",
          7395 => x"f8",
          7396 => x"3d",
          7397 => x"3d",
          7398 => x"08",
          7399 => x"57",
          7400 => x"80",
          7401 => x"39",
          7402 => x"85",
          7403 => x"80",
          7404 => x"15",
          7405 => x"33",
          7406 => x"a0",
          7407 => x"81",
          7408 => x"70",
          7409 => x"06",
          7410 => x"e6",
          7411 => x"53",
          7412 => x"09",
          7413 => x"38",
          7414 => x"81",
          7415 => x"80",
          7416 => x"29",
          7417 => x"05",
          7418 => x"70",
          7419 => x"fe",
          7420 => x"82",
          7421 => x"8b",
          7422 => x"33",
          7423 => x"2e",
          7424 => x"81",
          7425 => x"ff",
          7426 => x"bb",
          7427 => x"38",
          7428 => x"82",
          7429 => x"88",
          7430 => x"ce",
          7431 => x"70",
          7432 => x"72",
          7433 => x"5e",
          7434 => x"81",
          7435 => x"ff",
          7436 => x"82",
          7437 => x"81",
          7438 => x"78",
          7439 => x"81",
          7440 => x"82",
          7441 => x"96",
          7442 => x"59",
          7443 => x"3f",
          7444 => x"52",
          7445 => x"51",
          7446 => x"3f",
          7447 => x"08",
          7448 => x"2e",
          7449 => x"88",
          7450 => x"fd",
          7451 => x"39",
          7452 => x"5c",
          7453 => x"51",
          7454 => x"3f",
          7455 => x"43",
          7456 => x"70",
          7457 => x"52",
          7458 => x"e4",
          7459 => x"52",
          7460 => x"fd",
          7461 => x"3d",
          7462 => x"51",
          7463 => x"82",
          7464 => x"90",
          7465 => x"2c",
          7466 => x"81",
          7467 => x"af",
          7468 => x"10",
          7469 => x"05",
          7470 => x"04",
          7471 => x"f4",
          7472 => x"f8",
          7473 => x"fe",
          7474 => x"93",
          7475 => x"38",
          7476 => x"51",
          7477 => x"3f",
          7478 => x"b4",
          7479 => x"11",
          7480 => x"05",
          7481 => x"c3",
          7482 => x"c8",
          7483 => x"88",
          7484 => x"25",
          7485 => x"40",
          7486 => x"33",
          7487 => x"c3",
          7488 => x"ff",
          7489 => x"82",
          7490 => x"81",
          7491 => x"78",
          7492 => x"88",
          7493 => x"f6",
          7494 => x"5d",
          7495 => x"82",
          7496 => x"fe",
          7497 => x"fe",
          7498 => x"3d",
          7499 => x"53",
          7500 => x"51",
          7501 => x"3f",
          7502 => x"08",
          7503 => x"b4",
          7504 => x"80",
          7505 => x"c3",
          7506 => x"ff",
          7507 => x"82",
          7508 => x"52",
          7509 => x"51",
          7510 => x"3f",
          7511 => x"b4",
          7512 => x"11",
          7513 => x"05",
          7514 => x"bf",
          7515 => x"c8",
          7516 => x"87",
          7517 => x"26",
          7518 => x"b4",
          7519 => x"11",
          7520 => x"05",
          7521 => x"a3",
          7522 => x"c8",
          7523 => x"82",
          7524 => x"40",
          7525 => x"89",
          7526 => x"3d",
          7527 => x"fe",
          7528 => x"02",
          7529 => x"53",
          7530 => x"84",
          7531 => x"a0",
          7532 => x"ff",
          7533 => x"82",
          7534 => x"80",
          7535 => x"82",
          7536 => x"51",
          7537 => x"fd",
          7538 => x"88",
          7539 => x"f4",
          7540 => x"5c",
          7541 => x"b4",
          7542 => x"05",
          7543 => x"a4",
          7544 => x"c8",
          7545 => x"fe",
          7546 => x"5b",
          7547 => x"3f",
          7548 => x"93",
          7549 => x"7a",
          7550 => x"3f",
          7551 => x"08",
          7552 => x"f0",
          7553 => x"c8",
          7554 => x"d4",
          7555 => x"39",
          7556 => x"f8",
          7557 => x"e3",
          7558 => x"93",
          7559 => x"3d",
          7560 => x"52",
          7561 => x"c1",
          7562 => x"c8",
          7563 => x"fe",
          7564 => x"5a",
          7565 => x"3f",
          7566 => x"08",
          7567 => x"f8",
          7568 => x"fe",
          7569 => x"82",
          7570 => x"82",
          7571 => x"80",
          7572 => x"82",
          7573 => x"81",
          7574 => x"78",
          7575 => x"7a",
          7576 => x"3f",
          7577 => x"08",
          7578 => x"88",
          7579 => x"c8",
          7580 => x"ec",
          7581 => x"39",
          7582 => x"51",
          7583 => x"3f",
          7584 => x"f2",
          7585 => x"ec",
          7586 => x"b0",
          7587 => x"96",
          7588 => x"fe",
          7589 => x"fb",
          7590 => x"80",
          7591 => x"c0",
          7592 => x"84",
          7593 => x"87",
          7594 => x"0c",
          7595 => x"51",
          7596 => x"3f",
          7597 => x"82",
          7598 => x"fe",
          7599 => x"8c",
          7600 => x"87",
          7601 => x"0c",
          7602 => x"0b",
          7603 => x"94",
          7604 => x"39",
          7605 => x"f4",
          7606 => x"f8",
          7607 => x"fa",
          7608 => x"93",
          7609 => x"2e",
          7610 => x"60",
          7611 => x"f0",
          7612 => x"ac",
          7613 => x"78",
          7614 => x"fe",
          7615 => x"fe",
          7616 => x"fe",
          7617 => x"82",
          7618 => x"80",
          7619 => x"38",
          7620 => x"8a",
          7621 => x"f8",
          7622 => x"59",
          7623 => x"93",
          7624 => x"82",
          7625 => x"80",
          7626 => x"38",
          7627 => x"08",
          7628 => x"a8",
          7629 => x"e8",
          7630 => x"39",
          7631 => x"51",
          7632 => x"3f",
          7633 => x"3f",
          7634 => x"82",
          7635 => x"fe",
          7636 => x"80",
          7637 => x"39",
          7638 => x"3f",
          7639 => x"61",
          7640 => x"59",
          7641 => x"fa",
          7642 => x"7c",
          7643 => x"80",
          7644 => x"38",
          7645 => x"f8",
          7646 => x"e1",
          7647 => x"8a",
          7648 => x"93",
          7649 => x"82",
          7650 => x"80",
          7651 => x"fc",
          7652 => x"70",
          7653 => x"f7",
          7654 => x"8b",
          7655 => x"93",
          7656 => x"56",
          7657 => x"42",
          7658 => x"54",
          7659 => x"53",
          7660 => x"52",
          7661 => x"a6",
          7662 => x"c8",
          7663 => x"81",
          7664 => x"32",
          7665 => x"8a",
          7666 => x"2e",
          7667 => x"f9",
          7668 => x"8b",
          7669 => x"f6",
          7670 => x"98",
          7671 => x"0d",
          7672 => x"93",
          7673 => x"90",
          7674 => x"87",
          7675 => x"0c",
          7676 => x"e4",
          7677 => x"94",
          7678 => x"80",
          7679 => x"c0",
          7680 => x"8c",
          7681 => x"87",
          7682 => x"0c",
          7683 => x"0b",
          7684 => x"0c",
          7685 => x"0b",
          7686 => x"0c",
          7687 => x"3f",
          7688 => x"3f",
          7689 => x"51",
          7690 => x"3f",
          7691 => x"51",
          7692 => x"3f",
          7693 => x"51",
          7694 => x"3f",
          7695 => x"e5",
          7696 => x"3f",
          7697 => x"00",
          7698 => x"00",
          7699 => x"00",
          7700 => x"00",
          7701 => x"00",
          7702 => x"00",
          7703 => x"00",
          7704 => x"00",
          7705 => x"00",
          7706 => x"00",
          7707 => x"00",
          7708 => x"00",
          7709 => x"00",
          7710 => x"00",
          7711 => x"00",
          7712 => x"00",
          7713 => x"00",
          7714 => x"00",
          7715 => x"00",
          7716 => x"00",
          7717 => x"00",
          7718 => x"00",
          7719 => x"00",
          7720 => x"00",
          7721 => x"00",
          7722 => x"00",
          7723 => x"00",
          7724 => x"00",
          7725 => x"00",
          7726 => x"00",
          7727 => x"00",
          7728 => x"00",
          7729 => x"00",
          7730 => x"00",
          7731 => x"00",
          7732 => x"00",
          7733 => x"00",
          7734 => x"00",
          7735 => x"00",
          7736 => x"00",
          7737 => x"00",
          7738 => x"00",
          7739 => x"00",
          7740 => x"00",
          7741 => x"00",
          7742 => x"00",
          7743 => x"00",
          7744 => x"00",
          7745 => x"00",
          7746 => x"00",
          7747 => x"00",
          7748 => x"00",
          7749 => x"00",
          7750 => x"00",
          7751 => x"00",
          7752 => x"00",
          7753 => x"00",
          7754 => x"00",
          7755 => x"00",
          7756 => x"00",
          7757 => x"00",
          7758 => x"00",
          7759 => x"00",
          7760 => x"00",
          7761 => x"00",
          7762 => x"00",
          7763 => x"00",
          7764 => x"00",
          7765 => x"00",
          7766 => x"00",
          7767 => x"00",
          7768 => x"00",
          7769 => x"00",
          7770 => x"00",
          7771 => x"00",
          7772 => x"00",
          7773 => x"00",
          7774 => x"00",
          7775 => x"00",
          7776 => x"00",
          7777 => x"00",
          7778 => x"00",
          7779 => x"00",
          7780 => x"00",
          7781 => x"00",
          7782 => x"00",
          7783 => x"00",
          7784 => x"00",
          7785 => x"00",
          7786 => x"00",
          7787 => x"00",
          7788 => x"00",
          7789 => x"00",
          7790 => x"00",
          7791 => x"00",
          7792 => x"00",
          7793 => x"00",
          7794 => x"00",
          7795 => x"00",
          7796 => x"00",
          7797 => x"00",
          7798 => x"00",
          7799 => x"00",
          7800 => x"00",
          7801 => x"00",
          7802 => x"00",
          7803 => x"00",
          7804 => x"00",
          7805 => x"00",
          7806 => x"00",
          7807 => x"00",
          7808 => x"00",
          7809 => x"00",
          7810 => x"00",
          7811 => x"00",
          7812 => x"00",
          7813 => x"00",
          7814 => x"00",
          7815 => x"00",
          7816 => x"00",
          7817 => x"00",
          7818 => x"00",
          7819 => x"00",
          7820 => x"00",
          7821 => x"00",
          7822 => x"00",
          7823 => x"00",
          7824 => x"00",
          7825 => x"00",
          7826 => x"00",
          7827 => x"00",
          7828 => x"00",
          7829 => x"00",
          7830 => x"00",
          7831 => x"00",
          7832 => x"00",
          7833 => x"00",
          7834 => x"00",
          7835 => x"00",
          7836 => x"00",
          7837 => x"00",
          7838 => x"00",
          7839 => x"00",
          7840 => x"00",
          7841 => x"00",
          7842 => x"00",
          7843 => x"00",
          7844 => x"00",
          7845 => x"00",
          7846 => x"00",
          7847 => x"00",
          7848 => x"00",
          7849 => x"00",
          7850 => x"00",
          7851 => x"00",
          7852 => x"00",
          7853 => x"00",
          7854 => x"00",
          7855 => x"00",
          7856 => x"00",
          7857 => x"00",
          7858 => x"00",
          7859 => x"00",
          7860 => x"00",
          7861 => x"00",
          7862 => x"00",
          7863 => x"00",
          7864 => x"00",
          7865 => x"00",
          7866 => x"00",
          7867 => x"00",
          7868 => x"00",
          7869 => x"00",
          7870 => x"00",
          7871 => x"00",
          7872 => x"00",
          7873 => x"00",
          7874 => x"00",
          7875 => x"00",
          7876 => x"00",
          7877 => x"00",
          7878 => x"00",
          7879 => x"00",
          7880 => x"00",
          7881 => x"00",
          7882 => x"25",
          7883 => x"64",
          7884 => x"20",
          7885 => x"25",
          7886 => x"64",
          7887 => x"25",
          7888 => x"53",
          7889 => x"43",
          7890 => x"69",
          7891 => x"61",
          7892 => x"6e",
          7893 => x"20",
          7894 => x"6f",
          7895 => x"6f",
          7896 => x"6f",
          7897 => x"67",
          7898 => x"3a",
          7899 => x"76",
          7900 => x"73",
          7901 => x"70",
          7902 => x"65",
          7903 => x"64",
          7904 => x"20",
          7905 => x"49",
          7906 => x"20",
          7907 => x"4d",
          7908 => x"74",
          7909 => x"3d",
          7910 => x"58",
          7911 => x"69",
          7912 => x"25",
          7913 => x"29",
          7914 => x"20",
          7915 => x"42",
          7916 => x"20",
          7917 => x"61",
          7918 => x"25",
          7919 => x"2c",
          7920 => x"7a",
          7921 => x"30",
          7922 => x"2e",
          7923 => x"20",
          7924 => x"52",
          7925 => x"28",
          7926 => x"72",
          7927 => x"30",
          7928 => x"20",
          7929 => x"65",
          7930 => x"38",
          7931 => x"0a",
          7932 => x"20",
          7933 => x"49",
          7934 => x"4c",
          7935 => x"20",
          7936 => x"50",
          7937 => x"00",
          7938 => x"20",
          7939 => x"53",
          7940 => x"00",
          7941 => x"20",
          7942 => x"53",
          7943 => x"61",
          7944 => x"28",
          7945 => x"69",
          7946 => x"3d",
          7947 => x"58",
          7948 => x"00",
          7949 => x"20",
          7950 => x"49",
          7951 => x"52",
          7952 => x"54",
          7953 => x"4e",
          7954 => x"4c",
          7955 => x"0a",
          7956 => x"20",
          7957 => x"54",
          7958 => x"52",
          7959 => x"54",
          7960 => x"72",
          7961 => x"30",
          7962 => x"2e",
          7963 => x"41",
          7964 => x"65",
          7965 => x"73",
          7966 => x"20",
          7967 => x"43",
          7968 => x"52",
          7969 => x"74",
          7970 => x"63",
          7971 => x"20",
          7972 => x"72",
          7973 => x"20",
          7974 => x"30",
          7975 => x"00",
          7976 => x"20",
          7977 => x"43",
          7978 => x"4d",
          7979 => x"72",
          7980 => x"74",
          7981 => x"20",
          7982 => x"72",
          7983 => x"20",
          7984 => x"30",
          7985 => x"00",
          7986 => x"20",
          7987 => x"53",
          7988 => x"6b",
          7989 => x"61",
          7990 => x"41",
          7991 => x"65",
          7992 => x"20",
          7993 => x"20",
          7994 => x"30",
          7995 => x"00",
          7996 => x"20",
          7997 => x"5a",
          7998 => x"49",
          7999 => x"20",
          8000 => x"20",
          8001 => x"20",
          8002 => x"20",
          8003 => x"20",
          8004 => x"30",
          8005 => x"00",
          8006 => x"20",
          8007 => x"53",
          8008 => x"65",
          8009 => x"6c",
          8010 => x"20",
          8011 => x"71",
          8012 => x"20",
          8013 => x"20",
          8014 => x"30",
          8015 => x"00",
          8016 => x"53",
          8017 => x"6c",
          8018 => x"4d",
          8019 => x"75",
          8020 => x"46",
          8021 => x"00",
          8022 => x"45",
          8023 => x"45",
          8024 => x"69",
          8025 => x"55",
          8026 => x"6f",
          8027 => x"53",
          8028 => x"22",
          8029 => x"3a",
          8030 => x"3e",
          8031 => x"7c",
          8032 => x"46",
          8033 => x"46",
          8034 => x"32",
          8035 => x"30",
          8036 => x"31",
          8037 => x"32",
          8038 => x"33",
          8039 => x"35",
          8040 => x"36",
          8041 => x"37",
          8042 => x"38",
          8043 => x"39",
          8044 => x"31",
          8045 => x"eb",
          8046 => x"53",
          8047 => x"35",
          8048 => x"4e",
          8049 => x"41",
          8050 => x"20",
          8051 => x"41",
          8052 => x"20",
          8053 => x"4e",
          8054 => x"41",
          8055 => x"20",
          8056 => x"41",
          8057 => x"20",
          8058 => x"00",
          8059 => x"00",
          8060 => x"00",
          8061 => x"00",
          8062 => x"80",
          8063 => x"8e",
          8064 => x"45",
          8065 => x"49",
          8066 => x"90",
          8067 => x"99",
          8068 => x"59",
          8069 => x"9c",
          8070 => x"41",
          8071 => x"a5",
          8072 => x"a8",
          8073 => x"ac",
          8074 => x"b0",
          8075 => x"b4",
          8076 => x"b8",
          8077 => x"bc",
          8078 => x"c0",
          8079 => x"c4",
          8080 => x"c8",
          8081 => x"cc",
          8082 => x"d0",
          8083 => x"d4",
          8084 => x"d8",
          8085 => x"dc",
          8086 => x"e0",
          8087 => x"e4",
          8088 => x"e8",
          8089 => x"ec",
          8090 => x"f0",
          8091 => x"f4",
          8092 => x"f8",
          8093 => x"fc",
          8094 => x"2b",
          8095 => x"3d",
          8096 => x"5c",
          8097 => x"3c",
          8098 => x"7f",
          8099 => x"00",
          8100 => x"00",
          8101 => x"01",
          8102 => x"00",
          8103 => x"00",
          8104 => x"00",
          8105 => x"00",
          8106 => x"00",
          8107 => x"46",
          8108 => x"32",
          8109 => x"46",
          8110 => x"36",
          8111 => x"65",
          8112 => x"54",
          8113 => x"44",
          8114 => x"20",
          8115 => x"43",
          8116 => x"52",
          8117 => x"00",
          8118 => x"44",
          8119 => x"20",
          8120 => x"46",
          8121 => x"43",
          8122 => x"52",
          8123 => x"00",
          8124 => x"46",
          8125 => x"53",
          8126 => x"45",
          8127 => x"4f",
          8128 => x"4f",
          8129 => x"4d",
          8130 => x"52",
          8131 => x"48",
          8132 => x"57",
          8133 => x"00",
          8134 => x"54",
          8135 => x"49",
          8136 => x"45",
          8137 => x"55",
          8138 => x"4e",
          8139 => x"4d",
          8140 => x"20",
          8141 => x"4d",
          8142 => x"53",
          8143 => x"64",
          8144 => x"70",
          8145 => x"64",
          8146 => x"74",
          8147 => x"64",
          8148 => x"74",
          8149 => x"64",
          8150 => x"74",
          8151 => x"62",
          8152 => x"70",
          8153 => x"62",
          8154 => x"74",
          8155 => x"62",
          8156 => x"64",
          8157 => x"62",
          8158 => x"74",
          8159 => x"62",
          8160 => x"6c",
          8161 => x"62",
          8162 => x"00",
          8163 => x"66",
          8164 => x"74",
          8165 => x"66",
          8166 => x"6e",
          8167 => x"66",
          8168 => x"73",
          8169 => x"66",
          8170 => x"6b",
          8171 => x"66",
          8172 => x"64",
          8173 => x"66",
          8174 => x"70",
          8175 => x"00",
          8176 => x"66",
          8177 => x"74",
          8178 => x"66",
          8179 => x"6e",
          8180 => x"66",
          8181 => x"6f",
          8182 => x"66",
          8183 => x"72",
          8184 => x"66",
          8185 => x"65",
          8186 => x"66",
          8187 => x"61",
          8188 => x"66",
          8189 => x"00",
          8190 => x"66",
          8191 => x"69",
          8192 => x"66",
          8193 => x"74",
          8194 => x"66",
          8195 => x"00",
          8196 => x"66",
          8197 => x"00",
          8198 => x"66",
          8199 => x"66",
          8200 => x"63",
          8201 => x"66",
          8202 => x"61",
          8203 => x"66",
          8204 => x"64",
          8205 => x"66",
          8206 => x"63",
          8207 => x"66",
          8208 => x"65",
          8209 => x"66",
          8210 => x"70",
          8211 => x"66",
          8212 => x"66",
          8213 => x"76",
          8214 => x"66",
          8215 => x"77",
          8216 => x"00",
          8217 => x"66",
          8218 => x"65",
          8219 => x"66",
          8220 => x"73",
          8221 => x"6d",
          8222 => x"00",
          8223 => x"6d",
          8224 => x"70",
          8225 => x"6d",
          8226 => x"6d",
          8227 => x"6d",
          8228 => x"68",
          8229 => x"68",
          8230 => x"68",
          8231 => x"68",
          8232 => x"68",
          8233 => x"68",
          8234 => x"64",
          8235 => x"00",
          8236 => x"63",
          8237 => x"6d",
          8238 => x"00",
          8239 => x"63",
          8240 => x"00",
          8241 => x"6a",
          8242 => x"72",
          8243 => x"61",
          8244 => x"72",
          8245 => x"74",
          8246 => x"68",
          8247 => x"00",
          8248 => x"69",
          8249 => x"00",
          8250 => x"74",
          8251 => x"00",
          8252 => x"74",
          8253 => x"00",
          8254 => x"44",
          8255 => x"20",
          8256 => x"6f",
          8257 => x"49",
          8258 => x"72",
          8259 => x"20",
          8260 => x"6f",
          8261 => x"00",
          8262 => x"44",
          8263 => x"20",
          8264 => x"20",
          8265 => x"64",
          8266 => x"00",
          8267 => x"4e",
          8268 => x"69",
          8269 => x"66",
          8270 => x"64",
          8271 => x"4e",
          8272 => x"61",
          8273 => x"66",
          8274 => x"64",
          8275 => x"49",
          8276 => x"6c",
          8277 => x"66",
          8278 => x"6e",
          8279 => x"2e",
          8280 => x"41",
          8281 => x"73",
          8282 => x"65",
          8283 => x"64",
          8284 => x"46",
          8285 => x"20",
          8286 => x"65",
          8287 => x"20",
          8288 => x"73",
          8289 => x"0a",
          8290 => x"46",
          8291 => x"20",
          8292 => x"64",
          8293 => x"69",
          8294 => x"6c",
          8295 => x"0a",
          8296 => x"53",
          8297 => x"73",
          8298 => x"69",
          8299 => x"70",
          8300 => x"65",
          8301 => x"64",
          8302 => x"44",
          8303 => x"65",
          8304 => x"6d",
          8305 => x"20",
          8306 => x"69",
          8307 => x"6c",
          8308 => x"0a",
          8309 => x"44",
          8310 => x"20",
          8311 => x"20",
          8312 => x"62",
          8313 => x"2e",
          8314 => x"4e",
          8315 => x"6f",
          8316 => x"74",
          8317 => x"65",
          8318 => x"6c",
          8319 => x"73",
          8320 => x"20",
          8321 => x"6e",
          8322 => x"6e",
          8323 => x"73",
          8324 => x"00",
          8325 => x"46",
          8326 => x"61",
          8327 => x"62",
          8328 => x"65",
          8329 => x"00",
          8330 => x"54",
          8331 => x"6f",
          8332 => x"20",
          8333 => x"72",
          8334 => x"6f",
          8335 => x"61",
          8336 => x"6c",
          8337 => x"2e",
          8338 => x"46",
          8339 => x"20",
          8340 => x"6c",
          8341 => x"65",
          8342 => x"00",
          8343 => x"49",
          8344 => x"66",
          8345 => x"69",
          8346 => x"20",
          8347 => x"6f",
          8348 => x"0a",
          8349 => x"54",
          8350 => x"6d",
          8351 => x"20",
          8352 => x"6e",
          8353 => x"6c",
          8354 => x"0a",
          8355 => x"50",
          8356 => x"6d",
          8357 => x"72",
          8358 => x"6e",
          8359 => x"72",
          8360 => x"2e",
          8361 => x"53",
          8362 => x"65",
          8363 => x"0a",
          8364 => x"55",
          8365 => x"6f",
          8366 => x"65",
          8367 => x"72",
          8368 => x"0a",
          8369 => x"20",
          8370 => x"65",
          8371 => x"73",
          8372 => x"20",
          8373 => x"20",
          8374 => x"65",
          8375 => x"65",
          8376 => x"00",
          8377 => x"72",
          8378 => x"00",
          8379 => x"5a",
          8380 => x"41",
          8381 => x"0a",
          8382 => x"25",
          8383 => x"00",
          8384 => x"31",
          8385 => x"37",
          8386 => x"31",
          8387 => x"76",
          8388 => x"00",
          8389 => x"20",
          8390 => x"2c",
          8391 => x"76",
          8392 => x"32",
          8393 => x"25",
          8394 => x"73",
          8395 => x"0a",
          8396 => x"5a",
          8397 => x"41",
          8398 => x"74",
          8399 => x"75",
          8400 => x"48",
          8401 => x"6c",
          8402 => x"00",
          8403 => x"54",
          8404 => x"72",
          8405 => x"74",
          8406 => x"75",
          8407 => x"00",
          8408 => x"50",
          8409 => x"69",
          8410 => x"72",
          8411 => x"74",
          8412 => x"49",
          8413 => x"4c",
          8414 => x"20",
          8415 => x"65",
          8416 => x"70",
          8417 => x"49",
          8418 => x"4c",
          8419 => x"20",
          8420 => x"65",
          8421 => x"70",
          8422 => x"55",
          8423 => x"30",
          8424 => x"20",
          8425 => x"65",
          8426 => x"70",
          8427 => x"55",
          8428 => x"30",
          8429 => x"20",
          8430 => x"65",
          8431 => x"70",
          8432 => x"55",
          8433 => x"31",
          8434 => x"20",
          8435 => x"65",
          8436 => x"70",
          8437 => x"55",
          8438 => x"31",
          8439 => x"20",
          8440 => x"65",
          8441 => x"70",
          8442 => x"53",
          8443 => x"69",
          8444 => x"75",
          8445 => x"69",
          8446 => x"2e",
          8447 => x"00",
          8448 => x"45",
          8449 => x"6c",
          8450 => x"20",
          8451 => x"65",
          8452 => x"2e",
          8453 => x"30",
          8454 => x"46",
          8455 => x"65",
          8456 => x"6f",
          8457 => x"69",
          8458 => x"6c",
          8459 => x"20",
          8460 => x"63",
          8461 => x"20",
          8462 => x"70",
          8463 => x"73",
          8464 => x"6e",
          8465 => x"6d",
          8466 => x"61",
          8467 => x"2e",
          8468 => x"2a",
          8469 => x"42",
          8470 => x"64",
          8471 => x"20",
          8472 => x"0a",
          8473 => x"49",
          8474 => x"69",
          8475 => x"73",
          8476 => x"0a",
          8477 => x"46",
          8478 => x"65",
          8479 => x"6f",
          8480 => x"69",
          8481 => x"6c",
          8482 => x"2e",
          8483 => x"72",
          8484 => x"64",
          8485 => x"25",
          8486 => x"44",
          8487 => x"62",
          8488 => x"67",
          8489 => x"74",
          8490 => x"75",
          8491 => x"0a",
          8492 => x"45",
          8493 => x"6c",
          8494 => x"20",
          8495 => x"65",
          8496 => x"70",
          8497 => x"00",
          8498 => x"44",
          8499 => x"62",
          8500 => x"20",
          8501 => x"74",
          8502 => x"66",
          8503 => x"45",
          8504 => x"6c",
          8505 => x"20",
          8506 => x"74",
          8507 => x"66",
          8508 => x"45",
          8509 => x"75",
          8510 => x"67",
          8511 => x"64",
          8512 => x"20",
          8513 => x"78",
          8514 => x"2e",
          8515 => x"43",
          8516 => x"69",
          8517 => x"63",
          8518 => x"20",
          8519 => x"30",
          8520 => x"2e",
          8521 => x"00",
          8522 => x"43",
          8523 => x"20",
          8524 => x"75",
          8525 => x"64",
          8526 => x"64",
          8527 => x"25",
          8528 => x"0a",
          8529 => x"52",
          8530 => x"61",
          8531 => x"6e",
          8532 => x"70",
          8533 => x"63",
          8534 => x"6f",
          8535 => x"2e",
          8536 => x"43",
          8537 => x"20",
          8538 => x"6f",
          8539 => x"6e",
          8540 => x"2e",
          8541 => x"5a",
          8542 => x"62",
          8543 => x"25",
          8544 => x"25",
          8545 => x"73",
          8546 => x"00",
          8547 => x"42",
          8548 => x"63",
          8549 => x"61",
          8550 => x"0a",
          8551 => x"52",
          8552 => x"69",
          8553 => x"2e",
          8554 => x"45",
          8555 => x"6c",
          8556 => x"20",
          8557 => x"65",
          8558 => x"70",
          8559 => x"2e",
          8560 => x"00",
          8561 => x"00",
          8562 => x"00",
          8563 => x"00",
          8564 => x"00",
          8565 => x"00",
          8566 => x"00",
          8567 => x"00",
          8568 => x"00",
          8569 => x"00",
          8570 => x"00",
          8571 => x"05",
          8572 => x"00",
          8573 => x"01",
          8574 => x"80",
          8575 => x"01",
          8576 => x"00",
          8577 => x"01",
          8578 => x"00",
          8579 => x"00",
          8580 => x"00",
          8581 => x"00",
          8582 => x"00",
          8583 => x"01",
          8584 => x"00",
          8585 => x"00",
          8586 => x"00",
          8587 => x"00",
          8588 => x"00",
          8589 => x"00",
          8590 => x"00",
          8591 => x"01",
          8592 => x"00",
          8593 => x"00",
          8594 => x"00",
          8595 => x"00",
          8596 => x"00",
          8597 => x"00",
          8598 => x"00",
          8599 => x"00",
          8600 => x"00",
          8601 => x"00",
          8602 => x"00",
          8603 => x"00",
          8604 => x"00",
          8605 => x"00",
          8606 => x"00",
          8607 => x"00",
          8608 => x"00",
          8609 => x"00",
          8610 => x"00",
          8611 => x"00",
          8612 => x"00",
          8613 => x"00",
          8614 => x"00",
          8615 => x"00",
          8616 => x"00",
          8617 => x"00",
          8618 => x"00",
          8619 => x"01",
          8620 => x"00",
          8621 => x"00",
          8622 => x"00",
          8623 => x"00",
          8624 => x"00",
          8625 => x"00",
          8626 => x"00",
          8627 => x"00",
          8628 => x"00",
          8629 => x"00",
          8630 => x"00",
          8631 => x"00",
          8632 => x"00",
          8633 => x"00",
          8634 => x"00",
          8635 => x"00",
          8636 => x"00",
          8637 => x"00",
          8638 => x"00",
          8639 => x"00",
          8640 => x"00",
          8641 => x"00",
          8642 => x"00",
          8643 => x"00",
          8644 => x"00",
          8645 => x"00",
          8646 => x"00",
          8647 => x"00",
          8648 => x"00",
          8649 => x"00",
          8650 => x"00",
          8651 => x"00",
          8652 => x"00",
          8653 => x"00",
          8654 => x"00",
          8655 => x"00",
          8656 => x"00",
          8657 => x"00",
          8658 => x"00",
          8659 => x"00",
          8660 => x"00",
          8661 => x"00",
          8662 => x"00",
          8663 => x"00",
          8664 => x"00",
          8665 => x"00",
          8666 => x"00",
          8667 => x"00",
          8668 => x"00",
          8669 => x"00",
          8670 => x"00",
          8671 => x"00",
          8672 => x"00",
          8673 => x"00",
          8674 => x"00",
          8675 => x"00",
          8676 => x"00",
          8677 => x"00",
          8678 => x"00",
          8679 => x"00",
          8680 => x"00",
          8681 => x"00",
          8682 => x"00",
          8683 => x"00",
          8684 => x"00",
          8685 => x"00",
          8686 => x"00",
          8687 => x"00",
          8688 => x"00",
          8689 => x"00",
          8690 => x"00",
          8691 => x"00",
          8692 => x"00",
          8693 => x"00",
          8694 => x"00",
          8695 => x"00",
          8696 => x"00",
          8697 => x"00",
          8698 => x"00",
          8699 => x"01",
          8700 => x"00",
          8701 => x"00",
          8702 => x"00",
          8703 => x"01",
          8704 => x"00",
          8705 => x"00",
          8706 => x"00",
          8707 => x"00",
          8708 => x"00",
          8709 => x"00",
          8710 => x"00",
          8711 => x"00",
          8712 => x"00",
          8713 => x"00",
          8714 => x"00",
          8715 => x"00",
          8716 => x"00",
          8717 => x"00",
          8718 => x"00",
          8719 => x"00",
          8720 => x"00",
          8721 => x"00",
          8722 => x"00",
          8723 => x"00",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"01",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"01",
          8760 => x"00",
          8761 => x"00",
          8762 => x"00",
          8763 => x"00",
          8764 => x"00",
          8765 => x"00",
          8766 => x"00",
          8767 => x"00",
          8768 => x"00",
          8769 => x"00",
          8770 => x"00",
          8771 => x"01",
          8772 => x"00",
          8773 => x"00",
          8774 => x"00",
          8775 => x"01",
          8776 => x"00",
          8777 => x"00",
          8778 => x"00",
          8779 => x"00",
          8780 => x"00",
          8781 => x"00",
          8782 => x"00",
          8783 => x"00",
          8784 => x"00",
          8785 => x"00",
          8786 => x"00",
          8787 => x"01",
          8788 => x"00",
          8789 => x"00",
          8790 => x"00",
          8791 => x"01",
          8792 => x"00",
          8793 => x"00",
          8794 => x"00",
          8795 => x"01",
          8796 => x"00",
          8797 => x"00",
          8798 => x"00",
          8799 => x"01",
          8800 => x"00",
          8801 => x"00",
          8802 => x"00",
          8803 => x"00",
          8804 => x"00",
          8805 => x"00",
          8806 => x"00",
          8807 => x"01",
          8808 => x"00",
          8809 => x"00",
          8810 => x"00",
          8811 => x"00",
          8812 => x"00",
          8813 => x"00",
          8814 => x"00",
          8815 => x"01",
          8816 => x"00",
          8817 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
