-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8a",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"88",
           281 => x"00",
           282 => x"70",
           283 => x"8b",
           284 => x"70",
           285 => x"0c",
           286 => x"88",
           287 => x"99",
           288 => x"02",
           289 => x"3d",
           290 => x"94",
           291 => x"08",
           292 => x"88",
           293 => x"82",
           294 => x"08",
           295 => x"54",
           296 => x"94",
           297 => x"08",
           298 => x"fd",
           299 => x"53",
           300 => x"05",
           301 => x"08",
           302 => x"51",
           303 => x"88",
           304 => x"0c",
           305 => x"0d",
           306 => x"94",
           307 => x"0c",
           308 => x"80",
           309 => x"fc",
           310 => x"08",
           311 => x"80",
           312 => x"94",
           313 => x"08",
           314 => x"88",
           315 => x"0b",
           316 => x"05",
           317 => x"fc",
           318 => x"38",
           319 => x"08",
           320 => x"94",
           321 => x"08",
           322 => x"05",
           323 => x"8c",
           324 => x"25",
           325 => x"08",
           326 => x"30",
           327 => x"05",
           328 => x"94",
           329 => x"0c",
           330 => x"05",
           331 => x"81",
           332 => x"f0",
           333 => x"08",
           334 => x"94",
           335 => x"0c",
           336 => x"08",
           337 => x"52",
           338 => x"05",
           339 => x"a7",
           340 => x"70",
           341 => x"05",
           342 => x"08",
           343 => x"80",
           344 => x"94",
           345 => x"08",
           346 => x"f8",
           347 => x"08",
           348 => x"70",
           349 => x"89",
           350 => x"0c",
           351 => x"02",
           352 => x"3d",
           353 => x"94",
           354 => x"0c",
           355 => x"05",
           356 => x"93",
           357 => x"88",
           358 => x"94",
           359 => x"0c",
           360 => x"08",
           361 => x"94",
           362 => x"08",
           363 => x"38",
           364 => x"05",
           365 => x"08",
           366 => x"81",
           367 => x"8c",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"08",
           372 => x"54",
           373 => x"05",
           374 => x"8c",
           375 => x"f8",
           376 => x"94",
           377 => x"0c",
           378 => x"05",
           379 => x"0c",
           380 => x"0d",
           381 => x"94",
           382 => x"0c",
           383 => x"81",
           384 => x"fc",
           385 => x"0b",
           386 => x"05",
           387 => x"8c",
           388 => x"08",
           389 => x"27",
           390 => x"08",
           391 => x"80",
           392 => x"80",
           393 => x"8c",
           394 => x"99",
           395 => x"8c",
           396 => x"94",
           397 => x"0c",
           398 => x"05",
           399 => x"08",
           400 => x"c9",
           401 => x"fc",
           402 => x"2e",
           403 => x"94",
           404 => x"08",
           405 => x"05",
           406 => x"38",
           407 => x"05",
           408 => x"8c",
           409 => x"94",
           410 => x"0c",
           411 => x"05",
           412 => x"fc",
           413 => x"94",
           414 => x"0c",
           415 => x"05",
           416 => x"94",
           417 => x"0c",
           418 => x"05",
           419 => x"94",
           420 => x"0c",
           421 => x"94",
           422 => x"08",
           423 => x"38",
           424 => x"05",
           425 => x"08",
           426 => x"51",
           427 => x"08",
           428 => x"70",
           429 => x"05",
           430 => x"08",
           431 => x"88",
           432 => x"0d",
           433 => x"ff",
           434 => x"88",
           435 => x"92",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"8c",
           441 => x"06",
           442 => x"80",
           443 => x"87",
           444 => x"08",
           445 => x"38",
           446 => x"8c",
           447 => x"80",
           448 => x"93",
           449 => x"98",
           450 => x"70",
           451 => x"38",
           452 => x"0b",
           453 => x"0b",
           454 => x"a8",
           455 => x"83",
           456 => x"fa",
           457 => x"7b",
           458 => x"56",
           459 => x"0b",
           460 => x"33",
           461 => x"55",
           462 => x"75",
           463 => x"06",
           464 => x"85",
           465 => x"98",
           466 => x"87",
           467 => x"0c",
           468 => x"c0",
           469 => x"87",
           470 => x"08",
           471 => x"70",
           472 => x"52",
           473 => x"2e",
           474 => x"c0",
           475 => x"70",
           476 => x"76",
           477 => x"53",
           478 => x"2e",
           479 => x"80",
           480 => x"71",
           481 => x"05",
           482 => x"14",
           483 => x"55",
           484 => x"51",
           485 => x"8b",
           486 => x"98",
           487 => x"70",
           488 => x"87",
           489 => x"08",
           490 => x"38",
           491 => x"c0",
           492 => x"87",
           493 => x"08",
           494 => x"51",
           495 => x"38",
           496 => x"80",
           497 => x"52",
           498 => x"09",
           499 => x"38",
           500 => x"8c",
           501 => x"72",
           502 => x"06",
           503 => x"52",
           504 => x"88",
           505 => x"fe",
           506 => x"81",
           507 => x"33",
           508 => x"07",
           509 => x"51",
           510 => x"04",
           511 => x"75",
           512 => x"82",
           513 => x"90",
           514 => x"2b",
           515 => x"33",
           516 => x"88",
           517 => x"71",
           518 => x"52",
           519 => x"54",
           520 => x"0d",
           521 => x"0d",
           522 => x"0b",
           523 => x"57",
           524 => x"27",
           525 => x"76",
           526 => x"27",
           527 => x"75",
           528 => x"82",
           529 => x"74",
           530 => x"38",
           531 => x"74",
           532 => x"83",
           533 => x"76",
           534 => x"17",
           535 => x"88",
           536 => x"55",
           537 => x"88",
           538 => x"74",
           539 => x"3f",
           540 => x"ff",
           541 => x"ad",
           542 => x"76",
           543 => x"fc",
           544 => x"87",
           545 => x"08",
           546 => x"3d",
           547 => x"fd",
           548 => x"08",
           549 => x"51",
           550 => x"88",
           551 => x"06",
           552 => x"81",
           553 => x"0c",
           554 => x"04",
           555 => x"0b",
           556 => x"ac",
           557 => x"88",
           558 => x"05",
           559 => x"80",
           560 => x"27",
           561 => x"14",
           562 => x"29",
           563 => x"05",
           564 => x"88",
           565 => x"0d",
           566 => x"0d",
           567 => x"0b",
           568 => x"9f",
           569 => x"33",
           570 => x"71",
           571 => x"81",
           572 => x"94",
           573 => x"ef",
           574 => x"90",
           575 => x"14",
           576 => x"3f",
           577 => x"ff",
           578 => x"07",
           579 => x"3d",
           580 => x"3d",
           581 => x"0b",
           582 => x"08",
           583 => x"75",
           584 => x"08",
           585 => x"2e",
           586 => x"14",
           587 => x"85",
           588 => x"b0",
           589 => x"38",
           590 => x"71",
           591 => x"81",
           592 => x"90",
           593 => x"72",
           594 => x"72",
           595 => x"38",
           596 => x"d8",
           597 => x"52",
           598 => x"14",
           599 => x"90",
           600 => x"52",
           601 => x"86",
           602 => x"fa",
           603 => x"0b",
           604 => x"ac",
           605 => x"81",
           606 => x"ff",
           607 => x"54",
           608 => x"80",
           609 => x"90",
           610 => x"72",
           611 => x"52",
           612 => x"73",
           613 => x"71",
           614 => x"81",
           615 => x"0c",
           616 => x"53",
           617 => x"83",
           618 => x"22",
           619 => x"76",
           620 => x"b5",
           621 => x"33",
           622 => x"84",
           623 => x"71",
           624 => x"51",
           625 => x"81",
           626 => x"08",
           627 => x"83",
           628 => x"88",
           629 => x"96",
           630 => x"8c",
           631 => x"08",
           632 => x"3f",
           633 => x"16",
           634 => x"23",
           635 => x"88",
           636 => x"0d",
           637 => x"0d",
           638 => x"58",
           639 => x"33",
           640 => x"2e",
           641 => x"88",
           642 => x"70",
           643 => x"39",
           644 => x"56",
           645 => x"2e",
           646 => x"84",
           647 => x"43",
           648 => x"1d",
           649 => x"33",
           650 => x"9f",
           651 => x"7b",
           652 => x"3f",
           653 => x"80",
           654 => x"d3",
           655 => x"84",
           656 => x"58",
           657 => x"55",
           658 => x"81",
           659 => x"ff",
           660 => x"ff",
           661 => x"06",
           662 => x"70",
           663 => x"7f",
           664 => x"7a",
           665 => x"81",
           666 => x"13",
           667 => x"af",
           668 => x"a0",
           669 => x"80",
           670 => x"51",
           671 => x"5d",
           672 => x"80",
           673 => x"ae",
           674 => x"06",
           675 => x"55",
           676 => x"75",
           677 => x"80",
           678 => x"79",
           679 => x"30",
           680 => x"70",
           681 => x"07",
           682 => x"51",
           683 => x"75",
           684 => x"58",
           685 => x"ab",
           686 => x"19",
           687 => x"06",
           688 => x"5a",
           689 => x"75",
           690 => x"39",
           691 => x"0c",
           692 => x"a0",
           693 => x"81",
           694 => x"1a",
           695 => x"fc",
           696 => x"08",
           697 => x"a0",
           698 => x"70",
           699 => x"e0",
           700 => x"90",
           701 => x"7c",
           702 => x"3f",
           703 => x"88",
           704 => x"38",
           705 => x"74",
           706 => x"ee",
           707 => x"33",
           708 => x"70",
           709 => x"56",
           710 => x"38",
           711 => x"1e",
           712 => x"59",
           713 => x"ff",
           714 => x"ff",
           715 => x"79",
           716 => x"5b",
           717 => x"81",
           718 => x"71",
           719 => x"56",
           720 => x"2e",
           721 => x"39",
           722 => x"92",
           723 => x"fc",
           724 => x"8e",
           725 => x"56",
           726 => x"38",
           727 => x"56",
           728 => x"8b",
           729 => x"55",
           730 => x"8b",
           731 => x"84",
           732 => x"06",
           733 => x"74",
           734 => x"56",
           735 => x"56",
           736 => x"51",
           737 => x"88",
           738 => x"0c",
           739 => x"75",
           740 => x"3d",
           741 => x"3d",
           742 => x"59",
           743 => x"83",
           744 => x"52",
           745 => x"fb",
           746 => x"88",
           747 => x"38",
           748 => x"b3",
           749 => x"83",
           750 => x"55",
           751 => x"82",
           752 => x"09",
           753 => x"ce",
           754 => x"b6",
           755 => x"76",
           756 => x"3f",
           757 => x"88",
           758 => x"76",
           759 => x"3f",
           760 => x"ff",
           761 => x"74",
           762 => x"2e",
           763 => x"54",
           764 => x"77",
           765 => x"f6",
           766 => x"08",
           767 => x"94",
           768 => x"f7",
           769 => x"08",
           770 => x"06",
           771 => x"82",
           772 => x"38",
           773 => x"88",
           774 => x"0d",
           775 => x"0d",
           776 => x"0b",
           777 => x"9f",
           778 => x"9b",
           779 => x"81",
           780 => x"56",
           781 => x"38",
           782 => x"8d",
           783 => x"57",
           784 => x"3f",
           785 => x"ff",
           786 => x"81",
           787 => x"06",
           788 => x"54",
           789 => x"74",
           790 => x"f5",
           791 => x"08",
           792 => x"3d",
           793 => x"80",
           794 => x"95",
           795 => x"51",
           796 => x"88",
           797 => x"53",
           798 => x"fe",
           799 => x"08",
           800 => x"57",
           801 => x"09",
           802 => x"38",
           803 => x"99",
           804 => x"2e",
           805 => x"56",
           806 => x"a4",
           807 => x"79",
           808 => x"f4",
           809 => x"56",
           810 => x"fd",
           811 => x"e5",
           812 => x"b3",
           813 => x"83",
           814 => x"58",
           815 => x"95",
           816 => x"51",
           817 => x"88",
           818 => x"af",
           819 => x"71",
           820 => x"05",
           821 => x"54",
           822 => x"f6",
           823 => x"08",
           824 => x"06",
           825 => x"1a",
           826 => x"33",
           827 => x"95",
           828 => x"51",
           829 => x"88",
           830 => x"23",
           831 => x"05",
           832 => x"3f",
           833 => x"ff",
           834 => x"75",
           835 => x"3d",
           836 => x"f5",
           837 => x"08",
           838 => x"f5",
           839 => x"08",
           840 => x"06",
           841 => x"79",
           842 => x"22",
           843 => x"82",
           844 => x"72",
           845 => x"59",
           846 => x"ee",
           847 => x"08",
           848 => x"88",
           849 => x"08",
           850 => x"56",
           851 => x"df",
           852 => x"38",
           853 => x"ff",
           854 => x"85",
           855 => x"89",
           856 => x"76",
           857 => x"c1",
           858 => x"34",
           859 => x"09",
           860 => x"38",
           861 => x"05",
           862 => x"3f",
           863 => x"1a",
           864 => x"8c",
           865 => x"90",
           866 => x"83",
           867 => x"8c",
           868 => x"71",
           869 => x"94",
           870 => x"80",
           871 => x"34",
           872 => x"0b",
           873 => x"80",
           874 => x"0c",
           875 => x"04",
           876 => x"0b",
           877 => x"ac",
           878 => x"54",
           879 => x"80",
           880 => x"0b",
           881 => x"98",
           882 => x"45",
           883 => x"3d",
           884 => x"ec",
           885 => x"9d",
           886 => x"54",
           887 => x"c0",
           888 => x"33",
           889 => x"2e",
           890 => x"a7",
           891 => x"84",
           892 => x"06",
           893 => x"73",
           894 => x"38",
           895 => x"39",
           896 => x"d5",
           897 => x"a0",
           898 => x"3d",
           899 => x"f3",
           900 => x"08",
           901 => x"73",
           902 => x"81",
           903 => x"34",
           904 => x"98",
           905 => x"f6",
           906 => x"7f",
           907 => x"0b",
           908 => x"59",
           909 => x"80",
           910 => x"57",
           911 => x"81",
           912 => x"16",
           913 => x"55",
           914 => x"80",
           915 => x"38",
           916 => x"81",
           917 => x"39",
           918 => x"17",
           919 => x"81",
           920 => x"16",
           921 => x"08",
           922 => x"78",
           923 => x"74",
           924 => x"2e",
           925 => x"98",
           926 => x"83",
           927 => x"57",
           928 => x"38",
           929 => x"ff",
           930 => x"2a",
           931 => x"ff",
           932 => x"79",
           933 => x"87",
           934 => x"08",
           935 => x"a4",
           936 => x"f3",
           937 => x"08",
           938 => x"27",
           939 => x"74",
           940 => x"a4",
           941 => x"f3",
           942 => x"08",
           943 => x"80",
           944 => x"38",
           945 => x"a8",
           946 => x"16",
           947 => x"06",
           948 => x"31",
           949 => x"75",
           950 => x"77",
           951 => x"98",
           952 => x"ff",
           953 => x"16",
           954 => x"51",
           955 => x"88",
           956 => x"38",
           957 => x"15",
           958 => x"77",
           959 => x"08",
           960 => x"58",
           961 => x"fe",
           962 => x"19",
           963 => x"39",
           964 => x"88",
           965 => x"0d",
           966 => x"0d",
           967 => x"e4",
           968 => x"94",
           969 => x"90",
           970 => x"87",
           971 => x"0c",
           972 => x"0b",
           973 => x"84",
           974 => x"83",
           975 => x"94",
           976 => x"b0",
           977 => x"3f",
           978 => x"38",
           979 => x"fc",
           980 => x"08",
           981 => x"80",
           982 => x"87",
           983 => x"0c",
           984 => x"fc",
           985 => x"80",
           986 => x"fd",
           987 => x"08",
           988 => x"54",
           989 => x"86",
           990 => x"55",
           991 => x"80",
           992 => x"80",
           993 => x"00",
           994 => x"ff",
           995 => x"ff",
           996 => x"ff",
           997 => x"00",
           998 => x"54",
           999 => x"59",
          1000 => x"4d",
          1001 => x"00",
          1002 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"00",
           281 => x"00",
           282 => x"ac",
           283 => x"27",
           284 => x"71",
           285 => x"53",
           286 => x"04",
           287 => x"9e",
           288 => x"08",
           289 => x"fd",
           290 => x"53",
           291 => x"05",
           292 => x"08",
           293 => x"51",
           294 => x"88",
           295 => x"0c",
           296 => x"0d",
           297 => x"94",
           298 => x"0c",
           299 => x"81",
           300 => x"8c",
           301 => x"94",
           302 => x"08",
           303 => x"3f",
           304 => x"88",
           305 => x"3d",
           306 => x"04",
           307 => x"94",
           308 => x"0d",
           309 => x"08",
           310 => x"94",
           311 => x"08",
           312 => x"38",
           313 => x"05",
           314 => x"08",
           315 => x"80",
           316 => x"f4",
           317 => x"08",
           318 => x"88",
           319 => x"94",
           320 => x"0c",
           321 => x"05",
           322 => x"fc",
           323 => x"08",
           324 => x"80",
           325 => x"94",
           326 => x"08",
           327 => x"8c",
           328 => x"0b",
           329 => x"05",
           330 => x"fc",
           331 => x"38",
           332 => x"08",
           333 => x"94",
           334 => x"08",
           335 => x"05",
           336 => x"94",
           337 => x"08",
           338 => x"88",
           339 => x"81",
           340 => x"08",
           341 => x"f8",
           342 => x"94",
           343 => x"08",
           344 => x"38",
           345 => x"05",
           346 => x"08",
           347 => x"94",
           348 => x"08",
           349 => x"54",
           350 => x"94",
           351 => x"08",
           352 => x"fb",
           353 => x"0b",
           354 => x"05",
           355 => x"88",
           356 => x"25",
           357 => x"08",
           358 => x"30",
           359 => x"05",
           360 => x"94",
           361 => x"0c",
           362 => x"05",
           363 => x"8c",
           364 => x"8c",
           365 => x"94",
           366 => x"0c",
           367 => x"08",
           368 => x"52",
           369 => x"05",
           370 => x"3f",
           371 => x"94",
           372 => x"0c",
           373 => x"fc",
           374 => x"2e",
           375 => x"08",
           376 => x"30",
           377 => x"05",
           378 => x"f8",
           379 => x"88",
           380 => x"3d",
           381 => x"04",
           382 => x"94",
           383 => x"0d",
           384 => x"08",
           385 => x"80",
           386 => x"f8",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"94",
           391 => x"08",
           392 => x"38",
           393 => x"08",
           394 => x"24",
           395 => x"08",
           396 => x"10",
           397 => x"05",
           398 => x"fc",
           399 => x"94",
           400 => x"0c",
           401 => x"08",
           402 => x"80",
           403 => x"38",
           404 => x"05",
           405 => x"88",
           406 => x"a1",
           407 => x"88",
           408 => x"08",
           409 => x"31",
           410 => x"05",
           411 => x"f8",
           412 => x"08",
           413 => x"07",
           414 => x"05",
           415 => x"fc",
           416 => x"2a",
           417 => x"05",
           418 => x"8c",
           419 => x"2a",
           420 => x"05",
           421 => x"39",
           422 => x"05",
           423 => x"8f",
           424 => x"88",
           425 => x"94",
           426 => x"0c",
           427 => x"94",
           428 => x"08",
           429 => x"f4",
           430 => x"94",
           431 => x"08",
           432 => x"3d",
           433 => x"04",
           434 => x"81",
           435 => x"c0",
           436 => x"81",
           437 => x"92",
           438 => x"0b",
           439 => x"8c",
           440 => x"92",
           441 => x"82",
           442 => x"70",
           443 => x"38",
           444 => x"8c",
           445 => x"e9",
           446 => x"92",
           447 => x"80",
           448 => x"71",
           449 => x"c0",
           450 => x"51",
           451 => x"88",
           452 => x"0b",
           453 => x"34",
           454 => x"9f",
           455 => x"0c",
           456 => x"04",
           457 => x"78",
           458 => x"58",
           459 => x"0b",
           460 => x"a8",
           461 => x"52",
           462 => x"70",
           463 => x"81",
           464 => x"38",
           465 => x"c0",
           466 => x"79",
           467 => x"80",
           468 => x"87",
           469 => x"0c",
           470 => x"8c",
           471 => x"2a",
           472 => x"51",
           473 => x"80",
           474 => x"87",
           475 => x"08",
           476 => x"06",
           477 => x"52",
           478 => x"80",
           479 => x"70",
           480 => x"38",
           481 => x"81",
           482 => x"ff",
           483 => x"15",
           484 => x"06",
           485 => x"2e",
           486 => x"c0",
           487 => x"51",
           488 => x"38",
           489 => x"8c",
           490 => x"95",
           491 => x"87",
           492 => x"0c",
           493 => x"8c",
           494 => x"06",
           495 => x"f4",
           496 => x"fc",
           497 => x"52",
           498 => x"2e",
           499 => x"8f",
           500 => x"98",
           501 => x"70",
           502 => x"81",
           503 => x"81",
           504 => x"0c",
           505 => x"04",
           506 => x"74",
           507 => x"71",
           508 => x"2b",
           509 => x"53",
           510 => x"0d",
           511 => x"0d",
           512 => x"33",
           513 => x"71",
           514 => x"88",
           515 => x"14",
           516 => x"07",
           517 => x"33",
           518 => x"0c",
           519 => x"56",
           520 => x"3d",
           521 => x"3d",
           522 => x"0b",
           523 => x"08",
           524 => x"77",
           525 => x"38",
           526 => x"08",
           527 => x"38",
           528 => x"74",
           529 => x"38",
           530 => x"ae",
           531 => x"39",
           532 => x"10",
           533 => x"53",
           534 => x"8c",
           535 => x"52",
           536 => x"52",
           537 => x"3f",
           538 => x"38",
           539 => x"f8",
           540 => x"83",
           541 => x"55",
           542 => x"54",
           543 => x"83",
           544 => x"76",
           545 => x"17",
           546 => x"88",
           547 => x"55",
           548 => x"88",
           549 => x"74",
           550 => x"3f",
           551 => x"0a",
           552 => x"39",
           553 => x"88",
           554 => x"0d",
           555 => x"0d",
           556 => x"9f",
           557 => x"19",
           558 => x"fe",
           559 => x"54",
           560 => x"73",
           561 => x"82",
           562 => x"71",
           563 => x"08",
           564 => x"75",
           565 => x"3d",
           566 => x"3d",
           567 => x"80",
           568 => x"0b",
           569 => x"70",
           570 => x"53",
           571 => x"09",
           572 => x"38",
           573 => x"fd",
           574 => x"08",
           575 => x"9a",
           576 => x"e4",
           577 => x"83",
           578 => x"73",
           579 => x"85",
           580 => x"fc",
           581 => x"0b",
           582 => x"ac",
           583 => x"80",
           584 => x"15",
           585 => x"81",
           586 => x"88",
           587 => x"26",
           588 => x"52",
           589 => x"90",
           590 => x"52",
           591 => x"09",
           592 => x"38",
           593 => x"53",
           594 => x"0c",
           595 => x"8b",
           596 => x"fe",
           597 => x"08",
           598 => x"90",
           599 => x"71",
           600 => x"80",
           601 => x"0c",
           602 => x"04",
           603 => x"78",
           604 => x"9f",
           605 => x"22",
           606 => x"83",
           607 => x"57",
           608 => x"73",
           609 => x"38",
           610 => x"53",
           611 => x"83",
           612 => x"39",
           613 => x"52",
           614 => x"38",
           615 => x"16",
           616 => x"08",
           617 => x"38",
           618 => x"17",
           619 => x"73",
           620 => x"38",
           621 => x"16",
           622 => x"74",
           623 => x"52",
           624 => x"72",
           625 => x"3f",
           626 => x"88",
           627 => x"38",
           628 => x"08",
           629 => x"27",
           630 => x"08",
           631 => x"88",
           632 => x"c9",
           633 => x"90",
           634 => x"75",
           635 => x"71",
           636 => x"3d",
           637 => x"3d",
           638 => x"64",
           639 => x"75",
           640 => x"a0",
           641 => x"06",
           642 => x"16",
           643 => x"ef",
           644 => x"33",
           645 => x"af",
           646 => x"06",
           647 => x"16",
           648 => x"88",
           649 => x"70",
           650 => x"74",
           651 => x"38",
           652 => x"df",
           653 => x"56",
           654 => x"82",
           655 => x"3d",
           656 => x"70",
           657 => x"8a",
           658 => x"70",
           659 => x"34",
           660 => x"74",
           661 => x"81",
           662 => x"80",
           663 => x"88",
           664 => x"5a",
           665 => x"70",
           666 => x"60",
           667 => x"70",
           668 => x"30",
           669 => x"71",
           670 => x"51",
           671 => x"53",
           672 => x"74",
           673 => x"76",
           674 => x"81",
           675 => x"81",
           676 => x"27",
           677 => x"74",
           678 => x"38",
           679 => x"70",
           680 => x"32",
           681 => x"73",
           682 => x"53",
           683 => x"56",
           684 => x"88",
           685 => x"ff",
           686 => x"81",
           687 => x"ff",
           688 => x"53",
           689 => x"76",
           690 => x"98",
           691 => x"7f",
           692 => x"76",
           693 => x"38",
           694 => x"8b",
           695 => x"51",
           696 => x"88",
           697 => x"38",
           698 => x"22",
           699 => x"83",
           700 => x"55",
           701 => x"52",
           702 => x"a8",
           703 => x"57",
           704 => x"fb",
           705 => x"55",
           706 => x"80",
           707 => x"1d",
           708 => x"2a",
           709 => x"51",
           710 => x"b2",
           711 => x"84",
           712 => x"08",
           713 => x"58",
           714 => x"77",
           715 => x"38",
           716 => x"05",
           717 => x"70",
           718 => x"33",
           719 => x"52",
           720 => x"80",
           721 => x"86",
           722 => x"2e",
           723 => x"51",
           724 => x"ff",
           725 => x"08",
           726 => x"b4",
           727 => x"76",
           728 => x"08",
           729 => x"51",
           730 => x"38",
           731 => x"70",
           732 => x"81",
           733 => x"56",
           734 => x"83",
           735 => x"81",
           736 => x"7c",
           737 => x"3f",
           738 => x"1d",
           739 => x"39",
           740 => x"90",
           741 => x"f9",
           742 => x"7b",
           743 => x"54",
           744 => x"77",
           745 => x"f6",
           746 => x"56",
           747 => x"e7",
           748 => x"f8",
           749 => x"08",
           750 => x"06",
           751 => x"74",
           752 => x"2e",
           753 => x"80",
           754 => x"54",
           755 => x"52",
           756 => x"d0",
           757 => x"56",
           758 => x"38",
           759 => x"88",
           760 => x"83",
           761 => x"55",
           762 => x"c6",
           763 => x"82",
           764 => x"53",
           765 => x"51",
           766 => x"88",
           767 => x"08",
           768 => x"51",
           769 => x"88",
           770 => x"ff",
           771 => x"81",
           772 => x"83",
           773 => x"75",
           774 => x"3d",
           775 => x"3d",
           776 => x"80",
           777 => x"0b",
           778 => x"f5",
           779 => x"08",
           780 => x"82",
           781 => x"f2",
           782 => x"53",
           783 => x"53",
           784 => x"d3",
           785 => x"81",
           786 => x"76",
           787 => x"81",
           788 => x"90",
           789 => x"53",
           790 => x"51",
           791 => x"88",
           792 => x"8d",
           793 => x"74",
           794 => x"38",
           795 => x"05",
           796 => x"3f",
           797 => x"08",
           798 => x"5a",
           799 => x"88",
           800 => x"06",
           801 => x"2e",
           802 => x"86",
           803 => x"82",
           804 => x"80",
           805 => x"86",
           806 => x"39",
           807 => x"53",
           808 => x"51",
           809 => x"81",
           810 => x"81",
           811 => x"3d",
           812 => x"f6",
           813 => x"08",
           814 => x"06",
           815 => x"38",
           816 => x"05",
           817 => x"3f",
           818 => x"02",
           819 => x"78",
           820 => x"88",
           821 => x"70",
           822 => x"5b",
           823 => x"88",
           824 => x"ff",
           825 => x"8c",
           826 => x"3d",
           827 => x"34",
           828 => x"05",
           829 => x"3f",
           830 => x"1a",
           831 => x"e2",
           832 => x"e4",
           833 => x"83",
           834 => x"56",
           835 => x"95",
           836 => x"51",
           837 => x"88",
           838 => x"51",
           839 => x"88",
           840 => x"ff",
           841 => x"31",
           842 => x"1b",
           843 => x"2a",
           844 => x"56",
           845 => x"55",
           846 => x"55",
           847 => x"88",
           848 => x"70",
           849 => x"88",
           850 => x"05",
           851 => x"83",
           852 => x"83",
           853 => x"83",
           854 => x"27",
           855 => x"57",
           856 => x"56",
           857 => x"80",
           858 => x"79",
           859 => x"2e",
           860 => x"90",
           861 => x"fb",
           862 => x"81",
           863 => x"90",
           864 => x"39",
           865 => x"18",
           866 => x"79",
           867 => x"06",
           868 => x"19",
           869 => x"05",
           870 => x"55",
           871 => x"1a",
           872 => x"0b",
           873 => x"0c",
           874 => x"88",
           875 => x"0d",
           876 => x"0d",
           877 => x"9f",
           878 => x"85",
           879 => x"2e",
           880 => x"80",
           881 => x"34",
           882 => x"11",
           883 => x"89",
           884 => x"57",
           885 => x"f8",
           886 => x"08",
           887 => x"80",
           888 => x"3d",
           889 => x"80",
           890 => x"02",
           891 => x"70",
           892 => x"81",
           893 => x"57",
           894 => x"85",
           895 => x"a1",
           896 => x"f5",
           897 => x"08",
           898 => x"98",
           899 => x"51",
           900 => x"88",
           901 => x"0c",
           902 => x"0c",
           903 => x"16",
           904 => x"0c",
           905 => x"04",
           906 => x"7d",
           907 => x"0b",
           908 => x"08",
           909 => x"58",
           910 => x"85",
           911 => x"2e",
           912 => x"81",
           913 => x"06",
           914 => x"74",
           915 => x"c3",
           916 => x"74",
           917 => x"86",
           918 => x"81",
           919 => x"57",
           920 => x"9c",
           921 => x"17",
           922 => x"74",
           923 => x"38",
           924 => x"80",
           925 => x"38",
           926 => x"70",
           927 => x"56",
           928 => x"c7",
           929 => x"33",
           930 => x"89",
           931 => x"81",
           932 => x"55",
           933 => x"76",
           934 => x"16",
           935 => x"39",
           936 => x"51",
           937 => x"88",
           938 => x"75",
           939 => x"38",
           940 => x"0c",
           941 => x"51",
           942 => x"88",
           943 => x"08",
           944 => x"8f",
           945 => x"1a",
           946 => x"98",
           947 => x"ff",
           948 => x"71",
           949 => x"77",
           950 => x"38",
           951 => x"54",
           952 => x"83",
           953 => x"a8",
           954 => x"78",
           955 => x"3f",
           956 => x"e5",
           957 => x"08",
           958 => x"0c",
           959 => x"7b",
           960 => x"0c",
           961 => x"2e",
           962 => x"74",
           963 => x"e2",
           964 => x"76",
           965 => x"3d",
           966 => x"3d",
           967 => x"86",
           968 => x"c0",
           969 => x"9b",
           970 => x"0b",
           971 => x"9c",
           972 => x"83",
           973 => x"94",
           974 => x"80",
           975 => x"c0",
           976 => x"9f",
           977 => x"d6",
           978 => x"b8",
           979 => x"51",
           980 => x"88",
           981 => x"a0",
           982 => x"08",
           983 => x"88",
           984 => x"3d",
           985 => x"84",
           986 => x"51",
           987 => x"88",
           988 => x"75",
           989 => x"2e",
           990 => x"15",
           991 => x"a0",
           992 => x"04",
           993 => x"39",
           994 => x"ff",
           995 => x"ff",
           996 => x"00",
           997 => x"ff",
           998 => x"4f",
           999 => x"4e",
          1000 => x"4f",
          1001 => x"00",
          1002 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"04",
           281 => x"04",
           282 => x"9f",
           283 => x"dc",
           284 => x"80",
           285 => x"05",
           286 => x"eb",
           287 => x"51",
           288 => x"94",
           289 => x"0c",
           290 => x"80",
           291 => x"8c",
           292 => x"94",
           293 => x"08",
           294 => x"3f",
           295 => x"88",
           296 => x"3d",
           297 => x"04",
           298 => x"94",
           299 => x"0d",
           300 => x"08",
           301 => x"52",
           302 => x"05",
           303 => x"b9",
           304 => x"70",
           305 => x"85",
           306 => x"0c",
           307 => x"02",
           308 => x"3d",
           309 => x"94",
           310 => x"0c",
           311 => x"05",
           312 => x"ab",
           313 => x"88",
           314 => x"94",
           315 => x"0c",
           316 => x"08",
           317 => x"94",
           318 => x"08",
           319 => x"0b",
           320 => x"05",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"08",
           325 => x"38",
           326 => x"05",
           327 => x"08",
           328 => x"80",
           329 => x"f0",
           330 => x"08",
           331 => x"88",
           332 => x"94",
           333 => x"0c",
           334 => x"05",
           335 => x"fc",
           336 => x"53",
           337 => x"05",
           338 => x"08",
           339 => x"51",
           340 => x"88",
           341 => x"08",
           342 => x"54",
           343 => x"05",
           344 => x"8c",
           345 => x"f8",
           346 => x"94",
           347 => x"0c",
           348 => x"05",
           349 => x"0c",
           350 => x"0d",
           351 => x"94",
           352 => x"0c",
           353 => x"80",
           354 => x"fc",
           355 => x"08",
           356 => x"80",
           357 => x"94",
           358 => x"08",
           359 => x"88",
           360 => x"0b",
           361 => x"05",
           362 => x"8c",
           363 => x"25",
           364 => x"08",
           365 => x"30",
           366 => x"05",
           367 => x"94",
           368 => x"08",
           369 => x"88",
           370 => x"ad",
           371 => x"70",
           372 => x"05",
           373 => x"08",
           374 => x"80",
           375 => x"94",
           376 => x"08",
           377 => x"f8",
           378 => x"08",
           379 => x"70",
           380 => x"87",
           381 => x"0c",
           382 => x"02",
           383 => x"3d",
           384 => x"94",
           385 => x"0c",
           386 => x"08",
           387 => x"94",
           388 => x"08",
           389 => x"05",
           390 => x"38",
           391 => x"05",
           392 => x"a3",
           393 => x"94",
           394 => x"08",
           395 => x"94",
           396 => x"08",
           397 => x"8c",
           398 => x"08",
           399 => x"10",
           400 => x"05",
           401 => x"94",
           402 => x"08",
           403 => x"c9",
           404 => x"8c",
           405 => x"08",
           406 => x"26",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"88",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"f8",
           415 => x"08",
           416 => x"81",
           417 => x"fc",
           418 => x"08",
           419 => x"81",
           420 => x"8c",
           421 => x"af",
           422 => x"90",
           423 => x"2e",
           424 => x"08",
           425 => x"70",
           426 => x"05",
           427 => x"39",
           428 => x"05",
           429 => x"08",
           430 => x"51",
           431 => x"05",
           432 => x"85",
           433 => x"0c",
           434 => x"0d",
           435 => x"87",
           436 => x"0c",
           437 => x"c0",
           438 => x"85",
           439 => x"98",
           440 => x"c0",
           441 => x"70",
           442 => x"51",
           443 => x"8a",
           444 => x"98",
           445 => x"70",
           446 => x"c0",
           447 => x"fc",
           448 => x"52",
           449 => x"87",
           450 => x"08",
           451 => x"2e",
           452 => x"0b",
           453 => x"a8",
           454 => x"0b",
           455 => x"88",
           456 => x"0d",
           457 => x"0d",
           458 => x"56",
           459 => x"0b",
           460 => x"9f",
           461 => x"06",
           462 => x"52",
           463 => x"09",
           464 => x"9e",
           465 => x"87",
           466 => x"0c",
           467 => x"92",
           468 => x"0b",
           469 => x"8c",
           470 => x"92",
           471 => x"85",
           472 => x"06",
           473 => x"70",
           474 => x"38",
           475 => x"84",
           476 => x"ff",
           477 => x"27",
           478 => x"73",
           479 => x"38",
           480 => x"8b",
           481 => x"70",
           482 => x"34",
           483 => x"81",
           484 => x"a2",
           485 => x"80",
           486 => x"87",
           487 => x"08",
           488 => x"b5",
           489 => x"98",
           490 => x"70",
           491 => x"0b",
           492 => x"8c",
           493 => x"92",
           494 => x"82",
           495 => x"70",
           496 => x"73",
           497 => x"06",
           498 => x"72",
           499 => x"06",
           500 => x"c0",
           501 => x"51",
           502 => x"09",
           503 => x"38",
           504 => x"88",
           505 => x"0d",
           506 => x"0d",
           507 => x"33",
           508 => x"88",
           509 => x"0c",
           510 => x"3d",
           511 => x"3d",
           512 => x"11",
           513 => x"33",
           514 => x"71",
           515 => x"81",
           516 => x"72",
           517 => x"75",
           518 => x"88",
           519 => x"54",
           520 => x"85",
           521 => x"f9",
           522 => x"0b",
           523 => x"ac",
           524 => x"81",
           525 => x"ed",
           526 => x"17",
           527 => x"e5",
           528 => x"55",
           529 => x"89",
           530 => x"2e",
           531 => x"d5",
           532 => x"76",
           533 => x"06",
           534 => x"2a",
           535 => x"05",
           536 => x"70",
           537 => x"bd",
           538 => x"b9",
           539 => x"fe",
           540 => x"08",
           541 => x"06",
           542 => x"84",
           543 => x"2b",
           544 => x"53",
           545 => x"8c",
           546 => x"52",
           547 => x"52",
           548 => x"3f",
           549 => x"38",
           550 => x"e2",
           551 => x"f0",
           552 => x"83",
           553 => x"74",
           554 => x"3d",
           555 => x"3d",
           556 => x"0b",
           557 => x"fe",
           558 => x"08",
           559 => x"56",
           560 => x"74",
           561 => x"38",
           562 => x"75",
           563 => x"16",
           564 => x"53",
           565 => x"87",
           566 => x"fd",
           567 => x"54",
           568 => x"0b",
           569 => x"08",
           570 => x"53",
           571 => x"2e",
           572 => x"8c",
           573 => x"51",
           574 => x"88",
           575 => x"53",
           576 => x"fd",
           577 => x"08",
           578 => x"06",
           579 => x"0c",
           580 => x"04",
           581 => x"76",
           582 => x"9f",
           583 => x"55",
           584 => x"88",
           585 => x"72",
           586 => x"38",
           587 => x"73",
           588 => x"81",
           589 => x"72",
           590 => x"33",
           591 => x"2e",
           592 => x"85",
           593 => x"08",
           594 => x"16",
           595 => x"2e",
           596 => x"51",
           597 => x"88",
           598 => x"39",
           599 => x"52",
           600 => x"0c",
           601 => x"88",
           602 => x"0d",
           603 => x"0d",
           604 => x"0b",
           605 => x"71",
           606 => x"70",
           607 => x"06",
           608 => x"55",
           609 => x"88",
           610 => x"08",
           611 => x"38",
           612 => x"dc",
           613 => x"06",
           614 => x"cf",
           615 => x"90",
           616 => x"15",
           617 => x"8f",
           618 => x"84",
           619 => x"52",
           620 => x"bc",
           621 => x"82",
           622 => x"05",
           623 => x"06",
           624 => x"38",
           625 => x"df",
           626 => x"71",
           627 => x"a0",
           628 => x"88",
           629 => x"08",
           630 => x"88",
           631 => x"0c",
           632 => x"fd",
           633 => x"08",
           634 => x"73",
           635 => x"52",
           636 => x"88",
           637 => x"f2",
           638 => x"62",
           639 => x"5c",
           640 => x"74",
           641 => x"81",
           642 => x"81",
           643 => x"56",
           644 => x"70",
           645 => x"74",
           646 => x"81",
           647 => x"81",
           648 => x"0b",
           649 => x"62",
           650 => x"55",
           651 => x"8f",
           652 => x"fd",
           653 => x"08",
           654 => x"34",
           655 => x"93",
           656 => x"08",
           657 => x"5f",
           658 => x"76",
           659 => x"58",
           660 => x"55",
           661 => x"09",
           662 => x"38",
           663 => x"5b",
           664 => x"5f",
           665 => x"1c",
           666 => x"06",
           667 => x"33",
           668 => x"70",
           669 => x"27",
           670 => x"07",
           671 => x"5b",
           672 => x"55",
           673 => x"38",
           674 => x"09",
           675 => x"38",
           676 => x"7a",
           677 => x"55",
           678 => x"9f",
           679 => x"32",
           680 => x"ae",
           681 => x"70",
           682 => x"2a",
           683 => x"51",
           684 => x"38",
           685 => x"5a",
           686 => x"77",
           687 => x"81",
           688 => x"1c",
           689 => x"55",
           690 => x"ff",
           691 => x"1e",
           692 => x"55",
           693 => x"83",
           694 => x"74",
           695 => x"7b",
           696 => x"3f",
           697 => x"ef",
           698 => x"7b",
           699 => x"2b",
           700 => x"54",
           701 => x"08",
           702 => x"f8",
           703 => x"08",
           704 => x"80",
           705 => x"33",
           706 => x"2e",
           707 => x"8b",
           708 => x"83",
           709 => x"06",
           710 => x"74",
           711 => x"7d",
           712 => x"88",
           713 => x"5b",
           714 => x"58",
           715 => x"9a",
           716 => x"81",
           717 => x"79",
           718 => x"5b",
           719 => x"31",
           720 => x"75",
           721 => x"38",
           722 => x"80",
           723 => x"7b",
           724 => x"3f",
           725 => x"88",
           726 => x"08",
           727 => x"39",
           728 => x"1c",
           729 => x"33",
           730 => x"a5",
           731 => x"33",
           732 => x"70",
           733 => x"56",
           734 => x"38",
           735 => x"39",
           736 => x"39",
           737 => x"d3",
           738 => x"88",
           739 => x"af",
           740 => x"0c",
           741 => x"04",
           742 => x"79",
           743 => x"82",
           744 => x"53",
           745 => x"51",
           746 => x"83",
           747 => x"80",
           748 => x"51",
           749 => x"88",
           750 => x"ff",
           751 => x"56",
           752 => x"d5",
           753 => x"06",
           754 => x"75",
           755 => x"77",
           756 => x"f6",
           757 => x"08",
           758 => x"94",
           759 => x"f8",
           760 => x"08",
           761 => x"06",
           762 => x"82",
           763 => x"38",
           764 => x"d2",
           765 => x"76",
           766 => x"3f",
           767 => x"88",
           768 => x"76",
           769 => x"3f",
           770 => x"ff",
           771 => x"74",
           772 => x"2e",
           773 => x"56",
           774 => x"89",
           775 => x"ed",
           776 => x"59",
           777 => x"0b",
           778 => x"0c",
           779 => x"88",
           780 => x"55",
           781 => x"82",
           782 => x"75",
           783 => x"70",
           784 => x"fe",
           785 => x"08",
           786 => x"57",
           787 => x"09",
           788 => x"38",
           789 => x"be",
           790 => x"75",
           791 => x"3f",
           792 => x"38",
           793 => x"55",
           794 => x"ac",
           795 => x"e4",
           796 => x"8a",
           797 => x"88",
           798 => x"52",
           799 => x"3f",
           800 => x"ff",
           801 => x"83",
           802 => x"06",
           803 => x"56",
           804 => x"76",
           805 => x"38",
           806 => x"8f",
           807 => x"8d",
           808 => x"75",
           809 => x"3f",
           810 => x"08",
           811 => x"95",
           812 => x"51",
           813 => x"88",
           814 => x"ff",
           815 => x"8c",
           816 => x"f3",
           817 => x"b6",
           818 => x"58",
           819 => x"33",
           820 => x"02",
           821 => x"05",
           822 => x"59",
           823 => x"3f",
           824 => x"ff",
           825 => x"05",
           826 => x"8c",
           827 => x"1a",
           828 => x"e0",
           829 => x"f1",
           830 => x"84",
           831 => x"3d",
           832 => x"f5",
           833 => x"08",
           834 => x"06",
           835 => x"38",
           836 => x"05",
           837 => x"3f",
           838 => x"7a",
           839 => x"3f",
           840 => x"ff",
           841 => x"71",
           842 => x"84",
           843 => x"84",
           844 => x"33",
           845 => x"31",
           846 => x"51",
           847 => x"3f",
           848 => x"05",
           849 => x"0c",
           850 => x"8a",
           851 => x"74",
           852 => x"26",
           853 => x"57",
           854 => x"76",
           855 => x"83",
           856 => x"86",
           857 => x"2e",
           858 => x"76",
           859 => x"83",
           860 => x"06",
           861 => x"3d",
           862 => x"f5",
           863 => x"08",
           864 => x"88",
           865 => x"08",
           866 => x"0c",
           867 => x"ff",
           868 => x"08",
           869 => x"2a",
           870 => x"0c",
           871 => x"81",
           872 => x"0b",
           873 => x"ac",
           874 => x"75",
           875 => x"3d",
           876 => x"3d",
           877 => x"0b",
           878 => x"55",
           879 => x"80",
           880 => x"38",
           881 => x"16",
           882 => x"e0",
           883 => x"54",
           884 => x"54",
           885 => x"51",
           886 => x"88",
           887 => x"08",
           888 => x"88",
           889 => x"73",
           890 => x"38",
           891 => x"33",
           892 => x"70",
           893 => x"55",
           894 => x"2e",
           895 => x"54",
           896 => x"51",
           897 => x"88",
           898 => x"0c",
           899 => x"05",
           900 => x"3f",
           901 => x"16",
           902 => x"16",
           903 => x"81",
           904 => x"88",
           905 => x"0d",
           906 => x"0d",
           907 => x"0b",
           908 => x"ac",
           909 => x"5c",
           910 => x"0c",
           911 => x"80",
           912 => x"38",
           913 => x"81",
           914 => x"57",
           915 => x"81",
           916 => x"39",
           917 => x"34",
           918 => x"0b",
           919 => x"81",
           920 => x"39",
           921 => x"98",
           922 => x"55",
           923 => x"83",
           924 => x"77",
           925 => x"9a",
           926 => x"08",
           927 => x"06",
           928 => x"80",
           929 => x"16",
           930 => x"77",
           931 => x"70",
           932 => x"5b",
           933 => x"38",
           934 => x"a0",
           935 => x"8b",
           936 => x"08",
           937 => x"3f",
           938 => x"81",
           939 => x"aa",
           940 => x"17",
           941 => x"08",
           942 => x"3f",
           943 => x"88",
           944 => x"ff",
           945 => x"08",
           946 => x"0c",
           947 => x"83",
           948 => x"80",
           949 => x"55",
           950 => x"83",
           951 => x"74",
           952 => x"08",
           953 => x"53",
           954 => x"52",
           955 => x"b5",
           956 => x"fe",
           957 => x"16",
           958 => x"17",
           959 => x"31",
           960 => x"7c",
           961 => x"80",
           962 => x"38",
           963 => x"fe",
           964 => x"57",
           965 => x"8c",
           966 => x"fb",
           967 => x"90",
           968 => x"87",
           969 => x"0c",
           970 => x"e4",
           971 => x"94",
           972 => x"80",
           973 => x"c0",
           974 => x"8c",
           975 => x"87",
           976 => x"0c",
           977 => x"f9",
           978 => x"08",
           979 => x"98",
           980 => x"3f",
           981 => x"38",
           982 => x"88",
           983 => x"98",
           984 => x"87",
           985 => x"53",
           986 => x"74",
           987 => x"3f",
           988 => x"38",
           989 => x"80",
           990 => x"73",
           991 => x"39",
           992 => x"73",
           993 => x"fb",
           994 => x"ff",
           995 => x"00",
           996 => x"ff",
           997 => x"ff",
           998 => x"4f",
           999 => x"49",
          1000 => x"52",
          1001 => x"00",
          1002 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e9",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"88",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cb",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"fd",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"80",
           281 => x"e2",
           282 => x"00",
           283 => x"9f",
           284 => x"38",
           285 => x"84",
           286 => x"88",
           287 => x"e2",
           288 => x"04",
           289 => x"94",
           290 => x"0d",
           291 => x"08",
           292 => x"52",
           293 => x"05",
           294 => x"de",
           295 => x"70",
           296 => x"85",
           297 => x"0c",
           298 => x"02",
           299 => x"3d",
           300 => x"94",
           301 => x"08",
           302 => x"88",
           303 => x"82",
           304 => x"08",
           305 => x"54",
           306 => x"94",
           307 => x"08",
           308 => x"f9",
           309 => x"0b",
           310 => x"05",
           311 => x"88",
           312 => x"25",
           313 => x"08",
           314 => x"30",
           315 => x"05",
           316 => x"94",
           317 => x"0c",
           318 => x"05",
           319 => x"81",
           320 => x"f4",
           321 => x"08",
           322 => x"94",
           323 => x"0c",
           324 => x"05",
           325 => x"ab",
           326 => x"8c",
           327 => x"94",
           328 => x"0c",
           329 => x"08",
           330 => x"94",
           331 => x"08",
           332 => x"0b",
           333 => x"05",
           334 => x"f0",
           335 => x"08",
           336 => x"80",
           337 => x"8c",
           338 => x"94",
           339 => x"08",
           340 => x"3f",
           341 => x"94",
           342 => x"0c",
           343 => x"fc",
           344 => x"2e",
           345 => x"08",
           346 => x"30",
           347 => x"05",
           348 => x"f8",
           349 => x"88",
           350 => x"3d",
           351 => x"04",
           352 => x"94",
           353 => x"0d",
           354 => x"08",
           355 => x"94",
           356 => x"08",
           357 => x"38",
           358 => x"05",
           359 => x"08",
           360 => x"81",
           361 => x"fc",
           362 => x"08",
           363 => x"80",
           364 => x"94",
           365 => x"08",
           366 => x"8c",
           367 => x"53",
           368 => x"05",
           369 => x"08",
           370 => x"51",
           371 => x"08",
           372 => x"f8",
           373 => x"94",
           374 => x"08",
           375 => x"38",
           376 => x"05",
           377 => x"08",
           378 => x"94",
           379 => x"08",
           380 => x"54",
           381 => x"94",
           382 => x"08",
           383 => x"fd",
           384 => x"0b",
           385 => x"05",
           386 => x"94",
           387 => x"0c",
           388 => x"05",
           389 => x"88",
           390 => x"ac",
           391 => x"fc",
           392 => x"2e",
           393 => x"0b",
           394 => x"05",
           395 => x"38",
           396 => x"05",
           397 => x"08",
           398 => x"94",
           399 => x"08",
           400 => x"fc",
           401 => x"39",
           402 => x"05",
           403 => x"80",
           404 => x"08",
           405 => x"94",
           406 => x"08",
           407 => x"94",
           408 => x"08",
           409 => x"05",
           410 => x"08",
           411 => x"94",
           412 => x"08",
           413 => x"05",
           414 => x"08",
           415 => x"94",
           416 => x"08",
           417 => x"08",
           418 => x"94",
           419 => x"08",
           420 => x"08",
           421 => x"ff",
           422 => x"08",
           423 => x"80",
           424 => x"94",
           425 => x"08",
           426 => x"f4",
           427 => x"8d",
           428 => x"f8",
           429 => x"94",
           430 => x"0c",
           431 => x"f4",
           432 => x"0c",
           433 => x"94",
           434 => x"3d",
           435 => x"0b",
           436 => x"8c",
           437 => x"87",
           438 => x"0c",
           439 => x"c0",
           440 => x"87",
           441 => x"08",
           442 => x"51",
           443 => x"2e",
           444 => x"c0",
           445 => x"51",
           446 => x"87",
           447 => x"08",
           448 => x"06",
           449 => x"38",
           450 => x"8c",
           451 => x"80",
           452 => x"71",
           453 => x"9f",
           454 => x"0b",
           455 => x"33",
           456 => x"3d",
           457 => x"3d",
           458 => x"7d",
           459 => x"80",
           460 => x"0b",
           461 => x"81",
           462 => x"82",
           463 => x"2e",
           464 => x"81",
           465 => x"0b",
           466 => x"8c",
           467 => x"c0",
           468 => x"84",
           469 => x"92",
           470 => x"c0",
           471 => x"70",
           472 => x"81",
           473 => x"53",
           474 => x"a7",
           475 => x"92",
           476 => x"81",
           477 => x"79",
           478 => x"51",
           479 => x"90",
           480 => x"2e",
           481 => x"76",
           482 => x"58",
           483 => x"54",
           484 => x"72",
           485 => x"70",
           486 => x"38",
           487 => x"8c",
           488 => x"ff",
           489 => x"c0",
           490 => x"51",
           491 => x"81",
           492 => x"92",
           493 => x"c0",
           494 => x"70",
           495 => x"51",
           496 => x"80",
           497 => x"80",
           498 => x"70",
           499 => x"81",
           500 => x"87",
           501 => x"08",
           502 => x"2e",
           503 => x"83",
           504 => x"71",
           505 => x"3d",
           506 => x"3d",
           507 => x"11",
           508 => x"71",
           509 => x"88",
           510 => x"84",
           511 => x"fd",
           512 => x"83",
           513 => x"12",
           514 => x"2b",
           515 => x"07",
           516 => x"70",
           517 => x"2b",
           518 => x"07",
           519 => x"53",
           520 => x"52",
           521 => x"04",
           522 => x"79",
           523 => x"9f",
           524 => x"57",
           525 => x"80",
           526 => x"88",
           527 => x"80",
           528 => x"33",
           529 => x"2e",
           530 => x"83",
           531 => x"80",
           532 => x"54",
           533 => x"fe",
           534 => x"88",
           535 => x"08",
           536 => x"3d",
           537 => x"fd",
           538 => x"08",
           539 => x"51",
           540 => x"88",
           541 => x"ff",
           542 => x"39",
           543 => x"82",
           544 => x"06",
           545 => x"2a",
           546 => x"05",
           547 => x"70",
           548 => x"92",
           549 => x"8e",
           550 => x"fe",
           551 => x"08",
           552 => x"55",
           553 => x"55",
           554 => x"89",
           555 => x"fb",
           556 => x"0b",
           557 => x"08",
           558 => x"12",
           559 => x"55",
           560 => x"56",
           561 => x"8d",
           562 => x"33",
           563 => x"94",
           564 => x"57",
           565 => x"0c",
           566 => x"04",
           567 => x"75",
           568 => x"0b",
           569 => x"ac",
           570 => x"51",
           571 => x"83",
           572 => x"06",
           573 => x"14",
           574 => x"3f",
           575 => x"2b",
           576 => x"51",
           577 => x"88",
           578 => x"ff",
           579 => x"88",
           580 => x"0d",
           581 => x"0d",
           582 => x"0b",
           583 => x"55",
           584 => x"23",
           585 => x"53",
           586 => x"88",
           587 => x"08",
           588 => x"38",
           589 => x"39",
           590 => x"73",
           591 => x"83",
           592 => x"06",
           593 => x"14",
           594 => x"8c",
           595 => x"80",
           596 => x"72",
           597 => x"3f",
           598 => x"85",
           599 => x"08",
           600 => x"16",
           601 => x"71",
           602 => x"3d",
           603 => x"3d",
           604 => x"0b",
           605 => x"08",
           606 => x"05",
           607 => x"ff",
           608 => x"57",
           609 => x"2e",
           610 => x"15",
           611 => x"86",
           612 => x"80",
           613 => x"8f",
           614 => x"80",
           615 => x"13",
           616 => x"8c",
           617 => x"72",
           618 => x"0b",
           619 => x"57",
           620 => x"27",
           621 => x"39",
           622 => x"ff",
           623 => x"2a",
           624 => x"a8",
           625 => x"fc",
           626 => x"52",
           627 => x"27",
           628 => x"52",
           629 => x"17",
           630 => x"38",
           631 => x"16",
           632 => x"51",
           633 => x"88",
           634 => x"0c",
           635 => x"80",
           636 => x"0c",
           637 => x"04",
           638 => x"60",
           639 => x"5e",
           640 => x"55",
           641 => x"09",
           642 => x"38",
           643 => x"44",
           644 => x"62",
           645 => x"56",
           646 => x"09",
           647 => x"38",
           648 => x"80",
           649 => x"0c",
           650 => x"51",
           651 => x"26",
           652 => x"51",
           653 => x"88",
           654 => x"7d",
           655 => x"39",
           656 => x"1d",
           657 => x"5a",
           658 => x"a0",
           659 => x"05",
           660 => x"15",
           661 => x"2e",
           662 => x"ef",
           663 => x"59",
           664 => x"08",
           665 => x"81",
           666 => x"ff",
           667 => x"70",
           668 => x"32",
           669 => x"73",
           670 => x"25",
           671 => x"52",
           672 => x"57",
           673 => x"c7",
           674 => x"2e",
           675 => x"83",
           676 => x"77",
           677 => x"07",
           678 => x"2e",
           679 => x"88",
           680 => x"78",
           681 => x"30",
           682 => x"9f",
           683 => x"57",
           684 => x"9b",
           685 => x"8b",
           686 => x"39",
           687 => x"70",
           688 => x"72",
           689 => x"57",
           690 => x"34",
           691 => x"7a",
           692 => x"80",
           693 => x"26",
           694 => x"55",
           695 => x"34",
           696 => x"b1",
           697 => x"80",
           698 => x"54",
           699 => x"85",
           700 => x"06",
           701 => x"1c",
           702 => x"51",
           703 => x"88",
           704 => x"08",
           705 => x"7c",
           706 => x"80",
           707 => x"38",
           708 => x"70",
           709 => x"81",
           710 => x"56",
           711 => x"8b",
           712 => x"08",
           713 => x"5b",
           714 => x"18",
           715 => x"2e",
           716 => x"70",
           717 => x"33",
           718 => x"05",
           719 => x"71",
           720 => x"56",
           721 => x"e2",
           722 => x"75",
           723 => x"38",
           724 => x"9a",
           725 => x"39",
           726 => x"88",
           727 => x"83",
           728 => x"84",
           729 => x"11",
           730 => x"74",
           731 => x"1d",
           732 => x"2a",
           733 => x"51",
           734 => x"89",
           735 => x"92",
           736 => x"8e",
           737 => x"fa",
           738 => x"08",
           739 => x"fd",
           740 => x"88",
           741 => x"0d",
           742 => x"0d",
           743 => x"57",
           744 => x"fe",
           745 => x"76",
           746 => x"3f",
           747 => x"08",
           748 => x"76",
           749 => x"3f",
           750 => x"ff",
           751 => x"82",
           752 => x"d4",
           753 => x"81",
           754 => x"38",
           755 => x"53",
           756 => x"51",
           757 => x"88",
           758 => x"08",
           759 => x"51",
           760 => x"88",
           761 => x"ff",
           762 => x"81",
           763 => x"a9",
           764 => x"80",
           765 => x"52",
           766 => x"aa",
           767 => x"56",
           768 => x"38",
           769 => x"e2",
           770 => x"83",
           771 => x"55",
           772 => x"c6",
           773 => x"81",
           774 => x"0c",
           775 => x"04",
           776 => x"65",
           777 => x"0b",
           778 => x"ac",
           779 => x"3f",
           780 => x"06",
           781 => x"74",
           782 => x"74",
           783 => x"3d",
           784 => x"5a",
           785 => x"88",
           786 => x"06",
           787 => x"2e",
           788 => x"b3",
           789 => x"83",
           790 => x"52",
           791 => x"c6",
           792 => x"ab",
           793 => x"33",
           794 => x"2e",
           795 => x"3d",
           796 => x"f7",
           797 => x"08",
           798 => x"76",
           799 => x"99",
           800 => x"81",
           801 => x"76",
           802 => x"81",
           803 => x"81",
           804 => x"39",
           805 => x"86",
           806 => x"82",
           807 => x"54",
           808 => x"52",
           809 => x"fe",
           810 => x"88",
           811 => x"38",
           812 => x"05",
           813 => x"3f",
           814 => x"ff",
           815 => x"77",
           816 => x"3d",
           817 => x"f6",
           818 => x"08",
           819 => x"05",
           820 => x"29",
           821 => x"ad",
           822 => x"52",
           823 => x"8a",
           824 => x"83",
           825 => x"7a",
           826 => x"0c",
           827 => x"82",
           828 => x"3d",
           829 => x"f5",
           830 => x"08",
           831 => x"95",
           832 => x"51",
           833 => x"88",
           834 => x"ff",
           835 => x"8c",
           836 => x"ef",
           837 => x"e7",
           838 => x"56",
           839 => x"ca",
           840 => x"83",
           841 => x"76",
           842 => x"31",
           843 => x"70",
           844 => x"1d",
           845 => x"71",
           846 => x"5c",
           847 => x"c4",
           848 => x"82",
           849 => x"1b",
           850 => x"e0",
           851 => x"56",
           852 => x"fe",
           853 => x"82",
           854 => x"f6",
           855 => x"38",
           856 => x"39",
           857 => x"80",
           858 => x"38",
           859 => x"76",
           860 => x"81",
           861 => x"95",
           862 => x"51",
           863 => x"88",
           864 => x"0c",
           865 => x"19",
           866 => x"1a",
           867 => x"ff",
           868 => x"1a",
           869 => x"84",
           870 => x"1b",
           871 => x"0b",
           872 => x"78",
           873 => x"9f",
           874 => x"56",
           875 => x"95",
           876 => x"ea",
           877 => x"0b",
           878 => x"08",
           879 => x"74",
           880 => x"df",
           881 => x"81",
           882 => x"3d",
           883 => x"69",
           884 => x"70",
           885 => x"05",
           886 => x"3f",
           887 => x"88",
           888 => x"38",
           889 => x"54",
           890 => x"93",
           891 => x"05",
           892 => x"2a",
           893 => x"51",
           894 => x"80",
           895 => x"83",
           896 => x"75",
           897 => x"3f",
           898 => x"16",
           899 => x"dc",
           900 => x"eb",
           901 => x"9c",
           902 => x"98",
           903 => x"0b",
           904 => x"73",
           905 => x"3d",
           906 => x"3d",
           907 => x"7e",
           908 => x"9f",
           909 => x"5b",
           910 => x"7b",
           911 => x"75",
           912 => x"d1",
           913 => x"33",
           914 => x"84",
           915 => x"2e",
           916 => x"91",
           917 => x"17",
           918 => x"80",
           919 => x"34",
           920 => x"b1",
           921 => x"08",
           922 => x"31",
           923 => x"27",
           924 => x"58",
           925 => x"81",
           926 => x"16",
           927 => x"ff",
           928 => x"74",
           929 => x"82",
           930 => x"05",
           931 => x"06",
           932 => x"06",
           933 => x"9e",
           934 => x"38",
           935 => x"55",
           936 => x"16",
           937 => x"80",
           938 => x"55",
           939 => x"ff",
           940 => x"a4",
           941 => x"16",
           942 => x"f3",
           943 => x"55",
           944 => x"2e",
           945 => x"88",
           946 => x"17",
           947 => x"08",
           948 => x"84",
           949 => x"51",
           950 => x"27",
           951 => x"55",
           952 => x"16",
           953 => x"06",
           954 => x"08",
           955 => x"f0",
           956 => x"08",
           957 => x"98",
           958 => x"98",
           959 => x"75",
           960 => x"16",
           961 => x"78",
           962 => x"e8",
           963 => x"59",
           964 => x"80",
           965 => x"0c",
           966 => x"04",
           967 => x"9b",
           968 => x"0b",
           969 => x"8c",
           970 => x"86",
           971 => x"c0",
           972 => x"8c",
           973 => x"87",
           974 => x"0c",
           975 => x"0b",
           976 => x"94",
           977 => x"51",
           978 => x"88",
           979 => x"9f",
           980 => x"df",
           981 => x"ae",
           982 => x"0b",
           983 => x"c0",
           984 => x"55",
           985 => x"05",
           986 => x"52",
           987 => x"ba",
           988 => x"8d",
           989 => x"73",
           990 => x"38",
           991 => x"e4",
           992 => x"54",
           993 => x"54",
           994 => x"00",
           995 => x"ff",
           996 => x"ff",
           997 => x"ff",
           998 => x"42",
           999 => x"54",
          1000 => x"2e",
          1001 => x"00",
          1002 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
