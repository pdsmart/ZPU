-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b92",
             1 => x"d8040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b92",
            73 => x"bc040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b929f",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b81bd",
           162 => x"c0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"92a40400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b93",
           171 => x"dd2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b95",
           179 => x"c92d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"94040b0b",
           269 => x"0b8ca304",
           270 => x"0b0b0b8c",
           271 => x"b2040b0b",
           272 => x"0b8cc104",
           273 => x"0b0b0b8c",
           274 => x"d0040b0b",
           275 => x"0b8cdf04",
           276 => x"0b0b0b8c",
           277 => x"ee040b0b",
           278 => x"0b8cfd04",
           279 => x"0b0b0b8d",
           280 => x"8c040b0b",
           281 => x"0b8d9b04",
           282 => x"0b0b0b8d",
           283 => x"aa040b0b",
           284 => x"0b8db904",
           285 => x"0b0b0b8d",
           286 => x"c8040b0b",
           287 => x"0b8dd704",
           288 => x"0b0b0b8d",
           289 => x"e6040b0b",
           290 => x"0b8df504",
           291 => x"0b0b0b8e",
           292 => x"84040b0b",
           293 => x"0b8e9404",
           294 => x"0b0b0b8e",
           295 => x"a4040b0b",
           296 => x"0b8eb404",
           297 => x"0b0b0b8e",
           298 => x"c4040b0b",
           299 => x"0b8ed404",
           300 => x"0b0b0b8e",
           301 => x"e4040b0b",
           302 => x"0b8ef404",
           303 => x"0b0b0b8f",
           304 => x"84040b0b",
           305 => x"0b8f9404",
           306 => x"0b0b0b8f",
           307 => x"a4040b0b",
           308 => x"0b8fb404",
           309 => x"0b0b0b8f",
           310 => x"c4040b0b",
           311 => x"0b8fd404",
           312 => x"0b0b0b8f",
           313 => x"e4040b0b",
           314 => x"0b8ff404",
           315 => x"0b0b0b90",
           316 => x"84040b0b",
           317 => x"0b909404",
           318 => x"0b0b0b90",
           319 => x"a4040b0b",
           320 => x"0b90b404",
           321 => x"0b0b0b90",
           322 => x"c4040b0b",
           323 => x"0b90d404",
           324 => x"0b0b0b90",
           325 => x"e4040b0b",
           326 => x"0b90f404",
           327 => x"0b0b0b91",
           328 => x"84040b0b",
           329 => x"0b919404",
           330 => x"0b0b0b91",
           331 => x"a3040b0b",
           332 => x"0b91b204",
           333 => x"0b0b0b91",
           334 => x"c1040b0b",
           335 => x"0b91d004",
           336 => x"0b0b0b91",
           337 => x"df040b0b",
           338 => x"0b91ee04",
           339 => x"ffffffff",
           340 => x"ffffffff",
           341 => x"ffffffff",
           342 => x"ffffffff",
           343 => x"ffffffff",
           344 => x"ffffffff",
           345 => x"ffffffff",
           346 => x"ffffffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0481d3e4",
           386 => x"0ca0ae2d",
           387 => x"81d3e408",
           388 => x"82809004",
           389 => x"81d3e40c",
           390 => x"aadc2d81",
           391 => x"d3e40882",
           392 => x"80900481",
           393 => x"d3e40cab",
           394 => x"9b2d81d3",
           395 => x"e4088280",
           396 => x"900481d3",
           397 => x"e40cabb9",
           398 => x"2d81d3e4",
           399 => x"08828090",
           400 => x"0481d3e4",
           401 => x"0cb1f72d",
           402 => x"81d3e408",
           403 => x"82809004",
           404 => x"81d3e40c",
           405 => x"b2f52d81",
           406 => x"d3e40882",
           407 => x"80900481",
           408 => x"d3e40cab",
           409 => x"dc2d81d3",
           410 => x"e4088280",
           411 => x"900481d3",
           412 => x"e40cb392",
           413 => x"2d81d3e4",
           414 => x"08828090",
           415 => x"0481d3e4",
           416 => x"0cb5842d",
           417 => x"81d3e408",
           418 => x"82809004",
           419 => x"81d3e40c",
           420 => x"b19d2d81",
           421 => x"d3e40882",
           422 => x"80900481",
           423 => x"d3e40cb1",
           424 => x"b32d81d3",
           425 => x"e4088280",
           426 => x"900481d3",
           427 => x"e40cb1d7",
           428 => x"2d81d3e4",
           429 => x"08828090",
           430 => x"0481d3e4",
           431 => x"0ca2bb2d",
           432 => x"81d3e408",
           433 => x"82809004",
           434 => x"81d3e40c",
           435 => x"a38c2d81",
           436 => x"d3e40882",
           437 => x"80900481",
           438 => x"d3e40c9b",
           439 => x"a82d81d3",
           440 => x"e4088280",
           441 => x"900481d3",
           442 => x"e40c9cdd",
           443 => x"2d81d3e4",
           444 => x"08828090",
           445 => x"0481d3e4",
           446 => x"0c9e902d",
           447 => x"81d3e408",
           448 => x"82809004",
           449 => x"81d3e40c",
           450 => x"80e7b92d",
           451 => x"81d3e408",
           452 => x"82809004",
           453 => x"81d3e40c",
           454 => x"80f4aa2d",
           455 => x"81d3e408",
           456 => x"82809004",
           457 => x"81d3e40c",
           458 => x"80ec9e2d",
           459 => x"81d3e408",
           460 => x"82809004",
           461 => x"81d3e40c",
           462 => x"80ef9b2d",
           463 => x"81d3e408",
           464 => x"82809004",
           465 => x"81d3e40c",
           466 => x"80f9b92d",
           467 => x"81d3e408",
           468 => x"82809004",
           469 => x"81d3e40c",
           470 => x"8182992d",
           471 => x"81d3e408",
           472 => x"82809004",
           473 => x"81d3e40c",
           474 => x"80f38c2d",
           475 => x"81d3e408",
           476 => x"82809004",
           477 => x"81d3e40c",
           478 => x"80fcd82d",
           479 => x"81d3e408",
           480 => x"82809004",
           481 => x"81d3e40c",
           482 => x"80fdf72d",
           483 => x"81d3e408",
           484 => x"82809004",
           485 => x"81d3e40c",
           486 => x"80fe962d",
           487 => x"81d3e408",
           488 => x"82809004",
           489 => x"81d3e40c",
           490 => x"8186802d",
           491 => x"81d3e408",
           492 => x"82809004",
           493 => x"81d3e40c",
           494 => x"8183e62d",
           495 => x"81d3e408",
           496 => x"82809004",
           497 => x"81d3e40c",
           498 => x"8188d42d",
           499 => x"81d3e408",
           500 => x"82809004",
           501 => x"81d3e40c",
           502 => x"80ff9a2d",
           503 => x"81d3e408",
           504 => x"82809004",
           505 => x"81d3e40c",
           506 => x"818bd42d",
           507 => x"81d3e408",
           508 => x"82809004",
           509 => x"81d3e40c",
           510 => x"818cd52d",
           511 => x"81d3e408",
           512 => x"82809004",
           513 => x"81d3e40c",
           514 => x"80f58a2d",
           515 => x"81d3e408",
           516 => x"82809004",
           517 => x"81d3e40c",
           518 => x"80f4e32d",
           519 => x"81d3e408",
           520 => x"82809004",
           521 => x"81d3e40c",
           522 => x"80f68e2d",
           523 => x"81d3e408",
           524 => x"82809004",
           525 => x"81d3e40c",
           526 => x"80fff12d",
           527 => x"81d3e408",
           528 => x"82809004",
           529 => x"81d3e40c",
           530 => x"818dc62d",
           531 => x"81d3e408",
           532 => x"82809004",
           533 => x"81d3e40c",
           534 => x"818fd02d",
           535 => x"81d3e408",
           536 => x"82809004",
           537 => x"81d3e40c",
           538 => x"8193922d",
           539 => x"81d3e408",
           540 => x"82809004",
           541 => x"81d3e40c",
           542 => x"80e6d82d",
           543 => x"81d3e408",
           544 => x"82809004",
           545 => x"81d3e40c",
           546 => x"8195fe2d",
           547 => x"81d3e408",
           548 => x"82809004",
           549 => x"81d3e40c",
           550 => x"b8932d81",
           551 => x"d3e40882",
           552 => x"80900481",
           553 => x"d3e40cb9",
           554 => x"fd2d81d3",
           555 => x"e4088280",
           556 => x"900481d3",
           557 => x"e40cbbe1",
           558 => x"2d81d3e4",
           559 => x"08828090",
           560 => x"0481d3e4",
           561 => x"0c9bd12d",
           562 => x"81d3e408",
           563 => x"82809004",
           564 => x"81d3e40c",
           565 => x"9cb32d81",
           566 => x"d3e40882",
           567 => x"80900481",
           568 => x"d3e40c9f",
           569 => x"a02d81d3",
           570 => x"e4088280",
           571 => x"900481d3",
           572 => x"e40c81a2",
           573 => x"f92d81d3",
           574 => x"e4088280",
           575 => x"90043c04",
           576 => x"10101010",
           577 => x"10101010",
           578 => x"10101010",
           579 => x"10101010",
           580 => x"10101010",
           581 => x"10101010",
           582 => x"10101010",
           583 => x"10101053",
           584 => x"51040000",
           585 => x"7381ff06",
           586 => x"73830609",
           587 => x"81058305",
           588 => x"1010102b",
           589 => x"0772fc06",
           590 => x"0c515104",
           591 => x"72728072",
           592 => x"8106ff05",
           593 => x"09720605",
           594 => x"71105272",
           595 => x"0a100a53",
           596 => x"72ed3851",
           597 => x"51535104",
           598 => x"81d3d870",
           599 => x"81eb8427",
           600 => x"8e388071",
           601 => x"70840553",
           602 => x"0c0b0b0b",
           603 => x"92db048c",
           604 => x"815181bc",
           605 => x"d9040081",
           606 => x"d3e40802",
           607 => x"81d3e40c",
           608 => x"fd3d0d80",
           609 => x"5381d3e4",
           610 => x"088c0508",
           611 => x"5281d3e4",
           612 => x"08880508",
           613 => x"5183d43f",
           614 => x"81d3d808",
           615 => x"7081d3d8",
           616 => x"0c54853d",
           617 => x"0d81d3e4",
           618 => x"0c0481d3",
           619 => x"e4080281",
           620 => x"d3e40cfd",
           621 => x"3d0d8153",
           622 => x"81d3e408",
           623 => x"8c050852",
           624 => x"81d3e408",
           625 => x"88050851",
           626 => x"83a13f81",
           627 => x"d3d80870",
           628 => x"81d3d80c",
           629 => x"54853d0d",
           630 => x"81d3e40c",
           631 => x"0481d3e4",
           632 => x"080281d3",
           633 => x"e40cf93d",
           634 => x"0d800b81",
           635 => x"d3e408fc",
           636 => x"050c81d3",
           637 => x"e4088805",
           638 => x"088025b9",
           639 => x"3881d3e4",
           640 => x"08880508",
           641 => x"3081d3e4",
           642 => x"0888050c",
           643 => x"800b81d3",
           644 => x"e408f405",
           645 => x"0c81d3e4",
           646 => x"08fc0508",
           647 => x"8a38810b",
           648 => x"81d3e408",
           649 => x"f4050c81",
           650 => x"d3e408f4",
           651 => x"050881d3",
           652 => x"e408fc05",
           653 => x"0c81d3e4",
           654 => x"088c0508",
           655 => x"8025b938",
           656 => x"81d3e408",
           657 => x"8c050830",
           658 => x"81d3e408",
           659 => x"8c050c80",
           660 => x"0b81d3e4",
           661 => x"08f0050c",
           662 => x"81d3e408",
           663 => x"fc05088a",
           664 => x"38810b81",
           665 => x"d3e408f0",
           666 => x"050c81d3",
           667 => x"e408f005",
           668 => x"0881d3e4",
           669 => x"08fc050c",
           670 => x"805381d3",
           671 => x"e4088c05",
           672 => x"085281d3",
           673 => x"e4088805",
           674 => x"085181df",
           675 => x"3f81d3d8",
           676 => x"087081d3",
           677 => x"e408f805",
           678 => x"0c5481d3",
           679 => x"e408fc05",
           680 => x"08802e90",
           681 => x"3881d3e4",
           682 => x"08f80508",
           683 => x"3081d3e4",
           684 => x"08f8050c",
           685 => x"81d3e408",
           686 => x"f8050870",
           687 => x"81d3d80c",
           688 => x"54893d0d",
           689 => x"81d3e40c",
           690 => x"0481d3e4",
           691 => x"080281d3",
           692 => x"e40cfb3d",
           693 => x"0d800b81",
           694 => x"d3e408fc",
           695 => x"050c81d3",
           696 => x"e4088805",
           697 => x"08802599",
           698 => x"3881d3e4",
           699 => x"08880508",
           700 => x"3081d3e4",
           701 => x"0888050c",
           702 => x"810b81d3",
           703 => x"e408fc05",
           704 => x"0c81d3e4",
           705 => x"088c0508",
           706 => x"80259038",
           707 => x"81d3e408",
           708 => x"8c050830",
           709 => x"81d3e408",
           710 => x"8c050c81",
           711 => x"5381d3e4",
           712 => x"088c0508",
           713 => x"5281d3e4",
           714 => x"08880508",
           715 => x"51bd3f81",
           716 => x"d3d80870",
           717 => x"81d3e408",
           718 => x"f8050c54",
           719 => x"81d3e408",
           720 => x"fc050880",
           721 => x"2e903881",
           722 => x"d3e408f8",
           723 => x"05083081",
           724 => x"d3e408f8",
           725 => x"050c81d3",
           726 => x"e408f805",
           727 => x"087081d3",
           728 => x"d80c5487",
           729 => x"3d0d81d3",
           730 => x"e40c0481",
           731 => x"d3e40802",
           732 => x"81d3e40c",
           733 => x"fd3d0d81",
           734 => x"0b81d3e4",
           735 => x"08fc050c",
           736 => x"800b81d3",
           737 => x"e408f805",
           738 => x"0c81d3e4",
           739 => x"088c0508",
           740 => x"81d3e408",
           741 => x"88050827",
           742 => x"b93881d3",
           743 => x"e408fc05",
           744 => x"08802eae",
           745 => x"38800b81",
           746 => x"d3e4088c",
           747 => x"050824a2",
           748 => x"3881d3e4",
           749 => x"088c0508",
           750 => x"1081d3e4",
           751 => x"088c050c",
           752 => x"81d3e408",
           753 => x"fc050810",
           754 => x"81d3e408",
           755 => x"fc050cff",
           756 => x"b83981d3",
           757 => x"e408fc05",
           758 => x"08802e80",
           759 => x"e13881d3",
           760 => x"e4088c05",
           761 => x"0881d3e4",
           762 => x"08880508",
           763 => x"26ad3881",
           764 => x"d3e40888",
           765 => x"050881d3",
           766 => x"e4088c05",
           767 => x"083181d3",
           768 => x"e4088805",
           769 => x"0c81d3e4",
           770 => x"08f80508",
           771 => x"81d3e408",
           772 => x"fc050807",
           773 => x"81d3e408",
           774 => x"f8050c81",
           775 => x"d3e408fc",
           776 => x"0508812a",
           777 => x"81d3e408",
           778 => x"fc050c81",
           779 => x"d3e4088c",
           780 => x"0508812a",
           781 => x"81d3e408",
           782 => x"8c050cff",
           783 => x"953981d3",
           784 => x"e4089005",
           785 => x"08802e93",
           786 => x"3881d3e4",
           787 => x"08880508",
           788 => x"7081d3e4",
           789 => x"08f4050c",
           790 => x"51913981",
           791 => x"d3e408f8",
           792 => x"05087081",
           793 => x"d3e408f4",
           794 => x"050c5181",
           795 => x"d3e408f4",
           796 => x"050881d3",
           797 => x"d80c853d",
           798 => x"0d81d3e4",
           799 => x"0c04fc3d",
           800 => x"0d767971",
           801 => x"028c059f",
           802 => x"05335755",
           803 => x"53558372",
           804 => x"278a3874",
           805 => x"83065170",
           806 => x"802ea438",
           807 => x"ff125271",
           808 => x"ff2e9338",
           809 => x"73737081",
           810 => x"055534ff",
           811 => x"125271ff",
           812 => x"2e098106",
           813 => x"ef387481",
           814 => x"d3d80c86",
           815 => x"3d0d0474",
           816 => x"74882b75",
           817 => x"07707190",
           818 => x"2b075154",
           819 => x"518f7227",
           820 => x"a5387271",
           821 => x"70840553",
           822 => x"0c727170",
           823 => x"8405530c",
           824 => x"72717084",
           825 => x"05530c72",
           826 => x"71708405",
           827 => x"530cf012",
           828 => x"52718f26",
           829 => x"dd388372",
           830 => x"27903872",
           831 => x"71708405",
           832 => x"530cfc12",
           833 => x"52718326",
           834 => x"f2387053",
           835 => x"ff8e39fb",
           836 => x"3d0d7779",
           837 => x"70720783",
           838 => x"06535452",
           839 => x"70933871",
           840 => x"73730854",
           841 => x"56547173",
           842 => x"082e80c6",
           843 => x"38737554",
           844 => x"52713370",
           845 => x"81ff0652",
           846 => x"5470802e",
           847 => x"9d387233",
           848 => x"5570752e",
           849 => x"09810695",
           850 => x"38811281",
           851 => x"14713370",
           852 => x"81ff0654",
           853 => x"56545270",
           854 => x"e5387233",
           855 => x"557381ff",
           856 => x"067581ff",
           857 => x"06717131",
           858 => x"81d3d80c",
           859 => x"5252873d",
           860 => x"0d047109",
           861 => x"70f7fbfd",
           862 => x"ff140670",
           863 => x"f8848281",
           864 => x"80065151",
           865 => x"51709738",
           866 => x"84148416",
           867 => x"71085456",
           868 => x"54717508",
           869 => x"2edc3873",
           870 => x"755452ff",
           871 => x"9439800b",
           872 => x"81d3d80c",
           873 => x"873d0d04",
           874 => x"fe3d0d80",
           875 => x"52835371",
           876 => x"882b5287",
           877 => x"863f81d3",
           878 => x"d80881ff",
           879 => x"067207ff",
           880 => x"14545272",
           881 => x"8025e838",
           882 => x"7181d3d8",
           883 => x"0c843d0d",
           884 => x"04fb3d0d",
           885 => x"77700870",
           886 => x"53535671",
           887 => x"802e80ca",
           888 => x"38713351",
           889 => x"70a02e09",
           890 => x"81068638",
           891 => x"811252f1",
           892 => x"39715384",
           893 => x"39811353",
           894 => x"80733370",
           895 => x"81ff0653",
           896 => x"555570a0",
           897 => x"2e833881",
           898 => x"5570802e",
           899 => x"843874e5",
           900 => x"387381ff",
           901 => x"065170a0",
           902 => x"2e098106",
           903 => x"88388073",
           904 => x"70810555",
           905 => x"3472760c",
           906 => x"71517081",
           907 => x"d3d80c87",
           908 => x"3d0d04fc",
           909 => x"3d0d7653",
           910 => x"7208802e",
           911 => x"9138863d",
           912 => x"fc055272",
           913 => x"5198bd3f",
           914 => x"81d3d808",
           915 => x"85388053",
           916 => x"83397453",
           917 => x"7281d3d8",
           918 => x"0c863d0d",
           919 => x"04fc3d0d",
           920 => x"76821133",
           921 => x"ff055253",
           922 => x"8152708b",
           923 => x"26819838",
           924 => x"831333ff",
           925 => x"05518252",
           926 => x"709e2681",
           927 => x"8a388413",
           928 => x"33518352",
           929 => x"70972680",
           930 => x"fe388513",
           931 => x"33518452",
           932 => x"70bb2680",
           933 => x"f2388613",
           934 => x"33518552",
           935 => x"70bb2680",
           936 => x"e6388813",
           937 => x"22558652",
           938 => x"7487e726",
           939 => x"80d9388a",
           940 => x"13225487",
           941 => x"527387e7",
           942 => x"2680cc38",
           943 => x"810b87c0",
           944 => x"989c0c72",
           945 => x"2287c098",
           946 => x"bc0c8213",
           947 => x"3387c098",
           948 => x"b80c8313",
           949 => x"3387c098",
           950 => x"b40c8413",
           951 => x"3387c098",
           952 => x"b00c8513",
           953 => x"3387c098",
           954 => x"ac0c8613",
           955 => x"3387c098",
           956 => x"a80c7487",
           957 => x"c098a40c",
           958 => x"7387c098",
           959 => x"a00c800b",
           960 => x"87c0989c",
           961 => x"0c805271",
           962 => x"81d3d80c",
           963 => x"863d0d04",
           964 => x"f33d0d7f",
           965 => x"5b87c098",
           966 => x"9c5d817d",
           967 => x"0c87c098",
           968 => x"bc085e7d",
           969 => x"7b2387c0",
           970 => x"98b8085a",
           971 => x"79821c34",
           972 => x"87c098b4",
           973 => x"085a7983",
           974 => x"1c3487c0",
           975 => x"98b0085a",
           976 => x"79841c34",
           977 => x"87c098ac",
           978 => x"085a7985",
           979 => x"1c3487c0",
           980 => x"98a8085a",
           981 => x"79861c34",
           982 => x"87c098a4",
           983 => x"085c7b88",
           984 => x"1c2387c0",
           985 => x"98a0085a",
           986 => x"798a1c23",
           987 => x"807d0c79",
           988 => x"83ffff06",
           989 => x"597b83ff",
           990 => x"ff065886",
           991 => x"1b335785",
           992 => x"1b335684",
           993 => x"1b335583",
           994 => x"1b335482",
           995 => x"1b33537d",
           996 => x"83ffff06",
           997 => x"5281beb4",
           998 => x"5192823f",
           999 => x"8f3d0d04",
          1000 => x"ff3d0d02",
          1001 => x"8f053370",
          1002 => x"30709f2a",
          1003 => x"51525270",
          1004 => x"0b0b81d0",
          1005 => x"dc34833d",
          1006 => x"0d04fb3d",
          1007 => x"0d770b0b",
          1008 => x"81d0dc33",
          1009 => x"7081ff06",
          1010 => x"57555687",
          1011 => x"c0948451",
          1012 => x"74802e86",
          1013 => x"3887c094",
          1014 => x"94517008",
          1015 => x"70962a70",
          1016 => x"81065354",
          1017 => x"5270802e",
          1018 => x"8c387191",
          1019 => x"2a708106",
          1020 => x"515170d7",
          1021 => x"38728132",
          1022 => x"70810651",
          1023 => x"5170802e",
          1024 => x"8d387193",
          1025 => x"2a708106",
          1026 => x"515170ff",
          1027 => x"be387381",
          1028 => x"ff065187",
          1029 => x"c0948052",
          1030 => x"70802e86",
          1031 => x"3887c094",
          1032 => x"90527572",
          1033 => x"0c7581d3",
          1034 => x"d80c873d",
          1035 => x"0d04fb3d",
          1036 => x"0d029f05",
          1037 => x"330b0b81",
          1038 => x"d0dc3370",
          1039 => x"81ff0657",
          1040 => x"555687c0",
          1041 => x"94845174",
          1042 => x"802e8638",
          1043 => x"87c09494",
          1044 => x"51700870",
          1045 => x"962a7081",
          1046 => x"06535452",
          1047 => x"70802e8c",
          1048 => x"3871912a",
          1049 => x"70810651",
          1050 => x"5170d738",
          1051 => x"72813270",
          1052 => x"81065151",
          1053 => x"70802e8d",
          1054 => x"3871932a",
          1055 => x"70810651",
          1056 => x"5170ffbe",
          1057 => x"387381ff",
          1058 => x"065187c0",
          1059 => x"94805270",
          1060 => x"802e8638",
          1061 => x"87c09490",
          1062 => x"5275720c",
          1063 => x"873d0d04",
          1064 => x"f93d0d79",
          1065 => x"54807433",
          1066 => x"7081ff06",
          1067 => x"53535770",
          1068 => x"772e80fe",
          1069 => x"387181ff",
          1070 => x"0681150b",
          1071 => x"0b81d0dc",
          1072 => x"337081ff",
          1073 => x"06595755",
          1074 => x"5887c094",
          1075 => x"84517580",
          1076 => x"2e863887",
          1077 => x"c0949451",
          1078 => x"70087096",
          1079 => x"2a708106",
          1080 => x"53545270",
          1081 => x"802e8c38",
          1082 => x"71912a70",
          1083 => x"81065151",
          1084 => x"70d73872",
          1085 => x"81327081",
          1086 => x"06515170",
          1087 => x"802e8d38",
          1088 => x"71932a70",
          1089 => x"81065151",
          1090 => x"70ffbe38",
          1091 => x"7481ff06",
          1092 => x"5187c094",
          1093 => x"80527080",
          1094 => x"2e863887",
          1095 => x"c0949052",
          1096 => x"77720c81",
          1097 => x"17743370",
          1098 => x"81ff0653",
          1099 => x"535770ff",
          1100 => x"84387681",
          1101 => x"d3d80c89",
          1102 => x"3d0d04fe",
          1103 => x"3d0d0b0b",
          1104 => x"81d0dc33",
          1105 => x"7081ff06",
          1106 => x"545287c0",
          1107 => x"94845172",
          1108 => x"802e8638",
          1109 => x"87c09494",
          1110 => x"51700870",
          1111 => x"822a7081",
          1112 => x"06515151",
          1113 => x"70802ee2",
          1114 => x"387181ff",
          1115 => x"065187c0",
          1116 => x"94805270",
          1117 => x"802e8638",
          1118 => x"87c09490",
          1119 => x"52710870",
          1120 => x"81ff0681",
          1121 => x"d3d80c51",
          1122 => x"843d0d04",
          1123 => x"fe3d0d0b",
          1124 => x"0b81d0dc",
          1125 => x"337081ff",
          1126 => x"06525387",
          1127 => x"c0948452",
          1128 => x"70802e86",
          1129 => x"3887c094",
          1130 => x"94527108",
          1131 => x"70822a70",
          1132 => x"81065151",
          1133 => x"51ff5270",
          1134 => x"802ea038",
          1135 => x"7281ff06",
          1136 => x"5187c094",
          1137 => x"80527080",
          1138 => x"2e863887",
          1139 => x"c0949052",
          1140 => x"71087098",
          1141 => x"2b70982c",
          1142 => x"51535171",
          1143 => x"81d3d80c",
          1144 => x"843d0d04",
          1145 => x"ff3d0d87",
          1146 => x"c09e8008",
          1147 => x"709c2a8a",
          1148 => x"06515170",
          1149 => x"802e8393",
          1150 => x"3887c09e",
          1151 => x"9c0881d0",
          1152 => x"e00c87c0",
          1153 => x"9ea00881",
          1154 => x"d0e40c87",
          1155 => x"c09e8c08",
          1156 => x"81d0e80c",
          1157 => x"87c09e90",
          1158 => x"0881d0ec",
          1159 => x"0c87c09e",
          1160 => x"940881d0",
          1161 => x"f00c87c0",
          1162 => x"9e980881",
          1163 => x"d0f40c87",
          1164 => x"c09ea408",
          1165 => x"81d0f80c",
          1166 => x"87c09ea8",
          1167 => x"0881d0fc",
          1168 => x"0c87c09e",
          1169 => x"ac0881d1",
          1170 => x"800c87c0",
          1171 => x"9e800851",
          1172 => x"7081d184",
          1173 => x"2387c09e",
          1174 => x"840881d1",
          1175 => x"880c810b",
          1176 => x"81d18c34",
          1177 => x"800b87c0",
          1178 => x"9e880870",
          1179 => x"a0800651",
          1180 => x"52527080",
          1181 => x"2e833881",
          1182 => x"527181d1",
          1183 => x"8d34800b",
          1184 => x"87c09e88",
          1185 => x"08708180",
          1186 => x"80065152",
          1187 => x"5270802e",
          1188 => x"83388152",
          1189 => x"7181d18e",
          1190 => x"34800b87",
          1191 => x"c09e8808",
          1192 => x"7080c080",
          1193 => x"06515252",
          1194 => x"70802e83",
          1195 => x"38815271",
          1196 => x"81d18f34",
          1197 => x"800b87c0",
          1198 => x"9e880870",
          1199 => x"90800651",
          1200 => x"52527080",
          1201 => x"2e833881",
          1202 => x"527181d1",
          1203 => x"9034800b",
          1204 => x"87c09e88",
          1205 => x"08708880",
          1206 => x"06515252",
          1207 => x"70802e83",
          1208 => x"38815271",
          1209 => x"81d19134",
          1210 => x"800b87c0",
          1211 => x"9e880870",
          1212 => x"84800651",
          1213 => x"52527080",
          1214 => x"2e833881",
          1215 => x"527181d1",
          1216 => x"9234800b",
          1217 => x"87c09e88",
          1218 => x"08708280",
          1219 => x"06515252",
          1220 => x"70802e83",
          1221 => x"38815271",
          1222 => x"81d19334",
          1223 => x"800b87c0",
          1224 => x"9e880870",
          1225 => x"81800651",
          1226 => x"52527080",
          1227 => x"2e833881",
          1228 => x"527181d1",
          1229 => x"943487c0",
          1230 => x"9e880870",
          1231 => x"80e00670",
          1232 => x"862c5151",
          1233 => x"517081d1",
          1234 => x"9534800b",
          1235 => x"87c09e88",
          1236 => x"08709006",
          1237 => x"51525270",
          1238 => x"802e8338",
          1239 => x"81527181",
          1240 => x"d1963480",
          1241 => x"0b87c09e",
          1242 => x"88087088",
          1243 => x"06515252",
          1244 => x"70802e83",
          1245 => x"38815271",
          1246 => x"81d19734",
          1247 => x"87c09e88",
          1248 => x"08708706",
          1249 => x"51517081",
          1250 => x"d1983483",
          1251 => x"3d0d04fd",
          1252 => x"3d0d81be",
          1253 => x"cc5184a1",
          1254 => x"3f81d18c",
          1255 => x"33547380",
          1256 => x"2e883881",
          1257 => x"bee05184",
          1258 => x"903f81be",
          1259 => x"f4518489",
          1260 => x"3f81d18d",
          1261 => x"33547380",
          1262 => x"2e923881",
          1263 => x"d0e40853",
          1264 => x"81d0e008",
          1265 => x"5281bf8c",
          1266 => x"5189d23f",
          1267 => x"81d18e33",
          1268 => x"5473802e",
          1269 => x"923881d0",
          1270 => x"ec085381",
          1271 => x"d0e80852",
          1272 => x"81bfb451",
          1273 => x"89b73f81",
          1274 => x"d18f3354",
          1275 => x"738b3881",
          1276 => x"d1903354",
          1277 => x"73802e92",
          1278 => x"3881d0f4",
          1279 => x"085381d0",
          1280 => x"f0085281",
          1281 => x"bfd85189",
          1282 => x"943f81d1",
          1283 => x"91335473",
          1284 => x"802e8838",
          1285 => x"81bffc51",
          1286 => x"839f3f81",
          1287 => x"d1923354",
          1288 => x"73802e88",
          1289 => x"3881c088",
          1290 => x"51838e3f",
          1291 => x"81d19333",
          1292 => x"5473802e",
          1293 => x"883881c0",
          1294 => x"945182fd",
          1295 => x"3f81d194",
          1296 => x"33547380",
          1297 => x"2e8d3881",
          1298 => x"d1953352",
          1299 => x"81c0a051",
          1300 => x"88cb3f81",
          1301 => x"d1963354",
          1302 => x"73802e88",
          1303 => x"3881c0c0",
          1304 => x"5182d63f",
          1305 => x"81d19733",
          1306 => x"5473802e",
          1307 => x"8d3881d1",
          1308 => x"98335281",
          1309 => x"c0dc5188",
          1310 => x"a43f81c0",
          1311 => x"f85182b9",
          1312 => x"3f81d0f8",
          1313 => x"085281c1",
          1314 => x"84518891",
          1315 => x"3f81d0fc",
          1316 => x"085281c1",
          1317 => x"ac518885",
          1318 => x"3f81d180",
          1319 => x"085281c1",
          1320 => x"d45187f9",
          1321 => x"3f81d184",
          1322 => x"225281c1",
          1323 => x"fc5187ed",
          1324 => x"3f81d188",
          1325 => x"085281c2",
          1326 => x"a45187e1",
          1327 => x"3f853d0d",
          1328 => x"04fe3d0d",
          1329 => x"02920533",
          1330 => x"ff055271",
          1331 => x"8426aa38",
          1332 => x"71842981",
          1333 => x"bdd00552",
          1334 => x"71080481",
          1335 => x"c2cc519d",
          1336 => x"3981c2d4",
          1337 => x"51973981",
          1338 => x"c2dc5191",
          1339 => x"3981c2e4",
          1340 => x"518b3981",
          1341 => x"c2e85185",
          1342 => x"3981c2f0",
          1343 => x"51f7a13f",
          1344 => x"843d0d04",
          1345 => x"7188800c",
          1346 => x"04800b87",
          1347 => x"c096840c",
          1348 => x"04ff3d0d",
          1349 => x"87c09684",
          1350 => x"70085252",
          1351 => x"80720c70",
          1352 => x"74077081",
          1353 => x"d19c0c72",
          1354 => x"0c833d0d",
          1355 => x"04ff3d0d",
          1356 => x"87c09684",
          1357 => x"700881d1",
          1358 => x"9c0c5280",
          1359 => x"720c7309",
          1360 => x"7081d19c",
          1361 => x"08067081",
          1362 => x"d19c0c73",
          1363 => x"0c51833d",
          1364 => x"0d0481d1",
          1365 => x"9c0887c0",
          1366 => x"96840c04",
          1367 => x"fe3d0d02",
          1368 => x"93053353",
          1369 => x"728a2e09",
          1370 => x"81068538",
          1371 => x"8d51ed3f",
          1372 => x"81d3f008",
          1373 => x"5271802e",
          1374 => x"90387272",
          1375 => x"3481d3f0",
          1376 => x"08810581",
          1377 => x"d3f00c8f",
          1378 => x"3981d3e8",
          1379 => x"08527180",
          1380 => x"2e853872",
          1381 => x"51712d84",
          1382 => x"3d0d04fe",
          1383 => x"3d0d0297",
          1384 => x"053381d3",
          1385 => x"e8087681",
          1386 => x"d3e80c54",
          1387 => x"51ffad3f",
          1388 => x"7281d3e8",
          1389 => x"0c843d0d",
          1390 => x"04fd3d0d",
          1391 => x"75547333",
          1392 => x"7081ff06",
          1393 => x"53537180",
          1394 => x"2e8e3872",
          1395 => x"81ff0651",
          1396 => x"811454ff",
          1397 => x"873fe739",
          1398 => x"853d0d04",
          1399 => x"fc3d0d77",
          1400 => x"81d3e808",
          1401 => x"7881d3e8",
          1402 => x"0c565473",
          1403 => x"337081ff",
          1404 => x"06535371",
          1405 => x"802e8e38",
          1406 => x"7281ff06",
          1407 => x"51811454",
          1408 => x"feda3fe7",
          1409 => x"397481d3",
          1410 => x"e80c863d",
          1411 => x"0d04ec3d",
          1412 => x"0d666859",
          1413 => x"59787081",
          1414 => x"055a3356",
          1415 => x"75802e84",
          1416 => x"f83875a5",
          1417 => x"2e098106",
          1418 => x"82de3880",
          1419 => x"707a7081",
          1420 => x"055c3358",
          1421 => x"5b5b75b0",
          1422 => x"2e098106",
          1423 => x"8538815a",
          1424 => x"8b3975ad",
          1425 => x"2e098106",
          1426 => x"8a38825a",
          1427 => x"78708105",
          1428 => x"5a335675",
          1429 => x"aa2e0981",
          1430 => x"06923877",
          1431 => x"84197108",
          1432 => x"7b708105",
          1433 => x"5d33595d",
          1434 => x"59539d39",
          1435 => x"d0165372",
          1436 => x"89269538",
          1437 => x"7a88297b",
          1438 => x"10057605",
          1439 => x"d0057970",
          1440 => x"81055b33",
          1441 => x"575be539",
          1442 => x"7580ec32",
          1443 => x"70307072",
          1444 => x"07802578",
          1445 => x"80cc3270",
          1446 => x"30707207",
          1447 => x"80257307",
          1448 => x"53545851",
          1449 => x"55537380",
          1450 => x"2e8c3879",
          1451 => x"84077970",
          1452 => x"81055b33",
          1453 => x"575a7580",
          1454 => x"2e83de38",
          1455 => x"755480e0",
          1456 => x"76278938",
          1457 => x"e0167081",
          1458 => x"ff065553",
          1459 => x"7380cf2e",
          1460 => x"81aa3873",
          1461 => x"80cf24a2",
          1462 => x"387380c3",
          1463 => x"2e818e38",
          1464 => x"7380c324",
          1465 => x"8b387380",
          1466 => x"c22e818c",
          1467 => x"38819939",
          1468 => x"7380c42e",
          1469 => x"818a3881",
          1470 => x"8f397380",
          1471 => x"d52e8180",
          1472 => x"387380d5",
          1473 => x"248a3873",
          1474 => x"80d32e8e",
          1475 => x"3880f939",
          1476 => x"7380d82e",
          1477 => x"80ee3880",
          1478 => x"ef397784",
          1479 => x"19710856",
          1480 => x"59538074",
          1481 => x"33545572",
          1482 => x"752e8d38",
          1483 => x"81157015",
          1484 => x"70335154",
          1485 => x"5572f538",
          1486 => x"79812a56",
          1487 => x"90397481",
          1488 => x"16565372",
          1489 => x"7b278f38",
          1490 => x"a051fc90",
          1491 => x"3f758106",
          1492 => x"5372802e",
          1493 => x"e9387351",
          1494 => x"fcdf3f74",
          1495 => x"81165653",
          1496 => x"727b27fd",
          1497 => x"b038a051",
          1498 => x"fbf23fef",
          1499 => x"39778419",
          1500 => x"83123353",
          1501 => x"59539339",
          1502 => x"825c9539",
          1503 => x"885c9139",
          1504 => x"8a5c8d39",
          1505 => x"905c8939",
          1506 => x"7551fbd0",
          1507 => x"3ffd8639",
          1508 => x"79822a70",
          1509 => x"81065153",
          1510 => x"72802e88",
          1511 => x"38778419",
          1512 => x"59538639",
          1513 => x"84187854",
          1514 => x"58720874",
          1515 => x"80c43270",
          1516 => x"30707207",
          1517 => x"80255155",
          1518 => x"55557480",
          1519 => x"258d3872",
          1520 => x"802e8838",
          1521 => x"74307a90",
          1522 => x"075b5580",
          1523 => x"0b8f3d5e",
          1524 => x"577b5274",
          1525 => x"51e3d33f",
          1526 => x"81d3d808",
          1527 => x"81ff067c",
          1528 => x"53755254",
          1529 => x"e3913f81",
          1530 => x"d3d80855",
          1531 => x"89742792",
          1532 => x"38a71453",
          1533 => x"7580f82e",
          1534 => x"84388714",
          1535 => x"537281ff",
          1536 => x"0654b014",
          1537 => x"53727d70",
          1538 => x"81055f34",
          1539 => x"81177530",
          1540 => x"7077079f",
          1541 => x"2a515457",
          1542 => x"769f2685",
          1543 => x"3872ffb1",
          1544 => x"3879842a",
          1545 => x"70810651",
          1546 => x"5372802e",
          1547 => x"8e38963d",
          1548 => x"7705e005",
          1549 => x"53ad7334",
          1550 => x"81175776",
          1551 => x"7a810654",
          1552 => x"55b05472",
          1553 => x"8338a054",
          1554 => x"79812a70",
          1555 => x"81065456",
          1556 => x"729f3881",
          1557 => x"1755767b",
          1558 => x"27973873",
          1559 => x"51f9fd3f",
          1560 => x"75810653",
          1561 => x"728b3874",
          1562 => x"81165653",
          1563 => x"7a7326eb",
          1564 => x"38963d77",
          1565 => x"05e00553",
          1566 => x"ff17ff14",
          1567 => x"70335354",
          1568 => x"57f9d93f",
          1569 => x"76f23874",
          1570 => x"81165653",
          1571 => x"727b27fb",
          1572 => x"8438a051",
          1573 => x"f9c63fef",
          1574 => x"39963d0d",
          1575 => x"04fd3d0d",
          1576 => x"863d7070",
          1577 => x"84055208",
          1578 => x"55527351",
          1579 => x"fae03f85",
          1580 => x"3d0d04fe",
          1581 => x"3d0d7481",
          1582 => x"d3f00c85",
          1583 => x"3d880552",
          1584 => x"7551faca",
          1585 => x"3f81d3f0",
          1586 => x"08538073",
          1587 => x"34800b81",
          1588 => x"d3f00c84",
          1589 => x"3d0d04fd",
          1590 => x"3d0d81d3",
          1591 => x"e8087681",
          1592 => x"d3e80c87",
          1593 => x"3d880553",
          1594 => x"775253fa",
          1595 => x"a13f7281",
          1596 => x"d3e80c85",
          1597 => x"3d0d04fb",
          1598 => x"3d0d7779",
          1599 => x"81d3ec08",
          1600 => x"70565457",
          1601 => x"55805471",
          1602 => x"802e80e0",
          1603 => x"3881d3ec",
          1604 => x"0852712d",
          1605 => x"81d3d808",
          1606 => x"81ff0653",
          1607 => x"72802e80",
          1608 => x"cb38728d",
          1609 => x"2eb93872",
          1610 => x"88327030",
          1611 => x"70802551",
          1612 => x"51527380",
          1613 => x"2e8b3871",
          1614 => x"802e8638",
          1615 => x"ff145497",
          1616 => x"399f7325",
          1617 => x"c838ff16",
          1618 => x"52737225",
          1619 => x"c0387414",
          1620 => x"52727234",
          1621 => x"81145472",
          1622 => x"51f8813f",
          1623 => x"ffaf3973",
          1624 => x"15528072",
          1625 => x"348a51f7",
          1626 => x"f33f8153",
          1627 => x"7281d3d8",
          1628 => x"0c873d0d",
          1629 => x"04fe3d0d",
          1630 => x"81d3ec08",
          1631 => x"7581d3ec",
          1632 => x"0c775376",
          1633 => x"5253feef",
          1634 => x"3f7281d3",
          1635 => x"ec0c843d",
          1636 => x"0d04f83d",
          1637 => x"0d7a7c5a",
          1638 => x"5680707a",
          1639 => x"0c587508",
          1640 => x"70335553",
          1641 => x"73a02e09",
          1642 => x"81068738",
          1643 => x"8113760c",
          1644 => x"ed3973ad",
          1645 => x"2e098106",
          1646 => x"8e388176",
          1647 => x"0811770c",
          1648 => x"76087033",
          1649 => x"56545873",
          1650 => x"b02e0981",
          1651 => x"0680c238",
          1652 => x"75088105",
          1653 => x"760c7508",
          1654 => x"70335553",
          1655 => x"7380e22e",
          1656 => x"8b389057",
          1657 => x"7380f82e",
          1658 => x"85388f39",
          1659 => x"82578113",
          1660 => x"760c7508",
          1661 => x"70335553",
          1662 => x"ac398155",
          1663 => x"a0742780",
          1664 => x"fa38d014",
          1665 => x"53805588",
          1666 => x"57897327",
          1667 => x"983880eb",
          1668 => x"39d01453",
          1669 => x"80557289",
          1670 => x"2680e038",
          1671 => x"86398055",
          1672 => x"80d9398a",
          1673 => x"578055a0",
          1674 => x"742780c2",
          1675 => x"3880e074",
          1676 => x"278938e0",
          1677 => x"147081ff",
          1678 => x"065553d0",
          1679 => x"147081ff",
          1680 => x"06555390",
          1681 => x"74278e38",
          1682 => x"f9147081",
          1683 => x"ff065553",
          1684 => x"897427ca",
          1685 => x"38737727",
          1686 => x"c5387477",
          1687 => x"29147608",
          1688 => x"8105770c",
          1689 => x"76087033",
          1690 => x"565455ff",
          1691 => x"ba397780",
          1692 => x"2e843874",
          1693 => x"30557479",
          1694 => x"0c815574",
          1695 => x"81d3d80c",
          1696 => x"8a3d0d04",
          1697 => x"f83d0d7a",
          1698 => x"7c5a5680",
          1699 => x"707a0c58",
          1700 => x"75087033",
          1701 => x"555373a0",
          1702 => x"2e098106",
          1703 => x"87388113",
          1704 => x"760ced39",
          1705 => x"73ad2e09",
          1706 => x"81068e38",
          1707 => x"81760811",
          1708 => x"770c7608",
          1709 => x"70335654",
          1710 => x"5873b02e",
          1711 => x"09810680",
          1712 => x"c2387508",
          1713 => x"8105760c",
          1714 => x"75087033",
          1715 => x"55537380",
          1716 => x"e22e8b38",
          1717 => x"90577380",
          1718 => x"f82e8538",
          1719 => x"8f398257",
          1720 => x"8113760c",
          1721 => x"75087033",
          1722 => x"5553ac39",
          1723 => x"8155a074",
          1724 => x"2780fa38",
          1725 => x"d0145380",
          1726 => x"55885789",
          1727 => x"73279838",
          1728 => x"80eb39d0",
          1729 => x"14538055",
          1730 => x"72892680",
          1731 => x"e0388639",
          1732 => x"805580d9",
          1733 => x"398a5780",
          1734 => x"55a07427",
          1735 => x"80c23880",
          1736 => x"e0742789",
          1737 => x"38e01470",
          1738 => x"81ff0655",
          1739 => x"53d01470",
          1740 => x"81ff0655",
          1741 => x"53907427",
          1742 => x"8e38f914",
          1743 => x"7081ff06",
          1744 => x"55538974",
          1745 => x"27ca3873",
          1746 => x"7727c538",
          1747 => x"74772914",
          1748 => x"76088105",
          1749 => x"770c7608",
          1750 => x"70335654",
          1751 => x"55ffba39",
          1752 => x"77802e84",
          1753 => x"38743055",
          1754 => x"74790c81",
          1755 => x"557481d3",
          1756 => x"d80c8a3d",
          1757 => x"0d04ff3d",
          1758 => x"0d028f05",
          1759 => x"33518152",
          1760 => x"70722687",
          1761 => x"3881d1a0",
          1762 => x"11335271",
          1763 => x"81d3d80c",
          1764 => x"833d0d04",
          1765 => x"fc3d0d02",
          1766 => x"9b053302",
          1767 => x"84059f05",
          1768 => x"33565383",
          1769 => x"51728126",
          1770 => x"80e03872",
          1771 => x"842b87c0",
          1772 => x"928c1153",
          1773 => x"51885474",
          1774 => x"802e8438",
          1775 => x"81885473",
          1776 => x"720c87c0",
          1777 => x"928c1151",
          1778 => x"81710c85",
          1779 => x"0b87c098",
          1780 => x"8c0c7052",
          1781 => x"71087082",
          1782 => x"06515170",
          1783 => x"802e8a38",
          1784 => x"87c0988c",
          1785 => x"085170ec",
          1786 => x"387108fc",
          1787 => x"80800652",
          1788 => x"71923887",
          1789 => x"c0988c08",
          1790 => x"5170802e",
          1791 => x"87387181",
          1792 => x"d1a01434",
          1793 => x"81d1a013",
          1794 => x"33517081",
          1795 => x"d3d80c86",
          1796 => x"3d0d04f3",
          1797 => x"3d0d6062",
          1798 => x"64028c05",
          1799 => x"bf053357",
          1800 => x"40585b83",
          1801 => x"74525afe",
          1802 => x"cd3f81d3",
          1803 => x"d8088106",
          1804 => x"7a545271",
          1805 => x"81be3871",
          1806 => x"7275842b",
          1807 => x"87c09280",
          1808 => x"1187c092",
          1809 => x"8c1287c0",
          1810 => x"92841341",
          1811 => x"5a40575a",
          1812 => x"58850b87",
          1813 => x"c0988c0c",
          1814 => x"767d0c84",
          1815 => x"760c7508",
          1816 => x"70852a70",
          1817 => x"81065153",
          1818 => x"5471802e",
          1819 => x"8e387b08",
          1820 => x"52717b70",
          1821 => x"81055d34",
          1822 => x"81195980",
          1823 => x"74a20653",
          1824 => x"5371732e",
          1825 => x"83388153",
          1826 => x"7883ff26",
          1827 => x"8f387280",
          1828 => x"2e8a3887",
          1829 => x"c0988c08",
          1830 => x"5271c338",
          1831 => x"87c0988c",
          1832 => x"08527180",
          1833 => x"2e873878",
          1834 => x"84802e99",
          1835 => x"3881760c",
          1836 => x"87c0928c",
          1837 => x"15537208",
          1838 => x"70820651",
          1839 => x"5271f738",
          1840 => x"ff1a5a8d",
          1841 => x"39848017",
          1842 => x"81197081",
          1843 => x"ff065a53",
          1844 => x"5779802e",
          1845 => x"903873fc",
          1846 => x"80800652",
          1847 => x"7187387d",
          1848 => x"7826feed",
          1849 => x"3873fc80",
          1850 => x"80065271",
          1851 => x"802e8338",
          1852 => x"81527153",
          1853 => x"7281d3d8",
          1854 => x"0c8f3d0d",
          1855 => x"04f33d0d",
          1856 => x"60626402",
          1857 => x"8c05bf05",
          1858 => x"33574058",
          1859 => x"5b835980",
          1860 => x"745258fc",
          1861 => x"e13f81d3",
          1862 => x"d8088106",
          1863 => x"79545271",
          1864 => x"782e0981",
          1865 => x"0681b138",
          1866 => x"7774842b",
          1867 => x"87c09280",
          1868 => x"1187c092",
          1869 => x"8c1287c0",
          1870 => x"92841340",
          1871 => x"595f565a",
          1872 => x"850b87c0",
          1873 => x"988c0c76",
          1874 => x"7d0c8276",
          1875 => x"0c805875",
          1876 => x"0870842a",
          1877 => x"70810651",
          1878 => x"53547180",
          1879 => x"2e8c387a",
          1880 => x"7081055c",
          1881 => x"337c0c81",
          1882 => x"18587381",
          1883 => x"2a708106",
          1884 => x"51527180",
          1885 => x"2e8a3887",
          1886 => x"c0988c08",
          1887 => x"5271d038",
          1888 => x"87c0988c",
          1889 => x"08527180",
          1890 => x"2e873877",
          1891 => x"84802e99",
          1892 => x"3881760c",
          1893 => x"87c0928c",
          1894 => x"15537208",
          1895 => x"70820651",
          1896 => x"5271f738",
          1897 => x"ff19598d",
          1898 => x"39811a70",
          1899 => x"81ff0684",
          1900 => x"8019595b",
          1901 => x"5278802e",
          1902 => x"903873fc",
          1903 => x"80800652",
          1904 => x"7187387d",
          1905 => x"7a26fef8",
          1906 => x"3873fc80",
          1907 => x"80065271",
          1908 => x"802e8338",
          1909 => x"81527153",
          1910 => x"7281d3d8",
          1911 => x"0c8f3d0d",
          1912 => x"04f63d0d",
          1913 => x"7e028405",
          1914 => x"b3053302",
          1915 => x"8805b705",
          1916 => x"33715454",
          1917 => x"5657fafe",
          1918 => x"3f81d3d8",
          1919 => x"08810653",
          1920 => x"83547280",
          1921 => x"fe38850b",
          1922 => x"87c0988c",
          1923 => x"0c815671",
          1924 => x"762e80dc",
          1925 => x"38717624",
          1926 => x"93387484",
          1927 => x"2b87c092",
          1928 => x"8c115454",
          1929 => x"71802e8d",
          1930 => x"3880d439",
          1931 => x"71832e80",
          1932 => x"c63880cb",
          1933 => x"39720870",
          1934 => x"812a7081",
          1935 => x"06515152",
          1936 => x"71802e8a",
          1937 => x"3887c098",
          1938 => x"8c085271",
          1939 => x"e83887c0",
          1940 => x"988c0852",
          1941 => x"71963881",
          1942 => x"730c87c0",
          1943 => x"928c1453",
          1944 => x"72087082",
          1945 => x"06515271",
          1946 => x"f7389639",
          1947 => x"80569239",
          1948 => x"88800a77",
          1949 => x"0c853981",
          1950 => x"80770c72",
          1951 => x"56833984",
          1952 => x"56755473",
          1953 => x"81d3d80c",
          1954 => x"8c3d0d04",
          1955 => x"fe3d0d74",
          1956 => x"81113371",
          1957 => x"3371882b",
          1958 => x"0781d3d8",
          1959 => x"0c535184",
          1960 => x"3d0d04fd",
          1961 => x"3d0d7583",
          1962 => x"11338212",
          1963 => x"3371902b",
          1964 => x"71882b07",
          1965 => x"81143370",
          1966 => x"7207882b",
          1967 => x"75337107",
          1968 => x"81d3d80c",
          1969 => x"52535456",
          1970 => x"5452853d",
          1971 => x"0d04ff3d",
          1972 => x"0d730284",
          1973 => x"05920522",
          1974 => x"52527072",
          1975 => x"70810554",
          1976 => x"3470882a",
          1977 => x"51707234",
          1978 => x"833d0d04",
          1979 => x"ff3d0d73",
          1980 => x"75525270",
          1981 => x"72708105",
          1982 => x"54347088",
          1983 => x"2a517072",
          1984 => x"70810554",
          1985 => x"3470882a",
          1986 => x"51707270",
          1987 => x"81055434",
          1988 => x"70882a51",
          1989 => x"70723483",
          1990 => x"3d0d04fe",
          1991 => x"3d0d7675",
          1992 => x"77545451",
          1993 => x"70802e92",
          1994 => x"38717081",
          1995 => x"05533373",
          1996 => x"70810555",
          1997 => x"34ff1151",
          1998 => x"eb39843d",
          1999 => x"0d04fe3d",
          2000 => x"0d757776",
          2001 => x"54525372",
          2002 => x"72708105",
          2003 => x"5434ff11",
          2004 => x"5170f438",
          2005 => x"843d0d04",
          2006 => x"fc3d0d78",
          2007 => x"77795656",
          2008 => x"53747081",
          2009 => x"05563374",
          2010 => x"70810556",
          2011 => x"33717131",
          2012 => x"ff165652",
          2013 => x"52527280",
          2014 => x"2e863871",
          2015 => x"802ee238",
          2016 => x"7181d3d8",
          2017 => x"0c863d0d",
          2018 => x"04fe3d0d",
          2019 => x"74765451",
          2020 => x"89397173",
          2021 => x"2e8a3881",
          2022 => x"11517033",
          2023 => x"5271f338",
          2024 => x"703381d3",
          2025 => x"d80c843d",
          2026 => x"0d04800b",
          2027 => x"81d3d80c",
          2028 => x"04800b81",
          2029 => x"d3d80c04",
          2030 => x"f73d0d7b",
          2031 => x"56800b83",
          2032 => x"1733565a",
          2033 => x"747a2e80",
          2034 => x"d6388154",
          2035 => x"b0160853",
          2036 => x"b4167053",
          2037 => x"81173352",
          2038 => x"59faa23f",
          2039 => x"81d3d808",
          2040 => x"7a2e0981",
          2041 => x"06b73881",
          2042 => x"d3d80883",
          2043 => x"1734b016",
          2044 => x"0870a418",
          2045 => x"08319c18",
          2046 => x"08595658",
          2047 => x"7477279f",
          2048 => x"38821633",
          2049 => x"5574822e",
          2050 => x"09810693",
          2051 => x"38815476",
          2052 => x"18537852",
          2053 => x"81163351",
          2054 => x"f9e33f83",
          2055 => x"39815a79",
          2056 => x"81d3d80c",
          2057 => x"8b3d0d04",
          2058 => x"fa3d0d78",
          2059 => x"7a565680",
          2060 => x"5774b017",
          2061 => x"082eaf38",
          2062 => x"7551fefc",
          2063 => x"3f81d3d8",
          2064 => x"085781d3",
          2065 => x"d8089f38",
          2066 => x"81547453",
          2067 => x"b4165281",
          2068 => x"163351f7",
          2069 => x"be3f81d3",
          2070 => x"d808802e",
          2071 => x"8538ff55",
          2072 => x"815774b0",
          2073 => x"170c7681",
          2074 => x"d3d80c88",
          2075 => x"3d0d04f8",
          2076 => x"3d0d7a70",
          2077 => x"5257fec0",
          2078 => x"3f81d3d8",
          2079 => x"085881d3",
          2080 => x"d8088191",
          2081 => x"38763355",
          2082 => x"74832e09",
          2083 => x"810680f0",
          2084 => x"38841733",
          2085 => x"5978812e",
          2086 => x"09810680",
          2087 => x"e3388480",
          2088 => x"5381d3d8",
          2089 => x"0852b417",
          2090 => x"705256fd",
          2091 => x"913f82d4",
          2092 => x"d55284b2",
          2093 => x"1751fc96",
          2094 => x"3f848b85",
          2095 => x"a4d25275",
          2096 => x"51fca93f",
          2097 => x"868a85e4",
          2098 => x"f2528498",
          2099 => x"1751fc9c",
          2100 => x"3f901708",
          2101 => x"52849c17",
          2102 => x"51fc913f",
          2103 => x"8c170852",
          2104 => x"84a01751",
          2105 => x"fc863fa0",
          2106 => x"17088105",
          2107 => x"70b0190c",
          2108 => x"79555375",
          2109 => x"52811733",
          2110 => x"51f8823f",
          2111 => x"77841834",
          2112 => x"80538052",
          2113 => x"81173351",
          2114 => x"f9d73f81",
          2115 => x"d3d80880",
          2116 => x"2e833881",
          2117 => x"587781d3",
          2118 => x"d80c8a3d",
          2119 => x"0d04fb3d",
          2120 => x"0d77fe1a",
          2121 => x"981208fe",
          2122 => x"05555654",
          2123 => x"80567473",
          2124 => x"278d388a",
          2125 => x"14227571",
          2126 => x"29ac1608",
          2127 => x"05575375",
          2128 => x"81d3d80c",
          2129 => x"873d0d04",
          2130 => x"f93d0d7a",
          2131 => x"7a700856",
          2132 => x"54578177",
          2133 => x"2781df38",
          2134 => x"76981508",
          2135 => x"2781d738",
          2136 => x"ff743354",
          2137 => x"5872822e",
          2138 => x"80f53872",
          2139 => x"82248938",
          2140 => x"72812e8d",
          2141 => x"3881bf39",
          2142 => x"72832e81",
          2143 => x"8e3881b6",
          2144 => x"3976812a",
          2145 => x"1770892a",
          2146 => x"a4160805",
          2147 => x"53745255",
          2148 => x"fd963f81",
          2149 => x"d3d80881",
          2150 => x"9f387483",
          2151 => x"ff0614b4",
          2152 => x"11338117",
          2153 => x"70892aa4",
          2154 => x"18080555",
          2155 => x"76545757",
          2156 => x"53fcf53f",
          2157 => x"81d3d808",
          2158 => x"80fe3874",
          2159 => x"83ff0614",
          2160 => x"b4113370",
          2161 => x"882b7807",
          2162 => x"79810671",
          2163 => x"842a5c52",
          2164 => x"58515372",
          2165 => x"80e23875",
          2166 => x"9fff0658",
          2167 => x"80da3976",
          2168 => x"882aa415",
          2169 => x"08055273",
          2170 => x"51fcbd3f",
          2171 => x"81d3d808",
          2172 => x"80c63876",
          2173 => x"1083fe06",
          2174 => x"7405b405",
          2175 => x"51f98d3f",
          2176 => x"81d3d808",
          2177 => x"83ffff06",
          2178 => x"58ae3976",
          2179 => x"872aa415",
          2180 => x"08055273",
          2181 => x"51fc913f",
          2182 => x"81d3d808",
          2183 => x"9b387682",
          2184 => x"2b83fc06",
          2185 => x"7405b405",
          2186 => x"51f8f83f",
          2187 => x"81d3d808",
          2188 => x"f00a0658",
          2189 => x"83398158",
          2190 => x"7781d3d8",
          2191 => x"0c893d0d",
          2192 => x"04f83d0d",
          2193 => x"7a7c7e5a",
          2194 => x"58568259",
          2195 => x"81772782",
          2196 => x"9e387698",
          2197 => x"17082782",
          2198 => x"96387533",
          2199 => x"5372792e",
          2200 => x"819d3872",
          2201 => x"79248938",
          2202 => x"72812e8d",
          2203 => x"38828039",
          2204 => x"72832e81",
          2205 => x"b83881f7",
          2206 => x"3976812a",
          2207 => x"1770892a",
          2208 => x"a4180805",
          2209 => x"53765255",
          2210 => x"fb9e3f81",
          2211 => x"d3d80859",
          2212 => x"81d3d808",
          2213 => x"81d93874",
          2214 => x"83ff0616",
          2215 => x"b4058116",
          2216 => x"78810659",
          2217 => x"56547753",
          2218 => x"76802e8f",
          2219 => x"3877842b",
          2220 => x"9ff00674",
          2221 => x"338f0671",
          2222 => x"07515372",
          2223 => x"7434810b",
          2224 => x"83173474",
          2225 => x"892aa417",
          2226 => x"08055275",
          2227 => x"51fad93f",
          2228 => x"81d3d808",
          2229 => x"5981d3d8",
          2230 => x"08819438",
          2231 => x"7483ff06",
          2232 => x"16b40578",
          2233 => x"842a5454",
          2234 => x"768f3877",
          2235 => x"882a7433",
          2236 => x"81f00671",
          2237 => x"8f060751",
          2238 => x"53727434",
          2239 => x"80ec3976",
          2240 => x"882aa417",
          2241 => x"08055275",
          2242 => x"51fa9d3f",
          2243 => x"81d3d808",
          2244 => x"5981d3d8",
          2245 => x"0880d838",
          2246 => x"7783ffff",
          2247 => x"06527610",
          2248 => x"83fe0676",
          2249 => x"05b40551",
          2250 => x"f7a43fbe",
          2251 => x"3976872a",
          2252 => x"a4170805",
          2253 => x"527551f9",
          2254 => x"ef3f81d3",
          2255 => x"d8085981",
          2256 => x"d3d808ab",
          2257 => x"3877f00a",
          2258 => x"0677822b",
          2259 => x"83fc0670",
          2260 => x"18b40570",
          2261 => x"54515454",
          2262 => x"f6c93f81",
          2263 => x"d3d8088f",
          2264 => x"0a067407",
          2265 => x"527251f7",
          2266 => x"833f810b",
          2267 => x"83173478",
          2268 => x"81d3d80c",
          2269 => x"8a3d0d04",
          2270 => x"f83d0d7a",
          2271 => x"7c7e7208",
          2272 => x"59565659",
          2273 => x"817527a4",
          2274 => x"38749817",
          2275 => x"08279d38",
          2276 => x"73802eaa",
          2277 => x"38ff5373",
          2278 => x"527551fd",
          2279 => x"a43f81d3",
          2280 => x"d8085481",
          2281 => x"d3d80880",
          2282 => x"f2389339",
          2283 => x"825480eb",
          2284 => x"39815480",
          2285 => x"e63981d3",
          2286 => x"d8085480",
          2287 => x"de397452",
          2288 => x"7851fb84",
          2289 => x"3f81d3d8",
          2290 => x"085881d3",
          2291 => x"d808802e",
          2292 => x"80c73881",
          2293 => x"d3d80881",
          2294 => x"2ed23881",
          2295 => x"d3d808ff",
          2296 => x"2ecf3880",
          2297 => x"53745275",
          2298 => x"51fcd63f",
          2299 => x"81d3d808",
          2300 => x"c5389816",
          2301 => x"08fe1190",
          2302 => x"18085755",
          2303 => x"57747427",
          2304 => x"90388115",
          2305 => x"90170c84",
          2306 => x"16338107",
          2307 => x"54738417",
          2308 => x"34775576",
          2309 => x"7826ffa6",
          2310 => x"38805473",
          2311 => x"81d3d80c",
          2312 => x"8a3d0d04",
          2313 => x"f63d0d7c",
          2314 => x"7e710859",
          2315 => x"5b5b7995",
          2316 => x"388c1708",
          2317 => x"5877802e",
          2318 => x"88389817",
          2319 => x"087826b2",
          2320 => x"388158ae",
          2321 => x"3979527a",
          2322 => x"51f9fd3f",
          2323 => x"81557481",
          2324 => x"d3d80827",
          2325 => x"82e03881",
          2326 => x"d3d80855",
          2327 => x"81d3d808",
          2328 => x"ff2e82d2",
          2329 => x"38981708",
          2330 => x"81d3d808",
          2331 => x"2682c738",
          2332 => x"79589017",
          2333 => x"08705654",
          2334 => x"73802e82",
          2335 => x"b938777a",
          2336 => x"2e098106",
          2337 => x"80e23881",
          2338 => x"1a569817",
          2339 => x"08762683",
          2340 => x"38825675",
          2341 => x"527a51f9",
          2342 => x"af3f8059",
          2343 => x"81d3d808",
          2344 => x"812e0981",
          2345 => x"06863881",
          2346 => x"d3d80859",
          2347 => x"81d3d808",
          2348 => x"09703070",
          2349 => x"72078025",
          2350 => x"707c0781",
          2351 => x"d3d80854",
          2352 => x"51515555",
          2353 => x"7381ef38",
          2354 => x"81d3d808",
          2355 => x"802e9538",
          2356 => x"8c170854",
          2357 => x"81742790",
          2358 => x"38739818",
          2359 => x"08278938",
          2360 => x"73588539",
          2361 => x"7580db38",
          2362 => x"77568116",
          2363 => x"56981708",
          2364 => x"76268938",
          2365 => x"82567578",
          2366 => x"2681ac38",
          2367 => x"75527a51",
          2368 => x"f8c63f81",
          2369 => x"d3d80880",
          2370 => x"2eb83880",
          2371 => x"5981d3d8",
          2372 => x"08812e09",
          2373 => x"81068638",
          2374 => x"81d3d808",
          2375 => x"5981d3d8",
          2376 => x"08097030",
          2377 => x"70720780",
          2378 => x"25707c07",
          2379 => x"51515555",
          2380 => x"7380f838",
          2381 => x"75782e09",
          2382 => x"8106ffae",
          2383 => x"38735580",
          2384 => x"f539ff53",
          2385 => x"75527651",
          2386 => x"f9f73f81",
          2387 => x"d3d80881",
          2388 => x"d3d80830",
          2389 => x"7081d3d8",
          2390 => x"08078025",
          2391 => x"51555579",
          2392 => x"802e9438",
          2393 => x"73802e8f",
          2394 => x"38755379",
          2395 => x"527651f9",
          2396 => x"d03f81d3",
          2397 => x"d8085574",
          2398 => x"a538758c",
          2399 => x"180c9817",
          2400 => x"08fe0590",
          2401 => x"18085654",
          2402 => x"74742686",
          2403 => x"38ff1590",
          2404 => x"180c8417",
          2405 => x"33810754",
          2406 => x"73841834",
          2407 => x"9739ff56",
          2408 => x"74812e90",
          2409 => x"388c3980",
          2410 => x"558c3981",
          2411 => x"d3d80855",
          2412 => x"85398156",
          2413 => x"75557481",
          2414 => x"d3d80c8c",
          2415 => x"3d0d04f8",
          2416 => x"3d0d7a70",
          2417 => x"5255f3f0",
          2418 => x"3f81d3d8",
          2419 => x"08588156",
          2420 => x"81d3d808",
          2421 => x"80d8387b",
          2422 => x"527451f6",
          2423 => x"c13f81d3",
          2424 => x"d80881d3",
          2425 => x"d808b017",
          2426 => x"0c598480",
          2427 => x"537752b4",
          2428 => x"15705257",
          2429 => x"f2c83f77",
          2430 => x"56843981",
          2431 => x"16568a15",
          2432 => x"22587578",
          2433 => x"27973881",
          2434 => x"54751953",
          2435 => x"76528115",
          2436 => x"3351ede9",
          2437 => x"3f81d3d8",
          2438 => x"08802edf",
          2439 => x"388a1522",
          2440 => x"76327030",
          2441 => x"70720770",
          2442 => x"9f2a5351",
          2443 => x"56567581",
          2444 => x"d3d80c8a",
          2445 => x"3d0d04f8",
          2446 => x"3d0d7a7c",
          2447 => x"71085856",
          2448 => x"5774f080",
          2449 => x"0a2680f1",
          2450 => x"38749f06",
          2451 => x"537280e9",
          2452 => x"38749018",
          2453 => x"0c881708",
          2454 => x"5473aa38",
          2455 => x"75335382",
          2456 => x"73278838",
          2457 => x"a8160854",
          2458 => x"739b3874",
          2459 => x"852a5382",
          2460 => x"0b881722",
          2461 => x"5a587279",
          2462 => x"2780fe38",
          2463 => x"a8160898",
          2464 => x"180c80cd",
          2465 => x"398a1622",
          2466 => x"70892b54",
          2467 => x"58727526",
          2468 => x"b2387352",
          2469 => x"7651f5b0",
          2470 => x"3f81d3d8",
          2471 => x"085481d3",
          2472 => x"d808ff2e",
          2473 => x"bd38810b",
          2474 => x"81d3d808",
          2475 => x"278b3898",
          2476 => x"160881d3",
          2477 => x"d8082685",
          2478 => x"388258bd",
          2479 => x"39747331",
          2480 => x"55cb3973",
          2481 => x"527551f4",
          2482 => x"d53f81d3",
          2483 => x"d8089818",
          2484 => x"0c739418",
          2485 => x"0c981708",
          2486 => x"53825872",
          2487 => x"802e9a38",
          2488 => x"85398158",
          2489 => x"94397489",
          2490 => x"2a139818",
          2491 => x"0c7483ff",
          2492 => x"0616b405",
          2493 => x"9c180c80",
          2494 => x"587781d3",
          2495 => x"d80c8a3d",
          2496 => x"0d04f83d",
          2497 => x"0d7a7008",
          2498 => x"901208a0",
          2499 => x"05595754",
          2500 => x"f0800a77",
          2501 => x"27863880",
          2502 => x"0b98150c",
          2503 => x"98140853",
          2504 => x"84557280",
          2505 => x"2e81cb38",
          2506 => x"7683ff06",
          2507 => x"587781b5",
          2508 => x"38811398",
          2509 => x"150c9414",
          2510 => x"08557492",
          2511 => x"3876852a",
          2512 => x"88172256",
          2513 => x"53747326",
          2514 => x"819b3880",
          2515 => x"c0398a16",
          2516 => x"22ff0577",
          2517 => x"892a0653",
          2518 => x"72818a38",
          2519 => x"74527351",
          2520 => x"f3e63f81",
          2521 => x"d3d80853",
          2522 => x"8255810b",
          2523 => x"81d3d808",
          2524 => x"2780ff38",
          2525 => x"815581d3",
          2526 => x"d808ff2e",
          2527 => x"80f43898",
          2528 => x"160881d3",
          2529 => x"d8082680",
          2530 => x"ca387b8a",
          2531 => x"38779815",
          2532 => x"0c845580",
          2533 => x"dd399414",
          2534 => x"08527351",
          2535 => x"f9863f81",
          2536 => x"d3d80853",
          2537 => x"875581d3",
          2538 => x"d808802e",
          2539 => x"80c43882",
          2540 => x"5581d3d8",
          2541 => x"08812eba",
          2542 => x"38815581",
          2543 => x"d3d808ff",
          2544 => x"2eb03881",
          2545 => x"d3d80852",
          2546 => x"7551fbf3",
          2547 => x"3f81d3d8",
          2548 => x"08a03872",
          2549 => x"94150c72",
          2550 => x"527551f2",
          2551 => x"c13f81d3",
          2552 => x"d8089815",
          2553 => x"0c769015",
          2554 => x"0c7716b4",
          2555 => x"059c150c",
          2556 => x"80557481",
          2557 => x"d3d80c8a",
          2558 => x"3d0d04f7",
          2559 => x"3d0d7b7d",
          2560 => x"71085b5b",
          2561 => x"57805276",
          2562 => x"51fcac3f",
          2563 => x"81d3d808",
          2564 => x"5481d3d8",
          2565 => x"0880ec38",
          2566 => x"81d3d808",
          2567 => x"56981708",
          2568 => x"527851f0",
          2569 => x"833f81d3",
          2570 => x"d8085481",
          2571 => x"d3d80880",
          2572 => x"d23881d3",
          2573 => x"d8089c18",
          2574 => x"08703351",
          2575 => x"54587281",
          2576 => x"e52e0981",
          2577 => x"06833881",
          2578 => x"5881d3d8",
          2579 => x"08557283",
          2580 => x"38815577",
          2581 => x"75075372",
          2582 => x"802e8e38",
          2583 => x"81165675",
          2584 => x"7a2e0981",
          2585 => x"068838a5",
          2586 => x"3981d3d8",
          2587 => x"08568152",
          2588 => x"7651fd8e",
          2589 => x"3f81d3d8",
          2590 => x"085481d3",
          2591 => x"d808802e",
          2592 => x"ff9b3873",
          2593 => x"842e0981",
          2594 => x"06833887",
          2595 => x"547381d3",
          2596 => x"d80c8b3d",
          2597 => x"0d04fd3d",
          2598 => x"0d769a11",
          2599 => x"5254ebec",
          2600 => x"3f81d3d8",
          2601 => x"0883ffff",
          2602 => x"06767033",
          2603 => x"51535371",
          2604 => x"832e0981",
          2605 => x"06903894",
          2606 => x"1451ebd0",
          2607 => x"3f81d3d8",
          2608 => x"08902b73",
          2609 => x"07537281",
          2610 => x"d3d80c85",
          2611 => x"3d0d04fc",
          2612 => x"3d0d7779",
          2613 => x"7083ffff",
          2614 => x"06549a12",
          2615 => x"535555eb",
          2616 => x"ed3f7670",
          2617 => x"33515372",
          2618 => x"832e0981",
          2619 => x"068b3873",
          2620 => x"902a5294",
          2621 => x"1551ebd6",
          2622 => x"3f863d0d",
          2623 => x"04f73d0d",
          2624 => x"7b7d5b55",
          2625 => x"8475085a",
          2626 => x"58981508",
          2627 => x"802e818a",
          2628 => x"38981508",
          2629 => x"527851ee",
          2630 => x"8f3f81d3",
          2631 => x"d8085881",
          2632 => x"d3d80880",
          2633 => x"f5389c15",
          2634 => x"08703355",
          2635 => x"53738638",
          2636 => x"845880e6",
          2637 => x"398b1333",
          2638 => x"70bf0670",
          2639 => x"81ff0658",
          2640 => x"51537286",
          2641 => x"163481d3",
          2642 => x"d8085373",
          2643 => x"81e52e83",
          2644 => x"38815373",
          2645 => x"ae2ea938",
          2646 => x"81707406",
          2647 => x"54577280",
          2648 => x"2e9e3875",
          2649 => x"8f2e9938",
          2650 => x"81d3d808",
          2651 => x"76df0654",
          2652 => x"5472882e",
          2653 => x"09810683",
          2654 => x"38765473",
          2655 => x"7a2ea038",
          2656 => x"80527451",
          2657 => x"fafc3f81",
          2658 => x"d3d80858",
          2659 => x"81d3d808",
          2660 => x"89389815",
          2661 => x"08fefa38",
          2662 => x"8639800b",
          2663 => x"98160c77",
          2664 => x"81d3d80c",
          2665 => x"8b3d0d04",
          2666 => x"fb3d0d77",
          2667 => x"70085754",
          2668 => x"81527351",
          2669 => x"fcc53f81",
          2670 => x"d3d80855",
          2671 => x"81d3d808",
          2672 => x"b4389814",
          2673 => x"08527551",
          2674 => x"ecde3f81",
          2675 => x"d3d80855",
          2676 => x"81d3d808",
          2677 => x"a038a053",
          2678 => x"81d3d808",
          2679 => x"529c1408",
          2680 => x"51eadb3f",
          2681 => x"8b53a014",
          2682 => x"529c1408",
          2683 => x"51eaac3f",
          2684 => x"810b8317",
          2685 => x"347481d3",
          2686 => x"d80c873d",
          2687 => x"0d04fd3d",
          2688 => x"0d757008",
          2689 => x"98120854",
          2690 => x"70535553",
          2691 => x"ec9a3f81",
          2692 => x"d3d8088d",
          2693 => x"389c1308",
          2694 => x"53e57334",
          2695 => x"810b8315",
          2696 => x"34853d0d",
          2697 => x"04fa3d0d",
          2698 => x"787a5757",
          2699 => x"800b8917",
          2700 => x"34981708",
          2701 => x"802e8182",
          2702 => x"38807089",
          2703 => x"18555555",
          2704 => x"9c170814",
          2705 => x"70338116",
          2706 => x"56515271",
          2707 => x"a02ea838",
          2708 => x"71852e09",
          2709 => x"81068438",
          2710 => x"81e55273",
          2711 => x"892e0981",
          2712 => x"068b38ae",
          2713 => x"73708105",
          2714 => x"55348115",
          2715 => x"55717370",
          2716 => x"81055534",
          2717 => x"8115558a",
          2718 => x"7427c538",
          2719 => x"75158805",
          2720 => x"52800b81",
          2721 => x"13349c17",
          2722 => x"08528b12",
          2723 => x"33881734",
          2724 => x"9c17089c",
          2725 => x"115252e8",
          2726 => x"8a3f81d3",
          2727 => x"d808760c",
          2728 => x"961251e7",
          2729 => x"e73f81d3",
          2730 => x"d8088617",
          2731 => x"23981251",
          2732 => x"e7da3f81",
          2733 => x"d3d80884",
          2734 => x"1723883d",
          2735 => x"0d04f33d",
          2736 => x"0d7f7008",
          2737 => x"5e5b8061",
          2738 => x"70335155",
          2739 => x"5573af2e",
          2740 => x"83388155",
          2741 => x"7380dc2e",
          2742 => x"91387480",
          2743 => x"2e8c3894",
          2744 => x"1d08881c",
          2745 => x"0caa3981",
          2746 => x"15418061",
          2747 => x"70335656",
          2748 => x"5673af2e",
          2749 => x"09810683",
          2750 => x"38815673",
          2751 => x"80dc3270",
          2752 => x"30708025",
          2753 => x"78075151",
          2754 => x"5473dc38",
          2755 => x"73881c0c",
          2756 => x"60703351",
          2757 => x"54739f26",
          2758 => x"9638ff80",
          2759 => x"0bab1c34",
          2760 => x"80527a51",
          2761 => x"f6913f81",
          2762 => x"d3d80855",
          2763 => x"85983991",
          2764 => x"3d61a01d",
          2765 => x"5c5a5e8b",
          2766 => x"53a05279",
          2767 => x"51e7ff3f",
          2768 => x"80705957",
          2769 => x"88793355",
          2770 => x"5c73ae2e",
          2771 => x"09810680",
          2772 => x"d4387818",
          2773 => x"7033811a",
          2774 => x"71ae3270",
          2775 => x"30709f2a",
          2776 => x"73822607",
          2777 => x"5151535a",
          2778 => x"5754738c",
          2779 => x"38791754",
          2780 => x"75743481",
          2781 => x"1757db39",
          2782 => x"75af3270",
          2783 => x"30709f2a",
          2784 => x"51515475",
          2785 => x"80dc2e8c",
          2786 => x"3873802e",
          2787 => x"873875a0",
          2788 => x"2682bd38",
          2789 => x"77197e0c",
          2790 => x"a454a076",
          2791 => x"2782bd38",
          2792 => x"a05482b8",
          2793 => x"39781870",
          2794 => x"33811a5a",
          2795 => x"5754a076",
          2796 => x"2781fc38",
          2797 => x"75af3270",
          2798 => x"307780dc",
          2799 => x"32703072",
          2800 => x"80257180",
          2801 => x"25075151",
          2802 => x"56515573",
          2803 => x"802eac38",
          2804 => x"84398118",
          2805 => x"5880781a",
          2806 => x"70335155",
          2807 => x"5573af2e",
          2808 => x"09810683",
          2809 => x"38815573",
          2810 => x"80dc3270",
          2811 => x"30708025",
          2812 => x"77075151",
          2813 => x"5473db38",
          2814 => x"81b53975",
          2815 => x"ae2e0981",
          2816 => x"06833881",
          2817 => x"54767c27",
          2818 => x"74075473",
          2819 => x"802ea238",
          2820 => x"7b8b3270",
          2821 => x"3077ae32",
          2822 => x"70307280",
          2823 => x"25719f2a",
          2824 => x"07535156",
          2825 => x"51557481",
          2826 => x"a7388857",
          2827 => x"8b5cfef5",
          2828 => x"3975982b",
          2829 => x"54738025",
          2830 => x"8c387580",
          2831 => x"ff0681c3",
          2832 => x"dc113357",
          2833 => x"547551e6",
          2834 => x"e13f81d3",
          2835 => x"d808802e",
          2836 => x"b2387818",
          2837 => x"7033811a",
          2838 => x"71545a56",
          2839 => x"54e6d23f",
          2840 => x"81d3d808",
          2841 => x"802e80e8",
          2842 => x"38ff1c54",
          2843 => x"76742780",
          2844 => x"df387917",
          2845 => x"54757434",
          2846 => x"81177a11",
          2847 => x"55577474",
          2848 => x"34a73975",
          2849 => x"5281c2fc",
          2850 => x"51e5fe3f",
          2851 => x"81d3d808",
          2852 => x"bf38ff9f",
          2853 => x"16547399",
          2854 => x"268938e0",
          2855 => x"167081ff",
          2856 => x"06575479",
          2857 => x"17547574",
          2858 => x"34811757",
          2859 => x"fdf73977",
          2860 => x"197e0c76",
          2861 => x"802e9938",
          2862 => x"79335473",
          2863 => x"81e52e09",
          2864 => x"81068438",
          2865 => x"857a3484",
          2866 => x"54a07627",
          2867 => x"8f388b39",
          2868 => x"865581f2",
          2869 => x"39845680",
          2870 => x"f3398054",
          2871 => x"738b1b34",
          2872 => x"807b0858",
          2873 => x"527a51f2",
          2874 => x"ce3f81d3",
          2875 => x"d8085681",
          2876 => x"d3d80880",
          2877 => x"d738981b",
          2878 => x"08527651",
          2879 => x"e6aa3f81",
          2880 => x"d3d80856",
          2881 => x"81d3d808",
          2882 => x"80c2389c",
          2883 => x"1b087033",
          2884 => x"55557380",
          2885 => x"2effbe38",
          2886 => x"8b1533bf",
          2887 => x"06547386",
          2888 => x"1c348b15",
          2889 => x"3370832a",
          2890 => x"70810651",
          2891 => x"55587392",
          2892 => x"388b5379",
          2893 => x"527451e4",
          2894 => x"9f3f81d3",
          2895 => x"d808802e",
          2896 => x"8b387552",
          2897 => x"7a51f3ba",
          2898 => x"3fff9f39",
          2899 => x"75ab1c33",
          2900 => x"57557480",
          2901 => x"2ebb3874",
          2902 => x"842e0981",
          2903 => x"0680e738",
          2904 => x"75852a70",
          2905 => x"81067782",
          2906 => x"2a585154",
          2907 => x"73802e96",
          2908 => x"38758106",
          2909 => x"5473802e",
          2910 => x"fbb538ff",
          2911 => x"800bab1c",
          2912 => x"34805580",
          2913 => x"c1397581",
          2914 => x"065473ba",
          2915 => x"388555b6",
          2916 => x"3975822a",
          2917 => x"70810651",
          2918 => x"5473ab38",
          2919 => x"861b3370",
          2920 => x"842a7081",
          2921 => x"06515555",
          2922 => x"73802ee1",
          2923 => x"38901b08",
          2924 => x"83ff061d",
          2925 => x"b405527c",
          2926 => x"51f5db3f",
          2927 => x"81d3d808",
          2928 => x"881c0cfa",
          2929 => x"ea397481",
          2930 => x"d3d80c8f",
          2931 => x"3d0d04f6",
          2932 => x"3d0d7c5b",
          2933 => x"ff7b0870",
          2934 => x"71735559",
          2935 => x"5c555973",
          2936 => x"802e81c6",
          2937 => x"38757081",
          2938 => x"05573370",
          2939 => x"a0265252",
          2940 => x"71ba2e8d",
          2941 => x"3870ee38",
          2942 => x"71ba2e09",
          2943 => x"810681a5",
          2944 => x"387333d0",
          2945 => x"117081ff",
          2946 => x"06515253",
          2947 => x"70892691",
          2948 => x"38821473",
          2949 => x"81ff06d0",
          2950 => x"05565271",
          2951 => x"762e80f7",
          2952 => x"38800b81",
          2953 => x"c3cc5955",
          2954 => x"77087a55",
          2955 => x"57767081",
          2956 => x"05583374",
          2957 => x"70810556",
          2958 => x"33ff9f12",
          2959 => x"53535370",
          2960 => x"99268938",
          2961 => x"e0137081",
          2962 => x"ff065451",
          2963 => x"ff9f1251",
          2964 => x"70992689",
          2965 => x"38e01270",
          2966 => x"81ff0653",
          2967 => x"51723070",
          2968 => x"9f2a5151",
          2969 => x"72722e09",
          2970 => x"81068538",
          2971 => x"70ffbe38",
          2972 => x"72307477",
          2973 => x"32703070",
          2974 => x"72079f2a",
          2975 => x"739f2a07",
          2976 => x"53545451",
          2977 => x"70802e8f",
          2978 => x"38811584",
          2979 => x"19595583",
          2980 => x"7525ff94",
          2981 => x"388b3974",
          2982 => x"83248638",
          2983 => x"74767c0c",
          2984 => x"59785186",
          2985 => x"3981d488",
          2986 => x"33517081",
          2987 => x"d3d80c8c",
          2988 => x"3d0d04fa",
          2989 => x"3d0d7856",
          2990 => x"800b8317",
          2991 => x"34ff0bb0",
          2992 => x"170c7952",
          2993 => x"7551e2e0",
          2994 => x"3f845581",
          2995 => x"d3d80881",
          2996 => x"803884b2",
          2997 => x"1651dfb4",
          2998 => x"3f81d3d8",
          2999 => x"0883ffff",
          3000 => x"06548355",
          3001 => x"7382d4d5",
          3002 => x"2e098106",
          3003 => x"80e33880",
          3004 => x"0bb41733",
          3005 => x"56577481",
          3006 => x"e92e0981",
          3007 => x"06833881",
          3008 => x"577481eb",
          3009 => x"32703070",
          3010 => x"80257907",
          3011 => x"51515473",
          3012 => x"8a387481",
          3013 => x"e82e0981",
          3014 => x"06b53883",
          3015 => x"5381c38c",
          3016 => x"5280ea16",
          3017 => x"51e0b13f",
          3018 => x"81d3d808",
          3019 => x"5581d3d8",
          3020 => x"08802e9d",
          3021 => x"38855381",
          3022 => x"c3905281",
          3023 => x"861651e0",
          3024 => x"973f81d3",
          3025 => x"d8085581",
          3026 => x"d3d80880",
          3027 => x"2e833882",
          3028 => x"557481d3",
          3029 => x"d80c883d",
          3030 => x"0d04f23d",
          3031 => x"0d610284",
          3032 => x"0580cb05",
          3033 => x"33585580",
          3034 => x"750c6051",
          3035 => x"fce13f81",
          3036 => x"d3d80858",
          3037 => x"8b56800b",
          3038 => x"81d3d808",
          3039 => x"2486fc38",
          3040 => x"81d3d808",
          3041 => x"842981d3",
          3042 => x"f4057008",
          3043 => x"55538c56",
          3044 => x"73802e86",
          3045 => x"e6387375",
          3046 => x"0c7681fe",
          3047 => x"06743354",
          3048 => x"5772802e",
          3049 => x"ae388114",
          3050 => x"3351d7ca",
          3051 => x"3f81d3d8",
          3052 => x"0881ff06",
          3053 => x"70810654",
          3054 => x"55729838",
          3055 => x"76802e86",
          3056 => x"b8387482",
          3057 => x"2a708106",
          3058 => x"51538a56",
          3059 => x"7286ac38",
          3060 => x"86a73980",
          3061 => x"74347781",
          3062 => x"15348152",
          3063 => x"81143351",
          3064 => x"d7b23f81",
          3065 => x"d3d80881",
          3066 => x"ff067081",
          3067 => x"06545583",
          3068 => x"56728687",
          3069 => x"3876802e",
          3070 => x"8f387482",
          3071 => x"2a708106",
          3072 => x"51538a56",
          3073 => x"7285f438",
          3074 => x"80705374",
          3075 => x"525bfda3",
          3076 => x"3f81d3d8",
          3077 => x"0881ff06",
          3078 => x"5776822e",
          3079 => x"09810680",
          3080 => x"e2388c3d",
          3081 => x"74565883",
          3082 => x"5683f615",
          3083 => x"33705853",
          3084 => x"72802e8d",
          3085 => x"3883fa15",
          3086 => x"51dce83f",
          3087 => x"81d3d808",
          3088 => x"57767870",
          3089 => x"84055a0c",
          3090 => x"ff169016",
          3091 => x"56567580",
          3092 => x"25d73880",
          3093 => x"0b8d3d54",
          3094 => x"56727084",
          3095 => x"0554085b",
          3096 => x"83577a80",
          3097 => x"2e95387a",
          3098 => x"527351fc",
          3099 => x"c63f81d3",
          3100 => x"d80881ff",
          3101 => x"06578177",
          3102 => x"27893881",
          3103 => x"16568376",
          3104 => x"27d73881",
          3105 => x"5676842e",
          3106 => x"84f1388d",
          3107 => x"56768126",
          3108 => x"84e938bf",
          3109 => x"1451dbf4",
          3110 => x"3f81d3d8",
          3111 => x"0883ffff",
          3112 => x"06537284",
          3113 => x"802e0981",
          3114 => x"0684d038",
          3115 => x"80ca1451",
          3116 => x"dbda3f81",
          3117 => x"d3d80883",
          3118 => x"ffff0658",
          3119 => x"778d3880",
          3120 => x"d81451db",
          3121 => x"de3f81d3",
          3122 => x"d8085877",
          3123 => x"9c150c80",
          3124 => x"c4143382",
          3125 => x"153480c4",
          3126 => x"1433ff11",
          3127 => x"7081ff06",
          3128 => x"5154558d",
          3129 => x"56728126",
          3130 => x"84913874",
          3131 => x"81ff0678",
          3132 => x"712980c1",
          3133 => x"16335259",
          3134 => x"53728a15",
          3135 => x"2372802e",
          3136 => x"8b38ff13",
          3137 => x"73065372",
          3138 => x"802e8638",
          3139 => x"8d5683eb",
          3140 => x"3980c514",
          3141 => x"51daf53f",
          3142 => x"81d3d808",
          3143 => x"5381d3d8",
          3144 => x"08881523",
          3145 => x"728f0657",
          3146 => x"8d567683",
          3147 => x"ce3880c7",
          3148 => x"1451dad8",
          3149 => x"3f81d3d8",
          3150 => x"0883ffff",
          3151 => x"0655748d",
          3152 => x"3880d414",
          3153 => x"51dadc3f",
          3154 => x"81d3d808",
          3155 => x"5580c214",
          3156 => x"51dab93f",
          3157 => x"81d3d808",
          3158 => x"83ffff06",
          3159 => x"538d5672",
          3160 => x"802e8397",
          3161 => x"38881422",
          3162 => x"78147184",
          3163 => x"2a055a5a",
          3164 => x"78752683",
          3165 => x"86388a14",
          3166 => x"22527479",
          3167 => x"3151ffaf",
          3168 => x"f63f81d3",
          3169 => x"d8085581",
          3170 => x"d3d80880",
          3171 => x"2e82ec38",
          3172 => x"81d3d808",
          3173 => x"80ffffff",
          3174 => x"f5268338",
          3175 => x"83577483",
          3176 => x"fff52683",
          3177 => x"38825774",
          3178 => x"9ff52685",
          3179 => x"38815789",
          3180 => x"398d5676",
          3181 => x"802e82c3",
          3182 => x"38821570",
          3183 => x"98160c7b",
          3184 => x"a0160c73",
          3185 => x"1c70a417",
          3186 => x"0c7a1dac",
          3187 => x"170c5455",
          3188 => x"76832e09",
          3189 => x"8106af38",
          3190 => x"80de1451",
          3191 => x"d9ae3f81",
          3192 => x"d3d80883",
          3193 => x"ffff0653",
          3194 => x"8d567282",
          3195 => x"8e387982",
          3196 => x"8a3880e0",
          3197 => x"1451d9ab",
          3198 => x"3f81d3d8",
          3199 => x"08a8150c",
          3200 => x"74822b53",
          3201 => x"a2398d56",
          3202 => x"79802e81",
          3203 => x"ee387713",
          3204 => x"a8150c74",
          3205 => x"15537682",
          3206 => x"2e8d3874",
          3207 => x"10157081",
          3208 => x"2a768106",
          3209 => x"05515383",
          3210 => x"ff13892a",
          3211 => x"538d5672",
          3212 => x"9c150826",
          3213 => x"81c538ff",
          3214 => x"0b90150c",
          3215 => x"ff0b8c15",
          3216 => x"0cff800b",
          3217 => x"84153476",
          3218 => x"832e0981",
          3219 => x"06819238",
          3220 => x"80e41451",
          3221 => x"d8b63f81",
          3222 => x"d3d80883",
          3223 => x"ffff0653",
          3224 => x"72812e09",
          3225 => x"810680f9",
          3226 => x"38811b52",
          3227 => x"7351dbb8",
          3228 => x"3f81d3d8",
          3229 => x"0880ea38",
          3230 => x"81d3d808",
          3231 => x"84153484",
          3232 => x"b21451d8",
          3233 => x"873f81d3",
          3234 => x"d80883ff",
          3235 => x"ff065372",
          3236 => x"82d4d52e",
          3237 => x"09810680",
          3238 => x"c838b414",
          3239 => x"51d8843f",
          3240 => x"81d3d808",
          3241 => x"848b85a4",
          3242 => x"d22e0981",
          3243 => x"06b33884",
          3244 => x"981451d7",
          3245 => x"ee3f81d3",
          3246 => x"d808868a",
          3247 => x"85e4f22e",
          3248 => x"0981069d",
          3249 => x"38849c14",
          3250 => x"51d7d83f",
          3251 => x"81d3d808",
          3252 => x"90150c84",
          3253 => x"a01451d7",
          3254 => x"ca3f81d3",
          3255 => x"d8088c15",
          3256 => x"0c767434",
          3257 => x"81d48422",
          3258 => x"81055372",
          3259 => x"81d48423",
          3260 => x"72861523",
          3261 => x"800b9415",
          3262 => x"0c805675",
          3263 => x"81d3d80c",
          3264 => x"903d0d04",
          3265 => x"fb3d0d77",
          3266 => x"54895573",
          3267 => x"802eb938",
          3268 => x"73085372",
          3269 => x"802eb138",
          3270 => x"72335271",
          3271 => x"802ea938",
          3272 => x"86132284",
          3273 => x"15225752",
          3274 => x"71762e09",
          3275 => x"81069938",
          3276 => x"81133351",
          3277 => x"d0c03f81",
          3278 => x"d3d80881",
          3279 => x"06527188",
          3280 => x"38717408",
          3281 => x"54558339",
          3282 => x"80537873",
          3283 => x"710c5274",
          3284 => x"81d3d80c",
          3285 => x"873d0d04",
          3286 => x"fa3d0d02",
          3287 => x"ab05337a",
          3288 => x"58893dfc",
          3289 => x"055256f4",
          3290 => x"e63f8b54",
          3291 => x"800b81d3",
          3292 => x"d80824bc",
          3293 => x"3881d3d8",
          3294 => x"08842981",
          3295 => x"d3f40570",
          3296 => x"08555573",
          3297 => x"802e8438",
          3298 => x"80743478",
          3299 => x"5473802e",
          3300 => x"84388074",
          3301 => x"3478750c",
          3302 => x"75547580",
          3303 => x"2e923880",
          3304 => x"53893d70",
          3305 => x"53840551",
          3306 => x"f7b03f81",
          3307 => x"d3d80854",
          3308 => x"7381d3d8",
          3309 => x"0c883d0d",
          3310 => x"04eb3d0d",
          3311 => x"67028405",
          3312 => x"80e70533",
          3313 => x"59598954",
          3314 => x"78802e84",
          3315 => x"c83877bf",
          3316 => x"06705498",
          3317 => x"3dd00553",
          3318 => x"993d8405",
          3319 => x"5258f6fa",
          3320 => x"3f81d3d8",
          3321 => x"085581d3",
          3322 => x"d80884a4",
          3323 => x"387a5c68",
          3324 => x"528c3d70",
          3325 => x"5256edc6",
          3326 => x"3f81d3d8",
          3327 => x"085581d3",
          3328 => x"d8089238",
          3329 => x"0280d705",
          3330 => x"3370982b",
          3331 => x"55577380",
          3332 => x"25833886",
          3333 => x"55779c06",
          3334 => x"5473802e",
          3335 => x"81ab3874",
          3336 => x"802e9538",
          3337 => x"74842e09",
          3338 => x"8106aa38",
          3339 => x"7551eaf8",
          3340 => x"3f81d3d8",
          3341 => x"08559e39",
          3342 => x"02b20533",
          3343 => x"91065473",
          3344 => x"81b83877",
          3345 => x"822a7081",
          3346 => x"06515473",
          3347 => x"802e8e38",
          3348 => x"885583bc",
          3349 => x"39778807",
          3350 => x"587483b4",
          3351 => x"3877832a",
          3352 => x"70810651",
          3353 => x"5473802e",
          3354 => x"81af3862",
          3355 => x"527a51e8",
          3356 => x"a53f81d3",
          3357 => x"d8085682",
          3358 => x"88b20a52",
          3359 => x"628e0551",
          3360 => x"d4ea3f62",
          3361 => x"54a00b8b",
          3362 => x"15348053",
          3363 => x"62527a51",
          3364 => x"e8bd3f80",
          3365 => x"52629c05",
          3366 => x"51d4d13f",
          3367 => x"7a54810b",
          3368 => x"83153475",
          3369 => x"802e80f1",
          3370 => x"387ab011",
          3371 => x"08515480",
          3372 => x"53755297",
          3373 => x"3dd40551",
          3374 => x"ddbe3f81",
          3375 => x"d3d80855",
          3376 => x"81d3d808",
          3377 => x"82ca38b7",
          3378 => x"397482c4",
          3379 => x"3802b205",
          3380 => x"3370842a",
          3381 => x"70810651",
          3382 => x"55567380",
          3383 => x"2e863884",
          3384 => x"5582ad39",
          3385 => x"77812a70",
          3386 => x"81065154",
          3387 => x"73802ea9",
          3388 => x"38758106",
          3389 => x"5473802e",
          3390 => x"a0388755",
          3391 => x"82923973",
          3392 => x"527a51d6",
          3393 => x"a33f81d3",
          3394 => x"d8087bff",
          3395 => x"188c120c",
          3396 => x"555581d3",
          3397 => x"d80881f8",
          3398 => x"3877832a",
          3399 => x"70810651",
          3400 => x"5473802e",
          3401 => x"86387780",
          3402 => x"c007587a",
          3403 => x"b01108a0",
          3404 => x"1b0c63a4",
          3405 => x"1b0c6353",
          3406 => x"705257e6",
          3407 => x"d93f81d3",
          3408 => x"d80881d3",
          3409 => x"d808881b",
          3410 => x"0c639c05",
          3411 => x"525ad2d3",
          3412 => x"3f81d3d8",
          3413 => x"0881d3d8",
          3414 => x"088c1b0c",
          3415 => x"777a0c56",
          3416 => x"86172284",
          3417 => x"1a237790",
          3418 => x"1a34800b",
          3419 => x"911a3480",
          3420 => x"0b9c1a0c",
          3421 => x"800b941a",
          3422 => x"0c77852a",
          3423 => x"70810651",
          3424 => x"5473802e",
          3425 => x"818d3881",
          3426 => x"d3d80880",
          3427 => x"2e818438",
          3428 => x"81d3d808",
          3429 => x"941a0c8a",
          3430 => x"17227089",
          3431 => x"2b7b5259",
          3432 => x"57a83976",
          3433 => x"527851d7",
          3434 => x"9f3f81d3",
          3435 => x"d8085781",
          3436 => x"d3d80881",
          3437 => x"26833882",
          3438 => x"5581d3d8",
          3439 => x"08ff2e09",
          3440 => x"81068338",
          3441 => x"79557578",
          3442 => x"31567430",
          3443 => x"70760780",
          3444 => x"25515477",
          3445 => x"76278a38",
          3446 => x"81707506",
          3447 => x"555a73c3",
          3448 => x"3876981a",
          3449 => x"0c74a938",
          3450 => x"7583ff06",
          3451 => x"5473802e",
          3452 => x"a2387652",
          3453 => x"7a51d6a6",
          3454 => x"3f81d3d8",
          3455 => x"08853882",
          3456 => x"558e3975",
          3457 => x"892a81d3",
          3458 => x"d808059c",
          3459 => x"1a0c8439",
          3460 => x"80790c74",
          3461 => x"547381d3",
          3462 => x"d80c973d",
          3463 => x"0d04f23d",
          3464 => x"0d606365",
          3465 => x"6440405d",
          3466 => x"59807e0c",
          3467 => x"903dfc05",
          3468 => x"527851f9",
          3469 => x"cf3f81d3",
          3470 => x"d8085581",
          3471 => x"d3d8088a",
          3472 => x"38911933",
          3473 => x"5574802e",
          3474 => x"86387456",
          3475 => x"82c43990",
          3476 => x"19338106",
          3477 => x"55875674",
          3478 => x"802e82b6",
          3479 => x"38953982",
          3480 => x"0b911a34",
          3481 => x"825682aa",
          3482 => x"39810b91",
          3483 => x"1a348156",
          3484 => x"82a0398c",
          3485 => x"1908941a",
          3486 => x"08315574",
          3487 => x"7c278338",
          3488 => x"745c7b80",
          3489 => x"2e828938",
          3490 => x"94190870",
          3491 => x"83ff0656",
          3492 => x"567481b2",
          3493 => x"387e8a11",
          3494 => x"22ff0577",
          3495 => x"892a065b",
          3496 => x"5579a838",
          3497 => x"75873888",
          3498 => x"1908558f",
          3499 => x"39981908",
          3500 => x"527851d5",
          3501 => x"933f81d3",
          3502 => x"d8085581",
          3503 => x"7527ff9f",
          3504 => x"3874ff2e",
          3505 => x"ffa33874",
          3506 => x"981a0c98",
          3507 => x"1908527e",
          3508 => x"51d4cb3f",
          3509 => x"81d3d808",
          3510 => x"802eff83",
          3511 => x"3881d3d8",
          3512 => x"081a7c89",
          3513 => x"2a595777",
          3514 => x"802e80d6",
          3515 => x"38771a7f",
          3516 => x"8a112258",
          3517 => x"5c557575",
          3518 => x"27853875",
          3519 => x"7a315877",
          3520 => x"5476537c",
          3521 => x"52811b33",
          3522 => x"51ca883f",
          3523 => x"81d3d808",
          3524 => x"fed7387e",
          3525 => x"83113356",
          3526 => x"5674802e",
          3527 => x"9f38b016",
          3528 => x"08773155",
          3529 => x"74782794",
          3530 => x"38848053",
          3531 => x"b41652b0",
          3532 => x"16087731",
          3533 => x"892b7d05",
          3534 => x"51cfe03f",
          3535 => x"77892b56",
          3536 => x"b939769c",
          3537 => x"1a0c9419",
          3538 => x"0883ff06",
          3539 => x"84807131",
          3540 => x"57557b76",
          3541 => x"2783387b",
          3542 => x"569c1908",
          3543 => x"527e51d1",
          3544 => x"c73f81d3",
          3545 => x"d808fe81",
          3546 => x"38755394",
          3547 => x"190883ff",
          3548 => x"061fb405",
          3549 => x"527c51cf",
          3550 => x"a23f7b76",
          3551 => x"317e0817",
          3552 => x"7f0c761e",
          3553 => x"941b0818",
          3554 => x"941c0c5e",
          3555 => x"5cfdf339",
          3556 => x"80567581",
          3557 => x"d3d80c90",
          3558 => x"3d0d04f2",
          3559 => x"3d0d6063",
          3560 => x"65644040",
          3561 => x"5d58807e",
          3562 => x"0c903dfc",
          3563 => x"05527751",
          3564 => x"f6d23f81",
          3565 => x"d3d80855",
          3566 => x"81d3d808",
          3567 => x"8a389118",
          3568 => x"33557480",
          3569 => x"2e863874",
          3570 => x"5683b839",
          3571 => x"90183370",
          3572 => x"812a7081",
          3573 => x"06515656",
          3574 => x"87567480",
          3575 => x"2e83a438",
          3576 => x"9539820b",
          3577 => x"91193482",
          3578 => x"56839839",
          3579 => x"810b9119",
          3580 => x"34815683",
          3581 => x"8e399418",
          3582 => x"087c1156",
          3583 => x"56747627",
          3584 => x"84387509",
          3585 => x"5c7b802e",
          3586 => x"82ec3894",
          3587 => x"18087083",
          3588 => x"ff065656",
          3589 => x"7481fd38",
          3590 => x"7e8a1122",
          3591 => x"ff057789",
          3592 => x"2a065c55",
          3593 => x"7abf3875",
          3594 => x"8c388818",
          3595 => x"0855749c",
          3596 => x"387a5285",
          3597 => x"39981808",
          3598 => x"527751d7",
          3599 => x"e73f81d3",
          3600 => x"d8085581",
          3601 => x"d3d80880",
          3602 => x"2e82ab38",
          3603 => x"74812eff",
          3604 => x"913874ff",
          3605 => x"2eff9538",
          3606 => x"7498190c",
          3607 => x"88180885",
          3608 => x"38748819",
          3609 => x"0c7e55b0",
          3610 => x"15089c19",
          3611 => x"082e0981",
          3612 => x"068d3874",
          3613 => x"51cec13f",
          3614 => x"81d3d808",
          3615 => x"feee3898",
          3616 => x"1808527e",
          3617 => x"51d1973f",
          3618 => x"81d3d808",
          3619 => x"802efed2",
          3620 => x"3881d3d8",
          3621 => x"081b7c89",
          3622 => x"2a5a5778",
          3623 => x"802e80d5",
          3624 => x"38781b7f",
          3625 => x"8a112258",
          3626 => x"5b557575",
          3627 => x"27853875",
          3628 => x"7b315978",
          3629 => x"5476537c",
          3630 => x"52811a33",
          3631 => x"51c8be3f",
          3632 => x"81d3d808",
          3633 => x"fea6387e",
          3634 => x"b0110878",
          3635 => x"31565674",
          3636 => x"79279b38",
          3637 => x"848053b0",
          3638 => x"16087731",
          3639 => x"892b7d05",
          3640 => x"52b41651",
          3641 => x"ccb53f7e",
          3642 => x"55800b83",
          3643 => x"16347889",
          3644 => x"2b5680db",
          3645 => x"398c1808",
          3646 => x"94190826",
          3647 => x"93387e51",
          3648 => x"cdb63f81",
          3649 => x"d3d808fd",
          3650 => x"e3387e77",
          3651 => x"b0120c55",
          3652 => x"769c190c",
          3653 => x"94180883",
          3654 => x"ff068480",
          3655 => x"71315755",
          3656 => x"7b762783",
          3657 => x"387b569c",
          3658 => x"1808527e",
          3659 => x"51cdf93f",
          3660 => x"81d3d808",
          3661 => x"fdb63875",
          3662 => x"537c5294",
          3663 => x"180883ff",
          3664 => x"061fb405",
          3665 => x"51cbd43f",
          3666 => x"7e55810b",
          3667 => x"8316347b",
          3668 => x"76317e08",
          3669 => x"177f0c76",
          3670 => x"1e941a08",
          3671 => x"1870941c",
          3672 => x"0c8c1b08",
          3673 => x"58585e5c",
          3674 => x"74762783",
          3675 => x"38755574",
          3676 => x"8c190cfd",
          3677 => x"90399018",
          3678 => x"3380c007",
          3679 => x"55749019",
          3680 => x"34805675",
          3681 => x"81d3d80c",
          3682 => x"903d0d04",
          3683 => x"f83d0d7a",
          3684 => x"8b3dfc05",
          3685 => x"53705256",
          3686 => x"f2ea3f81",
          3687 => x"d3d80857",
          3688 => x"81d3d808",
          3689 => x"80fb3890",
          3690 => x"16337086",
          3691 => x"2a708106",
          3692 => x"51555573",
          3693 => x"802e80e9",
          3694 => x"38a01608",
          3695 => x"527851cc",
          3696 => x"e73f81d3",
          3697 => x"d8085781",
          3698 => x"d3d80880",
          3699 => x"d438a416",
          3700 => x"088b1133",
          3701 => x"a0075555",
          3702 => x"738b1634",
          3703 => x"88160853",
          3704 => x"74527508",
          3705 => x"51dde83f",
          3706 => x"8c160852",
          3707 => x"9c1551c9",
          3708 => x"fb3f8288",
          3709 => x"b20a5296",
          3710 => x"1551c9f0",
          3711 => x"3f765292",
          3712 => x"1551c9ca",
          3713 => x"3f785481",
          3714 => x"0b831534",
          3715 => x"7851ccdf",
          3716 => x"3f81d3d8",
          3717 => x"08901733",
          3718 => x"81bf0655",
          3719 => x"57739017",
          3720 => x"347681d3",
          3721 => x"d80c8a3d",
          3722 => x"0d04fc3d",
          3723 => x"0d767052",
          3724 => x"54fed93f",
          3725 => x"81d3d808",
          3726 => x"5381d3d8",
          3727 => x"089c3886",
          3728 => x"3dfc0552",
          3729 => x"7351f1bc",
          3730 => x"3f81d3d8",
          3731 => x"085381d3",
          3732 => x"d8088738",
          3733 => x"81d3d808",
          3734 => x"740c7281",
          3735 => x"d3d80c86",
          3736 => x"3d0d04ff",
          3737 => x"3d0d843d",
          3738 => x"51e6e43f",
          3739 => x"8b52800b",
          3740 => x"81d3d808",
          3741 => x"248b3881",
          3742 => x"d3d80881",
          3743 => x"d4883480",
          3744 => x"527181d3",
          3745 => x"d80c833d",
          3746 => x"0d04ef3d",
          3747 => x"0d805393",
          3748 => x"3dd00552",
          3749 => x"943d51e9",
          3750 => x"c13f81d3",
          3751 => x"d8085581",
          3752 => x"d3d80880",
          3753 => x"e0387658",
          3754 => x"6352933d",
          3755 => x"d40551e0",
          3756 => x"8d3f81d3",
          3757 => x"d8085581",
          3758 => x"d3d808bc",
          3759 => x"380280c7",
          3760 => x"05337098",
          3761 => x"2b555673",
          3762 => x"80258938",
          3763 => x"767a9412",
          3764 => x"0c54b239",
          3765 => x"02a20533",
          3766 => x"70842a70",
          3767 => x"81065155",
          3768 => x"5673802e",
          3769 => x"9e38767f",
          3770 => x"53705254",
          3771 => x"dba83f81",
          3772 => x"d3d80894",
          3773 => x"150c8e39",
          3774 => x"81d3d808",
          3775 => x"842e0981",
          3776 => x"06833885",
          3777 => x"557481d3",
          3778 => x"d80c933d",
          3779 => x"0d04e43d",
          3780 => x"0d6f6f5b",
          3781 => x"5b807a34",
          3782 => x"80539e3d",
          3783 => x"ffb80552",
          3784 => x"9f3d51e8",
          3785 => x"b53f81d3",
          3786 => x"d8085781",
          3787 => x"d3d80882",
          3788 => x"fc387b43",
          3789 => x"7a7c9411",
          3790 => x"08475558",
          3791 => x"64547380",
          3792 => x"2e81ed38",
          3793 => x"a052933d",
          3794 => x"705255d5",
          3795 => x"ea3f81d3",
          3796 => x"d8085781",
          3797 => x"d3d80882",
          3798 => x"d4386852",
          3799 => x"7b51c9c8",
          3800 => x"3f81d3d8",
          3801 => x"085781d3",
          3802 => x"d80882c1",
          3803 => x"3869527b",
          3804 => x"51daa33f",
          3805 => x"81d3d808",
          3806 => x"45765274",
          3807 => x"51d5b83f",
          3808 => x"81d3d808",
          3809 => x"5781d3d8",
          3810 => x"0882a238",
          3811 => x"80527451",
          3812 => x"daeb3f81",
          3813 => x"d3d80857",
          3814 => x"81d3d808",
          3815 => x"a4386952",
          3816 => x"7b51d9f2",
          3817 => x"3f7381d3",
          3818 => x"d8082ea6",
          3819 => x"38765274",
          3820 => x"51d6cf3f",
          3821 => x"81d3d808",
          3822 => x"5781d3d8",
          3823 => x"08802ecc",
          3824 => x"3876842e",
          3825 => x"09810686",
          3826 => x"38825781",
          3827 => x"e0397681",
          3828 => x"dc389e3d",
          3829 => x"ffbc0552",
          3830 => x"7451dcc9",
          3831 => x"3f76903d",
          3832 => x"78118111",
          3833 => x"3351565a",
          3834 => x"5673802e",
          3835 => x"913802b9",
          3836 => x"05558116",
          3837 => x"81167033",
          3838 => x"56565673",
          3839 => x"f5388116",
          3840 => x"54737826",
          3841 => x"81903875",
          3842 => x"802e9938",
          3843 => x"78168105",
          3844 => x"55ff186f",
          3845 => x"11ff18ff",
          3846 => x"18585855",
          3847 => x"58743374",
          3848 => x"3475ee38",
          3849 => x"ff186f11",
          3850 => x"5558af74",
          3851 => x"34fe8d39",
          3852 => x"777b2e09",
          3853 => x"81068a38",
          3854 => x"ff186f11",
          3855 => x"5558af74",
          3856 => x"34800b81",
          3857 => x"d4883370",
          3858 => x"842981c3",
          3859 => x"cc057008",
          3860 => x"7033525c",
          3861 => x"56565673",
          3862 => x"762e8d38",
          3863 => x"8116701a",
          3864 => x"70335155",
          3865 => x"5673f538",
          3866 => x"82165473",
          3867 => x"7826a738",
          3868 => x"80557476",
          3869 => x"27913874",
          3870 => x"19547333",
          3871 => x"7a708105",
          3872 => x"5c348115",
          3873 => x"55ec39ba",
          3874 => x"7a708105",
          3875 => x"5c3474ff",
          3876 => x"2e098106",
          3877 => x"85389157",
          3878 => x"94396e18",
          3879 => x"81195954",
          3880 => x"73337a70",
          3881 => x"81055c34",
          3882 => x"7a7826ee",
          3883 => x"38807a34",
          3884 => x"7681d3d8",
          3885 => x"0c9e3d0d",
          3886 => x"04f73d0d",
          3887 => x"7b7d8d3d",
          3888 => x"fc055471",
          3889 => x"535755ec",
          3890 => x"bb3f81d3",
          3891 => x"d8085381",
          3892 => x"d3d80882",
          3893 => x"fa389115",
          3894 => x"33537282",
          3895 => x"f2388c15",
          3896 => x"08547376",
          3897 => x"27923890",
          3898 => x"15337081",
          3899 => x"2a708106",
          3900 => x"51545772",
          3901 => x"83387356",
          3902 => x"94150854",
          3903 => x"80709417",
          3904 => x"0c587578",
          3905 => x"2e829738",
          3906 => x"798a1122",
          3907 => x"70892b59",
          3908 => x"51537378",
          3909 => x"2eb73876",
          3910 => x"52ff1651",
          3911 => x"ff98d83f",
          3912 => x"81d3d808",
          3913 => x"ff157854",
          3914 => x"70535553",
          3915 => x"ff98c83f",
          3916 => x"81d3d808",
          3917 => x"73269638",
          3918 => x"76307075",
          3919 => x"06709418",
          3920 => x"0c777131",
          3921 => x"98180857",
          3922 => x"585153b1",
          3923 => x"39881508",
          3924 => x"5473a638",
          3925 => x"73527451",
          3926 => x"cdca3f81",
          3927 => x"d3d80854",
          3928 => x"81d3d808",
          3929 => x"812e819a",
          3930 => x"3881d3d8",
          3931 => x"08ff2e81",
          3932 => x"9b3881d3",
          3933 => x"d8088816",
          3934 => x"0c739816",
          3935 => x"0c73802e",
          3936 => x"819c3876",
          3937 => x"762780dc",
          3938 => x"38757731",
          3939 => x"94160818",
          3940 => x"94170c90",
          3941 => x"16337081",
          3942 => x"2a708106",
          3943 => x"51555a56",
          3944 => x"72802e9a",
          3945 => x"38735274",
          3946 => x"51ccf93f",
          3947 => x"81d3d808",
          3948 => x"5481d3d8",
          3949 => x"08943881",
          3950 => x"d3d80856",
          3951 => x"a7397352",
          3952 => x"7451c784",
          3953 => x"3f81d3d8",
          3954 => x"085473ff",
          3955 => x"2ebe3881",
          3956 => x"7427af38",
          3957 => x"79537398",
          3958 => x"140827a6",
          3959 => x"38739816",
          3960 => x"0cffa039",
          3961 => x"94150816",
          3962 => x"94160c75",
          3963 => x"83ff0653",
          3964 => x"72802eaa",
          3965 => x"38735279",
          3966 => x"51c6a33f",
          3967 => x"81d3d808",
          3968 => x"9438820b",
          3969 => x"91163482",
          3970 => x"5380c439",
          3971 => x"810b9116",
          3972 => x"348153bb",
          3973 => x"3975892a",
          3974 => x"81d3d808",
          3975 => x"05589415",
          3976 => x"08548c15",
          3977 => x"08742790",
          3978 => x"38738c16",
          3979 => x"0c901533",
          3980 => x"80c00753",
          3981 => x"72901634",
          3982 => x"7383ff06",
          3983 => x"5372802e",
          3984 => x"8c38779c",
          3985 => x"16082e85",
          3986 => x"38779c16",
          3987 => x"0c805372",
          3988 => x"81d3d80c",
          3989 => x"8b3d0d04",
          3990 => x"f93d0d79",
          3991 => x"56895475",
          3992 => x"802e818a",
          3993 => x"38805389",
          3994 => x"3dfc0552",
          3995 => x"8a3d8405",
          3996 => x"51e1e73f",
          3997 => x"81d3d808",
          3998 => x"5581d3d8",
          3999 => x"0880ea38",
          4000 => x"77760c7a",
          4001 => x"527551d8",
          4002 => x"b53f81d3",
          4003 => x"d8085581",
          4004 => x"d3d80880",
          4005 => x"c338ab16",
          4006 => x"3370982b",
          4007 => x"55578074",
          4008 => x"24a23886",
          4009 => x"16337084",
          4010 => x"2a708106",
          4011 => x"51555773",
          4012 => x"802ead38",
          4013 => x"9c160852",
          4014 => x"7751d3da",
          4015 => x"3f81d3d8",
          4016 => x"0888170c",
          4017 => x"77548614",
          4018 => x"22841723",
          4019 => x"74527551",
          4020 => x"cee53f81",
          4021 => x"d3d80855",
          4022 => x"74842e09",
          4023 => x"81068538",
          4024 => x"85558639",
          4025 => x"74802e84",
          4026 => x"3880760c",
          4027 => x"74547381",
          4028 => x"d3d80c89",
          4029 => x"3d0d04fc",
          4030 => x"3d0d7687",
          4031 => x"3dfc0553",
          4032 => x"705253e7",
          4033 => x"ff3f81d3",
          4034 => x"d8088738",
          4035 => x"81d3d808",
          4036 => x"730c863d",
          4037 => x"0d04fb3d",
          4038 => x"0d777989",
          4039 => x"3dfc0554",
          4040 => x"71535654",
          4041 => x"e7de3f81",
          4042 => x"d3d80853",
          4043 => x"81d3d808",
          4044 => x"80df3874",
          4045 => x"933881d3",
          4046 => x"d8085273",
          4047 => x"51cdf83f",
          4048 => x"81d3d808",
          4049 => x"5380ca39",
          4050 => x"81d3d808",
          4051 => x"527351d3",
          4052 => x"ac3f81d3",
          4053 => x"d8085381",
          4054 => x"d3d80884",
          4055 => x"2e098106",
          4056 => x"85388053",
          4057 => x"873981d3",
          4058 => x"d808a638",
          4059 => x"74527351",
          4060 => x"d5b33f72",
          4061 => x"527351cf",
          4062 => x"893f81d3",
          4063 => x"d8088432",
          4064 => x"70307072",
          4065 => x"079f2c70",
          4066 => x"81d3d808",
          4067 => x"06515154",
          4068 => x"547281d3",
          4069 => x"d80c873d",
          4070 => x"0d04ee3d",
          4071 => x"0d655780",
          4072 => x"53893d70",
          4073 => x"53963d52",
          4074 => x"56dfaf3f",
          4075 => x"81d3d808",
          4076 => x"5581d3d8",
          4077 => x"08b23864",
          4078 => x"527551d6",
          4079 => x"813f81d3",
          4080 => x"d8085581",
          4081 => x"d3d808a0",
          4082 => x"380280cb",
          4083 => x"05337098",
          4084 => x"2b555873",
          4085 => x"80258538",
          4086 => x"86558d39",
          4087 => x"76802e88",
          4088 => x"38765275",
          4089 => x"51d4be3f",
          4090 => x"7481d3d8",
          4091 => x"0c943d0d",
          4092 => x"04f03d0d",
          4093 => x"6365555c",
          4094 => x"8053923d",
          4095 => x"ec055293",
          4096 => x"3d51ded6",
          4097 => x"3f81d3d8",
          4098 => x"085b81d3",
          4099 => x"d8088280",
          4100 => x"387c740c",
          4101 => x"73089811",
          4102 => x"08fe1190",
          4103 => x"13085956",
          4104 => x"58557574",
          4105 => x"26913875",
          4106 => x"7c0c81e4",
          4107 => x"39815b81",
          4108 => x"cc39825b",
          4109 => x"81c73981",
          4110 => x"d3d80875",
          4111 => x"33555973",
          4112 => x"812e0981",
          4113 => x"06bf3882",
          4114 => x"755f5776",
          4115 => x"52923df0",
          4116 => x"0551c1f4",
          4117 => x"3f81d3d8",
          4118 => x"08ff2ed1",
          4119 => x"3881d3d8",
          4120 => x"08812ece",
          4121 => x"3881d3d8",
          4122 => x"08307081",
          4123 => x"d3d80807",
          4124 => x"80257a05",
          4125 => x"81197f53",
          4126 => x"595a5498",
          4127 => x"14087726",
          4128 => x"ca3880f9",
          4129 => x"39a41508",
          4130 => x"81d3d808",
          4131 => x"57587598",
          4132 => x"38775281",
          4133 => x"187d5258",
          4134 => x"ffbf8d3f",
          4135 => x"81d3d808",
          4136 => x"5b81d3d8",
          4137 => x"0880d638",
          4138 => x"7c703377",
          4139 => x"12ff1a5d",
          4140 => x"52565474",
          4141 => x"822e0981",
          4142 => x"069e38b4",
          4143 => x"1451ffbb",
          4144 => x"cb3f81d3",
          4145 => x"d80883ff",
          4146 => x"ff067030",
          4147 => x"7080251b",
          4148 => x"8219595b",
          4149 => x"51549b39",
          4150 => x"b41451ff",
          4151 => x"bbc53f81",
          4152 => x"d3d808f0",
          4153 => x"0a067030",
          4154 => x"7080251b",
          4155 => x"8419595b",
          4156 => x"51547583",
          4157 => x"ff067a58",
          4158 => x"5679ff92",
          4159 => x"38787c0c",
          4160 => x"7c799012",
          4161 => x"0c841133",
          4162 => x"81075654",
          4163 => x"74841534",
          4164 => x"7a81d3d8",
          4165 => x"0c923d0d",
          4166 => x"04f93d0d",
          4167 => x"798a3dfc",
          4168 => x"05537052",
          4169 => x"57e3dd3f",
          4170 => x"81d3d808",
          4171 => x"5681d3d8",
          4172 => x"0881a838",
          4173 => x"91173356",
          4174 => x"7581a038",
          4175 => x"90173370",
          4176 => x"812a7081",
          4177 => x"06515555",
          4178 => x"87557380",
          4179 => x"2e818e38",
          4180 => x"94170854",
          4181 => x"738c1808",
          4182 => x"27818038",
          4183 => x"739b3881",
          4184 => x"d3d80853",
          4185 => x"88170852",
          4186 => x"7651c48c",
          4187 => x"3f81d3d8",
          4188 => x"08748819",
          4189 => x"0c5680c9",
          4190 => x"39981708",
          4191 => x"527651ff",
          4192 => x"bfc63f81",
          4193 => x"d3d808ff",
          4194 => x"2e098106",
          4195 => x"83388156",
          4196 => x"81d3d808",
          4197 => x"812e0981",
          4198 => x"06853882",
          4199 => x"56a33975",
          4200 => x"a0387754",
          4201 => x"81d3d808",
          4202 => x"98150827",
          4203 => x"94389817",
          4204 => x"085381d3",
          4205 => x"d8085276",
          4206 => x"51c3bd3f",
          4207 => x"81d3d808",
          4208 => x"56941708",
          4209 => x"8c180c90",
          4210 => x"173380c0",
          4211 => x"07547390",
          4212 => x"18347580",
          4213 => x"2e853875",
          4214 => x"91183475",
          4215 => x"557481d3",
          4216 => x"d80c893d",
          4217 => x"0d04e23d",
          4218 => x"0d8253a0",
          4219 => x"3dffa405",
          4220 => x"52a13d51",
          4221 => x"dae43f81",
          4222 => x"d3d80855",
          4223 => x"81d3d808",
          4224 => x"81f53878",
          4225 => x"45a13d08",
          4226 => x"52953d70",
          4227 => x"5258d1ae",
          4228 => x"3f81d3d8",
          4229 => x"085581d3",
          4230 => x"d80881db",
          4231 => x"380280fb",
          4232 => x"05337085",
          4233 => x"2a708106",
          4234 => x"51555686",
          4235 => x"557381c7",
          4236 => x"3875982b",
          4237 => x"54807424",
          4238 => x"81bd3802",
          4239 => x"80d60533",
          4240 => x"70810658",
          4241 => x"54875576",
          4242 => x"81ad386b",
          4243 => x"527851cc",
          4244 => x"c53f81d3",
          4245 => x"d8087484",
          4246 => x"2a708106",
          4247 => x"51555673",
          4248 => x"802e80d4",
          4249 => x"38785481",
          4250 => x"d3d80894",
          4251 => x"15082e81",
          4252 => x"8638735a",
          4253 => x"81d3d808",
          4254 => x"5c76528a",
          4255 => x"3d705254",
          4256 => x"c7b53f81",
          4257 => x"d3d80855",
          4258 => x"81d3d808",
          4259 => x"80e93881",
          4260 => x"d3d80852",
          4261 => x"7351cce5",
          4262 => x"3f81d3d8",
          4263 => x"085581d3",
          4264 => x"d8088638",
          4265 => x"875580cf",
          4266 => x"3981d3d8",
          4267 => x"08842e88",
          4268 => x"3881d3d8",
          4269 => x"0880c038",
          4270 => x"7751cec2",
          4271 => x"3f81d3d8",
          4272 => x"0881d3d8",
          4273 => x"08307081",
          4274 => x"d3d80807",
          4275 => x"80255155",
          4276 => x"5575802e",
          4277 => x"94387380",
          4278 => x"2e8f3880",
          4279 => x"53755277",
          4280 => x"51c1953f",
          4281 => x"81d3d808",
          4282 => x"55748c38",
          4283 => x"7851ffba",
          4284 => x"fe3f81d3",
          4285 => x"d8085574",
          4286 => x"81d3d80c",
          4287 => x"a03d0d04",
          4288 => x"e93d0d82",
          4289 => x"53993dc0",
          4290 => x"05529a3d",
          4291 => x"51d8cb3f",
          4292 => x"81d3d808",
          4293 => x"5481d3d8",
          4294 => x"0882b038",
          4295 => x"785e6952",
          4296 => x"8e3d7052",
          4297 => x"58cf973f",
          4298 => x"81d3d808",
          4299 => x"5481d3d8",
          4300 => x"08863888",
          4301 => x"54829439",
          4302 => x"81d3d808",
          4303 => x"842e0981",
          4304 => x"06828838",
          4305 => x"0280df05",
          4306 => x"3370852a",
          4307 => x"81065155",
          4308 => x"86547481",
          4309 => x"f638785a",
          4310 => x"74528a3d",
          4311 => x"705257c1",
          4312 => x"c33f81d3",
          4313 => x"d8087555",
          4314 => x"5681d3d8",
          4315 => x"08833887",
          4316 => x"5481d3d8",
          4317 => x"08812e09",
          4318 => x"81068338",
          4319 => x"825481d3",
          4320 => x"d808ff2e",
          4321 => x"09810686",
          4322 => x"38815481",
          4323 => x"b4397381",
          4324 => x"b03881d3",
          4325 => x"d8085278",
          4326 => x"51c4a43f",
          4327 => x"81d3d808",
          4328 => x"5481d3d8",
          4329 => x"08819a38",
          4330 => x"8b53a052",
          4331 => x"b41951ff",
          4332 => x"b78c3f78",
          4333 => x"54ae0bb4",
          4334 => x"15347854",
          4335 => x"900bbf15",
          4336 => x"348288b2",
          4337 => x"0a5280ca",
          4338 => x"1951ffb6",
          4339 => x"9f3f7553",
          4340 => x"78b41153",
          4341 => x"51c9f83f",
          4342 => x"a05378b4",
          4343 => x"115380d4",
          4344 => x"0551ffb6",
          4345 => x"b63f7854",
          4346 => x"ae0b80d5",
          4347 => x"15347f53",
          4348 => x"7880d411",
          4349 => x"5351c9d7",
          4350 => x"3f785481",
          4351 => x"0b831534",
          4352 => x"7751cba4",
          4353 => x"3f81d3d8",
          4354 => x"085481d3",
          4355 => x"d808b238",
          4356 => x"8288b20a",
          4357 => x"52649605",
          4358 => x"51ffb5d0",
          4359 => x"3f755364",
          4360 => x"527851c9",
          4361 => x"aa3f6454",
          4362 => x"900b8b15",
          4363 => x"34785481",
          4364 => x"0b831534",
          4365 => x"7851ffb8",
          4366 => x"b63f81d3",
          4367 => x"d808548b",
          4368 => x"39805375",
          4369 => x"527651ff",
          4370 => x"beae3f73",
          4371 => x"81d3d80c",
          4372 => x"993d0d04",
          4373 => x"da3d0da9",
          4374 => x"3d840551",
          4375 => x"d2f13f82",
          4376 => x"53a83dff",
          4377 => x"840552a9",
          4378 => x"3d51d5ee",
          4379 => x"3f81d3d8",
          4380 => x"085581d3",
          4381 => x"d80882d3",
          4382 => x"38784da9",
          4383 => x"3d08529d",
          4384 => x"3d705258",
          4385 => x"ccb83f81",
          4386 => x"d3d80855",
          4387 => x"81d3d808",
          4388 => x"82b93802",
          4389 => x"819b0533",
          4390 => x"81a00654",
          4391 => x"86557382",
          4392 => x"aa38a053",
          4393 => x"a43d0852",
          4394 => x"a83dff88",
          4395 => x"0551ffb4",
          4396 => x"ea3fac53",
          4397 => x"7752923d",
          4398 => x"705254ff",
          4399 => x"b4dd3faa",
          4400 => x"3d085273",
          4401 => x"51cbf73f",
          4402 => x"81d3d808",
          4403 => x"5581d3d8",
          4404 => x"08953863",
          4405 => x"6f2e0981",
          4406 => x"06883865",
          4407 => x"a23d082e",
          4408 => x"92388855",
          4409 => x"81e53981",
          4410 => x"d3d80884",
          4411 => x"2e098106",
          4412 => x"81b83873",
          4413 => x"51c9b13f",
          4414 => x"81d3d808",
          4415 => x"5581d3d8",
          4416 => x"0881c838",
          4417 => x"68569353",
          4418 => x"a83dff95",
          4419 => x"05528d16",
          4420 => x"51ffb487",
          4421 => x"3f02af05",
          4422 => x"338b1734",
          4423 => x"8b163370",
          4424 => x"842a7081",
          4425 => x"06515555",
          4426 => x"73893874",
          4427 => x"a0075473",
          4428 => x"8b173478",
          4429 => x"54810b83",
          4430 => x"15348b16",
          4431 => x"3370842a",
          4432 => x"70810651",
          4433 => x"55557380",
          4434 => x"2e80e538",
          4435 => x"6e642e80",
          4436 => x"df387552",
          4437 => x"7851c6be",
          4438 => x"3f81d3d8",
          4439 => x"08527851",
          4440 => x"ffb7bb3f",
          4441 => x"825581d3",
          4442 => x"d808802e",
          4443 => x"80dd3881",
          4444 => x"d3d80852",
          4445 => x"7851ffb5",
          4446 => x"af3f81d3",
          4447 => x"d8087980",
          4448 => x"d4115858",
          4449 => x"5581d3d8",
          4450 => x"0880c038",
          4451 => x"81163354",
          4452 => x"73ae2e09",
          4453 => x"81069938",
          4454 => x"63537552",
          4455 => x"7651c6af",
          4456 => x"3f785481",
          4457 => x"0b831534",
          4458 => x"873981d3",
          4459 => x"d8089c38",
          4460 => x"7751c8ca",
          4461 => x"3f81d3d8",
          4462 => x"085581d3",
          4463 => x"d8088c38",
          4464 => x"7851ffb5",
          4465 => x"aa3f81d3",
          4466 => x"d8085574",
          4467 => x"81d3d80c",
          4468 => x"a83d0d04",
          4469 => x"ed3d0d02",
          4470 => x"80db0533",
          4471 => x"02840580",
          4472 => x"df053357",
          4473 => x"57825395",
          4474 => x"3dd00552",
          4475 => x"963d51d2",
          4476 => x"e93f81d3",
          4477 => x"d8085581",
          4478 => x"d3d80880",
          4479 => x"cf38785a",
          4480 => x"6552953d",
          4481 => x"d40551c9",
          4482 => x"b53f81d3",
          4483 => x"d8085581",
          4484 => x"d3d808b8",
          4485 => x"380280cf",
          4486 => x"053381a0",
          4487 => x"06548655",
          4488 => x"73aa3875",
          4489 => x"a7066171",
          4490 => x"098b1233",
          4491 => x"71067a74",
          4492 => x"06075157",
          4493 => x"5556748b",
          4494 => x"15347854",
          4495 => x"810b8315",
          4496 => x"347851ff",
          4497 => x"b4a93f81",
          4498 => x"d3d80855",
          4499 => x"7481d3d8",
          4500 => x"0c953d0d",
          4501 => x"04ef3d0d",
          4502 => x"64568253",
          4503 => x"933dd005",
          4504 => x"52943d51",
          4505 => x"d1f43f81",
          4506 => x"d3d80855",
          4507 => x"81d3d808",
          4508 => x"80cb3876",
          4509 => x"58635293",
          4510 => x"3dd40551",
          4511 => x"c8c03f81",
          4512 => x"d3d80855",
          4513 => x"81d3d808",
          4514 => x"b4380280",
          4515 => x"c7053381",
          4516 => x"a0065486",
          4517 => x"5573a638",
          4518 => x"84162286",
          4519 => x"17227190",
          4520 => x"2b075354",
          4521 => x"961f51ff",
          4522 => x"b0c23f76",
          4523 => x"54810b83",
          4524 => x"15347651",
          4525 => x"ffb3b83f",
          4526 => x"81d3d808",
          4527 => x"557481d3",
          4528 => x"d80c933d",
          4529 => x"0d04ea3d",
          4530 => x"0d696b5c",
          4531 => x"5a805398",
          4532 => x"3dd00552",
          4533 => x"993d51d1",
          4534 => x"813f81d3",
          4535 => x"d80881d3",
          4536 => x"d8083070",
          4537 => x"81d3d808",
          4538 => x"07802551",
          4539 => x"55577980",
          4540 => x"2e818538",
          4541 => x"81707506",
          4542 => x"55557380",
          4543 => x"2e80f938",
          4544 => x"7b5d805f",
          4545 => x"80528d3d",
          4546 => x"705254ff",
          4547 => x"bea93f81",
          4548 => x"d3d80857",
          4549 => x"81d3d808",
          4550 => x"80d13874",
          4551 => x"527351c3",
          4552 => x"dc3f81d3",
          4553 => x"d8085781",
          4554 => x"d3d808bf",
          4555 => x"3881d3d8",
          4556 => x"0881d3d8",
          4557 => x"08655b59",
          4558 => x"56781881",
          4559 => x"197b1856",
          4560 => x"59557433",
          4561 => x"74348116",
          4562 => x"568a7827",
          4563 => x"ec388b56",
          4564 => x"751a5480",
          4565 => x"74347580",
          4566 => x"2e9e38ff",
          4567 => x"16701b70",
          4568 => x"33515556",
          4569 => x"73a02ee8",
          4570 => x"388e3976",
          4571 => x"842e0981",
          4572 => x"06863880",
          4573 => x"7a348057",
          4574 => x"76307078",
          4575 => x"07802551",
          4576 => x"547a802e",
          4577 => x"80c13873",
          4578 => x"802ebc38",
          4579 => x"7ba01108",
          4580 => x"5351ffb1",
          4581 => x"933f81d3",
          4582 => x"d8085781",
          4583 => x"d3d808a7",
          4584 => x"387b7033",
          4585 => x"555580c3",
          4586 => x"5673832e",
          4587 => x"8b3880e4",
          4588 => x"5673842e",
          4589 => x"8338a756",
          4590 => x"7515b405",
          4591 => x"51ffade3",
          4592 => x"3f81d3d8",
          4593 => x"087b0c76",
          4594 => x"81d3d80c",
          4595 => x"983d0d04",
          4596 => x"e63d0d82",
          4597 => x"539c3dff",
          4598 => x"b805529d",
          4599 => x"3d51cefa",
          4600 => x"3f81d3d8",
          4601 => x"0881d3d8",
          4602 => x"08565481",
          4603 => x"d3d80883",
          4604 => x"98388b53",
          4605 => x"a0528b3d",
          4606 => x"705259ff",
          4607 => x"aec03f73",
          4608 => x"6d703370",
          4609 => x"81ff0652",
          4610 => x"5755579f",
          4611 => x"742781bc",
          4612 => x"38785874",
          4613 => x"81ff066d",
          4614 => x"81054e70",
          4615 => x"5255ffaf",
          4616 => x"893f81d3",
          4617 => x"d808802e",
          4618 => x"a5386c70",
          4619 => x"33705357",
          4620 => x"54ffaefd",
          4621 => x"3f81d3d8",
          4622 => x"08802e8d",
          4623 => x"3874882b",
          4624 => x"76076d81",
          4625 => x"054e5586",
          4626 => x"3981d3d8",
          4627 => x"0855ff9f",
          4628 => x"157083ff",
          4629 => x"ff065154",
          4630 => x"7399268a",
          4631 => x"38e01570",
          4632 => x"83ffff06",
          4633 => x"565480ff",
          4634 => x"75278738",
          4635 => x"81c2dc15",
          4636 => x"33557480",
          4637 => x"2ea33874",
          4638 => x"5281c4dc",
          4639 => x"51ffae89",
          4640 => x"3f81d3d8",
          4641 => x"08933881",
          4642 => x"ff752788",
          4643 => x"38768926",
          4644 => x"88388b39",
          4645 => x"8a772786",
          4646 => x"38865581",
          4647 => x"ec3981ff",
          4648 => x"75278f38",
          4649 => x"74882a54",
          4650 => x"73787081",
          4651 => x"055a3481",
          4652 => x"17577478",
          4653 => x"7081055a",
          4654 => x"3481176d",
          4655 => x"70337081",
          4656 => x"ff065257",
          4657 => x"5557739f",
          4658 => x"26fec838",
          4659 => x"8b3d3354",
          4660 => x"86557381",
          4661 => x"e52e81b1",
          4662 => x"3876802e",
          4663 => x"993802a7",
          4664 => x"05557615",
          4665 => x"70335154",
          4666 => x"73a02e09",
          4667 => x"81068738",
          4668 => x"ff175776",
          4669 => x"ed387941",
          4670 => x"80438052",
          4671 => x"913d7052",
          4672 => x"55ffbab3",
          4673 => x"3f81d3d8",
          4674 => x"085481d3",
          4675 => x"d80880f7",
          4676 => x"38815274",
          4677 => x"51ffbfe5",
          4678 => x"3f81d3d8",
          4679 => x"085481d3",
          4680 => x"d8088d38",
          4681 => x"7680c438",
          4682 => x"6754e574",
          4683 => x"3480c639",
          4684 => x"81d3d808",
          4685 => x"842e0981",
          4686 => x"0680cc38",
          4687 => x"80547674",
          4688 => x"2e80c438",
          4689 => x"81527451",
          4690 => x"ffbdb03f",
          4691 => x"81d3d808",
          4692 => x"5481d3d8",
          4693 => x"08b138a0",
          4694 => x"5381d3d8",
          4695 => x"08526751",
          4696 => x"ffabdb3f",
          4697 => x"6754880b",
          4698 => x"8b15348b",
          4699 => x"53785267",
          4700 => x"51ffaba7",
          4701 => x"3f795481",
          4702 => x"0b831534",
          4703 => x"7951ffad",
          4704 => x"ee3f81d3",
          4705 => x"d8085473",
          4706 => x"557481d3",
          4707 => x"d80c9c3d",
          4708 => x"0d04f23d",
          4709 => x"0d606202",
          4710 => x"880580cb",
          4711 => x"0533933d",
          4712 => x"fc055572",
          4713 => x"54405e5a",
          4714 => x"d2da3f81",
          4715 => x"d3d80858",
          4716 => x"81d3d808",
          4717 => x"82bd3891",
          4718 => x"1a335877",
          4719 => x"82b5387c",
          4720 => x"802e9738",
          4721 => x"8c1a0859",
          4722 => x"78903890",
          4723 => x"1a337081",
          4724 => x"2a708106",
          4725 => x"51555573",
          4726 => x"90388754",
          4727 => x"82973982",
          4728 => x"58829039",
          4729 => x"8158828b",
          4730 => x"397e8a11",
          4731 => x"2270892b",
          4732 => x"70557f54",
          4733 => x"565656fe",
          4734 => x"fefd3fff",
          4735 => x"147d0670",
          4736 => x"30707207",
          4737 => x"9f2a81d3",
          4738 => x"d808058c",
          4739 => x"19087c40",
          4740 => x"5a5d5555",
          4741 => x"81772788",
          4742 => x"38981608",
          4743 => x"77268338",
          4744 => x"82577677",
          4745 => x"56598056",
          4746 => x"74527951",
          4747 => x"ffae993f",
          4748 => x"81157f55",
          4749 => x"55981408",
          4750 => x"75268338",
          4751 => x"825581d3",
          4752 => x"d808812e",
          4753 => x"ff993881",
          4754 => x"d3d808ff",
          4755 => x"2eff9538",
          4756 => x"81d3d808",
          4757 => x"8e388116",
          4758 => x"56757b2e",
          4759 => x"09810687",
          4760 => x"38933974",
          4761 => x"59805674",
          4762 => x"772e0981",
          4763 => x"06ffb938",
          4764 => x"875880ff",
          4765 => x"397d802e",
          4766 => x"ba38787b",
          4767 => x"55557a80",
          4768 => x"2eb43881",
          4769 => x"15567381",
          4770 => x"2e098106",
          4771 => x"8338ff56",
          4772 => x"75537452",
          4773 => x"7e51ffaf",
          4774 => x"a83f81d3",
          4775 => x"d8085881",
          4776 => x"d3d80880",
          4777 => x"ce387481",
          4778 => x"16ff1656",
          4779 => x"565c73d3",
          4780 => x"388439ff",
          4781 => x"195c7e7c",
          4782 => x"8c120c55",
          4783 => x"7d802eb3",
          4784 => x"3878881b",
          4785 => x"0c7c8c1b",
          4786 => x"0c901a33",
          4787 => x"80c00754",
          4788 => x"73901b34",
          4789 => x"981508fe",
          4790 => x"05901608",
          4791 => x"57547574",
          4792 => x"26913875",
          4793 => x"7b319016",
          4794 => x"0c841533",
          4795 => x"81075473",
          4796 => x"84163477",
          4797 => x"547381d3",
          4798 => x"d80c903d",
          4799 => x"0d04e93d",
          4800 => x"0d6b6d02",
          4801 => x"880580eb",
          4802 => x"05339d3d",
          4803 => x"545a5c59",
          4804 => x"c5bd3f8b",
          4805 => x"56800b81",
          4806 => x"d3d80824",
          4807 => x"8bf83881",
          4808 => x"d3d80884",
          4809 => x"2981d3f4",
          4810 => x"05700851",
          4811 => x"5574802e",
          4812 => x"84388075",
          4813 => x"3481d3d8",
          4814 => x"0881ff06",
          4815 => x"5f81527e",
          4816 => x"51ffa0d0",
          4817 => x"3f81d3d8",
          4818 => x"0881ff06",
          4819 => x"70810656",
          4820 => x"57835674",
          4821 => x"8bc03876",
          4822 => x"822a7081",
          4823 => x"0651558a",
          4824 => x"56748bb2",
          4825 => x"38993dfc",
          4826 => x"05538352",
          4827 => x"7e51ffa4",
          4828 => x"f03f81d3",
          4829 => x"d8089938",
          4830 => x"67557480",
          4831 => x"2e923874",
          4832 => x"82808026",
          4833 => x"8b38ff15",
          4834 => x"75065574",
          4835 => x"802e8338",
          4836 => x"81487880",
          4837 => x"2e873884",
          4838 => x"80792692",
          4839 => x"38788180",
          4840 => x"0a268b38",
          4841 => x"ff197906",
          4842 => x"5574802e",
          4843 => x"86389356",
          4844 => x"8ae43978",
          4845 => x"892a6e89",
          4846 => x"2a70892b",
          4847 => x"77594843",
          4848 => x"597a8338",
          4849 => x"81566130",
          4850 => x"70802577",
          4851 => x"07515591",
          4852 => x"56748ac2",
          4853 => x"38993df8",
          4854 => x"05538152",
          4855 => x"7e51ffa4",
          4856 => x"803f8156",
          4857 => x"81d3d808",
          4858 => x"8aac3877",
          4859 => x"832a7077",
          4860 => x"0681d3d8",
          4861 => x"08435645",
          4862 => x"748338bf",
          4863 => x"4166558e",
          4864 => x"56607526",
          4865 => x"8a903874",
          4866 => x"61317048",
          4867 => x"5580ff75",
          4868 => x"278a8338",
          4869 => x"93567881",
          4870 => x"802689fa",
          4871 => x"3877812a",
          4872 => x"70810656",
          4873 => x"4374802e",
          4874 => x"95387787",
          4875 => x"06557482",
          4876 => x"2e838d38",
          4877 => x"77810655",
          4878 => x"74802e83",
          4879 => x"83387781",
          4880 => x"06559356",
          4881 => x"825e7480",
          4882 => x"2e89cb38",
          4883 => x"785a7d83",
          4884 => x"2e098106",
          4885 => x"80e13878",
          4886 => x"ae386691",
          4887 => x"2a57810b",
          4888 => x"81c58022",
          4889 => x"565a7480",
          4890 => x"2e9d3874",
          4891 => x"77269838",
          4892 => x"81c58056",
          4893 => x"79108217",
          4894 => x"70225757",
          4895 => x"5a74802e",
          4896 => x"86387675",
          4897 => x"27ee3879",
          4898 => x"526651fe",
          4899 => x"f9e93f81",
          4900 => x"d3d80884",
          4901 => x"29848705",
          4902 => x"70892a5e",
          4903 => x"55a05c80",
          4904 => x"0b81d3d8",
          4905 => x"08fc808a",
          4906 => x"055644fd",
          4907 => x"fff00a75",
          4908 => x"2780ec38",
          4909 => x"88d33978",
          4910 => x"ae38668c",
          4911 => x"2a57810b",
          4912 => x"81c4f022",
          4913 => x"565a7480",
          4914 => x"2e9d3874",
          4915 => x"77269838",
          4916 => x"81c4f056",
          4917 => x"79108217",
          4918 => x"70225757",
          4919 => x"5a74802e",
          4920 => x"86387675",
          4921 => x"27ee3879",
          4922 => x"526651fe",
          4923 => x"f9893f81",
          4924 => x"d3d80810",
          4925 => x"84055781",
          4926 => x"d3d8089f",
          4927 => x"f5269638",
          4928 => x"810b81d3",
          4929 => x"d8081081",
          4930 => x"d3d80805",
          4931 => x"7111722a",
          4932 => x"83055956",
          4933 => x"5e83ff17",
          4934 => x"892a5d81",
          4935 => x"5ca04460",
          4936 => x"1c7d1165",
          4937 => x"05697012",
          4938 => x"ff057130",
          4939 => x"70720674",
          4940 => x"315c5259",
          4941 => x"5759407d",
          4942 => x"832e0981",
          4943 => x"06893876",
          4944 => x"1c601841",
          4945 => x"5c843976",
          4946 => x"1d5d7990",
          4947 => x"29187062",
          4948 => x"31685851",
          4949 => x"55747626",
          4950 => x"87af3875",
          4951 => x"7c317d31",
          4952 => x"7a537065",
          4953 => x"315255fe",
          4954 => x"f88d3f81",
          4955 => x"d3d80858",
          4956 => x"7d832e09",
          4957 => x"81069b38",
          4958 => x"81d3d808",
          4959 => x"83fff526",
          4960 => x"80dd3878",
          4961 => x"87833879",
          4962 => x"812a5978",
          4963 => x"fdbe3886",
          4964 => x"f8397d82",
          4965 => x"2e098106",
          4966 => x"80c53883",
          4967 => x"fff50b81",
          4968 => x"d3d80827",
          4969 => x"a038788f",
          4970 => x"38791a55",
          4971 => x"7480c026",
          4972 => x"86387459",
          4973 => x"fd963962",
          4974 => x"81065574",
          4975 => x"802e8f38",
          4976 => x"835efd88",
          4977 => x"3981d3d8",
          4978 => x"089ff526",
          4979 => x"92387886",
          4980 => x"b838791a",
          4981 => x"59818079",
          4982 => x"27fcf138",
          4983 => x"86ab3980",
          4984 => x"557d812e",
          4985 => x"09810683",
          4986 => x"387d559f",
          4987 => x"f578278b",
          4988 => x"38748106",
          4989 => x"558e5674",
          4990 => x"869c3884",
          4991 => x"80538052",
          4992 => x"7a51ffa2",
          4993 => x"b93f8b53",
          4994 => x"81c39852",
          4995 => x"7a51ffa2",
          4996 => x"8a3f8480",
          4997 => x"528b1b51",
          4998 => x"ffa1b33f",
          4999 => x"798d1c34",
          5000 => x"7b83ffff",
          5001 => x"06528e1b",
          5002 => x"51ffa1a2",
          5003 => x"3f810b90",
          5004 => x"1c347d83",
          5005 => x"32703070",
          5006 => x"962a8480",
          5007 => x"06545155",
          5008 => x"911b51ff",
          5009 => x"a1883f66",
          5010 => x"557483ff",
          5011 => x"ff269038",
          5012 => x"7483ffff",
          5013 => x"0652931b",
          5014 => x"51ffa0f2",
          5015 => x"3f8a3974",
          5016 => x"52a01b51",
          5017 => x"ffa1853f",
          5018 => x"f80b951c",
          5019 => x"34bf5298",
          5020 => x"1b51ffa0",
          5021 => x"d93f81ff",
          5022 => x"529a1b51",
          5023 => x"ffa0cf3f",
          5024 => x"60529c1b",
          5025 => x"51ffa0e4",
          5026 => x"3f7d832e",
          5027 => x"09810680",
          5028 => x"cb388288",
          5029 => x"b20a5280",
          5030 => x"c31b51ff",
          5031 => x"a0ce3f7c",
          5032 => x"52a41b51",
          5033 => x"ffa0c53f",
          5034 => x"8252ac1b",
          5035 => x"51ffa0bc",
          5036 => x"3f8152b0",
          5037 => x"1b51ffa0",
          5038 => x"953f8652",
          5039 => x"b21b51ff",
          5040 => x"a08c3fff",
          5041 => x"800b80c0",
          5042 => x"1c34a90b",
          5043 => x"80c21c34",
          5044 => x"935381c3",
          5045 => x"a45280c7",
          5046 => x"1b51ae39",
          5047 => x"8288b20a",
          5048 => x"52a71b51",
          5049 => x"ffa0853f",
          5050 => x"7c83ffff",
          5051 => x"0652961b",
          5052 => x"51ff9fda",
          5053 => x"3fff800b",
          5054 => x"a41c34a9",
          5055 => x"0ba61c34",
          5056 => x"935381c3",
          5057 => x"b852ab1b",
          5058 => x"51ffa08f",
          5059 => x"3f82d4d5",
          5060 => x"5283fe1b",
          5061 => x"705259ff",
          5062 => x"9fb43f81",
          5063 => x"5460537a",
          5064 => x"527e51ff",
          5065 => x"9bd73f81",
          5066 => x"5681d3d8",
          5067 => x"0883e738",
          5068 => x"7d832e09",
          5069 => x"810680ee",
          5070 => x"38755460",
          5071 => x"8605537a",
          5072 => x"527e51ff",
          5073 => x"9bb73f84",
          5074 => x"80538052",
          5075 => x"7a51ff9f",
          5076 => x"ed3f848b",
          5077 => x"85a4d252",
          5078 => x"7a51ff9f",
          5079 => x"8f3f868a",
          5080 => x"85e4f252",
          5081 => x"83e41b51",
          5082 => x"ff9f813f",
          5083 => x"ff185283",
          5084 => x"e81b51ff",
          5085 => x"9ef63f82",
          5086 => x"5283ec1b",
          5087 => x"51ff9eec",
          5088 => x"3f82d4d5",
          5089 => x"527851ff",
          5090 => x"9ec43f75",
          5091 => x"54608705",
          5092 => x"537a527e",
          5093 => x"51ff9ae5",
          5094 => x"3f755460",
          5095 => x"16537a52",
          5096 => x"7e51ff9a",
          5097 => x"d83f6553",
          5098 => x"80527a51",
          5099 => x"ff9f8f3f",
          5100 => x"7f568058",
          5101 => x"7d832e09",
          5102 => x"81069a38",
          5103 => x"f8527a51",
          5104 => x"ff9ea93f",
          5105 => x"ff52841b",
          5106 => x"51ff9ea0",
          5107 => x"3ff00a52",
          5108 => x"881b5191",
          5109 => x"3987ffff",
          5110 => x"f8557d81",
          5111 => x"2e8338f8",
          5112 => x"5574527a",
          5113 => x"51ff9e84",
          5114 => x"3f7c5561",
          5115 => x"57746226",
          5116 => x"83387457",
          5117 => x"76547553",
          5118 => x"7a527e51",
          5119 => x"ff99fe3f",
          5120 => x"81d3d808",
          5121 => x"82873884",
          5122 => x"805381d3",
          5123 => x"d808527a",
          5124 => x"51ff9eaa",
          5125 => x"3f761675",
          5126 => x"78315656",
          5127 => x"74cd3881",
          5128 => x"18587780",
          5129 => x"2eff8d38",
          5130 => x"79557d83",
          5131 => x"2e833863",
          5132 => x"55615774",
          5133 => x"62268338",
          5134 => x"74577654",
          5135 => x"75537a52",
          5136 => x"7e51ff99",
          5137 => x"b83f81d3",
          5138 => x"d80881c1",
          5139 => x"38761675",
          5140 => x"78315656",
          5141 => x"74db388c",
          5142 => x"567d832e",
          5143 => x"93388656",
          5144 => x"6683ffff",
          5145 => x"268a3884",
          5146 => x"567d822e",
          5147 => x"83388156",
          5148 => x"64810658",
          5149 => x"7780fe38",
          5150 => x"84805377",
          5151 => x"527a51ff",
          5152 => x"9dbc3f82",
          5153 => x"d4d55278",
          5154 => x"51ff9cc2",
          5155 => x"3f83be1b",
          5156 => x"55777534",
          5157 => x"810b8116",
          5158 => x"34810b82",
          5159 => x"16347783",
          5160 => x"16347584",
          5161 => x"16346067",
          5162 => x"055680fd",
          5163 => x"c1527551",
          5164 => x"fef1c43f",
          5165 => x"fe0b8516",
          5166 => x"3481d3d8",
          5167 => x"08822abf",
          5168 => x"07567586",
          5169 => x"163481d3",
          5170 => x"d8088716",
          5171 => x"34605283",
          5172 => x"c61b51ff",
          5173 => x"9c963f66",
          5174 => x"5283ca1b",
          5175 => x"51ff9c8c",
          5176 => x"3f815477",
          5177 => x"537a527e",
          5178 => x"51ff9891",
          5179 => x"3f815681",
          5180 => x"d3d808a2",
          5181 => x"38805380",
          5182 => x"527e51ff",
          5183 => x"99e33f81",
          5184 => x"5681d3d8",
          5185 => x"08903889",
          5186 => x"398e568a",
          5187 => x"39815686",
          5188 => x"3981d3d8",
          5189 => x"08567581",
          5190 => x"d3d80c99",
          5191 => x"3d0d04f5",
          5192 => x"3d0d7d60",
          5193 => x"5b598079",
          5194 => x"60ff055a",
          5195 => x"57577678",
          5196 => x"25b4388d",
          5197 => x"3df81155",
          5198 => x"558153fc",
          5199 => x"15527951",
          5200 => x"c9dc3f7a",
          5201 => x"812e0981",
          5202 => x"069c388c",
          5203 => x"3d335574",
          5204 => x"8d2edb38",
          5205 => x"74767081",
          5206 => x"05583481",
          5207 => x"1757748a",
          5208 => x"2e098106",
          5209 => x"c9388076",
          5210 => x"34785576",
          5211 => x"83387655",
          5212 => x"7481d3d8",
          5213 => x"0c8d3d0d",
          5214 => x"04ff3d0d",
          5215 => x"73527193",
          5216 => x"26818e38",
          5217 => x"71842981",
          5218 => x"bde40552",
          5219 => x"71080481",
          5220 => x"c6885181",
          5221 => x"803981c6",
          5222 => x"945180f9",
          5223 => x"3981c6a8",
          5224 => x"5180f239",
          5225 => x"81c6bc51",
          5226 => x"80eb3981",
          5227 => x"c6cc5180",
          5228 => x"e43981c6",
          5229 => x"dc5180dd",
          5230 => x"3981c6f0",
          5231 => x"5180d639",
          5232 => x"81c78051",
          5233 => x"80cf3981",
          5234 => x"c7985180",
          5235 => x"c83981c7",
          5236 => x"b05180c1",
          5237 => x"3981c7c8",
          5238 => x"51bb3981",
          5239 => x"c7e451b5",
          5240 => x"3981c7f8",
          5241 => x"51af3981",
          5242 => x"c8a451a9",
          5243 => x"3981c8b8",
          5244 => x"51a33981",
          5245 => x"c8d8519d",
          5246 => x"3981c8ec",
          5247 => x"51973981",
          5248 => x"c9845191",
          5249 => x"3981c99c",
          5250 => x"518b3981",
          5251 => x"c9b45185",
          5252 => x"3981c9c0",
          5253 => x"51ff87a1",
          5254 => x"3f833d0d",
          5255 => x"04fb3d0d",
          5256 => x"77795656",
          5257 => x"7487e726",
          5258 => x"8a387452",
          5259 => x"7587e829",
          5260 => x"51913987",
          5261 => x"e8527451",
          5262 => x"feeebc3f",
          5263 => x"81d3d808",
          5264 => x"527551fe",
          5265 => x"eeb13f81",
          5266 => x"d3d80854",
          5267 => x"79537552",
          5268 => x"81c9d051",
          5269 => x"ff8cc63f",
          5270 => x"873d0d04",
          5271 => x"f53d0d7d",
          5272 => x"7f61028c",
          5273 => x"0580c705",
          5274 => x"33737315",
          5275 => x"665f5d5a",
          5276 => x"5a5c5c5c",
          5277 => x"785281c9",
          5278 => x"f451ff8c",
          5279 => x"a03f81c9",
          5280 => x"fc51ff86",
          5281 => x"b43f8055",
          5282 => x"74772780",
          5283 => x"fc387990",
          5284 => x"2e893879",
          5285 => x"a02ea738",
          5286 => x"80c63974",
          5287 => x"16537278",
          5288 => x"278e3872",
          5289 => x"225281ca",
          5290 => x"8051ff8b",
          5291 => x"f03f8939",
          5292 => x"81ca8c51",
          5293 => x"ff86823f",
          5294 => x"82155580",
          5295 => x"c3397416",
          5296 => x"53727827",
          5297 => x"8e387208",
          5298 => x"5281c9f4",
          5299 => x"51ff8bcd",
          5300 => x"3f893981",
          5301 => x"ca8851ff",
          5302 => x"85df3f84",
          5303 => x"1555a139",
          5304 => x"74165372",
          5305 => x"78278e38",
          5306 => x"72335281",
          5307 => x"ca9451ff",
          5308 => x"8bab3f89",
          5309 => x"3981ca9c",
          5310 => x"51ff85bd",
          5311 => x"3f811555",
          5312 => x"a051fef9",
          5313 => x"b53fff80",
          5314 => x"3981caa0",
          5315 => x"51ff85a9",
          5316 => x"3f805574",
          5317 => x"7727aa38",
          5318 => x"74167033",
          5319 => x"79722652",
          5320 => x"55539f74",
          5321 => x"27903872",
          5322 => x"802e8b38",
          5323 => x"7380fe26",
          5324 => x"85387351",
          5325 => x"8339a051",
          5326 => x"fef8ff3f",
          5327 => x"811555d3",
          5328 => x"3981caa4",
          5329 => x"51ff84f1",
          5330 => x"3f761677",
          5331 => x"1a5a56fe",
          5332 => x"fcba3f81",
          5333 => x"d3d80898",
          5334 => x"2b70982c",
          5335 => x"515574a0",
          5336 => x"2e098106",
          5337 => x"a538fefc",
          5338 => x"a33f81d3",
          5339 => x"d808982b",
          5340 => x"70982c70",
          5341 => x"a0327030",
          5342 => x"7072079f",
          5343 => x"2a515656",
          5344 => x"5155749b",
          5345 => x"2e8c3872",
          5346 => x"dd38749b",
          5347 => x"2e098106",
          5348 => x"85388053",
          5349 => x"8c397a1c",
          5350 => x"53727626",
          5351 => x"fdd638ff",
          5352 => x"537281d3",
          5353 => x"d80c8d3d",
          5354 => x"0d04ec3d",
          5355 => x"0d660284",
          5356 => x"0580e305",
          5357 => x"33697230",
          5358 => x"70740780",
          5359 => x"257087ff",
          5360 => x"74270751",
          5361 => x"51585a5b",
          5362 => x"56935774",
          5363 => x"80fc3881",
          5364 => x"5375528c",
          5365 => x"3d705257",
          5366 => x"ffbfde3f",
          5367 => x"81d3d808",
          5368 => x"5681d3d8",
          5369 => x"08b83881",
          5370 => x"d3d80887",
          5371 => x"c098880c",
          5372 => x"81d3d808",
          5373 => x"59963dd4",
          5374 => x"05548480",
          5375 => x"53775276",
          5376 => x"51c49b3f",
          5377 => x"81d3d808",
          5378 => x"5681d3d8",
          5379 => x"0890387a",
          5380 => x"5574802e",
          5381 => x"89387419",
          5382 => x"75195959",
          5383 => x"d839963d",
          5384 => x"d80551cc",
          5385 => x"853f7530",
          5386 => x"70770780",
          5387 => x"25515579",
          5388 => x"802e9538",
          5389 => x"74802e90",
          5390 => x"3881caa8",
          5391 => x"5387c098",
          5392 => x"88085278",
          5393 => x"51fbd63f",
          5394 => x"75577681",
          5395 => x"d3d80c96",
          5396 => x"3d0d04f9",
          5397 => x"3d0d7b02",
          5398 => x"8405b305",
          5399 => x"335758ff",
          5400 => x"5780537a",
          5401 => x"527951fe",
          5402 => x"c13f81d3",
          5403 => x"d808a438",
          5404 => x"75802e88",
          5405 => x"3875812e",
          5406 => x"98389839",
          5407 => x"60557f54",
          5408 => x"81d3d853",
          5409 => x"7e527d51",
          5410 => x"772d81d3",
          5411 => x"d8085783",
          5412 => x"39770476",
          5413 => x"81d3d80c",
          5414 => x"893d0d04",
          5415 => x"fc3d0d02",
          5416 => x"9b053381",
          5417 => x"cab05381",
          5418 => x"cab85255",
          5419 => x"ff87ee3f",
          5420 => x"81d18422",
          5421 => x"51ff8089",
          5422 => x"3f81cac4",
          5423 => x"5481cad0",
          5424 => x"5381d185",
          5425 => x"335281ca",
          5426 => x"d851ff87",
          5427 => x"d03f7480",
          5428 => x"2e8538fe",
          5429 => x"fdb93f86",
          5430 => x"3d0d04fe",
          5431 => x"3d0d87c0",
          5432 => x"96800853",
          5433 => x"ff80a23f",
          5434 => x"8151fef5",
          5435 => x"b33f81ca",
          5436 => x"f451fef7",
          5437 => x"ab3f8051",
          5438 => x"fef5a53f",
          5439 => x"72812a70",
          5440 => x"81065152",
          5441 => x"71802e95",
          5442 => x"388151fe",
          5443 => x"f5923f81",
          5444 => x"cb9051fe",
          5445 => x"f78a3f80",
          5446 => x"51fef584",
          5447 => x"3f72822a",
          5448 => x"70810651",
          5449 => x"5271802e",
          5450 => x"95388151",
          5451 => x"fef4f13f",
          5452 => x"81cba451",
          5453 => x"fef6e93f",
          5454 => x"8051fef4",
          5455 => x"e33f7283",
          5456 => x"2a708106",
          5457 => x"51527180",
          5458 => x"2e953881",
          5459 => x"51fef4d0",
          5460 => x"3f81cbb4",
          5461 => x"51fef6c8",
          5462 => x"3f8051fe",
          5463 => x"f4c23f72",
          5464 => x"842a7081",
          5465 => x"06515271",
          5466 => x"802e9538",
          5467 => x"8151fef4",
          5468 => x"af3f81cb",
          5469 => x"c851fef6",
          5470 => x"a73f8051",
          5471 => x"fef4a13f",
          5472 => x"72852a70",
          5473 => x"81065152",
          5474 => x"71802e95",
          5475 => x"388151fe",
          5476 => x"f48e3f81",
          5477 => x"cbdc51fe",
          5478 => x"f6863f80",
          5479 => x"51fef480",
          5480 => x"3f72862a",
          5481 => x"70810651",
          5482 => x"5271802e",
          5483 => x"95388151",
          5484 => x"fef3ed3f",
          5485 => x"81cbf051",
          5486 => x"fef5e53f",
          5487 => x"8051fef3",
          5488 => x"df3f7287",
          5489 => x"2a708106",
          5490 => x"51527180",
          5491 => x"2e953881",
          5492 => x"51fef3cc",
          5493 => x"3f81cc84",
          5494 => x"51fef5c4",
          5495 => x"3f8051fe",
          5496 => x"f3be3f72",
          5497 => x"882a7081",
          5498 => x"06515271",
          5499 => x"802e9538",
          5500 => x"8151fef3",
          5501 => x"ab3f81cc",
          5502 => x"9851fef5",
          5503 => x"a33f8051",
          5504 => x"fef39d3f",
          5505 => x"fefecb3f",
          5506 => x"843d0d04",
          5507 => x"fa3d0d78",
          5508 => x"70087055",
          5509 => x"55577380",
          5510 => x"2e80f038",
          5511 => x"8e397377",
          5512 => x"0c851533",
          5513 => x"5380e439",
          5514 => x"81145480",
          5515 => x"74337081",
          5516 => x"ff065757",
          5517 => x"5374a02e",
          5518 => x"83388153",
          5519 => x"74802e84",
          5520 => x"3872e538",
          5521 => x"7581ff06",
          5522 => x"5372a02e",
          5523 => x"09810688",
          5524 => x"38807470",
          5525 => x"81055634",
          5526 => x"80567590",
          5527 => x"2981d1a8",
          5528 => x"05770853",
          5529 => x"70085255",
          5530 => x"feeda43f",
          5531 => x"81d3d808",
          5532 => x"8b388415",
          5533 => x"33537281",
          5534 => x"2effa338",
          5535 => x"81167081",
          5536 => x"ff065753",
          5537 => x"927627d2",
          5538 => x"38ff5372",
          5539 => x"81d3d80c",
          5540 => x"883d0d04",
          5541 => x"fb3d0d77",
          5542 => x"79705556",
          5543 => x"56805275",
          5544 => x"51feebda",
          5545 => x"3f81d1a4",
          5546 => x"335473a7",
          5547 => x"38815381",
          5548 => x"ccd85281",
          5549 => x"eadc51ff",
          5550 => x"b9ff3f81",
          5551 => x"d3d80830",
          5552 => x"7081d3d8",
          5553 => x"08078025",
          5554 => x"82713151",
          5555 => x"51547381",
          5556 => x"d1a43481",
          5557 => x"d1a43354",
          5558 => x"73812e09",
          5559 => x"8106ac38",
          5560 => x"81eadc53",
          5561 => x"74527551",
          5562 => x"f4b53f81",
          5563 => x"d3d80880",
          5564 => x"2e8c3881",
          5565 => x"d3d80851",
          5566 => x"fefdbe3f",
          5567 => x"8e3981ea",
          5568 => x"dc51c6a6",
          5569 => x"3f820b81",
          5570 => x"d1a43481",
          5571 => x"d1a43354",
          5572 => x"73822e09",
          5573 => x"81068938",
          5574 => x"74527551",
          5575 => x"ff83d83f",
          5576 => x"800b81d3",
          5577 => x"d80c873d",
          5578 => x"0d04cb3d",
          5579 => x"0d807071",
          5580 => x"81ead80c",
          5581 => x"5e5c8152",
          5582 => x"7b51ff88",
          5583 => x"d73f81d3",
          5584 => x"d80881ff",
          5585 => x"0659787c",
          5586 => x"2e098106",
          5587 => x"a23881cc",
          5588 => x"e852993d",
          5589 => x"705259ff",
          5590 => x"82d93f7b",
          5591 => x"53785281",
          5592 => x"d58851ff",
          5593 => x"b7f23f81",
          5594 => x"d3d8087c",
          5595 => x"2e883881",
          5596 => x"ccec518d",
          5597 => x"dd398170",
          5598 => x"5e5c81cd",
          5599 => x"a451fefc",
          5600 => x"b83f993d",
          5601 => x"70465a80",
          5602 => x"f8527951",
          5603 => x"fe863fb7",
          5604 => x"3dfef805",
          5605 => x"51fcf53f",
          5606 => x"81d3d808",
          5607 => x"902b7090",
          5608 => x"2c515978",
          5609 => x"80c32e89",
          5610 => x"a8387880",
          5611 => x"c32480d6",
          5612 => x"3878ab2e",
          5613 => x"83b63878",
          5614 => x"ab24a438",
          5615 => x"78822e81",
          5616 => x"a9387882",
          5617 => x"248a3878",
          5618 => x"802effae",
          5619 => x"388c8939",
          5620 => x"78842e81",
          5621 => x"fc387894",
          5622 => x"2e82a738",
          5623 => x"8bfa3978",
          5624 => x"80c02e84",
          5625 => x"97387880",
          5626 => x"c0248a38",
          5627 => x"78b02e83",
          5628 => x"a3388be4",
          5629 => x"397880c1",
          5630 => x"2e85fe38",
          5631 => x"7880c22e",
          5632 => x"879f388b",
          5633 => x"d3397880",
          5634 => x"f82e8ac1",
          5635 => x"387880f8",
          5636 => x"24a93878",
          5637 => x"80d12e89",
          5638 => x"e9387880",
          5639 => x"d1248b38",
          5640 => x"7880d02e",
          5641 => x"89cb388b",
          5642 => x"af397880",
          5643 => x"d42e89e3",
          5644 => x"387880d5",
          5645 => x"2e89f938",
          5646 => x"8b9e3978",
          5647 => x"81832e8b",
          5648 => x"83387881",
          5649 => x"83249238",
          5650 => x"7880f92e",
          5651 => x"8aa43878",
          5652 => x"81822e8a",
          5653 => x"e0388b80",
          5654 => x"39788185",
          5655 => x"2e8af238",
          5656 => x"7881872e",
          5657 => x"fe94388a",
          5658 => x"ef39b73d",
          5659 => x"fef41153",
          5660 => x"fef80551",
          5661 => x"ff829b3f",
          5662 => x"81d3d808",
          5663 => x"883881cd",
          5664 => x"a8518bce",
          5665 => x"39b73dfe",
          5666 => x"f01153fe",
          5667 => x"f80551ff",
          5668 => x"82803f81",
          5669 => x"d3d80880",
          5670 => x"2e883881",
          5671 => x"63258338",
          5672 => x"80430280",
          5673 => x"cb053352",
          5674 => x"0280cf05",
          5675 => x"3351ff85",
          5676 => x"e33f81d3",
          5677 => x"d80881ff",
          5678 => x"0659788e",
          5679 => x"3881cdb8",
          5680 => x"51fef9f5",
          5681 => x"3f815dfd",
          5682 => x"b13981cd",
          5683 => x"c85188d9",
          5684 => x"39b73dfe",
          5685 => x"f41153fe",
          5686 => x"f80551ff",
          5687 => x"81b43f81",
          5688 => x"d3d80880",
          5689 => x"2efd9338",
          5690 => x"80538052",
          5691 => x"0280cf05",
          5692 => x"3351ff89",
          5693 => x"ec3f81d3",
          5694 => x"d8085281",
          5695 => x"cde05189",
          5696 => x"ad39b73d",
          5697 => x"fef41153",
          5698 => x"fef80551",
          5699 => x"ff81833f",
          5700 => x"81d3d808",
          5701 => x"802e8738",
          5702 => x"638926fc",
          5703 => x"dd38b73d",
          5704 => x"fef01153",
          5705 => x"fef80551",
          5706 => x"ff80e73f",
          5707 => x"81d3d808",
          5708 => x"863881d3",
          5709 => x"d8084363",
          5710 => x"5381cde8",
          5711 => x"527951fe",
          5712 => x"fef13f02",
          5713 => x"80cb0533",
          5714 => x"53795263",
          5715 => x"84b42981",
          5716 => x"d5880551",
          5717 => x"ffb4813f",
          5718 => x"81d3d808",
          5719 => x"81933881",
          5720 => x"cdb851fe",
          5721 => x"f8d33f81",
          5722 => x"5cfc8f39",
          5723 => x"b73dfef8",
          5724 => x"0551fee8",
          5725 => x"dc3f81d3",
          5726 => x"d808b83d",
          5727 => x"fef80552",
          5728 => x"5bfee9af",
          5729 => x"3f815381",
          5730 => x"d3d80852",
          5731 => x"7a51f49a",
          5732 => x"3f80d539",
          5733 => x"b73dfef8",
          5734 => x"0551fee8",
          5735 => x"b43f81d3",
          5736 => x"d808b83d",
          5737 => x"fef80552",
          5738 => x"5bfee987",
          5739 => x"3f81d3d8",
          5740 => x"08b83dfe",
          5741 => x"f805525a",
          5742 => x"fee8f83f",
          5743 => x"81d3d808",
          5744 => x"b83dfef8",
          5745 => x"055259fe",
          5746 => x"e8e93f81",
          5747 => x"d0e05881",
          5748 => x"d48c5780",
          5749 => x"56805581",
          5750 => x"d3d80881",
          5751 => x"ff065478",
          5752 => x"5379527a",
          5753 => x"51f4ec3f",
          5754 => x"81d3d808",
          5755 => x"802efb8a",
          5756 => x"3881d3d8",
          5757 => x"0851ef81",
          5758 => x"3ffaff39",
          5759 => x"b73dfef4",
          5760 => x"1153fef8",
          5761 => x"0551feff",
          5762 => x"893f81d3",
          5763 => x"d80880c4",
          5764 => x"3881d18d",
          5765 => x"33597880",
          5766 => x"2e883881",
          5767 => x"d0e00844",
          5768 => x"b33981d1",
          5769 => x"8e335978",
          5770 => x"802e8838",
          5771 => x"81d0e808",
          5772 => x"44a23981",
          5773 => x"d18f3359",
          5774 => x"788b3881",
          5775 => x"d1903359",
          5776 => x"78802e88",
          5777 => x"3881d0f0",
          5778 => x"08448939",
          5779 => x"81d18008",
          5780 => x"fc800544",
          5781 => x"b73dfef0",
          5782 => x"1153fef8",
          5783 => x"0551fefe",
          5784 => x"b13f81d3",
          5785 => x"d80880c3",
          5786 => x"3881d18d",
          5787 => x"33597880",
          5788 => x"2e883881",
          5789 => x"d0e40843",
          5790 => x"b23981d1",
          5791 => x"8e335978",
          5792 => x"802e8838",
          5793 => x"81d0ec08",
          5794 => x"43a13981",
          5795 => x"d18f3359",
          5796 => x"788b3881",
          5797 => x"d1903359",
          5798 => x"78802e88",
          5799 => x"3881d0f4",
          5800 => x"08438839",
          5801 => x"81d18008",
          5802 => x"880543b7",
          5803 => x"3dfeec11",
          5804 => x"53fef805",
          5805 => x"51fefdda",
          5806 => x"3f81d3d8",
          5807 => x"08802e9b",
          5808 => x"3880625b",
          5809 => x"5979882e",
          5810 => x"83388159",
          5811 => x"79902e8d",
          5812 => x"3878802e",
          5813 => x"883879a0",
          5814 => x"2e833888",
          5815 => x"4281cdec",
          5816 => x"51fef5d5",
          5817 => x"3fa05563",
          5818 => x"54615362",
          5819 => x"526351ee",
          5820 => x"eb3f81cd",
          5821 => x"fc5184b1",
          5822 => x"39b73dfe",
          5823 => x"f41153fe",
          5824 => x"f80551fe",
          5825 => x"fd8c3f81",
          5826 => x"d3d80880",
          5827 => x"2ef8eb38",
          5828 => x"b73dfef0",
          5829 => x"1153fef8",
          5830 => x"0551fefc",
          5831 => x"f53f81d3",
          5832 => x"d808802e",
          5833 => x"a5386359",
          5834 => x"0280cb05",
          5835 => x"33793463",
          5836 => x"810544b7",
          5837 => x"3dfef011",
          5838 => x"53fef805",
          5839 => x"51fefcd2",
          5840 => x"3f81d3d8",
          5841 => x"08e038f8",
          5842 => x"b1396370",
          5843 => x"33545281",
          5844 => x"ce8851fe",
          5845 => x"fac73f80",
          5846 => x"f8527951",
          5847 => x"fefb983f",
          5848 => x"79457933",
          5849 => x"5978ae2e",
          5850 => x"f890389f",
          5851 => x"7927a038",
          5852 => x"b73dfef0",
          5853 => x"1153fef8",
          5854 => x"0551fefc",
          5855 => x"953f81d3",
          5856 => x"d808802e",
          5857 => x"91386359",
          5858 => x"0280cb05",
          5859 => x"33793463",
          5860 => x"810544ff",
          5861 => x"b53981ce",
          5862 => x"9451fef4",
          5863 => x"9c3fffaa",
          5864 => x"39b73dfe",
          5865 => x"e81153fe",
          5866 => x"f80551fe",
          5867 => x"fdd63f81",
          5868 => x"d3d80880",
          5869 => x"2ef7c338",
          5870 => x"b73dfee4",
          5871 => x"1153fef8",
          5872 => x"0551fefd",
          5873 => x"bf3f81d3",
          5874 => x"d808802e",
          5875 => x"a6386059",
          5876 => x"02be0522",
          5877 => x"79708205",
          5878 => x"5b237841",
          5879 => x"b73dfee4",
          5880 => x"1153fef8",
          5881 => x"0551fefd",
          5882 => x"9b3f81d3",
          5883 => x"d808df38",
          5884 => x"f7883960",
          5885 => x"70225452",
          5886 => x"81ce9c51",
          5887 => x"fef99e3f",
          5888 => x"80f85279",
          5889 => x"51fef9ef",
          5890 => x"3f794579",
          5891 => x"335978ae",
          5892 => x"2ef6e738",
          5893 => x"789f2687",
          5894 => x"38608405",
          5895 => x"41d539b7",
          5896 => x"3dfee411",
          5897 => x"53fef805",
          5898 => x"51fefcd8",
          5899 => x"3f81d3d8",
          5900 => x"08802e92",
          5901 => x"38605902",
          5902 => x"be052279",
          5903 => x"7082055b",
          5904 => x"237841ff",
          5905 => x"ae3981ce",
          5906 => x"9451fef2",
          5907 => x"ec3fffa3",
          5908 => x"39b73dfe",
          5909 => x"e81153fe",
          5910 => x"f80551fe",
          5911 => x"fca63f81",
          5912 => x"d3d80880",
          5913 => x"2ef69338",
          5914 => x"b73dfee4",
          5915 => x"1153fef8",
          5916 => x"0551fefc",
          5917 => x"8f3f81d3",
          5918 => x"d808802e",
          5919 => x"a1386060",
          5920 => x"710c5960",
          5921 => x"840541b7",
          5922 => x"3dfee411",
          5923 => x"53fef805",
          5924 => x"51fefbf0",
          5925 => x"3f81d3d8",
          5926 => x"08e438f5",
          5927 => x"dd396070",
          5928 => x"08545281",
          5929 => x"cea851fe",
          5930 => x"f7f33f80",
          5931 => x"f8527951",
          5932 => x"fef8c43f",
          5933 => x"79457933",
          5934 => x"5978ae2e",
          5935 => x"f5bc389f",
          5936 => x"79279c38",
          5937 => x"b73dfee4",
          5938 => x"1153fef8",
          5939 => x"0551fefb",
          5940 => x"b33f81d3",
          5941 => x"d808802e",
          5942 => x"8d386060",
          5943 => x"710c5960",
          5944 => x"840541ff",
          5945 => x"b93981ce",
          5946 => x"9451fef1",
          5947 => x"cc3fffae",
          5948 => x"3981ceb4",
          5949 => x"51fef1c1",
          5950 => x"3f8251fe",
          5951 => x"f0af3ff4",
          5952 => x"f93981ce",
          5953 => x"cc51fef1",
          5954 => x"b03fa251",
          5955 => x"fef0823f",
          5956 => x"f4e83984",
          5957 => x"80810b87",
          5958 => x"c094840c",
          5959 => x"8480810b",
          5960 => x"87c09494",
          5961 => x"0c81cee4",
          5962 => x"51fef18d",
          5963 => x"3ff4cb39",
          5964 => x"81cef851",
          5965 => x"fef1823f",
          5966 => x"8c80830b",
          5967 => x"87c09484",
          5968 => x"0c8c8083",
          5969 => x"0b87c094",
          5970 => x"940cf4ae",
          5971 => x"39b73dfe",
          5972 => x"f41153fe",
          5973 => x"f80551fe",
          5974 => x"f8b83f81",
          5975 => x"d3d80880",
          5976 => x"2ef49738",
          5977 => x"635281cf",
          5978 => x"8c51fef6",
          5979 => x"b03f6359",
          5980 => x"7804b73d",
          5981 => x"fef41153",
          5982 => x"fef80551",
          5983 => x"fef8933f",
          5984 => x"81d3d808",
          5985 => x"802ef3f2",
          5986 => x"38635281",
          5987 => x"cfa851fe",
          5988 => x"f68b3f63",
          5989 => x"59782d81",
          5990 => x"d3d8085e",
          5991 => x"81d3d808",
          5992 => x"802ef3d6",
          5993 => x"3881d3d8",
          5994 => x"085281cf",
          5995 => x"c451fef5",
          5996 => x"ec3ff3c6",
          5997 => x"3981cfe0",
          5998 => x"51feeffd",
          5999 => x"3ffec4c0",
          6000 => x"3ff3b739",
          6001 => x"81cffc51",
          6002 => x"feefee3f",
          6003 => x"8059ffa0",
          6004 => x"39feebbb",
          6005 => x"3ff3a339",
          6006 => x"64703351",
          6007 => x"5978802e",
          6008 => x"f398387b",
          6009 => x"802e80d2",
          6010 => x"387c802e",
          6011 => x"80cc38b7",
          6012 => x"3dfef805",
          6013 => x"51fedfd9",
          6014 => x"3f81d090",
          6015 => x"5681d3d8",
          6016 => x"085581d0",
          6017 => x"94548053",
          6018 => x"81d09852",
          6019 => x"a33d7052",
          6020 => x"5afef59f",
          6021 => x"3f81d0e0",
          6022 => x"5881d48c",
          6023 => x"57805664",
          6024 => x"81114681",
          6025 => x"05558054",
          6026 => x"82808053",
          6027 => x"82808052",
          6028 => x"7951ec9f",
          6029 => x"3f81d3d8",
          6030 => x"085e7c81",
          6031 => x"327c8132",
          6032 => x"0759788a",
          6033 => x"387dff2e",
          6034 => x"098106f2",
          6035 => x"ad3881d0",
          6036 => x"a851fef4",
          6037 => x"c83ff2a2",
          6038 => x"39803d0d",
          6039 => x"800b81d4",
          6040 => x"8c349b90",
          6041 => x"86e40b87",
          6042 => x"c0948c0c",
          6043 => x"9b9086e4",
          6044 => x"0b87c094",
          6045 => x"9c0c8c80",
          6046 => x"830b87c0",
          6047 => x"94840c8c",
          6048 => x"80830b87",
          6049 => x"c094940c",
          6050 => x"9fba0b81",
          6051 => x"d3e80ca2",
          6052 => x"bb0b81d3",
          6053 => x"ec0cfee6",
          6054 => x"cb3ffeec",
          6055 => x"ec3f81d0",
          6056 => x"b851fee3",
          6057 => x"fb3f81d0",
          6058 => x"c451feee",
          6059 => x"8c3f81a9",
          6060 => x"db51feec",
          6061 => x"cf3f8151",
          6062 => x"ebe23ff0",
          6063 => x"ed3f8004",
          6064 => x"00ffffff",
          6065 => x"ff00ffff",
          6066 => x"ffff00ff",
          6067 => x"ffffff00",
          6068 => x"000014db",
          6069 => x"000014e1",
          6070 => x"000014e7",
          6071 => x"000014ed",
          6072 => x"000014f3",
          6073 => x"0000520b",
          6074 => x"0000518f",
          6075 => x"00005196",
          6076 => x"0000519d",
          6077 => x"000051a4",
          6078 => x"000051ab",
          6079 => x"000051b2",
          6080 => x"000051b9",
          6081 => x"000051c0",
          6082 => x"000051c7",
          6083 => x"000051ce",
          6084 => x"000051d5",
          6085 => x"000051db",
          6086 => x"000051e1",
          6087 => x"000051e7",
          6088 => x"000051ed",
          6089 => x"000051f3",
          6090 => x"000051f9",
          6091 => x"000051ff",
          6092 => x"00005205",
          6093 => x"25642f25",
          6094 => x"642f2564",
          6095 => x"2025643a",
          6096 => x"25643a25",
          6097 => x"642e2564",
          6098 => x"25640a00",
          6099 => x"536f4320",
          6100 => x"436f6e66",
          6101 => x"69677572",
          6102 => x"6174696f",
          6103 => x"6e000000",
          6104 => x"20286672",
          6105 => x"6f6d2053",
          6106 => x"6f432063",
          6107 => x"6f6e6669",
          6108 => x"67290000",
          6109 => x"3a0a4465",
          6110 => x"76696365",
          6111 => x"7320696d",
          6112 => x"706c656d",
          6113 => x"656e7465",
          6114 => x"643a0a00",
          6115 => x"20202020",
          6116 => x"494e534e",
          6117 => x"20425241",
          6118 => x"4d202853",
          6119 => x"74617274",
          6120 => x"3d253038",
          6121 => x"582c2053",
          6122 => x"697a653d",
          6123 => x"25303858",
          6124 => x"292e0a00",
          6125 => x"20202020",
          6126 => x"4252414d",
          6127 => x"20285374",
          6128 => x"6172743d",
          6129 => x"25303858",
          6130 => x"2c205369",
          6131 => x"7a653d25",
          6132 => x"30385829",
          6133 => x"2e0a0000",
          6134 => x"20202020",
          6135 => x"52414d20",
          6136 => x"28537461",
          6137 => x"72743d25",
          6138 => x"3038582c",
          6139 => x"2053697a",
          6140 => x"653d2530",
          6141 => x"3858292e",
          6142 => x"0a000000",
          6143 => x"20202020",
          6144 => x"494f4354",
          6145 => x"4c0a0000",
          6146 => x"20202020",
          6147 => x"5053320a",
          6148 => x"00000000",
          6149 => x"20202020",
          6150 => x"5350490a",
          6151 => x"00000000",
          6152 => x"20202020",
          6153 => x"53442043",
          6154 => x"61726420",
          6155 => x"28446576",
          6156 => x"69636573",
          6157 => x"3d253032",
          6158 => x"58292e0a",
          6159 => x"00000000",
          6160 => x"20202020",
          6161 => x"494e5445",
          6162 => x"52525550",
          6163 => x"5420434f",
          6164 => x"4e54524f",
          6165 => x"4c4c4552",
          6166 => x"0a000000",
          6167 => x"20202020",
          6168 => x"54494d45",
          6169 => x"52312028",
          6170 => x"54696d65",
          6171 => x"72733d25",
          6172 => x"30315829",
          6173 => x"2e0a0000",
          6174 => x"41646472",
          6175 => x"65737365",
          6176 => x"733a0a00",
          6177 => x"20202020",
          6178 => x"43505520",
          6179 => x"52657365",
          6180 => x"74205665",
          6181 => x"63746f72",
          6182 => x"20416464",
          6183 => x"72657373",
          6184 => x"203d2025",
          6185 => x"3038580a",
          6186 => x"00000000",
          6187 => x"20202020",
          6188 => x"43505520",
          6189 => x"4d656d6f",
          6190 => x"72792053",
          6191 => x"74617274",
          6192 => x"20416464",
          6193 => x"72657373",
          6194 => x"203d2025",
          6195 => x"3038580a",
          6196 => x"00000000",
          6197 => x"20202020",
          6198 => x"53746163",
          6199 => x"6b205374",
          6200 => x"61727420",
          6201 => x"41646472",
          6202 => x"65737320",
          6203 => x"20202020",
          6204 => x"203d2025",
          6205 => x"3038580a",
          6206 => x"00000000",
          6207 => x"20202020",
          6208 => x"5a505520",
          6209 => x"49642020",
          6210 => x"20202020",
          6211 => x"20202020",
          6212 => x"20202020",
          6213 => x"20202020",
          6214 => x"203d2025",
          6215 => x"3038580a",
          6216 => x"00000000",
          6217 => x"20202020",
          6218 => x"53797374",
          6219 => x"656d2043",
          6220 => x"6c6f636b",
          6221 => x"20467265",
          6222 => x"71202020",
          6223 => x"20202020",
          6224 => x"203d2025",
          6225 => x"3038580a",
          6226 => x"00000000",
          6227 => x"536d616c",
          6228 => x"6c000000",
          6229 => x"4d656469",
          6230 => x"756d0000",
          6231 => x"466c6578",
          6232 => x"00000000",
          6233 => x"45564f00",
          6234 => x"45564f6d",
          6235 => x"696e0000",
          6236 => x"556e6b6e",
          6237 => x"6f776e00",
          6238 => x"53440000",
          6239 => x"222a2b2c",
          6240 => x"3a3b3c3d",
          6241 => x"3e3f5b5d",
          6242 => x"7c7f0000",
          6243 => x"46415400",
          6244 => x"46415433",
          6245 => x"32000000",
          6246 => x"ebfe904d",
          6247 => x"53444f53",
          6248 => x"352e3000",
          6249 => x"4e4f204e",
          6250 => x"414d4520",
          6251 => x"20202046",
          6252 => x"41543332",
          6253 => x"20202000",
          6254 => x"4e4f204e",
          6255 => x"414d4520",
          6256 => x"20202046",
          6257 => x"41542020",
          6258 => x"20202000",
          6259 => x"00006178",
          6260 => x"00000000",
          6261 => x"00000000",
          6262 => x"00000000",
          6263 => x"809a4541",
          6264 => x"8e418f80",
          6265 => x"45454549",
          6266 => x"49498e8f",
          6267 => x"9092924f",
          6268 => x"994f5555",
          6269 => x"59999a9b",
          6270 => x"9c9d9e9f",
          6271 => x"41494f55",
          6272 => x"a5a5a6a7",
          6273 => x"a8a9aaab",
          6274 => x"acadaeaf",
          6275 => x"b0b1b2b3",
          6276 => x"b4b5b6b7",
          6277 => x"b8b9babb",
          6278 => x"bcbdbebf",
          6279 => x"c0c1c2c3",
          6280 => x"c4c5c6c7",
          6281 => x"c8c9cacb",
          6282 => x"cccdcecf",
          6283 => x"d0d1d2d3",
          6284 => x"d4d5d6d7",
          6285 => x"d8d9dadb",
          6286 => x"dcdddedf",
          6287 => x"e0e1e2e3",
          6288 => x"e4e5e6e7",
          6289 => x"e8e9eaeb",
          6290 => x"ecedeeef",
          6291 => x"f0f1f2f3",
          6292 => x"f4f5f6f7",
          6293 => x"f8f9fafb",
          6294 => x"fcfdfeff",
          6295 => x"2b2e2c3b",
          6296 => x"3d5b5d2f",
          6297 => x"5c222a3a",
          6298 => x"3c3e3f7c",
          6299 => x"7f000000",
          6300 => x"00010004",
          6301 => x"00100040",
          6302 => x"01000200",
          6303 => x"00000000",
          6304 => x"00010002",
          6305 => x"00040008",
          6306 => x"00100020",
          6307 => x"00000000",
          6308 => x"64696e69",
          6309 => x"74000000",
          6310 => x"64696f63",
          6311 => x"746c0000",
          6312 => x"66696e69",
          6313 => x"74000000",
          6314 => x"666c6f61",
          6315 => x"64000000",
          6316 => x"66657865",
          6317 => x"63000000",
          6318 => x"6d64756d",
          6319 => x"70000000",
          6320 => x"6d656200",
          6321 => x"6d656800",
          6322 => x"6d657700",
          6323 => x"68696400",
          6324 => x"68696500",
          6325 => x"68666400",
          6326 => x"68666500",
          6327 => x"63616c6c",
          6328 => x"00000000",
          6329 => x"6a6d7000",
          6330 => x"72657374",
          6331 => x"61727400",
          6332 => x"72657365",
          6333 => x"74000000",
          6334 => x"696e666f",
          6335 => x"00000000",
          6336 => x"74657374",
          6337 => x"00000000",
          6338 => x"4469736b",
          6339 => x"20457272",
          6340 => x"6f720a00",
          6341 => x"496e7465",
          6342 => x"726e616c",
          6343 => x"20657272",
          6344 => x"6f722e0a",
          6345 => x"00000000",
          6346 => x"4469736b",
          6347 => x"206e6f74",
          6348 => x"20726561",
          6349 => x"64792e0a",
          6350 => x"00000000",
          6351 => x"4e6f2066",
          6352 => x"696c6520",
          6353 => x"666f756e",
          6354 => x"642e0a00",
          6355 => x"4e6f2070",
          6356 => x"61746820",
          6357 => x"666f756e",
          6358 => x"642e0a00",
          6359 => x"496e7661",
          6360 => x"6c696420",
          6361 => x"66696c65",
          6362 => x"6e616d65",
          6363 => x"2e0a0000",
          6364 => x"41636365",
          6365 => x"73732064",
          6366 => x"656e6965",
          6367 => x"642e0a00",
          6368 => x"46696c65",
          6369 => x"20616c72",
          6370 => x"65616479",
          6371 => x"20657869",
          6372 => x"7374732e",
          6373 => x"0a000000",
          6374 => x"46696c65",
          6375 => x"2068616e",
          6376 => x"646c6520",
          6377 => x"696e7661",
          6378 => x"6c69642e",
          6379 => x"0a000000",
          6380 => x"53442069",
          6381 => x"73207772",
          6382 => x"69746520",
          6383 => x"70726f74",
          6384 => x"65637465",
          6385 => x"642e0a00",
          6386 => x"44726976",
          6387 => x"65206e75",
          6388 => x"6d626572",
          6389 => x"20697320",
          6390 => x"696e7661",
          6391 => x"6c69642e",
          6392 => x"0a000000",
          6393 => x"4469736b",
          6394 => x"206e6f74",
          6395 => x"20656e61",
          6396 => x"626c6564",
          6397 => x"2e0a0000",
          6398 => x"4e6f2063",
          6399 => x"6f6d7061",
          6400 => x"7469626c",
          6401 => x"65206669",
          6402 => x"6c657379",
          6403 => x"7374656d",
          6404 => x"20666f75",
          6405 => x"6e64206f",
          6406 => x"6e206469",
          6407 => x"736b2e0a",
          6408 => x"00000000",
          6409 => x"466f726d",
          6410 => x"61742061",
          6411 => x"626f7274",
          6412 => x"65642e0a",
          6413 => x"00000000",
          6414 => x"54696d65",
          6415 => x"6f75742c",
          6416 => x"206f7065",
          6417 => x"72617469",
          6418 => x"6f6e2063",
          6419 => x"616e6365",
          6420 => x"6c6c6564",
          6421 => x"2e0a0000",
          6422 => x"46696c65",
          6423 => x"20697320",
          6424 => x"6c6f636b",
          6425 => x"65642e0a",
          6426 => x"00000000",
          6427 => x"496e7375",
          6428 => x"66666963",
          6429 => x"69656e74",
          6430 => x"206d656d",
          6431 => x"6f72792e",
          6432 => x"0a000000",
          6433 => x"546f6f20",
          6434 => x"6d616e79",
          6435 => x"206f7065",
          6436 => x"6e206669",
          6437 => x"6c65732e",
          6438 => x"0a000000",
          6439 => x"50617261",
          6440 => x"6d657465",
          6441 => x"72732069",
          6442 => x"6e636f72",
          6443 => x"72656374",
          6444 => x"2e0a0000",
          6445 => x"53756363",
          6446 => x"6573732e",
          6447 => x"0a000000",
          6448 => x"556e6b6e",
          6449 => x"6f776e20",
          6450 => x"6572726f",
          6451 => x"722e0a00",
          6452 => x"0a256c75",
          6453 => x"20627974",
          6454 => x"65732025",
          6455 => x"73206174",
          6456 => x"20256c75",
          6457 => x"20627974",
          6458 => x"65732f73",
          6459 => x"65632e0a",
          6460 => x"00000000",
          6461 => x"25303858",
          6462 => x"00000000",
          6463 => x"3a202000",
          6464 => x"25303458",
          6465 => x"00000000",
          6466 => x"20202020",
          6467 => x"20202020",
          6468 => x"00000000",
          6469 => x"25303258",
          6470 => x"00000000",
          6471 => x"20200000",
          6472 => x"207c0000",
          6473 => x"7c0d0a00",
          6474 => x"72656164",
          6475 => x"00000000",
          6476 => x"5a505554",
          6477 => x"41000000",
          6478 => x"0a2a2a20",
          6479 => x"25732028",
          6480 => x"00000000",
          6481 => x"31382f30",
          6482 => x"372f3230",
          6483 => x"31390000",
          6484 => x"76312e33",
          6485 => x"00000000",
          6486 => x"205a5055",
          6487 => x"2c207265",
          6488 => x"76202530",
          6489 => x"32782920",
          6490 => x"25732025",
          6491 => x"73202a2a",
          6492 => x"0a0a0000",
          6493 => x"5a505554",
          6494 => x"4120496e",
          6495 => x"74657272",
          6496 => x"75707420",
          6497 => x"48616e64",
          6498 => x"6c65720a",
          6499 => x"00000000",
          6500 => x"54696d65",
          6501 => x"7220696e",
          6502 => x"74657272",
          6503 => x"7570740a",
          6504 => x"00000000",
          6505 => x"50533220",
          6506 => x"696e7465",
          6507 => x"72727570",
          6508 => x"740a0000",
          6509 => x"494f4354",
          6510 => x"4c205244",
          6511 => x"20696e74",
          6512 => x"65727275",
          6513 => x"70740a00",
          6514 => x"494f4354",
          6515 => x"4c205752",
          6516 => x"20696e74",
          6517 => x"65727275",
          6518 => x"70740a00",
          6519 => x"55415254",
          6520 => x"30205258",
          6521 => x"20696e74",
          6522 => x"65727275",
          6523 => x"70740a00",
          6524 => x"55415254",
          6525 => x"30205458",
          6526 => x"20696e74",
          6527 => x"65727275",
          6528 => x"70740a00",
          6529 => x"55415254",
          6530 => x"31205258",
          6531 => x"20696e74",
          6532 => x"65727275",
          6533 => x"70740a00",
          6534 => x"55415254",
          6535 => x"31205458",
          6536 => x"20696e74",
          6537 => x"65727275",
          6538 => x"70740a00",
          6539 => x"53657474",
          6540 => x"696e6720",
          6541 => x"75702074",
          6542 => x"696d6572",
          6543 => x"2e2e2e0a",
          6544 => x"00000000",
          6545 => x"456e6162",
          6546 => x"6c696e67",
          6547 => x"2074696d",
          6548 => x"65722e2e",
          6549 => x"2e0a0000",
          6550 => x"6175746f",
          6551 => x"65786563",
          6552 => x"2e626174",
          6553 => x"00000000",
          6554 => x"303a0000",
          6555 => x"4661696c",
          6556 => x"65642074",
          6557 => x"6f20696e",
          6558 => x"69746961",
          6559 => x"6c697365",
          6560 => x"20736420",
          6561 => x"63617264",
          6562 => x"20302c20",
          6563 => x"706c6561",
          6564 => x"73652069",
          6565 => x"6e697420",
          6566 => x"6d616e75",
          6567 => x"616c6c79",
          6568 => x"2e0a0000",
          6569 => x"2a200000",
          6570 => x"42616420",
          6571 => x"6469736b",
          6572 => x"20696421",
          6573 => x"0a000000",
          6574 => x"496e6974",
          6575 => x"69616c69",
          6576 => x"7365642e",
          6577 => x"0a000000",
          6578 => x"4661696c",
          6579 => x"65642074",
          6580 => x"6f20696e",
          6581 => x"69746961",
          6582 => x"6c697365",
          6583 => x"2e0a0000",
          6584 => x"72633d25",
          6585 => x"640a0000",
          6586 => x"25753a00",
          6587 => x"44756d70",
          6588 => x"204d656d",
          6589 => x"6f72790a",
          6590 => x"00000000",
          6591 => x"0a436f6d",
          6592 => x"706c6574",
          6593 => x"652e0a00",
          6594 => x"25303858",
          6595 => x"20253032",
          6596 => x"582d0000",
          6597 => x"3f3f3f0a",
          6598 => x"00000000",
          6599 => x"25303858",
          6600 => x"20253034",
          6601 => x"582d0000",
          6602 => x"25303858",
          6603 => x"20253038",
          6604 => x"582d0000",
          6605 => x"44697361",
          6606 => x"626c696e",
          6607 => x"6720696e",
          6608 => x"74657272",
          6609 => x"75707473",
          6610 => x"0a000000",
          6611 => x"456e6162",
          6612 => x"6c696e67",
          6613 => x"20696e74",
          6614 => x"65727275",
          6615 => x"7074730a",
          6616 => x"00000000",
          6617 => x"44697361",
          6618 => x"626c6564",
          6619 => x"20756172",
          6620 => x"74206669",
          6621 => x"666f0a00",
          6622 => x"456e6162",
          6623 => x"6c696e67",
          6624 => x"20756172",
          6625 => x"74206669",
          6626 => x"666f0a00",
          6627 => x"45786563",
          6628 => x"7574696e",
          6629 => x"6720636f",
          6630 => x"64652040",
          6631 => x"20253038",
          6632 => x"78202e2e",
          6633 => x"2e0a0000",
          6634 => x"43616c6c",
          6635 => x"696e6720",
          6636 => x"636f6465",
          6637 => x"20402025",
          6638 => x"30387820",
          6639 => x"2e2e2e0a",
          6640 => x"00000000",
          6641 => x"43616c6c",
          6642 => x"20726574",
          6643 => x"75726e65",
          6644 => x"6420636f",
          6645 => x"64652028",
          6646 => x"2564292e",
          6647 => x"0a000000",
          6648 => x"52657374",
          6649 => x"61727469",
          6650 => x"6e672061",
          6651 => x"70706c69",
          6652 => x"63617469",
          6653 => x"6f6e2e2e",
          6654 => x"2e0a0000",
          6655 => x"436f6c64",
          6656 => x"20726562",
          6657 => x"6f6f7469",
          6658 => x"6e672e2e",
          6659 => x"2e0a0000",
          6660 => x"5a505500",
          6661 => x"62696e00",
          6662 => x"25643a5c",
          6663 => x"25735c25",
          6664 => x"732e2573",
          6665 => x"00000000",
          6666 => x"42616420",
          6667 => x"636f6d6d",
          6668 => x"616e642e",
          6669 => x"0a000000",
          6670 => x"52756e6e",
          6671 => x"696e672e",
          6672 => x"2e2e0a00",
          6673 => x"456e6162",
          6674 => x"6c696e67",
          6675 => x"20696e74",
          6676 => x"65727275",
          6677 => x"7074732e",
          6678 => x"2e2e0a00",
          6679 => x"00000000",
          6680 => x"00000000",
          6681 => x"00007fff",
          6682 => x"00000000",
          6683 => x"00007fff",
          6684 => x"00010000",
          6685 => x"00007fff",
          6686 => x"00000000",
          6687 => x"00000000",
          6688 => x"00007800",
          6689 => x"00000000",
          6690 => x"05f5e100",
          6691 => x"00010101",
          6692 => x"01010101",
          6693 => x"80010101",
          6694 => x"01000000",
          6695 => x"00000000",
          6696 => x"01000000",
          6697 => x"00000000",
          6698 => x"00006290",
          6699 => x"01020100",
          6700 => x"00000000",
          6701 => x"00000000",
          6702 => x"00006298",
          6703 => x"01040100",
          6704 => x"00000000",
          6705 => x"00000000",
          6706 => x"000062a0",
          6707 => x"01140300",
          6708 => x"00000000",
          6709 => x"00000000",
          6710 => x"000062a8",
          6711 => x"012b0300",
          6712 => x"00000000",
          6713 => x"00000000",
          6714 => x"000062b0",
          6715 => x"01300300",
          6716 => x"00000000",
          6717 => x"00000000",
          6718 => x"000062b8",
          6719 => x"01400400",
          6720 => x"00000000",
          6721 => x"00000000",
          6722 => x"000062c0",
          6723 => x"01410400",
          6724 => x"00000000",
          6725 => x"00000000",
          6726 => x"000062c4",
          6727 => x"01420400",
          6728 => x"00000000",
          6729 => x"00000000",
          6730 => x"000062c8",
          6731 => x"01430400",
          6732 => x"00000000",
          6733 => x"00000000",
          6734 => x"000062cc",
          6735 => x"01500500",
          6736 => x"00000000",
          6737 => x"00000000",
          6738 => x"000062d0",
          6739 => x"01510500",
          6740 => x"00000000",
          6741 => x"00000000",
          6742 => x"000062d4",
          6743 => x"01540500",
          6744 => x"00000000",
          6745 => x"00000000",
          6746 => x"000062d8",
          6747 => x"01550500",
          6748 => x"00000000",
          6749 => x"00000000",
          6750 => x"000062dc",
          6751 => x"01790700",
          6752 => x"00000000",
          6753 => x"00000000",
          6754 => x"000062e4",
          6755 => x"01780700",
          6756 => x"00000000",
          6757 => x"00000000",
          6758 => x"000062e8",
          6759 => x"01820800",
          6760 => x"00000000",
          6761 => x"00000000",
          6762 => x"000062f0",
          6763 => x"01830800",
          6764 => x"00000000",
          6765 => x"00000000",
          6766 => x"000062f8",
          6767 => x"01850800",
          6768 => x"00000000",
          6769 => x"00000000",
          6770 => x"00006300",
          6771 => x"01870800",
          6772 => x"00000000",
          6773 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

