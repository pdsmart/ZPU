-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8b",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"a0",
           281 => x"38",
           282 => x"84",
           283 => x"0b",
           284 => x"e2",
           285 => x"51",
           286 => x"00",
           287 => x"88",
           288 => x"00",
           289 => x"02",
           290 => x"3d",
           291 => x"94",
           292 => x"08",
           293 => x"88",
           294 => x"82",
           295 => x"08",
           296 => x"54",
           297 => x"94",
           298 => x"08",
           299 => x"fd",
           300 => x"53",
           301 => x"05",
           302 => x"08",
           303 => x"51",
           304 => x"88",
           305 => x"0c",
           306 => x"0d",
           307 => x"94",
           308 => x"0c",
           309 => x"80",
           310 => x"fc",
           311 => x"08",
           312 => x"80",
           313 => x"94",
           314 => x"08",
           315 => x"88",
           316 => x"0b",
           317 => x"05",
           318 => x"fc",
           319 => x"38",
           320 => x"08",
           321 => x"94",
           322 => x"08",
           323 => x"05",
           324 => x"8c",
           325 => x"25",
           326 => x"08",
           327 => x"30",
           328 => x"05",
           329 => x"94",
           330 => x"0c",
           331 => x"05",
           332 => x"81",
           333 => x"f0",
           334 => x"08",
           335 => x"94",
           336 => x"0c",
           337 => x"08",
           338 => x"52",
           339 => x"05",
           340 => x"a7",
           341 => x"70",
           342 => x"05",
           343 => x"08",
           344 => x"80",
           345 => x"94",
           346 => x"08",
           347 => x"f8",
           348 => x"08",
           349 => x"70",
           350 => x"89",
           351 => x"0c",
           352 => x"02",
           353 => x"3d",
           354 => x"94",
           355 => x"0c",
           356 => x"05",
           357 => x"93",
           358 => x"88",
           359 => x"94",
           360 => x"0c",
           361 => x"08",
           362 => x"94",
           363 => x"08",
           364 => x"38",
           365 => x"05",
           366 => x"08",
           367 => x"81",
           368 => x"8c",
           369 => x"94",
           370 => x"08",
           371 => x"88",
           372 => x"08",
           373 => x"54",
           374 => x"05",
           375 => x"8c",
           376 => x"f8",
           377 => x"94",
           378 => x"0c",
           379 => x"05",
           380 => x"0c",
           381 => x"0d",
           382 => x"94",
           383 => x"0c",
           384 => x"81",
           385 => x"fc",
           386 => x"0b",
           387 => x"05",
           388 => x"8c",
           389 => x"08",
           390 => x"27",
           391 => x"08",
           392 => x"80",
           393 => x"80",
           394 => x"8c",
           395 => x"99",
           396 => x"8c",
           397 => x"94",
           398 => x"0c",
           399 => x"05",
           400 => x"08",
           401 => x"c9",
           402 => x"fc",
           403 => x"2e",
           404 => x"94",
           405 => x"08",
           406 => x"05",
           407 => x"38",
           408 => x"05",
           409 => x"8c",
           410 => x"94",
           411 => x"0c",
           412 => x"05",
           413 => x"fc",
           414 => x"94",
           415 => x"0c",
           416 => x"05",
           417 => x"94",
           418 => x"0c",
           419 => x"05",
           420 => x"94",
           421 => x"0c",
           422 => x"94",
           423 => x"08",
           424 => x"38",
           425 => x"05",
           426 => x"08",
           427 => x"51",
           428 => x"08",
           429 => x"70",
           430 => x"05",
           431 => x"08",
           432 => x"88",
           433 => x"0d",
           434 => x"ff",
           435 => x"88",
           436 => x"92",
           437 => x"0b",
           438 => x"8c",
           439 => x"87",
           440 => x"0c",
           441 => x"8c",
           442 => x"06",
           443 => x"80",
           444 => x"87",
           445 => x"08",
           446 => x"38",
           447 => x"8c",
           448 => x"80",
           449 => x"93",
           450 => x"98",
           451 => x"70",
           452 => x"38",
           453 => x"0b",
           454 => x"0b",
           455 => x"f0",
           456 => x"83",
           457 => x"fa",
           458 => x"7b",
           459 => x"56",
           460 => x"0b",
           461 => x"33",
           462 => x"55",
           463 => x"75",
           464 => x"06",
           465 => x"85",
           466 => x"98",
           467 => x"87",
           468 => x"0c",
           469 => x"c0",
           470 => x"87",
           471 => x"08",
           472 => x"70",
           473 => x"52",
           474 => x"2e",
           475 => x"c0",
           476 => x"70",
           477 => x"76",
           478 => x"53",
           479 => x"2e",
           480 => x"80",
           481 => x"71",
           482 => x"05",
           483 => x"14",
           484 => x"55",
           485 => x"51",
           486 => x"8b",
           487 => x"98",
           488 => x"70",
           489 => x"87",
           490 => x"08",
           491 => x"38",
           492 => x"c0",
           493 => x"87",
           494 => x"08",
           495 => x"51",
           496 => x"38",
           497 => x"80",
           498 => x"52",
           499 => x"09",
           500 => x"38",
           501 => x"8c",
           502 => x"72",
           503 => x"06",
           504 => x"52",
           505 => x"88",
           506 => x"fe",
           507 => x"81",
           508 => x"33",
           509 => x"07",
           510 => x"51",
           511 => x"04",
           512 => x"75",
           513 => x"82",
           514 => x"90",
           515 => x"2b",
           516 => x"33",
           517 => x"88",
           518 => x"71",
           519 => x"52",
           520 => x"54",
           521 => x"0d",
           522 => x"0d",
           523 => x"0b",
           524 => x"57",
           525 => x"27",
           526 => x"76",
           527 => x"27",
           528 => x"75",
           529 => x"82",
           530 => x"74",
           531 => x"38",
           532 => x"74",
           533 => x"83",
           534 => x"76",
           535 => x"17",
           536 => x"88",
           537 => x"55",
           538 => x"88",
           539 => x"74",
           540 => x"3f",
           541 => x"ff",
           542 => x"ad",
           543 => x"76",
           544 => x"fc",
           545 => x"87",
           546 => x"08",
           547 => x"3d",
           548 => x"fd",
           549 => x"08",
           550 => x"51",
           551 => x"88",
           552 => x"06",
           553 => x"81",
           554 => x"0c",
           555 => x"04",
           556 => x"0b",
           557 => x"f4",
           558 => x"88",
           559 => x"05",
           560 => x"80",
           561 => x"27",
           562 => x"14",
           563 => x"29",
           564 => x"05",
           565 => x"88",
           566 => x"0d",
           567 => x"0d",
           568 => x"0b",
           569 => x"9f",
           570 => x"33",
           571 => x"71",
           572 => x"81",
           573 => x"94",
           574 => x"ef",
           575 => x"90",
           576 => x"14",
           577 => x"3f",
           578 => x"ff",
           579 => x"07",
           580 => x"3d",
           581 => x"3d",
           582 => x"0b",
           583 => x"08",
           584 => x"75",
           585 => x"08",
           586 => x"2e",
           587 => x"14",
           588 => x"85",
           589 => x"b0",
           590 => x"38",
           591 => x"71",
           592 => x"81",
           593 => x"90",
           594 => x"72",
           595 => x"72",
           596 => x"38",
           597 => x"d8",
           598 => x"52",
           599 => x"14",
           600 => x"90",
           601 => x"52",
           602 => x"86",
           603 => x"fa",
           604 => x"0b",
           605 => x"f4",
           606 => x"81",
           607 => x"ff",
           608 => x"54",
           609 => x"80",
           610 => x"90",
           611 => x"72",
           612 => x"52",
           613 => x"73",
           614 => x"71",
           615 => x"81",
           616 => x"0c",
           617 => x"53",
           618 => x"83",
           619 => x"22",
           620 => x"76",
           621 => x"b5",
           622 => x"33",
           623 => x"84",
           624 => x"71",
           625 => x"51",
           626 => x"81",
           627 => x"08",
           628 => x"83",
           629 => x"88",
           630 => x"96",
           631 => x"8c",
           632 => x"08",
           633 => x"3f",
           634 => x"16",
           635 => x"23",
           636 => x"88",
           637 => x"0d",
           638 => x"0d",
           639 => x"58",
           640 => x"33",
           641 => x"2e",
           642 => x"88",
           643 => x"70",
           644 => x"39",
           645 => x"56",
           646 => x"2e",
           647 => x"84",
           648 => x"43",
           649 => x"1d",
           650 => x"33",
           651 => x"9f",
           652 => x"7b",
           653 => x"3f",
           654 => x"80",
           655 => x"d3",
           656 => x"84",
           657 => x"58",
           658 => x"55",
           659 => x"81",
           660 => x"ff",
           661 => x"ff",
           662 => x"06",
           663 => x"70",
           664 => x"7f",
           665 => x"7a",
           666 => x"81",
           667 => x"13",
           668 => x"af",
           669 => x"a0",
           670 => x"80",
           671 => x"51",
           672 => x"5d",
           673 => x"80",
           674 => x"ae",
           675 => x"06",
           676 => x"55",
           677 => x"75",
           678 => x"80",
           679 => x"79",
           680 => x"30",
           681 => x"70",
           682 => x"07",
           683 => x"51",
           684 => x"75",
           685 => x"58",
           686 => x"ab",
           687 => x"19",
           688 => x"06",
           689 => x"5a",
           690 => x"75",
           691 => x"39",
           692 => x"0c",
           693 => x"a0",
           694 => x"81",
           695 => x"1a",
           696 => x"fc",
           697 => x"08",
           698 => x"a0",
           699 => x"70",
           700 => x"e0",
           701 => x"90",
           702 => x"7c",
           703 => x"3f",
           704 => x"88",
           705 => x"38",
           706 => x"74",
           707 => x"ee",
           708 => x"33",
           709 => x"70",
           710 => x"56",
           711 => x"38",
           712 => x"1e",
           713 => x"59",
           714 => x"ff",
           715 => x"ff",
           716 => x"79",
           717 => x"5b",
           718 => x"81",
           719 => x"71",
           720 => x"56",
           721 => x"2e",
           722 => x"39",
           723 => x"92",
           724 => x"fc",
           725 => x"8e",
           726 => x"56",
           727 => x"38",
           728 => x"56",
           729 => x"8b",
           730 => x"55",
           731 => x"8b",
           732 => x"84",
           733 => x"06",
           734 => x"74",
           735 => x"56",
           736 => x"56",
           737 => x"51",
           738 => x"88",
           739 => x"0c",
           740 => x"75",
           741 => x"3d",
           742 => x"3d",
           743 => x"59",
           744 => x"83",
           745 => x"52",
           746 => x"fb",
           747 => x"88",
           748 => x"38",
           749 => x"b3",
           750 => x"83",
           751 => x"55",
           752 => x"82",
           753 => x"09",
           754 => x"ce",
           755 => x"b6",
           756 => x"76",
           757 => x"3f",
           758 => x"88",
           759 => x"76",
           760 => x"3f",
           761 => x"ff",
           762 => x"74",
           763 => x"2e",
           764 => x"54",
           765 => x"77",
           766 => x"f6",
           767 => x"08",
           768 => x"94",
           769 => x"f7",
           770 => x"08",
           771 => x"06",
           772 => x"82",
           773 => x"38",
           774 => x"88",
           775 => x"0d",
           776 => x"0d",
           777 => x"0b",
           778 => x"9f",
           779 => x"9b",
           780 => x"81",
           781 => x"56",
           782 => x"38",
           783 => x"8d",
           784 => x"57",
           785 => x"3f",
           786 => x"ff",
           787 => x"81",
           788 => x"06",
           789 => x"54",
           790 => x"74",
           791 => x"f5",
           792 => x"08",
           793 => x"3d",
           794 => x"80",
           795 => x"95",
           796 => x"51",
           797 => x"88",
           798 => x"53",
           799 => x"fe",
           800 => x"08",
           801 => x"57",
           802 => x"09",
           803 => x"38",
           804 => x"99",
           805 => x"2e",
           806 => x"56",
           807 => x"a4",
           808 => x"79",
           809 => x"f4",
           810 => x"56",
           811 => x"fd",
           812 => x"e5",
           813 => x"b3",
           814 => x"83",
           815 => x"58",
           816 => x"95",
           817 => x"51",
           818 => x"88",
           819 => x"af",
           820 => x"71",
           821 => x"05",
           822 => x"54",
           823 => x"f6",
           824 => x"08",
           825 => x"06",
           826 => x"1a",
           827 => x"33",
           828 => x"95",
           829 => x"51",
           830 => x"88",
           831 => x"23",
           832 => x"05",
           833 => x"3f",
           834 => x"ff",
           835 => x"75",
           836 => x"3d",
           837 => x"f5",
           838 => x"08",
           839 => x"f5",
           840 => x"08",
           841 => x"06",
           842 => x"79",
           843 => x"22",
           844 => x"82",
           845 => x"72",
           846 => x"59",
           847 => x"ee",
           848 => x"08",
           849 => x"88",
           850 => x"08",
           851 => x"56",
           852 => x"df",
           853 => x"38",
           854 => x"ff",
           855 => x"85",
           856 => x"89",
           857 => x"76",
           858 => x"c1",
           859 => x"34",
           860 => x"09",
           861 => x"38",
           862 => x"05",
           863 => x"3f",
           864 => x"1a",
           865 => x"8c",
           866 => x"90",
           867 => x"83",
           868 => x"8c",
           869 => x"71",
           870 => x"94",
           871 => x"80",
           872 => x"34",
           873 => x"0b",
           874 => x"80",
           875 => x"0c",
           876 => x"04",
           877 => x"0b",
           878 => x"f4",
           879 => x"54",
           880 => x"80",
           881 => x"0b",
           882 => x"98",
           883 => x"45",
           884 => x"3d",
           885 => x"ec",
           886 => x"9d",
           887 => x"54",
           888 => x"c0",
           889 => x"33",
           890 => x"2e",
           891 => x"a7",
           892 => x"84",
           893 => x"06",
           894 => x"73",
           895 => x"38",
           896 => x"39",
           897 => x"d5",
           898 => x"a0",
           899 => x"3d",
           900 => x"f3",
           901 => x"08",
           902 => x"73",
           903 => x"81",
           904 => x"34",
           905 => x"98",
           906 => x"f6",
           907 => x"7f",
           908 => x"0b",
           909 => x"59",
           910 => x"80",
           911 => x"57",
           912 => x"81",
           913 => x"16",
           914 => x"55",
           915 => x"80",
           916 => x"38",
           917 => x"81",
           918 => x"39",
           919 => x"17",
           920 => x"81",
           921 => x"16",
           922 => x"08",
           923 => x"78",
           924 => x"74",
           925 => x"2e",
           926 => x"98",
           927 => x"83",
           928 => x"57",
           929 => x"38",
           930 => x"ff",
           931 => x"2a",
           932 => x"ff",
           933 => x"79",
           934 => x"87",
           935 => x"08",
           936 => x"a4",
           937 => x"f3",
           938 => x"08",
           939 => x"27",
           940 => x"74",
           941 => x"a4",
           942 => x"f3",
           943 => x"08",
           944 => x"80",
           945 => x"38",
           946 => x"a8",
           947 => x"16",
           948 => x"06",
           949 => x"31",
           950 => x"75",
           951 => x"77",
           952 => x"98",
           953 => x"ff",
           954 => x"16",
           955 => x"51",
           956 => x"88",
           957 => x"38",
           958 => x"15",
           959 => x"77",
           960 => x"08",
           961 => x"58",
           962 => x"fe",
           963 => x"19",
           964 => x"39",
           965 => x"88",
           966 => x"0d",
           967 => x"0d",
           968 => x"8c",
           969 => x"84",
           970 => x"51",
           971 => x"88",
           972 => x"87",
           973 => x"08",
           974 => x"84",
           975 => x"51",
           976 => x"73",
           977 => x"87",
           978 => x"0c",
           979 => x"9c",
           980 => x"84",
           981 => x"51",
           982 => x"88",
           983 => x"87",
           984 => x"08",
           985 => x"84",
           986 => x"51",
           987 => x"73",
           988 => x"87",
           989 => x"0c",
           990 => x"0b",
           991 => x"84",
           992 => x"83",
           993 => x"94",
           994 => x"f8",
           995 => x"3f",
           996 => x"38",
           997 => x"fc",
           998 => x"08",
           999 => x"80",
          1000 => x"87",
          1001 => x"0c",
          1002 => x"fc",
          1003 => x"80",
          1004 => x"fc",
          1005 => x"08",
          1006 => x"54",
          1007 => x"86",
          1008 => x"55",
          1009 => x"80",
          1010 => x"80",
          1011 => x"00",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"00",
          1016 => x"54",
          1017 => x"59",
          1018 => x"4d",
          1019 => x"00",
          1020 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"70",
           281 => x"8e",
           282 => x"70",
           283 => x"0c",
           284 => x"88",
           285 => x"fe",
           286 => x"04",
           287 => x"00",
           288 => x"00",
           289 => x"08",
           290 => x"fd",
           291 => x"53",
           292 => x"05",
           293 => x"08",
           294 => x"51",
           295 => x"88",
           296 => x"0c",
           297 => x"0d",
           298 => x"94",
           299 => x"0c",
           300 => x"81",
           301 => x"8c",
           302 => x"94",
           303 => x"08",
           304 => x"3f",
           305 => x"88",
           306 => x"3d",
           307 => x"04",
           308 => x"94",
           309 => x"0d",
           310 => x"08",
           311 => x"94",
           312 => x"08",
           313 => x"38",
           314 => x"05",
           315 => x"08",
           316 => x"80",
           317 => x"f4",
           318 => x"08",
           319 => x"88",
           320 => x"94",
           321 => x"0c",
           322 => x"05",
           323 => x"fc",
           324 => x"08",
           325 => x"80",
           326 => x"94",
           327 => x"08",
           328 => x"8c",
           329 => x"0b",
           330 => x"05",
           331 => x"fc",
           332 => x"38",
           333 => x"08",
           334 => x"94",
           335 => x"08",
           336 => x"05",
           337 => x"94",
           338 => x"08",
           339 => x"88",
           340 => x"81",
           341 => x"08",
           342 => x"f8",
           343 => x"94",
           344 => x"08",
           345 => x"38",
           346 => x"05",
           347 => x"08",
           348 => x"94",
           349 => x"08",
           350 => x"54",
           351 => x"94",
           352 => x"08",
           353 => x"fb",
           354 => x"0b",
           355 => x"05",
           356 => x"88",
           357 => x"25",
           358 => x"08",
           359 => x"30",
           360 => x"05",
           361 => x"94",
           362 => x"0c",
           363 => x"05",
           364 => x"8c",
           365 => x"8c",
           366 => x"94",
           367 => x"0c",
           368 => x"08",
           369 => x"52",
           370 => x"05",
           371 => x"3f",
           372 => x"94",
           373 => x"0c",
           374 => x"fc",
           375 => x"2e",
           376 => x"08",
           377 => x"30",
           378 => x"05",
           379 => x"f8",
           380 => x"88",
           381 => x"3d",
           382 => x"04",
           383 => x"94",
           384 => x"0d",
           385 => x"08",
           386 => x"80",
           387 => x"f8",
           388 => x"08",
           389 => x"94",
           390 => x"08",
           391 => x"94",
           392 => x"08",
           393 => x"38",
           394 => x"08",
           395 => x"24",
           396 => x"08",
           397 => x"10",
           398 => x"05",
           399 => x"fc",
           400 => x"94",
           401 => x"0c",
           402 => x"08",
           403 => x"80",
           404 => x"38",
           405 => x"05",
           406 => x"88",
           407 => x"a1",
           408 => x"88",
           409 => x"08",
           410 => x"31",
           411 => x"05",
           412 => x"f8",
           413 => x"08",
           414 => x"07",
           415 => x"05",
           416 => x"fc",
           417 => x"2a",
           418 => x"05",
           419 => x"8c",
           420 => x"2a",
           421 => x"05",
           422 => x"39",
           423 => x"05",
           424 => x"8f",
           425 => x"88",
           426 => x"94",
           427 => x"0c",
           428 => x"94",
           429 => x"08",
           430 => x"f4",
           431 => x"94",
           432 => x"08",
           433 => x"3d",
           434 => x"04",
           435 => x"81",
           436 => x"c0",
           437 => x"81",
           438 => x"92",
           439 => x"0b",
           440 => x"8c",
           441 => x"92",
           442 => x"82",
           443 => x"70",
           444 => x"38",
           445 => x"8c",
           446 => x"e9",
           447 => x"92",
           448 => x"80",
           449 => x"71",
           450 => x"c0",
           451 => x"51",
           452 => x"88",
           453 => x"0b",
           454 => x"34",
           455 => x"9f",
           456 => x"0c",
           457 => x"04",
           458 => x"78",
           459 => x"58",
           460 => x"0b",
           461 => x"f0",
           462 => x"52",
           463 => x"70",
           464 => x"81",
           465 => x"38",
           466 => x"c0",
           467 => x"79",
           468 => x"80",
           469 => x"87",
           470 => x"0c",
           471 => x"8c",
           472 => x"2a",
           473 => x"51",
           474 => x"80",
           475 => x"87",
           476 => x"08",
           477 => x"06",
           478 => x"52",
           479 => x"80",
           480 => x"70",
           481 => x"38",
           482 => x"81",
           483 => x"ff",
           484 => x"15",
           485 => x"06",
           486 => x"2e",
           487 => x"c0",
           488 => x"51",
           489 => x"38",
           490 => x"8c",
           491 => x"95",
           492 => x"87",
           493 => x"0c",
           494 => x"8c",
           495 => x"06",
           496 => x"f4",
           497 => x"fc",
           498 => x"52",
           499 => x"2e",
           500 => x"8f",
           501 => x"98",
           502 => x"70",
           503 => x"81",
           504 => x"81",
           505 => x"0c",
           506 => x"04",
           507 => x"74",
           508 => x"71",
           509 => x"2b",
           510 => x"53",
           511 => x"0d",
           512 => x"0d",
           513 => x"33",
           514 => x"71",
           515 => x"88",
           516 => x"14",
           517 => x"07",
           518 => x"33",
           519 => x"0c",
           520 => x"56",
           521 => x"3d",
           522 => x"3d",
           523 => x"0b",
           524 => x"08",
           525 => x"77",
           526 => x"38",
           527 => x"08",
           528 => x"38",
           529 => x"74",
           530 => x"38",
           531 => x"ae",
           532 => x"39",
           533 => x"10",
           534 => x"53",
           535 => x"8c",
           536 => x"52",
           537 => x"52",
           538 => x"3f",
           539 => x"38",
           540 => x"f8",
           541 => x"83",
           542 => x"55",
           543 => x"54",
           544 => x"83",
           545 => x"76",
           546 => x"17",
           547 => x"88",
           548 => x"55",
           549 => x"88",
           550 => x"74",
           551 => x"3f",
           552 => x"0a",
           553 => x"39",
           554 => x"88",
           555 => x"0d",
           556 => x"0d",
           557 => x"9f",
           558 => x"19",
           559 => x"fe",
           560 => x"54",
           561 => x"73",
           562 => x"82",
           563 => x"71",
           564 => x"08",
           565 => x"75",
           566 => x"3d",
           567 => x"3d",
           568 => x"80",
           569 => x"0b",
           570 => x"70",
           571 => x"53",
           572 => x"09",
           573 => x"38",
           574 => x"fd",
           575 => x"08",
           576 => x"9a",
           577 => x"e4",
           578 => x"83",
           579 => x"73",
           580 => x"85",
           581 => x"fc",
           582 => x"0b",
           583 => x"f4",
           584 => x"80",
           585 => x"15",
           586 => x"81",
           587 => x"88",
           588 => x"26",
           589 => x"52",
           590 => x"90",
           591 => x"52",
           592 => x"09",
           593 => x"38",
           594 => x"53",
           595 => x"0c",
           596 => x"8b",
           597 => x"fe",
           598 => x"08",
           599 => x"90",
           600 => x"71",
           601 => x"80",
           602 => x"0c",
           603 => x"04",
           604 => x"78",
           605 => x"9f",
           606 => x"22",
           607 => x"83",
           608 => x"57",
           609 => x"73",
           610 => x"38",
           611 => x"53",
           612 => x"83",
           613 => x"39",
           614 => x"52",
           615 => x"38",
           616 => x"16",
           617 => x"08",
           618 => x"38",
           619 => x"17",
           620 => x"73",
           621 => x"38",
           622 => x"16",
           623 => x"74",
           624 => x"52",
           625 => x"72",
           626 => x"3f",
           627 => x"88",
           628 => x"38",
           629 => x"08",
           630 => x"27",
           631 => x"08",
           632 => x"88",
           633 => x"c9",
           634 => x"90",
           635 => x"75",
           636 => x"71",
           637 => x"3d",
           638 => x"3d",
           639 => x"64",
           640 => x"75",
           641 => x"a0",
           642 => x"06",
           643 => x"16",
           644 => x"ef",
           645 => x"33",
           646 => x"af",
           647 => x"06",
           648 => x"16",
           649 => x"88",
           650 => x"70",
           651 => x"74",
           652 => x"38",
           653 => x"df",
           654 => x"56",
           655 => x"82",
           656 => x"3d",
           657 => x"70",
           658 => x"8a",
           659 => x"70",
           660 => x"34",
           661 => x"74",
           662 => x"81",
           663 => x"80",
           664 => x"88",
           665 => x"5a",
           666 => x"70",
           667 => x"60",
           668 => x"70",
           669 => x"30",
           670 => x"71",
           671 => x"51",
           672 => x"53",
           673 => x"74",
           674 => x"76",
           675 => x"81",
           676 => x"81",
           677 => x"27",
           678 => x"74",
           679 => x"38",
           680 => x"70",
           681 => x"32",
           682 => x"73",
           683 => x"53",
           684 => x"56",
           685 => x"88",
           686 => x"ff",
           687 => x"81",
           688 => x"ff",
           689 => x"53",
           690 => x"76",
           691 => x"98",
           692 => x"7f",
           693 => x"76",
           694 => x"38",
           695 => x"8b",
           696 => x"51",
           697 => x"88",
           698 => x"38",
           699 => x"22",
           700 => x"83",
           701 => x"55",
           702 => x"52",
           703 => x"a8",
           704 => x"57",
           705 => x"fb",
           706 => x"55",
           707 => x"80",
           708 => x"1d",
           709 => x"2a",
           710 => x"51",
           711 => x"b2",
           712 => x"84",
           713 => x"08",
           714 => x"58",
           715 => x"77",
           716 => x"38",
           717 => x"05",
           718 => x"70",
           719 => x"33",
           720 => x"52",
           721 => x"80",
           722 => x"86",
           723 => x"2e",
           724 => x"51",
           725 => x"ff",
           726 => x"08",
           727 => x"b4",
           728 => x"76",
           729 => x"08",
           730 => x"51",
           731 => x"38",
           732 => x"70",
           733 => x"81",
           734 => x"56",
           735 => x"83",
           736 => x"81",
           737 => x"7c",
           738 => x"3f",
           739 => x"1d",
           740 => x"39",
           741 => x"90",
           742 => x"f9",
           743 => x"7b",
           744 => x"54",
           745 => x"77",
           746 => x"f6",
           747 => x"56",
           748 => x"e7",
           749 => x"f8",
           750 => x"08",
           751 => x"06",
           752 => x"74",
           753 => x"2e",
           754 => x"80",
           755 => x"54",
           756 => x"52",
           757 => x"d0",
           758 => x"56",
           759 => x"38",
           760 => x"88",
           761 => x"83",
           762 => x"55",
           763 => x"c6",
           764 => x"82",
           765 => x"53",
           766 => x"51",
           767 => x"88",
           768 => x"08",
           769 => x"51",
           770 => x"88",
           771 => x"ff",
           772 => x"81",
           773 => x"83",
           774 => x"75",
           775 => x"3d",
           776 => x"3d",
           777 => x"80",
           778 => x"0b",
           779 => x"f5",
           780 => x"08",
           781 => x"82",
           782 => x"f2",
           783 => x"53",
           784 => x"53",
           785 => x"d3",
           786 => x"81",
           787 => x"76",
           788 => x"81",
           789 => x"90",
           790 => x"53",
           791 => x"51",
           792 => x"88",
           793 => x"8d",
           794 => x"74",
           795 => x"38",
           796 => x"05",
           797 => x"3f",
           798 => x"08",
           799 => x"5a",
           800 => x"88",
           801 => x"06",
           802 => x"2e",
           803 => x"86",
           804 => x"82",
           805 => x"80",
           806 => x"86",
           807 => x"39",
           808 => x"53",
           809 => x"51",
           810 => x"81",
           811 => x"81",
           812 => x"3d",
           813 => x"f6",
           814 => x"08",
           815 => x"06",
           816 => x"38",
           817 => x"05",
           818 => x"3f",
           819 => x"02",
           820 => x"78",
           821 => x"88",
           822 => x"70",
           823 => x"5b",
           824 => x"88",
           825 => x"ff",
           826 => x"8c",
           827 => x"3d",
           828 => x"34",
           829 => x"05",
           830 => x"3f",
           831 => x"1a",
           832 => x"e2",
           833 => x"e4",
           834 => x"83",
           835 => x"56",
           836 => x"95",
           837 => x"51",
           838 => x"88",
           839 => x"51",
           840 => x"88",
           841 => x"ff",
           842 => x"31",
           843 => x"1b",
           844 => x"2a",
           845 => x"56",
           846 => x"55",
           847 => x"55",
           848 => x"88",
           849 => x"70",
           850 => x"88",
           851 => x"05",
           852 => x"83",
           853 => x"83",
           854 => x"83",
           855 => x"27",
           856 => x"57",
           857 => x"56",
           858 => x"80",
           859 => x"79",
           860 => x"2e",
           861 => x"90",
           862 => x"fb",
           863 => x"81",
           864 => x"90",
           865 => x"39",
           866 => x"18",
           867 => x"79",
           868 => x"06",
           869 => x"19",
           870 => x"05",
           871 => x"55",
           872 => x"1a",
           873 => x"0b",
           874 => x"0c",
           875 => x"88",
           876 => x"0d",
           877 => x"0d",
           878 => x"9f",
           879 => x"85",
           880 => x"2e",
           881 => x"80",
           882 => x"34",
           883 => x"11",
           884 => x"89",
           885 => x"57",
           886 => x"f8",
           887 => x"08",
           888 => x"80",
           889 => x"3d",
           890 => x"80",
           891 => x"02",
           892 => x"70",
           893 => x"81",
           894 => x"57",
           895 => x"85",
           896 => x"a1",
           897 => x"f5",
           898 => x"08",
           899 => x"98",
           900 => x"51",
           901 => x"88",
           902 => x"0c",
           903 => x"0c",
           904 => x"16",
           905 => x"0c",
           906 => x"04",
           907 => x"7d",
           908 => x"0b",
           909 => x"08",
           910 => x"58",
           911 => x"85",
           912 => x"2e",
           913 => x"81",
           914 => x"06",
           915 => x"74",
           916 => x"c3",
           917 => x"74",
           918 => x"86",
           919 => x"81",
           920 => x"57",
           921 => x"9c",
           922 => x"17",
           923 => x"74",
           924 => x"38",
           925 => x"80",
           926 => x"38",
           927 => x"70",
           928 => x"56",
           929 => x"c7",
           930 => x"33",
           931 => x"89",
           932 => x"81",
           933 => x"55",
           934 => x"76",
           935 => x"16",
           936 => x"39",
           937 => x"51",
           938 => x"88",
           939 => x"75",
           940 => x"38",
           941 => x"0c",
           942 => x"51",
           943 => x"88",
           944 => x"08",
           945 => x"8f",
           946 => x"1a",
           947 => x"98",
           948 => x"ff",
           949 => x"71",
           950 => x"77",
           951 => x"38",
           952 => x"54",
           953 => x"83",
           954 => x"a8",
           955 => x"78",
           956 => x"3f",
           957 => x"e5",
           958 => x"08",
           959 => x"0c",
           960 => x"7b",
           961 => x"0c",
           962 => x"2e",
           963 => x"74",
           964 => x"e2",
           965 => x"76",
           966 => x"3d",
           967 => x"3d",
           968 => x"94",
           969 => x"87",
           970 => x"73",
           971 => x"3f",
           972 => x"2b",
           973 => x"8c",
           974 => x"87",
           975 => x"74",
           976 => x"3f",
           977 => x"07",
           978 => x"8c",
           979 => x"94",
           980 => x"87",
           981 => x"73",
           982 => x"3f",
           983 => x"2b",
           984 => x"9c",
           985 => x"87",
           986 => x"74",
           987 => x"3f",
           988 => x"07",
           989 => x"9c",
           990 => x"83",
           991 => x"94",
           992 => x"80",
           993 => x"c0",
           994 => x"9f",
           995 => x"92",
           996 => x"b8",
           997 => x"51",
           998 => x"88",
           999 => x"a0",
          1000 => x"08",
          1001 => x"88",
          1002 => x"3d",
          1003 => x"84",
          1004 => x"51",
          1005 => x"88",
          1006 => x"75",
          1007 => x"2e",
          1008 => x"15",
          1009 => x"a0",
          1010 => x"04",
          1011 => x"39",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"00",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"4e",
          1018 => x"4f",
          1019 => x"00",
          1020 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"f4",
           281 => x"27",
           282 => x"71",
           283 => x"53",
           284 => x"0b",
           285 => x"88",
           286 => x"9d",
           287 => x"04",
           288 => x"04",
           289 => x"94",
           290 => x"0c",
           291 => x"80",
           292 => x"8c",
           293 => x"94",
           294 => x"08",
           295 => x"3f",
           296 => x"88",
           297 => x"3d",
           298 => x"04",
           299 => x"94",
           300 => x"0d",
           301 => x"08",
           302 => x"52",
           303 => x"05",
           304 => x"b9",
           305 => x"70",
           306 => x"85",
           307 => x"0c",
           308 => x"02",
           309 => x"3d",
           310 => x"94",
           311 => x"0c",
           312 => x"05",
           313 => x"ab",
           314 => x"88",
           315 => x"94",
           316 => x"0c",
           317 => x"08",
           318 => x"94",
           319 => x"08",
           320 => x"0b",
           321 => x"05",
           322 => x"f4",
           323 => x"08",
           324 => x"94",
           325 => x"08",
           326 => x"38",
           327 => x"05",
           328 => x"08",
           329 => x"80",
           330 => x"f0",
           331 => x"08",
           332 => x"88",
           333 => x"94",
           334 => x"0c",
           335 => x"05",
           336 => x"fc",
           337 => x"53",
           338 => x"05",
           339 => x"08",
           340 => x"51",
           341 => x"88",
           342 => x"08",
           343 => x"54",
           344 => x"05",
           345 => x"8c",
           346 => x"f8",
           347 => x"94",
           348 => x"0c",
           349 => x"05",
           350 => x"0c",
           351 => x"0d",
           352 => x"94",
           353 => x"0c",
           354 => x"80",
           355 => x"fc",
           356 => x"08",
           357 => x"80",
           358 => x"94",
           359 => x"08",
           360 => x"88",
           361 => x"0b",
           362 => x"05",
           363 => x"8c",
           364 => x"25",
           365 => x"08",
           366 => x"30",
           367 => x"05",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"ad",
           372 => x"70",
           373 => x"05",
           374 => x"08",
           375 => x"80",
           376 => x"94",
           377 => x"08",
           378 => x"f8",
           379 => x"08",
           380 => x"70",
           381 => x"87",
           382 => x"0c",
           383 => x"02",
           384 => x"3d",
           385 => x"94",
           386 => x"0c",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"05",
           391 => x"38",
           392 => x"05",
           393 => x"a3",
           394 => x"94",
           395 => x"08",
           396 => x"94",
           397 => x"08",
           398 => x"8c",
           399 => x"08",
           400 => x"10",
           401 => x"05",
           402 => x"94",
           403 => x"08",
           404 => x"c9",
           405 => x"8c",
           406 => x"08",
           407 => x"26",
           408 => x"08",
           409 => x"94",
           410 => x"08",
           411 => x"88",
           412 => x"08",
           413 => x"94",
           414 => x"08",
           415 => x"f8",
           416 => x"08",
           417 => x"81",
           418 => x"fc",
           419 => x"08",
           420 => x"81",
           421 => x"8c",
           422 => x"af",
           423 => x"90",
           424 => x"2e",
           425 => x"08",
           426 => x"70",
           427 => x"05",
           428 => x"39",
           429 => x"05",
           430 => x"08",
           431 => x"51",
           432 => x"05",
           433 => x"85",
           434 => x"0c",
           435 => x"0d",
           436 => x"87",
           437 => x"0c",
           438 => x"c0",
           439 => x"85",
           440 => x"98",
           441 => x"c0",
           442 => x"70",
           443 => x"51",
           444 => x"8a",
           445 => x"98",
           446 => x"70",
           447 => x"c0",
           448 => x"fc",
           449 => x"52",
           450 => x"87",
           451 => x"08",
           452 => x"2e",
           453 => x"0b",
           454 => x"f0",
           455 => x"0b",
           456 => x"88",
           457 => x"0d",
           458 => x"0d",
           459 => x"56",
           460 => x"0b",
           461 => x"9f",
           462 => x"06",
           463 => x"52",
           464 => x"09",
           465 => x"9e",
           466 => x"87",
           467 => x"0c",
           468 => x"92",
           469 => x"0b",
           470 => x"8c",
           471 => x"92",
           472 => x"85",
           473 => x"06",
           474 => x"70",
           475 => x"38",
           476 => x"84",
           477 => x"ff",
           478 => x"27",
           479 => x"73",
           480 => x"38",
           481 => x"8b",
           482 => x"70",
           483 => x"34",
           484 => x"81",
           485 => x"a2",
           486 => x"80",
           487 => x"87",
           488 => x"08",
           489 => x"b5",
           490 => x"98",
           491 => x"70",
           492 => x"0b",
           493 => x"8c",
           494 => x"92",
           495 => x"82",
           496 => x"70",
           497 => x"73",
           498 => x"06",
           499 => x"72",
           500 => x"06",
           501 => x"c0",
           502 => x"51",
           503 => x"09",
           504 => x"38",
           505 => x"88",
           506 => x"0d",
           507 => x"0d",
           508 => x"33",
           509 => x"88",
           510 => x"0c",
           511 => x"3d",
           512 => x"3d",
           513 => x"11",
           514 => x"33",
           515 => x"71",
           516 => x"81",
           517 => x"72",
           518 => x"75",
           519 => x"88",
           520 => x"54",
           521 => x"85",
           522 => x"f9",
           523 => x"0b",
           524 => x"f4",
           525 => x"81",
           526 => x"ed",
           527 => x"17",
           528 => x"e5",
           529 => x"55",
           530 => x"89",
           531 => x"2e",
           532 => x"d5",
           533 => x"76",
           534 => x"06",
           535 => x"2a",
           536 => x"05",
           537 => x"70",
           538 => x"bd",
           539 => x"b9",
           540 => x"fe",
           541 => x"08",
           542 => x"06",
           543 => x"84",
           544 => x"2b",
           545 => x"53",
           546 => x"8c",
           547 => x"52",
           548 => x"52",
           549 => x"3f",
           550 => x"38",
           551 => x"e2",
           552 => x"f0",
           553 => x"83",
           554 => x"74",
           555 => x"3d",
           556 => x"3d",
           557 => x"0b",
           558 => x"fe",
           559 => x"08",
           560 => x"56",
           561 => x"74",
           562 => x"38",
           563 => x"75",
           564 => x"16",
           565 => x"53",
           566 => x"87",
           567 => x"fd",
           568 => x"54",
           569 => x"0b",
           570 => x"08",
           571 => x"53",
           572 => x"2e",
           573 => x"8c",
           574 => x"51",
           575 => x"88",
           576 => x"53",
           577 => x"fd",
           578 => x"08",
           579 => x"06",
           580 => x"0c",
           581 => x"04",
           582 => x"76",
           583 => x"9f",
           584 => x"55",
           585 => x"88",
           586 => x"72",
           587 => x"38",
           588 => x"73",
           589 => x"81",
           590 => x"72",
           591 => x"33",
           592 => x"2e",
           593 => x"85",
           594 => x"08",
           595 => x"16",
           596 => x"2e",
           597 => x"51",
           598 => x"88",
           599 => x"39",
           600 => x"52",
           601 => x"0c",
           602 => x"88",
           603 => x"0d",
           604 => x"0d",
           605 => x"0b",
           606 => x"71",
           607 => x"70",
           608 => x"06",
           609 => x"55",
           610 => x"88",
           611 => x"08",
           612 => x"38",
           613 => x"dc",
           614 => x"06",
           615 => x"cf",
           616 => x"90",
           617 => x"15",
           618 => x"8f",
           619 => x"84",
           620 => x"52",
           621 => x"bc",
           622 => x"82",
           623 => x"05",
           624 => x"06",
           625 => x"38",
           626 => x"df",
           627 => x"71",
           628 => x"a0",
           629 => x"88",
           630 => x"08",
           631 => x"88",
           632 => x"0c",
           633 => x"fd",
           634 => x"08",
           635 => x"73",
           636 => x"52",
           637 => x"88",
           638 => x"f2",
           639 => x"62",
           640 => x"5c",
           641 => x"74",
           642 => x"81",
           643 => x"81",
           644 => x"56",
           645 => x"70",
           646 => x"74",
           647 => x"81",
           648 => x"81",
           649 => x"0b",
           650 => x"62",
           651 => x"55",
           652 => x"8f",
           653 => x"fd",
           654 => x"08",
           655 => x"34",
           656 => x"93",
           657 => x"08",
           658 => x"5f",
           659 => x"76",
           660 => x"58",
           661 => x"55",
           662 => x"09",
           663 => x"38",
           664 => x"5b",
           665 => x"5f",
           666 => x"1c",
           667 => x"06",
           668 => x"33",
           669 => x"70",
           670 => x"27",
           671 => x"07",
           672 => x"5b",
           673 => x"55",
           674 => x"38",
           675 => x"09",
           676 => x"38",
           677 => x"7a",
           678 => x"55",
           679 => x"9f",
           680 => x"32",
           681 => x"ae",
           682 => x"70",
           683 => x"2a",
           684 => x"51",
           685 => x"38",
           686 => x"5a",
           687 => x"77",
           688 => x"81",
           689 => x"1c",
           690 => x"55",
           691 => x"ff",
           692 => x"1e",
           693 => x"55",
           694 => x"83",
           695 => x"74",
           696 => x"7b",
           697 => x"3f",
           698 => x"ef",
           699 => x"7b",
           700 => x"2b",
           701 => x"54",
           702 => x"08",
           703 => x"f8",
           704 => x"08",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"8b",
           709 => x"83",
           710 => x"06",
           711 => x"74",
           712 => x"7d",
           713 => x"88",
           714 => x"5b",
           715 => x"58",
           716 => x"9a",
           717 => x"81",
           718 => x"79",
           719 => x"5b",
           720 => x"31",
           721 => x"75",
           722 => x"38",
           723 => x"80",
           724 => x"7b",
           725 => x"3f",
           726 => x"88",
           727 => x"08",
           728 => x"39",
           729 => x"1c",
           730 => x"33",
           731 => x"a5",
           732 => x"33",
           733 => x"70",
           734 => x"56",
           735 => x"38",
           736 => x"39",
           737 => x"39",
           738 => x"d3",
           739 => x"88",
           740 => x"af",
           741 => x"0c",
           742 => x"04",
           743 => x"79",
           744 => x"82",
           745 => x"53",
           746 => x"51",
           747 => x"83",
           748 => x"80",
           749 => x"51",
           750 => x"88",
           751 => x"ff",
           752 => x"56",
           753 => x"d5",
           754 => x"06",
           755 => x"75",
           756 => x"77",
           757 => x"f6",
           758 => x"08",
           759 => x"94",
           760 => x"f8",
           761 => x"08",
           762 => x"06",
           763 => x"82",
           764 => x"38",
           765 => x"d2",
           766 => x"76",
           767 => x"3f",
           768 => x"88",
           769 => x"76",
           770 => x"3f",
           771 => x"ff",
           772 => x"74",
           773 => x"2e",
           774 => x"56",
           775 => x"89",
           776 => x"ed",
           777 => x"59",
           778 => x"0b",
           779 => x"0c",
           780 => x"88",
           781 => x"55",
           782 => x"82",
           783 => x"75",
           784 => x"70",
           785 => x"fe",
           786 => x"08",
           787 => x"57",
           788 => x"09",
           789 => x"38",
           790 => x"be",
           791 => x"75",
           792 => x"3f",
           793 => x"38",
           794 => x"55",
           795 => x"ac",
           796 => x"e4",
           797 => x"8a",
           798 => x"88",
           799 => x"52",
           800 => x"3f",
           801 => x"ff",
           802 => x"83",
           803 => x"06",
           804 => x"56",
           805 => x"76",
           806 => x"38",
           807 => x"8f",
           808 => x"8d",
           809 => x"75",
           810 => x"3f",
           811 => x"08",
           812 => x"95",
           813 => x"51",
           814 => x"88",
           815 => x"ff",
           816 => x"8c",
           817 => x"f3",
           818 => x"b6",
           819 => x"58",
           820 => x"33",
           821 => x"02",
           822 => x"05",
           823 => x"59",
           824 => x"3f",
           825 => x"ff",
           826 => x"05",
           827 => x"8c",
           828 => x"1a",
           829 => x"e0",
           830 => x"f1",
           831 => x"84",
           832 => x"3d",
           833 => x"f5",
           834 => x"08",
           835 => x"06",
           836 => x"38",
           837 => x"05",
           838 => x"3f",
           839 => x"7a",
           840 => x"3f",
           841 => x"ff",
           842 => x"71",
           843 => x"84",
           844 => x"84",
           845 => x"33",
           846 => x"31",
           847 => x"51",
           848 => x"3f",
           849 => x"05",
           850 => x"0c",
           851 => x"8a",
           852 => x"74",
           853 => x"26",
           854 => x"57",
           855 => x"76",
           856 => x"83",
           857 => x"86",
           858 => x"2e",
           859 => x"76",
           860 => x"83",
           861 => x"06",
           862 => x"3d",
           863 => x"f5",
           864 => x"08",
           865 => x"88",
           866 => x"08",
           867 => x"0c",
           868 => x"ff",
           869 => x"08",
           870 => x"2a",
           871 => x"0c",
           872 => x"81",
           873 => x"0b",
           874 => x"f4",
           875 => x"75",
           876 => x"3d",
           877 => x"3d",
           878 => x"0b",
           879 => x"55",
           880 => x"80",
           881 => x"38",
           882 => x"16",
           883 => x"e0",
           884 => x"54",
           885 => x"54",
           886 => x"51",
           887 => x"88",
           888 => x"08",
           889 => x"88",
           890 => x"73",
           891 => x"38",
           892 => x"33",
           893 => x"70",
           894 => x"55",
           895 => x"2e",
           896 => x"54",
           897 => x"51",
           898 => x"88",
           899 => x"0c",
           900 => x"05",
           901 => x"3f",
           902 => x"16",
           903 => x"16",
           904 => x"81",
           905 => x"88",
           906 => x"0d",
           907 => x"0d",
           908 => x"0b",
           909 => x"f4",
           910 => x"5c",
           911 => x"0c",
           912 => x"80",
           913 => x"38",
           914 => x"81",
           915 => x"57",
           916 => x"81",
           917 => x"39",
           918 => x"34",
           919 => x"0b",
           920 => x"81",
           921 => x"39",
           922 => x"98",
           923 => x"55",
           924 => x"83",
           925 => x"77",
           926 => x"9a",
           927 => x"08",
           928 => x"06",
           929 => x"80",
           930 => x"16",
           931 => x"77",
           932 => x"70",
           933 => x"5b",
           934 => x"38",
           935 => x"a0",
           936 => x"8b",
           937 => x"08",
           938 => x"3f",
           939 => x"81",
           940 => x"aa",
           941 => x"17",
           942 => x"08",
           943 => x"3f",
           944 => x"88",
           945 => x"ff",
           946 => x"08",
           947 => x"0c",
           948 => x"83",
           949 => x"80",
           950 => x"55",
           951 => x"83",
           952 => x"74",
           953 => x"08",
           954 => x"53",
           955 => x"52",
           956 => x"b5",
           957 => x"fe",
           958 => x"16",
           959 => x"17",
           960 => x"31",
           961 => x"7c",
           962 => x"80",
           963 => x"38",
           964 => x"fe",
           965 => x"57",
           966 => x"8c",
           967 => x"fb",
           968 => x"c0",
           969 => x"54",
           970 => x"52",
           971 => x"d7",
           972 => x"90",
           973 => x"94",
           974 => x"54",
           975 => x"52",
           976 => x"c3",
           977 => x"08",
           978 => x"94",
           979 => x"c0",
           980 => x"54",
           981 => x"52",
           982 => x"ab",
           983 => x"90",
           984 => x"94",
           985 => x"54",
           986 => x"52",
           987 => x"97",
           988 => x"08",
           989 => x"94",
           990 => x"80",
           991 => x"c0",
           992 => x"8c",
           993 => x"87",
           994 => x"0c",
           995 => x"f9",
           996 => x"08",
           997 => x"e0",
           998 => x"3f",
           999 => x"38",
          1000 => x"88",
          1001 => x"98",
          1002 => x"87",
          1003 => x"53",
          1004 => x"74",
          1005 => x"3f",
          1006 => x"38",
          1007 => x"80",
          1008 => x"73",
          1009 => x"39",
          1010 => x"73",
          1011 => x"fb",
          1012 => x"ff",
          1013 => x"00",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"49",
          1018 => x"52",
          1019 => x"00",
          1020 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e0",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"d0",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cf",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"81",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"9f",
           281 => x"a4",
           282 => x"80",
           283 => x"05",
           284 => x"0b",
           285 => x"04",
           286 => x"9e",
           287 => x"80",
           288 => x"fe",
           289 => x"00",
           290 => x"94",
           291 => x"0d",
           292 => x"08",
           293 => x"52",
           294 => x"05",
           295 => x"de",
           296 => x"70",
           297 => x"85",
           298 => x"0c",
           299 => x"02",
           300 => x"3d",
           301 => x"94",
           302 => x"08",
           303 => x"88",
           304 => x"82",
           305 => x"08",
           306 => x"54",
           307 => x"94",
           308 => x"08",
           309 => x"f9",
           310 => x"0b",
           311 => x"05",
           312 => x"88",
           313 => x"25",
           314 => x"08",
           315 => x"30",
           316 => x"05",
           317 => x"94",
           318 => x"0c",
           319 => x"05",
           320 => x"81",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"0c",
           325 => x"05",
           326 => x"ab",
           327 => x"8c",
           328 => x"94",
           329 => x"0c",
           330 => x"08",
           331 => x"94",
           332 => x"08",
           333 => x"0b",
           334 => x"05",
           335 => x"f0",
           336 => x"08",
           337 => x"80",
           338 => x"8c",
           339 => x"94",
           340 => x"08",
           341 => x"3f",
           342 => x"94",
           343 => x"0c",
           344 => x"fc",
           345 => x"2e",
           346 => x"08",
           347 => x"30",
           348 => x"05",
           349 => x"f8",
           350 => x"88",
           351 => x"3d",
           352 => x"04",
           353 => x"94",
           354 => x"0d",
           355 => x"08",
           356 => x"94",
           357 => x"08",
           358 => x"38",
           359 => x"05",
           360 => x"08",
           361 => x"81",
           362 => x"fc",
           363 => x"08",
           364 => x"80",
           365 => x"94",
           366 => x"08",
           367 => x"8c",
           368 => x"53",
           369 => x"05",
           370 => x"08",
           371 => x"51",
           372 => x"08",
           373 => x"f8",
           374 => x"94",
           375 => x"08",
           376 => x"38",
           377 => x"05",
           378 => x"08",
           379 => x"94",
           380 => x"08",
           381 => x"54",
           382 => x"94",
           383 => x"08",
           384 => x"fd",
           385 => x"0b",
           386 => x"05",
           387 => x"94",
           388 => x"0c",
           389 => x"05",
           390 => x"88",
           391 => x"ac",
           392 => x"fc",
           393 => x"2e",
           394 => x"0b",
           395 => x"05",
           396 => x"38",
           397 => x"05",
           398 => x"08",
           399 => x"94",
           400 => x"08",
           401 => x"fc",
           402 => x"39",
           403 => x"05",
           404 => x"80",
           405 => x"08",
           406 => x"94",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"05",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"05",
           415 => x"08",
           416 => x"94",
           417 => x"08",
           418 => x"08",
           419 => x"94",
           420 => x"08",
           421 => x"08",
           422 => x"ff",
           423 => x"08",
           424 => x"80",
           425 => x"94",
           426 => x"08",
           427 => x"f4",
           428 => x"8d",
           429 => x"f8",
           430 => x"94",
           431 => x"0c",
           432 => x"f4",
           433 => x"0c",
           434 => x"94",
           435 => x"3d",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"c0",
           441 => x"87",
           442 => x"08",
           443 => x"51",
           444 => x"2e",
           445 => x"c0",
           446 => x"51",
           447 => x"87",
           448 => x"08",
           449 => x"06",
           450 => x"38",
           451 => x"8c",
           452 => x"80",
           453 => x"71",
           454 => x"9f",
           455 => x"0b",
           456 => x"33",
           457 => x"3d",
           458 => x"3d",
           459 => x"7d",
           460 => x"80",
           461 => x"0b",
           462 => x"81",
           463 => x"82",
           464 => x"2e",
           465 => x"81",
           466 => x"0b",
           467 => x"8c",
           468 => x"c0",
           469 => x"84",
           470 => x"92",
           471 => x"c0",
           472 => x"70",
           473 => x"81",
           474 => x"53",
           475 => x"a7",
           476 => x"92",
           477 => x"81",
           478 => x"79",
           479 => x"51",
           480 => x"90",
           481 => x"2e",
           482 => x"76",
           483 => x"58",
           484 => x"54",
           485 => x"72",
           486 => x"70",
           487 => x"38",
           488 => x"8c",
           489 => x"ff",
           490 => x"c0",
           491 => x"51",
           492 => x"81",
           493 => x"92",
           494 => x"c0",
           495 => x"70",
           496 => x"51",
           497 => x"80",
           498 => x"80",
           499 => x"70",
           500 => x"81",
           501 => x"87",
           502 => x"08",
           503 => x"2e",
           504 => x"83",
           505 => x"71",
           506 => x"3d",
           507 => x"3d",
           508 => x"11",
           509 => x"71",
           510 => x"88",
           511 => x"84",
           512 => x"fd",
           513 => x"83",
           514 => x"12",
           515 => x"2b",
           516 => x"07",
           517 => x"70",
           518 => x"2b",
           519 => x"07",
           520 => x"53",
           521 => x"52",
           522 => x"04",
           523 => x"79",
           524 => x"9f",
           525 => x"57",
           526 => x"80",
           527 => x"88",
           528 => x"80",
           529 => x"33",
           530 => x"2e",
           531 => x"83",
           532 => x"80",
           533 => x"54",
           534 => x"fe",
           535 => x"88",
           536 => x"08",
           537 => x"3d",
           538 => x"fd",
           539 => x"08",
           540 => x"51",
           541 => x"88",
           542 => x"ff",
           543 => x"39",
           544 => x"82",
           545 => x"06",
           546 => x"2a",
           547 => x"05",
           548 => x"70",
           549 => x"92",
           550 => x"8e",
           551 => x"fe",
           552 => x"08",
           553 => x"55",
           554 => x"55",
           555 => x"89",
           556 => x"fb",
           557 => x"0b",
           558 => x"08",
           559 => x"12",
           560 => x"55",
           561 => x"56",
           562 => x"8d",
           563 => x"33",
           564 => x"94",
           565 => x"57",
           566 => x"0c",
           567 => x"04",
           568 => x"75",
           569 => x"0b",
           570 => x"f4",
           571 => x"51",
           572 => x"83",
           573 => x"06",
           574 => x"14",
           575 => x"3f",
           576 => x"2b",
           577 => x"51",
           578 => x"88",
           579 => x"ff",
           580 => x"88",
           581 => x"0d",
           582 => x"0d",
           583 => x"0b",
           584 => x"55",
           585 => x"23",
           586 => x"53",
           587 => x"88",
           588 => x"08",
           589 => x"38",
           590 => x"39",
           591 => x"73",
           592 => x"83",
           593 => x"06",
           594 => x"14",
           595 => x"8c",
           596 => x"80",
           597 => x"72",
           598 => x"3f",
           599 => x"85",
           600 => x"08",
           601 => x"16",
           602 => x"71",
           603 => x"3d",
           604 => x"3d",
           605 => x"0b",
           606 => x"08",
           607 => x"05",
           608 => x"ff",
           609 => x"57",
           610 => x"2e",
           611 => x"15",
           612 => x"86",
           613 => x"80",
           614 => x"8f",
           615 => x"80",
           616 => x"13",
           617 => x"8c",
           618 => x"72",
           619 => x"0b",
           620 => x"57",
           621 => x"27",
           622 => x"39",
           623 => x"ff",
           624 => x"2a",
           625 => x"a8",
           626 => x"fc",
           627 => x"52",
           628 => x"27",
           629 => x"52",
           630 => x"17",
           631 => x"38",
           632 => x"16",
           633 => x"51",
           634 => x"88",
           635 => x"0c",
           636 => x"80",
           637 => x"0c",
           638 => x"04",
           639 => x"60",
           640 => x"5e",
           641 => x"55",
           642 => x"09",
           643 => x"38",
           644 => x"44",
           645 => x"62",
           646 => x"56",
           647 => x"09",
           648 => x"38",
           649 => x"80",
           650 => x"0c",
           651 => x"51",
           652 => x"26",
           653 => x"51",
           654 => x"88",
           655 => x"7d",
           656 => x"39",
           657 => x"1d",
           658 => x"5a",
           659 => x"a0",
           660 => x"05",
           661 => x"15",
           662 => x"2e",
           663 => x"ef",
           664 => x"59",
           665 => x"08",
           666 => x"81",
           667 => x"ff",
           668 => x"70",
           669 => x"32",
           670 => x"73",
           671 => x"25",
           672 => x"52",
           673 => x"57",
           674 => x"c7",
           675 => x"2e",
           676 => x"83",
           677 => x"77",
           678 => x"07",
           679 => x"2e",
           680 => x"88",
           681 => x"78",
           682 => x"30",
           683 => x"9f",
           684 => x"57",
           685 => x"9b",
           686 => x"8b",
           687 => x"39",
           688 => x"70",
           689 => x"72",
           690 => x"57",
           691 => x"34",
           692 => x"7a",
           693 => x"80",
           694 => x"26",
           695 => x"55",
           696 => x"34",
           697 => x"b1",
           698 => x"80",
           699 => x"54",
           700 => x"85",
           701 => x"06",
           702 => x"1c",
           703 => x"51",
           704 => x"88",
           705 => x"08",
           706 => x"7c",
           707 => x"80",
           708 => x"38",
           709 => x"70",
           710 => x"81",
           711 => x"56",
           712 => x"8b",
           713 => x"08",
           714 => x"5b",
           715 => x"18",
           716 => x"2e",
           717 => x"70",
           718 => x"33",
           719 => x"05",
           720 => x"71",
           721 => x"56",
           722 => x"e2",
           723 => x"75",
           724 => x"38",
           725 => x"9a",
           726 => x"39",
           727 => x"88",
           728 => x"83",
           729 => x"84",
           730 => x"11",
           731 => x"74",
           732 => x"1d",
           733 => x"2a",
           734 => x"51",
           735 => x"89",
           736 => x"92",
           737 => x"8e",
           738 => x"fa",
           739 => x"08",
           740 => x"fd",
           741 => x"88",
           742 => x"0d",
           743 => x"0d",
           744 => x"57",
           745 => x"fe",
           746 => x"76",
           747 => x"3f",
           748 => x"08",
           749 => x"76",
           750 => x"3f",
           751 => x"ff",
           752 => x"82",
           753 => x"d4",
           754 => x"81",
           755 => x"38",
           756 => x"53",
           757 => x"51",
           758 => x"88",
           759 => x"08",
           760 => x"51",
           761 => x"88",
           762 => x"ff",
           763 => x"81",
           764 => x"a9",
           765 => x"80",
           766 => x"52",
           767 => x"aa",
           768 => x"56",
           769 => x"38",
           770 => x"e2",
           771 => x"83",
           772 => x"55",
           773 => x"c6",
           774 => x"81",
           775 => x"0c",
           776 => x"04",
           777 => x"65",
           778 => x"0b",
           779 => x"f4",
           780 => x"3f",
           781 => x"06",
           782 => x"74",
           783 => x"74",
           784 => x"3d",
           785 => x"5a",
           786 => x"88",
           787 => x"06",
           788 => x"2e",
           789 => x"b3",
           790 => x"83",
           791 => x"52",
           792 => x"c6",
           793 => x"ab",
           794 => x"33",
           795 => x"2e",
           796 => x"3d",
           797 => x"f7",
           798 => x"08",
           799 => x"76",
           800 => x"99",
           801 => x"81",
           802 => x"76",
           803 => x"81",
           804 => x"81",
           805 => x"39",
           806 => x"86",
           807 => x"82",
           808 => x"54",
           809 => x"52",
           810 => x"fe",
           811 => x"88",
           812 => x"38",
           813 => x"05",
           814 => x"3f",
           815 => x"ff",
           816 => x"77",
           817 => x"3d",
           818 => x"f6",
           819 => x"08",
           820 => x"05",
           821 => x"29",
           822 => x"ad",
           823 => x"52",
           824 => x"8a",
           825 => x"83",
           826 => x"7a",
           827 => x"0c",
           828 => x"82",
           829 => x"3d",
           830 => x"f5",
           831 => x"08",
           832 => x"95",
           833 => x"51",
           834 => x"88",
           835 => x"ff",
           836 => x"8c",
           837 => x"ef",
           838 => x"e7",
           839 => x"56",
           840 => x"ca",
           841 => x"83",
           842 => x"76",
           843 => x"31",
           844 => x"70",
           845 => x"1d",
           846 => x"71",
           847 => x"5c",
           848 => x"c4",
           849 => x"82",
           850 => x"1b",
           851 => x"e0",
           852 => x"56",
           853 => x"fe",
           854 => x"82",
           855 => x"f6",
           856 => x"38",
           857 => x"39",
           858 => x"80",
           859 => x"38",
           860 => x"76",
           861 => x"81",
           862 => x"95",
           863 => x"51",
           864 => x"88",
           865 => x"0c",
           866 => x"19",
           867 => x"1a",
           868 => x"ff",
           869 => x"1a",
           870 => x"84",
           871 => x"1b",
           872 => x"0b",
           873 => x"78",
           874 => x"9f",
           875 => x"56",
           876 => x"95",
           877 => x"ea",
           878 => x"0b",
           879 => x"08",
           880 => x"74",
           881 => x"df",
           882 => x"81",
           883 => x"3d",
           884 => x"69",
           885 => x"70",
           886 => x"05",
           887 => x"3f",
           888 => x"88",
           889 => x"38",
           890 => x"54",
           891 => x"93",
           892 => x"05",
           893 => x"2a",
           894 => x"51",
           895 => x"80",
           896 => x"83",
           897 => x"75",
           898 => x"3f",
           899 => x"16",
           900 => x"dc",
           901 => x"eb",
           902 => x"9c",
           903 => x"98",
           904 => x"0b",
           905 => x"73",
           906 => x"3d",
           907 => x"3d",
           908 => x"7e",
           909 => x"9f",
           910 => x"5b",
           911 => x"7b",
           912 => x"75",
           913 => x"d1",
           914 => x"33",
           915 => x"84",
           916 => x"2e",
           917 => x"91",
           918 => x"17",
           919 => x"80",
           920 => x"34",
           921 => x"b1",
           922 => x"08",
           923 => x"31",
           924 => x"27",
           925 => x"58",
           926 => x"81",
           927 => x"16",
           928 => x"ff",
           929 => x"74",
           930 => x"82",
           931 => x"05",
           932 => x"06",
           933 => x"06",
           934 => x"9e",
           935 => x"38",
           936 => x"55",
           937 => x"16",
           938 => x"80",
           939 => x"55",
           940 => x"ff",
           941 => x"a4",
           942 => x"16",
           943 => x"f3",
           944 => x"55",
           945 => x"2e",
           946 => x"88",
           947 => x"17",
           948 => x"08",
           949 => x"84",
           950 => x"51",
           951 => x"27",
           952 => x"55",
           953 => x"16",
           954 => x"06",
           955 => x"08",
           956 => x"f0",
           957 => x"08",
           958 => x"98",
           959 => x"98",
           960 => x"75",
           961 => x"16",
           962 => x"78",
           963 => x"e8",
           964 => x"59",
           965 => x"80",
           966 => x"0c",
           967 => x"04",
           968 => x"87",
           969 => x"08",
           970 => x"80",
           971 => x"ea",
           972 => x"08",
           973 => x"c0",
           974 => x"56",
           975 => x"80",
           976 => x"ea",
           977 => x"88",
           978 => x"c0",
           979 => x"87",
           980 => x"08",
           981 => x"80",
           982 => x"ea",
           983 => x"08",
           984 => x"c0",
           985 => x"56",
           986 => x"80",
           987 => x"ea",
           988 => x"88",
           989 => x"c0",
           990 => x"8c",
           991 => x"87",
           992 => x"0c",
           993 => x"0b",
           994 => x"94",
           995 => x"51",
           996 => x"88",
           997 => x"9f",
           998 => x"9b",
           999 => x"ae",
          1000 => x"0b",
          1001 => x"c0",
          1002 => x"55",
          1003 => x"05",
          1004 => x"52",
          1005 => x"f6",
          1006 => x"8d",
          1007 => x"73",
          1008 => x"38",
          1009 => x"e4",
          1010 => x"54",
          1011 => x"54",
          1012 => x"00",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"42",
          1017 => x"54",
          1018 => x"2e",
          1019 => x"00",
          1020 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
