-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBRAM;

architecture arch of SinglePortBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"a4",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"a4",
             9 => x"0b",
            10 => x"04",
            11 => x"a4",
            12 => x"0b",
            13 => x"04",
            14 => x"a4",
            15 => x"0b",
            16 => x"04",
            17 => x"a4",
            18 => x"0b",
            19 => x"04",
            20 => x"a4",
            21 => x"0b",
            22 => x"04",
            23 => x"a5",
            24 => x"0b",
            25 => x"04",
            26 => x"a5",
            27 => x"0b",
            28 => x"04",
            29 => x"a5",
            30 => x"0b",
            31 => x"04",
            32 => x"a5",
            33 => x"0b",
            34 => x"04",
            35 => x"a6",
            36 => x"0b",
            37 => x"04",
            38 => x"a6",
            39 => x"0b",
            40 => x"04",
            41 => x"a6",
            42 => x"0b",
            43 => x"04",
            44 => x"a6",
            45 => x"0b",
            46 => x"04",
            47 => x"a7",
            48 => x"0b",
            49 => x"04",
            50 => x"a7",
            51 => x"0b",
            52 => x"04",
            53 => x"a7",
            54 => x"0b",
            55 => x"04",
            56 => x"a7",
            57 => x"0b",
            58 => x"04",
            59 => x"a8",
            60 => x"0b",
            61 => x"04",
            62 => x"a8",
            63 => x"0b",
            64 => x"04",
            65 => x"a8",
            66 => x"0b",
            67 => x"04",
            68 => x"a8",
            69 => x"0b",
            70 => x"04",
            71 => x"a9",
            72 => x"0b",
            73 => x"04",
            74 => x"a9",
            75 => x"0b",
            76 => x"04",
            77 => x"a9",
            78 => x"0b",
            79 => x"04",
            80 => x"a9",
            81 => x"0b",
            82 => x"04",
            83 => x"aa",
            84 => x"0b",
            85 => x"04",
            86 => x"aa",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"04",
           129 => x"0c",
           130 => x"82",
           131 => x"83",
           132 => x"82",
           133 => x"80",
           134 => x"82",
           135 => x"83",
           136 => x"82",
           137 => x"80",
           138 => x"82",
           139 => x"83",
           140 => x"82",
           141 => x"80",
           142 => x"82",
           143 => x"83",
           144 => x"82",
           145 => x"80",
           146 => x"82",
           147 => x"83",
           148 => x"82",
           149 => x"80",
           150 => x"82",
           151 => x"83",
           152 => x"82",
           153 => x"80",
           154 => x"82",
           155 => x"83",
           156 => x"82",
           157 => x"80",
           158 => x"82",
           159 => x"83",
           160 => x"82",
           161 => x"80",
           162 => x"82",
           163 => x"83",
           164 => x"82",
           165 => x"80",
           166 => x"82",
           167 => x"83",
           168 => x"82",
           169 => x"80",
           170 => x"82",
           171 => x"83",
           172 => x"82",
           173 => x"80",
           174 => x"82",
           175 => x"83",
           176 => x"82",
           177 => x"80",
           178 => x"82",
           179 => x"83",
           180 => x"82",
           181 => x"ba",
           182 => x"8c",
           183 => x"80",
           184 => x"8c",
           185 => x"fe",
           186 => x"e8",
           187 => x"90",
           188 => x"e8",
           189 => x"2d",
           190 => x"08",
           191 => x"04",
           192 => x"0c",
           193 => x"82",
           194 => x"83",
           195 => x"82",
           196 => x"b6",
           197 => x"8c",
           198 => x"80",
           199 => x"8c",
           200 => x"98",
           201 => x"8c",
           202 => x"80",
           203 => x"8c",
           204 => x"a5",
           205 => x"8c",
           206 => x"80",
           207 => x"8c",
           208 => x"9d",
           209 => x"8c",
           210 => x"80",
           211 => x"8c",
           212 => x"a0",
           213 => x"8c",
           214 => x"80",
           215 => x"8c",
           216 => x"aa",
           217 => x"8c",
           218 => x"80",
           219 => x"8c",
           220 => x"b3",
           221 => x"8c",
           222 => x"80",
           223 => x"8c",
           224 => x"a3",
           225 => x"8c",
           226 => x"80",
           227 => x"8c",
           228 => x"ad",
           229 => x"8c",
           230 => x"80",
           231 => x"8c",
           232 => x"ae",
           233 => x"8c",
           234 => x"80",
           235 => x"8c",
           236 => x"af",
           237 => x"8c",
           238 => x"80",
           239 => x"8c",
           240 => x"b6",
           241 => x"8c",
           242 => x"80",
           243 => x"8c",
           244 => x"b4",
           245 => x"8c",
           246 => x"80",
           247 => x"8c",
           248 => x"b9",
           249 => x"8c",
           250 => x"80",
           251 => x"8c",
           252 => x"b0",
           253 => x"8c",
           254 => x"80",
           255 => x"8c",
           256 => x"bc",
           257 => x"8c",
           258 => x"80",
           259 => x"8c",
           260 => x"bd",
           261 => x"8c",
           262 => x"80",
           263 => x"8c",
           264 => x"a5",
           265 => x"8c",
           266 => x"80",
           267 => x"8c",
           268 => x"a5",
           269 => x"8c",
           270 => x"80",
           271 => x"8c",
           272 => x"a6",
           273 => x"8c",
           274 => x"80",
           275 => x"8c",
           276 => x"b0",
           277 => x"8c",
           278 => x"80",
           279 => x"8c",
           280 => x"be",
           281 => x"8c",
           282 => x"80",
           283 => x"8c",
           284 => x"c0",
           285 => x"8c",
           286 => x"80",
           287 => x"8c",
           288 => x"c3",
           289 => x"8c",
           290 => x"80",
           291 => x"8c",
           292 => x"97",
           293 => x"8c",
           294 => x"80",
           295 => x"8c",
           296 => x"c6",
           297 => x"8c",
           298 => x"80",
           299 => x"8c",
           300 => x"d5",
           301 => x"8c",
           302 => x"80",
           303 => x"8c",
           304 => x"d3",
           305 => x"8c",
           306 => x"80",
           307 => x"8c",
           308 => x"e8",
           309 => x"8c",
           310 => x"80",
           311 => x"8c",
           312 => x"ea",
           313 => x"8c",
           314 => x"80",
           315 => x"8c",
           316 => x"ec",
           317 => x"8c",
           318 => x"80",
           319 => x"8c",
           320 => x"c3",
           321 => x"e8",
           322 => x"90",
           323 => x"e8",
           324 => x"2d",
           325 => x"08",
           326 => x"04",
           327 => x"0c",
           328 => x"82",
           329 => x"83",
           330 => x"82",
           331 => x"81",
           332 => x"82",
           333 => x"83",
           334 => x"82",
           335 => x"82",
           336 => x"8e",
           337 => x"70",
           338 => x"0c",
           339 => x"aa",
           340 => x"80",
           341 => x"a0",
           342 => x"82",
           343 => x"02",
           344 => x"0c",
           345 => x"80",
           346 => x"e8",
           347 => x"08",
           348 => x"e8",
           349 => x"08",
           350 => x"3f",
           351 => x"08",
           352 => x"dc",
           353 => x"3d",
           354 => x"e8",
           355 => x"8c",
           356 => x"82",
           357 => x"fd",
           358 => x"53",
           359 => x"08",
           360 => x"52",
           361 => x"08",
           362 => x"51",
           363 => x"8c",
           364 => x"82",
           365 => x"54",
           366 => x"82",
           367 => x"04",
           368 => x"08",
           369 => x"e8",
           370 => x"0d",
           371 => x"8c",
           372 => x"05",
           373 => x"82",
           374 => x"f8",
           375 => x"8c",
           376 => x"05",
           377 => x"e8",
           378 => x"08",
           379 => x"82",
           380 => x"fc",
           381 => x"2e",
           382 => x"0b",
           383 => x"08",
           384 => x"24",
           385 => x"8c",
           386 => x"05",
           387 => x"8c",
           388 => x"05",
           389 => x"e8",
           390 => x"08",
           391 => x"e8",
           392 => x"0c",
           393 => x"82",
           394 => x"fc",
           395 => x"2e",
           396 => x"82",
           397 => x"8c",
           398 => x"8c",
           399 => x"05",
           400 => x"38",
           401 => x"08",
           402 => x"82",
           403 => x"8c",
           404 => x"82",
           405 => x"88",
           406 => x"8c",
           407 => x"05",
           408 => x"e8",
           409 => x"08",
           410 => x"e8",
           411 => x"0c",
           412 => x"08",
           413 => x"81",
           414 => x"e8",
           415 => x"0c",
           416 => x"08",
           417 => x"81",
           418 => x"e8",
           419 => x"0c",
           420 => x"82",
           421 => x"90",
           422 => x"2e",
           423 => x"8c",
           424 => x"05",
           425 => x"8c",
           426 => x"05",
           427 => x"39",
           428 => x"08",
           429 => x"70",
           430 => x"08",
           431 => x"51",
           432 => x"08",
           433 => x"82",
           434 => x"85",
           435 => x"8c",
           436 => x"fc",
           437 => x"70",
           438 => x"55",
           439 => x"72",
           440 => x"72",
           441 => x"06",
           442 => x"2e",
           443 => x"12",
           444 => x"2e",
           445 => x"70",
           446 => x"33",
           447 => x"05",
           448 => x"12",
           449 => x"2e",
           450 => x"ea",
           451 => x"8c",
           452 => x"3d",
           453 => x"51",
           454 => x"05",
           455 => x"70",
           456 => x"0c",
           457 => x"05",
           458 => x"70",
           459 => x"0c",
           460 => x"05",
           461 => x"70",
           462 => x"0c",
           463 => x"05",
           464 => x"70",
           465 => x"0c",
           466 => x"71",
           467 => x"38",
           468 => x"95",
           469 => x"84",
           470 => x"71",
           471 => x"53",
           472 => x"52",
           473 => x"ed",
           474 => x"ff",
           475 => x"3d",
           476 => x"71",
           477 => x"9f",
           478 => x"55",
           479 => x"72",
           480 => x"74",
           481 => x"70",
           482 => x"38",
           483 => x"71",
           484 => x"38",
           485 => x"81",
           486 => x"ff",
           487 => x"ff",
           488 => x"06",
           489 => x"82",
           490 => x"86",
           491 => x"74",
           492 => x"75",
           493 => x"90",
           494 => x"54",
           495 => x"27",
           496 => x"71",
           497 => x"53",
           498 => x"70",
           499 => x"0c",
           500 => x"84",
           501 => x"72",
           502 => x"05",
           503 => x"12",
           504 => x"26",
           505 => x"72",
           506 => x"72",
           507 => x"05",
           508 => x"12",
           509 => x"26",
           510 => x"53",
           511 => x"fc",
           512 => x"70",
           513 => x"07",
           514 => x"54",
           515 => x"80",
           516 => x"70",
           517 => x"70",
           518 => x"ff",
           519 => x"f8",
           520 => x"80",
           521 => x"53",
           522 => x"a6",
           523 => x"72",
           524 => x"05",
           525 => x"08",
           526 => x"f7",
           527 => x"13",
           528 => x"84",
           529 => x"06",
           530 => x"53",
           531 => x"2e",
           532 => x"52",
           533 => x"05",
           534 => x"70",
           535 => x"05",
           536 => x"f0",
           537 => x"8c",
           538 => x"3d",
           539 => x"3d",
           540 => x"71",
           541 => x"55",
           542 => x"38",
           543 => x"70",
           544 => x"fd",
           545 => x"70",
           546 => x"81",
           547 => x"51",
           548 => x"9d",
           549 => x"70",
           550 => x"f7",
           551 => x"12",
           552 => x"84",
           553 => x"06",
           554 => x"53",
           555 => x"e5",
           556 => x"71",
           557 => x"80",
           558 => x"81",
           559 => x"52",
           560 => x"38",
           561 => x"82",
           562 => x"85",
           563 => x"fa",
           564 => x"7a",
           565 => x"55",
           566 => x"80",
           567 => x"38",
           568 => x"83",
           569 => x"80",
           570 => x"38",
           571 => x"72",
           572 => x"38",
           573 => x"33",
           574 => x"71",
           575 => x"06",
           576 => x"80",
           577 => x"38",
           578 => x"06",
           579 => x"2e",
           580 => x"81",
           581 => x"ff",
           582 => x"52",
           583 => x"09",
           584 => x"38",
           585 => x"33",
           586 => x"81",
           587 => x"81",
           588 => x"71",
           589 => x"52",
           590 => x"dc",
           591 => x"0d",
           592 => x"57",
           593 => x"27",
           594 => x"08",
           595 => x"88",
           596 => x"55",
           597 => x"39",
           598 => x"72",
           599 => x"38",
           600 => x"09",
           601 => x"ff",
           602 => x"f8",
           603 => x"80",
           604 => x"51",
           605 => x"84",
           606 => x"57",
           607 => x"27",
           608 => x"08",
           609 => x"d0",
           610 => x"55",
           611 => x"39",
           612 => x"8c",
           613 => x"3d",
           614 => x"3d",
           615 => x"83",
           616 => x"2b",
           617 => x"3f",
           618 => x"08",
           619 => x"72",
           620 => x"54",
           621 => x"25",
           622 => x"82",
           623 => x"84",
           624 => x"fb",
           625 => x"70",
           626 => x"53",
           627 => x"2e",
           628 => x"71",
           629 => x"a0",
           630 => x"06",
           631 => x"12",
           632 => x"71",
           633 => x"81",
           634 => x"73",
           635 => x"ff",
           636 => x"55",
           637 => x"83",
           638 => x"70",
           639 => x"38",
           640 => x"73",
           641 => x"51",
           642 => x"09",
           643 => x"38",
           644 => x"81",
           645 => x"72",
           646 => x"51",
           647 => x"dc",
           648 => x"0d",
           649 => x"0d",
           650 => x"08",
           651 => x"38",
           652 => x"05",
           653 => x"9f",
           654 => x"8c",
           655 => x"38",
           656 => x"39",
           657 => x"82",
           658 => x"86",
           659 => x"fc",
           660 => x"82",
           661 => x"05",
           662 => x"52",
           663 => x"81",
           664 => x"13",
           665 => x"51",
           666 => x"9e",
           667 => x"38",
           668 => x"51",
           669 => x"97",
           670 => x"38",
           671 => x"51",
           672 => x"bb",
           673 => x"38",
           674 => x"51",
           675 => x"bb",
           676 => x"38",
           677 => x"55",
           678 => x"87",
           679 => x"d9",
           680 => x"22",
           681 => x"73",
           682 => x"80",
           683 => x"0b",
           684 => x"9c",
           685 => x"87",
           686 => x"0c",
           687 => x"87",
           688 => x"0c",
           689 => x"87",
           690 => x"0c",
           691 => x"87",
           692 => x"0c",
           693 => x"87",
           694 => x"0c",
           695 => x"87",
           696 => x"0c",
           697 => x"98",
           698 => x"87",
           699 => x"0c",
           700 => x"c0",
           701 => x"80",
           702 => x"8c",
           703 => x"3d",
           704 => x"3d",
           705 => x"87",
           706 => x"5d",
           707 => x"87",
           708 => x"08",
           709 => x"23",
           710 => x"b8",
           711 => x"82",
           712 => x"c0",
           713 => x"5a",
           714 => x"34",
           715 => x"b0",
           716 => x"84",
           717 => x"c0",
           718 => x"5a",
           719 => x"34",
           720 => x"a8",
           721 => x"86",
           722 => x"c0",
           723 => x"5c",
           724 => x"23",
           725 => x"a0",
           726 => x"8a",
           727 => x"7d",
           728 => x"ff",
           729 => x"7b",
           730 => x"06",
           731 => x"33",
           732 => x"33",
           733 => x"33",
           734 => x"33",
           735 => x"33",
           736 => x"ff",
           737 => x"81",
           738 => x"98",
           739 => x"3d",
           740 => x"3d",
           741 => x"05",
           742 => x"70",
           743 => x"52",
           744 => x"0b",
           745 => x"34",
           746 => x"04",
           747 => x"77",
           748 => x"87",
           749 => x"81",
           750 => x"55",
           751 => x"94",
           752 => x"80",
           753 => x"87",
           754 => x"51",
           755 => x"96",
           756 => x"06",
           757 => x"70",
           758 => x"38",
           759 => x"70",
           760 => x"51",
           761 => x"72",
           762 => x"81",
           763 => x"70",
           764 => x"38",
           765 => x"70",
           766 => x"51",
           767 => x"38",
           768 => x"06",
           769 => x"94",
           770 => x"80",
           771 => x"87",
           772 => x"52",
           773 => x"75",
           774 => x"0c",
           775 => x"04",
           776 => x"02",
           777 => x"0b",
           778 => x"d4",
           779 => x"ff",
           780 => x"56",
           781 => x"84",
           782 => x"2e",
           783 => x"c0",
           784 => x"70",
           785 => x"2a",
           786 => x"53",
           787 => x"80",
           788 => x"71",
           789 => x"81",
           790 => x"70",
           791 => x"81",
           792 => x"06",
           793 => x"80",
           794 => x"71",
           795 => x"81",
           796 => x"70",
           797 => x"73",
           798 => x"51",
           799 => x"80",
           800 => x"2e",
           801 => x"c0",
           802 => x"75",
           803 => x"3d",
           804 => x"3d",
           805 => x"80",
           806 => x"81",
           807 => x"53",
           808 => x"2e",
           809 => x"71",
           810 => x"81",
           811 => x"82",
           812 => x"70",
           813 => x"59",
           814 => x"87",
           815 => x"51",
           816 => x"86",
           817 => x"94",
           818 => x"08",
           819 => x"70",
           820 => x"54",
           821 => x"2e",
           822 => x"91",
           823 => x"06",
           824 => x"d7",
           825 => x"32",
           826 => x"51",
           827 => x"2e",
           828 => x"93",
           829 => x"06",
           830 => x"ff",
           831 => x"81",
           832 => x"87",
           833 => x"52",
           834 => x"86",
           835 => x"94",
           836 => x"72",
           837 => x"74",
           838 => x"ff",
           839 => x"57",
           840 => x"38",
           841 => x"dc",
           842 => x"0d",
           843 => x"0d",
           844 => x"87",
           845 => x"81",
           846 => x"52",
           847 => x"84",
           848 => x"2e",
           849 => x"c0",
           850 => x"70",
           851 => x"2a",
           852 => x"51",
           853 => x"80",
           854 => x"71",
           855 => x"51",
           856 => x"80",
           857 => x"2e",
           858 => x"c0",
           859 => x"71",
           860 => x"ff",
           861 => x"dc",
           862 => x"3d",
           863 => x"3d",
           864 => x"82",
           865 => x"70",
           866 => x"52",
           867 => x"94",
           868 => x"80",
           869 => x"87",
           870 => x"52",
           871 => x"82",
           872 => x"06",
           873 => x"ff",
           874 => x"2e",
           875 => x"81",
           876 => x"87",
           877 => x"52",
           878 => x"86",
           879 => x"94",
           880 => x"08",
           881 => x"70",
           882 => x"53",
           883 => x"8c",
           884 => x"3d",
           885 => x"3d",
           886 => x"9e",
           887 => x"9c",
           888 => x"51",
           889 => x"2e",
           890 => x"87",
           891 => x"08",
           892 => x"0c",
           893 => x"a8",
           894 => x"dc",
           895 => x"9e",
           896 => x"87",
           897 => x"c0",
           898 => x"82",
           899 => x"87",
           900 => x"08",
           901 => x"0c",
           902 => x"a0",
           903 => x"ec",
           904 => x"9e",
           905 => x"87",
           906 => x"c0",
           907 => x"82",
           908 => x"87",
           909 => x"08",
           910 => x"0c",
           911 => x"b8",
           912 => x"fc",
           913 => x"9e",
           914 => x"88",
           915 => x"c0",
           916 => x"82",
           917 => x"87",
           918 => x"08",
           919 => x"0c",
           920 => x"80",
           921 => x"82",
           922 => x"87",
           923 => x"08",
           924 => x"0c",
           925 => x"88",
           926 => x"94",
           927 => x"9e",
           928 => x"88",
           929 => x"0b",
           930 => x"34",
           931 => x"c0",
           932 => x"70",
           933 => x"06",
           934 => x"70",
           935 => x"38",
           936 => x"82",
           937 => x"80",
           938 => x"9e",
           939 => x"88",
           940 => x"51",
           941 => x"80",
           942 => x"81",
           943 => x"88",
           944 => x"0b",
           945 => x"90",
           946 => x"80",
           947 => x"52",
           948 => x"2e",
           949 => x"52",
           950 => x"9f",
           951 => x"87",
           952 => x"08",
           953 => x"80",
           954 => x"52",
           955 => x"83",
           956 => x"71",
           957 => x"34",
           958 => x"c0",
           959 => x"70",
           960 => x"06",
           961 => x"70",
           962 => x"38",
           963 => x"82",
           964 => x"80",
           965 => x"9e",
           966 => x"90",
           967 => x"51",
           968 => x"80",
           969 => x"81",
           970 => x"88",
           971 => x"0b",
           972 => x"90",
           973 => x"80",
           974 => x"52",
           975 => x"2e",
           976 => x"52",
           977 => x"a3",
           978 => x"87",
           979 => x"08",
           980 => x"80",
           981 => x"52",
           982 => x"83",
           983 => x"71",
           984 => x"34",
           985 => x"c0",
           986 => x"70",
           987 => x"06",
           988 => x"70",
           989 => x"38",
           990 => x"82",
           991 => x"80",
           992 => x"9e",
           993 => x"80",
           994 => x"51",
           995 => x"80",
           996 => x"81",
           997 => x"88",
           998 => x"0b",
           999 => x"90",
          1000 => x"80",
          1001 => x"52",
          1002 => x"83",
          1003 => x"71",
          1004 => x"34",
          1005 => x"90",
          1006 => x"80",
          1007 => x"2a",
          1008 => x"70",
          1009 => x"34",
          1010 => x"c0",
          1011 => x"70",
          1012 => x"51",
          1013 => x"80",
          1014 => x"81",
          1015 => x"88",
          1016 => x"c0",
          1017 => x"70",
          1018 => x"70",
          1019 => x"51",
          1020 => x"88",
          1021 => x"0b",
          1022 => x"90",
          1023 => x"06",
          1024 => x"70",
          1025 => x"38",
          1026 => x"82",
          1027 => x"87",
          1028 => x"08",
          1029 => x"51",
          1030 => x"88",
          1031 => x"3d",
          1032 => x"3d",
          1033 => x"fc",
          1034 => x"3f",
          1035 => x"33",
          1036 => x"2e",
          1037 => x"f2",
          1038 => x"cb",
          1039 => x"a4",
          1040 => x"3f",
          1041 => x"33",
          1042 => x"2e",
          1043 => x"87",
          1044 => x"87",
          1045 => x"54",
          1046 => x"bc",
          1047 => x"3f",
          1048 => x"33",
          1049 => x"2e",
          1050 => x"87",
          1051 => x"87",
          1052 => x"54",
          1053 => x"d8",
          1054 => x"3f",
          1055 => x"33",
          1056 => x"2e",
          1057 => x"87",
          1058 => x"87",
          1059 => x"54",
          1060 => x"f4",
          1061 => x"3f",
          1062 => x"33",
          1063 => x"2e",
          1064 => x"87",
          1065 => x"87",
          1066 => x"54",
          1067 => x"90",
          1068 => x"3f",
          1069 => x"33",
          1070 => x"2e",
          1071 => x"87",
          1072 => x"87",
          1073 => x"54",
          1074 => x"ac",
          1075 => x"3f",
          1076 => x"33",
          1077 => x"2e",
          1078 => x"88",
          1079 => x"81",
          1080 => x"8e",
          1081 => x"88",
          1082 => x"73",
          1083 => x"38",
          1084 => x"33",
          1085 => x"e8",
          1086 => x"3f",
          1087 => x"33",
          1088 => x"2e",
          1089 => x"88",
          1090 => x"81",
          1091 => x"8d",
          1092 => x"88",
          1093 => x"73",
          1094 => x"38",
          1095 => x"51",
          1096 => x"82",
          1097 => x"54",
          1098 => x"88",
          1099 => x"bc",
          1100 => x"3f",
          1101 => x"33",
          1102 => x"2e",
          1103 => x"f4",
          1104 => x"c3",
          1105 => x"a5",
          1106 => x"80",
          1107 => x"81",
          1108 => x"87",
          1109 => x"88",
          1110 => x"73",
          1111 => x"38",
          1112 => x"51",
          1113 => x"81",
          1114 => x"87",
          1115 => x"88",
          1116 => x"81",
          1117 => x"8c",
          1118 => x"88",
          1119 => x"81",
          1120 => x"8c",
          1121 => x"88",
          1122 => x"81",
          1123 => x"8c",
          1124 => x"f5",
          1125 => x"ef",
          1126 => x"8c",
          1127 => x"f5",
          1128 => x"c7",
          1129 => x"90",
          1130 => x"84",
          1131 => x"51",
          1132 => x"82",
          1133 => x"bd",
          1134 => x"76",
          1135 => x"54",
          1136 => x"08",
          1137 => x"a0",
          1138 => x"3f",
          1139 => x"33",
          1140 => x"2e",
          1141 => x"88",
          1142 => x"bd",
          1143 => x"75",
          1144 => x"3f",
          1145 => x"08",
          1146 => x"29",
          1147 => x"54",
          1148 => x"dc",
          1149 => x"f6",
          1150 => x"ef",
          1151 => x"9e",
          1152 => x"80",
          1153 => x"82",
          1154 => x"56",
          1155 => x"52",
          1156 => x"c7",
          1157 => x"dc",
          1158 => x"c0",
          1159 => x"31",
          1160 => x"8c",
          1161 => x"81",
          1162 => x"8b",
          1163 => x"85",
          1164 => x"d3",
          1165 => x"0d",
          1166 => x"0d",
          1167 => x"33",
          1168 => x"71",
          1169 => x"38",
          1170 => x"0b",
          1171 => x"d0",
          1172 => x"08",
          1173 => x"a4",
          1174 => x"81",
          1175 => x"97",
          1176 => x"b4",
          1177 => x"81",
          1178 => x"8b",
          1179 => x"c0",
          1180 => x"81",
          1181 => x"85",
          1182 => x"3d",
          1183 => x"88",
          1184 => x"80",
          1185 => x"96",
          1186 => x"82",
          1187 => x"87",
          1188 => x"0c",
          1189 => x"0d",
          1190 => x"08",
          1191 => x"a4",
          1192 => x"8c",
          1193 => x"8c",
          1194 => x"11",
          1195 => x"53",
          1196 => x"f8",
          1197 => x"70",
          1198 => x"0c",
          1199 => x"82",
          1200 => x"84",
          1201 => x"f9",
          1202 => x"7b",
          1203 => x"a0",
          1204 => x"08",
          1205 => x"90",
          1206 => x"58",
          1207 => x"53",
          1208 => x"ba",
          1209 => x"88",
          1210 => x"51",
          1211 => x"76",
          1212 => x"12",
          1213 => x"0c",
          1214 => x"0c",
          1215 => x"0c",
          1216 => x"0c",
          1217 => x"0c",
          1218 => x"0c",
          1219 => x"0c",
          1220 => x"0c",
          1221 => x"0c",
          1222 => x"0c",
          1223 => x"73",
          1224 => x"16",
          1225 => x"15",
          1226 => x"8c",
          1227 => x"3d",
          1228 => x"3d",
          1229 => x"11",
          1230 => x"08",
          1231 => x"71",
          1232 => x"09",
          1233 => x"38",
          1234 => x"70",
          1235 => x"70",
          1236 => x"81",
          1237 => x"84",
          1238 => x"84",
          1239 => x"88",
          1240 => x"8c",
          1241 => x"53",
          1242 => x"73",
          1243 => x"c4",
          1244 => x"0c",
          1245 => x"0b",
          1246 => x"72",
          1247 => x"0c",
          1248 => x"73",
          1249 => x"51",
          1250 => x"2e",
          1251 => x"b3",
          1252 => x"08",
          1253 => x"52",
          1254 => x"09",
          1255 => x"38",
          1256 => x"12",
          1257 => x"94",
          1258 => x"15",
          1259 => x"13",
          1260 => x"12",
          1261 => x"08",
          1262 => x"70",
          1263 => x"52",
          1264 => x"72",
          1265 => x"0c",
          1266 => x"04",
          1267 => x"79",
          1268 => x"76",
          1269 => x"b5",
          1270 => x"f0",
          1271 => x"c4",
          1272 => x"75",
          1273 => x"8f",
          1274 => x"08",
          1275 => x"c7",
          1276 => x"08",
          1277 => x"83",
          1278 => x"fc",
          1279 => x"70",
          1280 => x"91",
          1281 => x"dc",
          1282 => x"dc",
          1283 => x"82",
          1284 => x"07",
          1285 => x"8c",
          1286 => x"70",
          1287 => x"07",
          1288 => x"07",
          1289 => x"51",
          1290 => x"54",
          1291 => x"09",
          1292 => x"d9",
          1293 => x"76",
          1294 => x"80",
          1295 => x"0b",
          1296 => x"08",
          1297 => x"8c",
          1298 => x"05",
          1299 => x"c0",
          1300 => x"08",
          1301 => x"38",
          1302 => x"87",
          1303 => x"08",
          1304 => x"88",
          1305 => x"17",
          1306 => x"17",
          1307 => x"14",
          1308 => x"08",
          1309 => x"0c",
          1310 => x"fd",
          1311 => x"52",
          1312 => x"08",
          1313 => x"3f",
          1314 => x"08",
          1315 => x"8c",
          1316 => x"3d",
          1317 => x"3d",
          1318 => x"71",
          1319 => x"38",
          1320 => x"fd",
          1321 => x"3d",
          1322 => x"3d",
          1323 => x"05",
          1324 => x"8a",
          1325 => x"06",
          1326 => x"51",
          1327 => x"8c",
          1328 => x"71",
          1329 => x"38",
          1330 => x"82",
          1331 => x"81",
          1332 => x"f8",
          1333 => x"82",
          1334 => x"52",
          1335 => x"85",
          1336 => x"71",
          1337 => x"0d",
          1338 => x"0d",
          1339 => x"33",
          1340 => x"08",
          1341 => x"f0",
          1342 => x"ff",
          1343 => x"82",
          1344 => x"84",
          1345 => x"fd",
          1346 => x"54",
          1347 => x"81",
          1348 => x"53",
          1349 => x"8e",
          1350 => x"ff",
          1351 => x"14",
          1352 => x"3f",
          1353 => x"3d",
          1354 => x"3d",
          1355 => x"8c",
          1356 => x"82",
          1357 => x"56",
          1358 => x"70",
          1359 => x"53",
          1360 => x"2e",
          1361 => x"81",
          1362 => x"81",
          1363 => x"da",
          1364 => x"74",
          1365 => x"0c",
          1366 => x"04",
          1367 => x"66",
          1368 => x"78",
          1369 => x"5a",
          1370 => x"80",
          1371 => x"38",
          1372 => x"09",
          1373 => x"de",
          1374 => x"7a",
          1375 => x"5c",
          1376 => x"5b",
          1377 => x"09",
          1378 => x"38",
          1379 => x"39",
          1380 => x"09",
          1381 => x"38",
          1382 => x"70",
          1383 => x"33",
          1384 => x"2e",
          1385 => x"92",
          1386 => x"19",
          1387 => x"70",
          1388 => x"33",
          1389 => x"53",
          1390 => x"16",
          1391 => x"26",
          1392 => x"88",
          1393 => x"05",
          1394 => x"05",
          1395 => x"05",
          1396 => x"5b",
          1397 => x"80",
          1398 => x"30",
          1399 => x"80",
          1400 => x"cc",
          1401 => x"70",
          1402 => x"25",
          1403 => x"54",
          1404 => x"53",
          1405 => x"8c",
          1406 => x"07",
          1407 => x"05",
          1408 => x"5a",
          1409 => x"83",
          1410 => x"54",
          1411 => x"27",
          1412 => x"16",
          1413 => x"06",
          1414 => x"80",
          1415 => x"aa",
          1416 => x"cf",
          1417 => x"73",
          1418 => x"81",
          1419 => x"80",
          1420 => x"38",
          1421 => x"2e",
          1422 => x"81",
          1423 => x"80",
          1424 => x"8a",
          1425 => x"39",
          1426 => x"2e",
          1427 => x"73",
          1428 => x"8a",
          1429 => x"d3",
          1430 => x"80",
          1431 => x"80",
          1432 => x"ee",
          1433 => x"39",
          1434 => x"71",
          1435 => x"53",
          1436 => x"54",
          1437 => x"2e",
          1438 => x"15",
          1439 => x"33",
          1440 => x"72",
          1441 => x"81",
          1442 => x"39",
          1443 => x"56",
          1444 => x"27",
          1445 => x"51",
          1446 => x"75",
          1447 => x"72",
          1448 => x"38",
          1449 => x"df",
          1450 => x"16",
          1451 => x"7b",
          1452 => x"38",
          1453 => x"f2",
          1454 => x"77",
          1455 => x"12",
          1456 => x"53",
          1457 => x"5c",
          1458 => x"5c",
          1459 => x"5c",
          1460 => x"5c",
          1461 => x"51",
          1462 => x"fd",
          1463 => x"82",
          1464 => x"06",
          1465 => x"80",
          1466 => x"77",
          1467 => x"53",
          1468 => x"18",
          1469 => x"72",
          1470 => x"c4",
          1471 => x"70",
          1472 => x"25",
          1473 => x"55",
          1474 => x"8d",
          1475 => x"2e",
          1476 => x"30",
          1477 => x"5b",
          1478 => x"8f",
          1479 => x"7b",
          1480 => x"dc",
          1481 => x"8c",
          1482 => x"ff",
          1483 => x"75",
          1484 => x"a7",
          1485 => x"dc",
          1486 => x"74",
          1487 => x"a7",
          1488 => x"80",
          1489 => x"38",
          1490 => x"72",
          1491 => x"54",
          1492 => x"72",
          1493 => x"05",
          1494 => x"17",
          1495 => x"77",
          1496 => x"51",
          1497 => x"9f",
          1498 => x"72",
          1499 => x"79",
          1500 => x"81",
          1501 => x"72",
          1502 => x"38",
          1503 => x"05",
          1504 => x"ad",
          1505 => x"17",
          1506 => x"81",
          1507 => x"b0",
          1508 => x"38",
          1509 => x"81",
          1510 => x"06",
          1511 => x"9f",
          1512 => x"55",
          1513 => x"97",
          1514 => x"f9",
          1515 => x"81",
          1516 => x"8b",
          1517 => x"16",
          1518 => x"73",
          1519 => x"96",
          1520 => x"e0",
          1521 => x"17",
          1522 => x"33",
          1523 => x"f9",
          1524 => x"f2",
          1525 => x"16",
          1526 => x"7b",
          1527 => x"38",
          1528 => x"c6",
          1529 => x"96",
          1530 => x"fd",
          1531 => x"3d",
          1532 => x"05",
          1533 => x"52",
          1534 => x"e0",
          1535 => x"0d",
          1536 => x"0d",
          1537 => x"f8",
          1538 => x"88",
          1539 => x"51",
          1540 => x"82",
          1541 => x"53",
          1542 => x"80",
          1543 => x"f8",
          1544 => x"0d",
          1545 => x"0d",
          1546 => x"08",
          1547 => x"f0",
          1548 => x"88",
          1549 => x"52",
          1550 => x"3f",
          1551 => x"f0",
          1552 => x"0d",
          1553 => x"0d",
          1554 => x"8c",
          1555 => x"56",
          1556 => x"80",
          1557 => x"2e",
          1558 => x"82",
          1559 => x"52",
          1560 => x"8c",
          1561 => x"ff",
          1562 => x"80",
          1563 => x"38",
          1564 => x"b9",
          1565 => x"32",
          1566 => x"80",
          1567 => x"52",
          1568 => x"8b",
          1569 => x"2e",
          1570 => x"14",
          1571 => x"9f",
          1572 => x"38",
          1573 => x"73",
          1574 => x"38",
          1575 => x"72",
          1576 => x"14",
          1577 => x"f8",
          1578 => x"af",
          1579 => x"52",
          1580 => x"8a",
          1581 => x"3f",
          1582 => x"82",
          1583 => x"87",
          1584 => x"fe",
          1585 => x"8c",
          1586 => x"82",
          1587 => x"77",
          1588 => x"53",
          1589 => x"72",
          1590 => x"0c",
          1591 => x"04",
          1592 => x"7a",
          1593 => x"80",
          1594 => x"58",
          1595 => x"33",
          1596 => x"a0",
          1597 => x"06",
          1598 => x"13",
          1599 => x"39",
          1600 => x"09",
          1601 => x"38",
          1602 => x"11",
          1603 => x"08",
          1604 => x"54",
          1605 => x"2e",
          1606 => x"80",
          1607 => x"08",
          1608 => x"0c",
          1609 => x"33",
          1610 => x"80",
          1611 => x"38",
          1612 => x"80",
          1613 => x"38",
          1614 => x"57",
          1615 => x"0c",
          1616 => x"33",
          1617 => x"39",
          1618 => x"74",
          1619 => x"38",
          1620 => x"80",
          1621 => x"89",
          1622 => x"38",
          1623 => x"d0",
          1624 => x"55",
          1625 => x"80",
          1626 => x"39",
          1627 => x"d9",
          1628 => x"80",
          1629 => x"27",
          1630 => x"80",
          1631 => x"89",
          1632 => x"70",
          1633 => x"55",
          1634 => x"70",
          1635 => x"55",
          1636 => x"27",
          1637 => x"14",
          1638 => x"06",
          1639 => x"74",
          1640 => x"73",
          1641 => x"38",
          1642 => x"14",
          1643 => x"05",
          1644 => x"08",
          1645 => x"54",
          1646 => x"39",
          1647 => x"84",
          1648 => x"55",
          1649 => x"81",
          1650 => x"8c",
          1651 => x"3d",
          1652 => x"3d",
          1653 => x"5a",
          1654 => x"7a",
          1655 => x"08",
          1656 => x"53",
          1657 => x"09",
          1658 => x"38",
          1659 => x"0c",
          1660 => x"ad",
          1661 => x"06",
          1662 => x"76",
          1663 => x"0c",
          1664 => x"33",
          1665 => x"73",
          1666 => x"81",
          1667 => x"38",
          1668 => x"05",
          1669 => x"08",
          1670 => x"53",
          1671 => x"2e",
          1672 => x"57",
          1673 => x"2e",
          1674 => x"39",
          1675 => x"13",
          1676 => x"08",
          1677 => x"53",
          1678 => x"55",
          1679 => x"80",
          1680 => x"14",
          1681 => x"88",
          1682 => x"27",
          1683 => x"eb",
          1684 => x"53",
          1685 => x"89",
          1686 => x"38",
          1687 => x"55",
          1688 => x"8a",
          1689 => x"a0",
          1690 => x"c2",
          1691 => x"74",
          1692 => x"e0",
          1693 => x"ff",
          1694 => x"d0",
          1695 => x"ff",
          1696 => x"90",
          1697 => x"38",
          1698 => x"81",
          1699 => x"53",
          1700 => x"ca",
          1701 => x"27",
          1702 => x"77",
          1703 => x"08",
          1704 => x"0c",
          1705 => x"33",
          1706 => x"ff",
          1707 => x"80",
          1708 => x"74",
          1709 => x"79",
          1710 => x"74",
          1711 => x"0c",
          1712 => x"04",
          1713 => x"76",
          1714 => x"98",
          1715 => x"2b",
          1716 => x"72",
          1717 => x"82",
          1718 => x"51",
          1719 => x"80",
          1720 => x"dc",
          1721 => x"53",
          1722 => x"9c",
          1723 => x"d8",
          1724 => x"02",
          1725 => x"05",
          1726 => x"52",
          1727 => x"72",
          1728 => x"06",
          1729 => x"53",
          1730 => x"dc",
          1731 => x"0d",
          1732 => x"0d",
          1733 => x"05",
          1734 => x"71",
          1735 => x"53",
          1736 => x"9f",
          1737 => x"f3",
          1738 => x"51",
          1739 => x"88",
          1740 => x"3f",
          1741 => x"05",
          1742 => x"34",
          1743 => x"06",
          1744 => x"76",
          1745 => x"3f",
          1746 => x"86",
          1747 => x"f6",
          1748 => x"02",
          1749 => x"05",
          1750 => x"05",
          1751 => x"82",
          1752 => x"70",
          1753 => x"88",
          1754 => x"08",
          1755 => x"5a",
          1756 => x"80",
          1757 => x"74",
          1758 => x"3f",
          1759 => x"33",
          1760 => x"82",
          1761 => x"81",
          1762 => x"58",
          1763 => x"bc",
          1764 => x"dc",
          1765 => x"82",
          1766 => x"70",
          1767 => x"88",
          1768 => x"08",
          1769 => x"74",
          1770 => x"38",
          1771 => x"52",
          1772 => x"9f",
          1773 => x"a8",
          1774 => x"55",
          1775 => x"a8",
          1776 => x"ff",
          1777 => x"75",
          1778 => x"80",
          1779 => x"a8",
          1780 => x"2e",
          1781 => x"89",
          1782 => x"75",
          1783 => x"38",
          1784 => x"33",
          1785 => x"38",
          1786 => x"05",
          1787 => x"78",
          1788 => x"80",
          1789 => x"82",
          1790 => x"52",
          1791 => x"fd",
          1792 => x"89",
          1793 => x"80",
          1794 => x"8c",
          1795 => x"dc",
          1796 => x"57",
          1797 => x"89",
          1798 => x"80",
          1799 => x"82",
          1800 => x"80",
          1801 => x"89",
          1802 => x"80",
          1803 => x"3d",
          1804 => x"80",
          1805 => x"82",
          1806 => x"80",
          1807 => x"75",
          1808 => x"3f",
          1809 => x"08",
          1810 => x"82",
          1811 => x"25",
          1812 => x"8c",
          1813 => x"05",
          1814 => x"55",
          1815 => x"75",
          1816 => x"81",
          1817 => x"f0",
          1818 => x"ff",
          1819 => x"2e",
          1820 => x"ff",
          1821 => x"3d",
          1822 => x"3d",
          1823 => x"08",
          1824 => x"5a",
          1825 => x"58",
          1826 => x"82",
          1827 => x"51",
          1828 => x"3f",
          1829 => x"08",
          1830 => x"ff",
          1831 => x"a4",
          1832 => x"80",
          1833 => x"3d",
          1834 => x"80",
          1835 => x"82",
          1836 => x"80",
          1837 => x"75",
          1838 => x"3f",
          1839 => x"08",
          1840 => x"55",
          1841 => x"8c",
          1842 => x"8e",
          1843 => x"dc",
          1844 => x"70",
          1845 => x"80",
          1846 => x"09",
          1847 => x"72",
          1848 => x"51",
          1849 => x"77",
          1850 => x"73",
          1851 => x"82",
          1852 => x"8c",
          1853 => x"51",
          1854 => x"3f",
          1855 => x"08",
          1856 => x"38",
          1857 => x"51",
          1858 => x"78",
          1859 => x"81",
          1860 => x"75",
          1861 => x"d5",
          1862 => x"51",
          1863 => x"ab",
          1864 => x"82",
          1865 => x"74",
          1866 => x"77",
          1867 => x"0c",
          1868 => x"04",
          1869 => x"7c",
          1870 => x"71",
          1871 => x"59",
          1872 => x"a0",
          1873 => x"06",
          1874 => x"33",
          1875 => x"77",
          1876 => x"38",
          1877 => x"5b",
          1878 => x"56",
          1879 => x"a0",
          1880 => x"06",
          1881 => x"75",
          1882 => x"80",
          1883 => x"29",
          1884 => x"05",
          1885 => x"55",
          1886 => x"82",
          1887 => x"53",
          1888 => x"08",
          1889 => x"3f",
          1890 => x"08",
          1891 => x"84",
          1892 => x"74",
          1893 => x"38",
          1894 => x"88",
          1895 => x"fc",
          1896 => x"39",
          1897 => x"8c",
          1898 => x"53",
          1899 => x"f6",
          1900 => x"8c",
          1901 => x"2e",
          1902 => x"53",
          1903 => x"51",
          1904 => x"82",
          1905 => x"81",
          1906 => x"74",
          1907 => x"54",
          1908 => x"14",
          1909 => x"06",
          1910 => x"74",
          1911 => x"38",
          1912 => x"82",
          1913 => x"8c",
          1914 => x"d3",
          1915 => x"3d",
          1916 => x"05",
          1917 => x"33",
          1918 => x"0b",
          1919 => x"82",
          1920 => x"5b",
          1921 => x"08",
          1922 => x"82",
          1923 => x"54",
          1924 => x"38",
          1925 => x"b4",
          1926 => x"dc",
          1927 => x"a4",
          1928 => x"dc",
          1929 => x"80",
          1930 => x"53",
          1931 => x"08",
          1932 => x"dc",
          1933 => x"ed",
          1934 => x"dc",
          1935 => x"8b",
          1936 => x"a8",
          1937 => x"3f",
          1938 => x"82",
          1939 => x"53",
          1940 => x"90",
          1941 => x"54",
          1942 => x"3f",
          1943 => x"08",
          1944 => x"dc",
          1945 => x"09",
          1946 => x"c1",
          1947 => x"dc",
          1948 => x"fa",
          1949 => x"dc",
          1950 => x"0b",
          1951 => x"08",
          1952 => x"82",
          1953 => x"ff",
          1954 => x"55",
          1955 => x"34",
          1956 => x"81",
          1957 => x"75",
          1958 => x"3f",
          1959 => x"09",
          1960 => x"a7",
          1961 => x"81",
          1962 => x"a0",
          1963 => x"5d",
          1964 => x"82",
          1965 => x"98",
          1966 => x"2c",
          1967 => x"ff",
          1968 => x"78",
          1969 => x"82",
          1970 => x"70",
          1971 => x"98",
          1972 => x"fc",
          1973 => x"2b",
          1974 => x"71",
          1975 => x"70",
          1976 => x"f8",
          1977 => x"08",
          1978 => x"51",
          1979 => x"59",
          1980 => x"5d",
          1981 => x"73",
          1982 => x"e9",
          1983 => x"27",
          1984 => x"81",
          1985 => x"81",
          1986 => x"70",
          1987 => x"55",
          1988 => x"80",
          1989 => x"53",
          1990 => x"51",
          1991 => x"82",
          1992 => x"81",
          1993 => x"73",
          1994 => x"38",
          1995 => x"fc",
          1996 => x"b1",
          1997 => x"80",
          1998 => x"80",
          1999 => x"98",
          2000 => x"ff",
          2001 => x"55",
          2002 => x"97",
          2003 => x"74",
          2004 => x"f6",
          2005 => x"8c",
          2006 => x"ff",
          2007 => x"cc",
          2008 => x"80",
          2009 => x"2e",
          2010 => x"81",
          2011 => x"82",
          2012 => x"74",
          2013 => x"98",
          2014 => x"fc",
          2015 => x"2b",
          2016 => x"70",
          2017 => x"82",
          2018 => x"dc",
          2019 => x"51",
          2020 => x"58",
          2021 => x"77",
          2022 => x"06",
          2023 => x"81",
          2024 => x"08",
          2025 => x"0b",
          2026 => x"34",
          2027 => x"8c",
          2028 => x"39",
          2029 => x"80",
          2030 => x"8c",
          2031 => x"af",
          2032 => x"7d",
          2033 => x"73",
          2034 => x"e1",
          2035 => x"29",
          2036 => x"05",
          2037 => x"04",
          2038 => x"33",
          2039 => x"2e",
          2040 => x"82",
          2041 => x"55",
          2042 => x"ab",
          2043 => x"2b",
          2044 => x"51",
          2045 => x"24",
          2046 => x"1a",
          2047 => x"81",
          2048 => x"81",
          2049 => x"81",
          2050 => x"70",
          2051 => x"8d",
          2052 => x"51",
          2053 => x"82",
          2054 => x"81",
          2055 => x"74",
          2056 => x"34",
          2057 => x"ae",
          2058 => x"34",
          2059 => x"33",
          2060 => x"27",
          2061 => x"14",
          2062 => x"8d",
          2063 => x"8d",
          2064 => x"81",
          2065 => x"81",
          2066 => x"70",
          2067 => x"8d",
          2068 => x"51",
          2069 => x"77",
          2070 => x"74",
          2071 => x"52",
          2072 => x"3f",
          2073 => x"0a",
          2074 => x"0a",
          2075 => x"2c",
          2076 => x"33",
          2077 => x"73",
          2078 => x"38",
          2079 => x"33",
          2080 => x"70",
          2081 => x"8d",
          2082 => x"51",
          2083 => x"77",
          2084 => x"38",
          2085 => x"92",
          2086 => x"80",
          2087 => x"80",
          2088 => x"98",
          2089 => x"84",
          2090 => x"55",
          2091 => x"e4",
          2092 => x"39",
          2093 => x"33",
          2094 => x"06",
          2095 => x"80",
          2096 => x"38",
          2097 => x"33",
          2098 => x"73",
          2099 => x"34",
          2100 => x"73",
          2101 => x"34",
          2102 => x"ce",
          2103 => x"88",
          2104 => x"2b",
          2105 => x"82",
          2106 => x"57",
          2107 => x"74",
          2108 => x"38",
          2109 => x"81",
          2110 => x"34",
          2111 => x"e7",
          2112 => x"81",
          2113 => x"81",
          2114 => x"70",
          2115 => x"8d",
          2116 => x"51",
          2117 => x"24",
          2118 => x"51",
          2119 => x"82",
          2120 => x"70",
          2121 => x"98",
          2122 => x"84",
          2123 => x"56",
          2124 => x"24",
          2125 => x"88",
          2126 => x"3f",
          2127 => x"0a",
          2128 => x"0a",
          2129 => x"2c",
          2130 => x"33",
          2131 => x"75",
          2132 => x"38",
          2133 => x"82",
          2134 => x"7a",
          2135 => x"74",
          2136 => x"e6",
          2137 => x"8d",
          2138 => x"51",
          2139 => x"82",
          2140 => x"81",
          2141 => x"73",
          2142 => x"8d",
          2143 => x"73",
          2144 => x"c9",
          2145 => x"73",
          2146 => x"f3",
          2147 => x"bd",
          2148 => x"34",
          2149 => x"82",
          2150 => x"54",
          2151 => x"fa",
          2152 => x"51",
          2153 => x"82",
          2154 => x"ff",
          2155 => x"82",
          2156 => x"73",
          2157 => x"54",
          2158 => x"8d",
          2159 => x"8d",
          2160 => x"55",
          2161 => x"f9",
          2162 => x"14",
          2163 => x"8d",
          2164 => x"98",
          2165 => x"2c",
          2166 => x"06",
          2167 => x"74",
          2168 => x"38",
          2169 => x"81",
          2170 => x"34",
          2171 => x"e5",
          2172 => x"81",
          2173 => x"81",
          2174 => x"70",
          2175 => x"8d",
          2176 => x"51",
          2177 => x"24",
          2178 => x"51",
          2179 => x"82",
          2180 => x"70",
          2181 => x"98",
          2182 => x"84",
          2183 => x"56",
          2184 => x"24",
          2185 => x"88",
          2186 => x"3f",
          2187 => x"0a",
          2188 => x"0a",
          2189 => x"2c",
          2190 => x"33",
          2191 => x"75",
          2192 => x"38",
          2193 => x"82",
          2194 => x"70",
          2195 => x"82",
          2196 => x"59",
          2197 => x"77",
          2198 => x"38",
          2199 => x"73",
          2200 => x"34",
          2201 => x"33",
          2202 => x"be",
          2203 => x"88",
          2204 => x"ff",
          2205 => x"84",
          2206 => x"54",
          2207 => x"dc",
          2208 => x"39",
          2209 => x"82",
          2210 => x"55",
          2211 => x"a4",
          2212 => x"cb",
          2213 => x"8c",
          2214 => x"8d",
          2215 => x"8c",
          2216 => x"ff",
          2217 => x"53",
          2218 => x"51",
          2219 => x"93",
          2220 => x"39",
          2221 => x"82",
          2222 => x"fc",
          2223 => x"54",
          2224 => x"a5",
          2225 => x"cb",
          2226 => x"8c",
          2227 => x"8d",
          2228 => x"8c",
          2229 => x"ff",
          2230 => x"53",
          2231 => x"51",
          2232 => x"ff",
          2233 => x"de",
          2234 => x"55",
          2235 => x"f7",
          2236 => x"51",
          2237 => x"80",
          2238 => x"93",
          2239 => x"06",
          2240 => x"88",
          2241 => x"74",
          2242 => x"38",
          2243 => x"de",
          2244 => x"39",
          2245 => x"82",
          2246 => x"84",
          2247 => x"54",
          2248 => x"a9",
          2249 => x"ca",
          2250 => x"8c",
          2251 => x"8d",
          2252 => x"8c",
          2253 => x"ff",
          2254 => x"53",
          2255 => x"51",
          2256 => x"81",
          2257 => x"81",
          2258 => x"a8",
          2259 => x"55",
          2260 => x"f6",
          2261 => x"51",
          2262 => x"82",
          2263 => x"82",
          2264 => x"82",
          2265 => x"81",
          2266 => x"05",
          2267 => x"79",
          2268 => x"3f",
          2269 => x"53",
          2270 => x"33",
          2271 => x"ef",
          2272 => x"a9",
          2273 => x"88",
          2274 => x"ff",
          2275 => x"84",
          2276 => x"54",
          2277 => x"f6",
          2278 => x"14",
          2279 => x"8d",
          2280 => x"1a",
          2281 => x"54",
          2282 => x"f6",
          2283 => x"8d",
          2284 => x"73",
          2285 => x"f5",
          2286 => x"e1",
          2287 => x"8d",
          2288 => x"05",
          2289 => x"8d",
          2290 => x"e1",
          2291 => x"82",
          2292 => x"80",
          2293 => x"84",
          2294 => x"8c",
          2295 => x"3d",
          2296 => x"3d",
          2297 => x"05",
          2298 => x"52",
          2299 => x"87",
          2300 => x"c4",
          2301 => x"71",
          2302 => x"0c",
          2303 => x"04",
          2304 => x"02",
          2305 => x"02",
          2306 => x"05",
          2307 => x"83",
          2308 => x"26",
          2309 => x"72",
          2310 => x"c0",
          2311 => x"53",
          2312 => x"74",
          2313 => x"38",
          2314 => x"73",
          2315 => x"c0",
          2316 => x"51",
          2317 => x"85",
          2318 => x"98",
          2319 => x"52",
          2320 => x"82",
          2321 => x"70",
          2322 => x"38",
          2323 => x"8c",
          2324 => x"ec",
          2325 => x"fc",
          2326 => x"52",
          2327 => x"87",
          2328 => x"08",
          2329 => x"2e",
          2330 => x"82",
          2331 => x"34",
          2332 => x"13",
          2333 => x"82",
          2334 => x"86",
          2335 => x"f3",
          2336 => x"62",
          2337 => x"05",
          2338 => x"57",
          2339 => x"83",
          2340 => x"fe",
          2341 => x"8c",
          2342 => x"06",
          2343 => x"71",
          2344 => x"71",
          2345 => x"2b",
          2346 => x"80",
          2347 => x"92",
          2348 => x"c0",
          2349 => x"41",
          2350 => x"5a",
          2351 => x"87",
          2352 => x"0c",
          2353 => x"84",
          2354 => x"08",
          2355 => x"70",
          2356 => x"53",
          2357 => x"2e",
          2358 => x"08",
          2359 => x"70",
          2360 => x"34",
          2361 => x"80",
          2362 => x"53",
          2363 => x"2e",
          2364 => x"53",
          2365 => x"26",
          2366 => x"80",
          2367 => x"87",
          2368 => x"08",
          2369 => x"38",
          2370 => x"8c",
          2371 => x"80",
          2372 => x"78",
          2373 => x"99",
          2374 => x"0c",
          2375 => x"8c",
          2376 => x"08",
          2377 => x"51",
          2378 => x"38",
          2379 => x"8d",
          2380 => x"17",
          2381 => x"81",
          2382 => x"53",
          2383 => x"2e",
          2384 => x"fc",
          2385 => x"52",
          2386 => x"7d",
          2387 => x"ed",
          2388 => x"80",
          2389 => x"71",
          2390 => x"38",
          2391 => x"53",
          2392 => x"dc",
          2393 => x"0d",
          2394 => x"0d",
          2395 => x"02",
          2396 => x"05",
          2397 => x"58",
          2398 => x"80",
          2399 => x"fc",
          2400 => x"8c",
          2401 => x"06",
          2402 => x"71",
          2403 => x"81",
          2404 => x"38",
          2405 => x"2b",
          2406 => x"80",
          2407 => x"92",
          2408 => x"c0",
          2409 => x"40",
          2410 => x"5a",
          2411 => x"c0",
          2412 => x"76",
          2413 => x"76",
          2414 => x"75",
          2415 => x"2a",
          2416 => x"51",
          2417 => x"80",
          2418 => x"7a",
          2419 => x"5c",
          2420 => x"81",
          2421 => x"81",
          2422 => x"06",
          2423 => x"80",
          2424 => x"87",
          2425 => x"08",
          2426 => x"38",
          2427 => x"8c",
          2428 => x"80",
          2429 => x"77",
          2430 => x"99",
          2431 => x"0c",
          2432 => x"8c",
          2433 => x"08",
          2434 => x"51",
          2435 => x"38",
          2436 => x"8d",
          2437 => x"70",
          2438 => x"84",
          2439 => x"5b",
          2440 => x"2e",
          2441 => x"fc",
          2442 => x"52",
          2443 => x"7d",
          2444 => x"f8",
          2445 => x"80",
          2446 => x"71",
          2447 => x"38",
          2448 => x"53",
          2449 => x"dc",
          2450 => x"0d",
          2451 => x"0d",
          2452 => x"05",
          2453 => x"02",
          2454 => x"05",
          2455 => x"54",
          2456 => x"fe",
          2457 => x"dc",
          2458 => x"53",
          2459 => x"80",
          2460 => x"0b",
          2461 => x"8c",
          2462 => x"71",
          2463 => x"dc",
          2464 => x"24",
          2465 => x"84",
          2466 => x"92",
          2467 => x"54",
          2468 => x"8d",
          2469 => x"39",
          2470 => x"80",
          2471 => x"cb",
          2472 => x"70",
          2473 => x"81",
          2474 => x"52",
          2475 => x"8a",
          2476 => x"98",
          2477 => x"71",
          2478 => x"c0",
          2479 => x"52",
          2480 => x"81",
          2481 => x"c0",
          2482 => x"53",
          2483 => x"82",
          2484 => x"71",
          2485 => x"39",
          2486 => x"39",
          2487 => x"77",
          2488 => x"81",
          2489 => x"72",
          2490 => x"84",
          2491 => x"73",
          2492 => x"0c",
          2493 => x"04",
          2494 => x"74",
          2495 => x"71",
          2496 => x"2b",
          2497 => x"dc",
          2498 => x"84",
          2499 => x"fd",
          2500 => x"83",
          2501 => x"12",
          2502 => x"2b",
          2503 => x"07",
          2504 => x"70",
          2505 => x"2b",
          2506 => x"07",
          2507 => x"0c",
          2508 => x"56",
          2509 => x"3d",
          2510 => x"3d",
          2511 => x"84",
          2512 => x"22",
          2513 => x"72",
          2514 => x"54",
          2515 => x"2a",
          2516 => x"34",
          2517 => x"04",
          2518 => x"73",
          2519 => x"70",
          2520 => x"05",
          2521 => x"88",
          2522 => x"72",
          2523 => x"54",
          2524 => x"2a",
          2525 => x"70",
          2526 => x"34",
          2527 => x"51",
          2528 => x"83",
          2529 => x"fe",
          2530 => x"75",
          2531 => x"51",
          2532 => x"92",
          2533 => x"81",
          2534 => x"73",
          2535 => x"55",
          2536 => x"51",
          2537 => x"3d",
          2538 => x"3d",
          2539 => x"76",
          2540 => x"72",
          2541 => x"05",
          2542 => x"11",
          2543 => x"38",
          2544 => x"04",
          2545 => x"78",
          2546 => x"56",
          2547 => x"81",
          2548 => x"74",
          2549 => x"56",
          2550 => x"31",
          2551 => x"52",
          2552 => x"80",
          2553 => x"71",
          2554 => x"38",
          2555 => x"dc",
          2556 => x"0d",
          2557 => x"0d",
          2558 => x"51",
          2559 => x"73",
          2560 => x"81",
          2561 => x"33",
          2562 => x"38",
          2563 => x"8c",
          2564 => x"3d",
          2565 => x"0b",
          2566 => x"0c",
          2567 => x"82",
          2568 => x"04",
          2569 => x"7b",
          2570 => x"83",
          2571 => x"5a",
          2572 => x"80",
          2573 => x"54",
          2574 => x"53",
          2575 => x"53",
          2576 => x"52",
          2577 => x"3f",
          2578 => x"08",
          2579 => x"81",
          2580 => x"82",
          2581 => x"83",
          2582 => x"16",
          2583 => x"18",
          2584 => x"18",
          2585 => x"58",
          2586 => x"9f",
          2587 => x"33",
          2588 => x"2e",
          2589 => x"93",
          2590 => x"76",
          2591 => x"52",
          2592 => x"51",
          2593 => x"83",
          2594 => x"79",
          2595 => x"0c",
          2596 => x"04",
          2597 => x"78",
          2598 => x"80",
          2599 => x"17",
          2600 => x"38",
          2601 => x"fc",
          2602 => x"dc",
          2603 => x"8c",
          2604 => x"38",
          2605 => x"53",
          2606 => x"81",
          2607 => x"f7",
          2608 => x"8c",
          2609 => x"2e",
          2610 => x"55",
          2611 => x"b0",
          2612 => x"82",
          2613 => x"88",
          2614 => x"f8",
          2615 => x"70",
          2616 => x"c0",
          2617 => x"dc",
          2618 => x"8c",
          2619 => x"91",
          2620 => x"55",
          2621 => x"09",
          2622 => x"f0",
          2623 => x"33",
          2624 => x"2e",
          2625 => x"80",
          2626 => x"80",
          2627 => x"dc",
          2628 => x"17",
          2629 => x"fd",
          2630 => x"d4",
          2631 => x"b2",
          2632 => x"96",
          2633 => x"85",
          2634 => x"75",
          2635 => x"3f",
          2636 => x"e4",
          2637 => x"98",
          2638 => x"9c",
          2639 => x"08",
          2640 => x"17",
          2641 => x"3f",
          2642 => x"52",
          2643 => x"51",
          2644 => x"a0",
          2645 => x"05",
          2646 => x"0c",
          2647 => x"75",
          2648 => x"33",
          2649 => x"3f",
          2650 => x"34",
          2651 => x"52",
          2652 => x"51",
          2653 => x"82",
          2654 => x"80",
          2655 => x"81",
          2656 => x"8c",
          2657 => x"3d",
          2658 => x"3d",
          2659 => x"1a",
          2660 => x"fe",
          2661 => x"54",
          2662 => x"73",
          2663 => x"8a",
          2664 => x"71",
          2665 => x"08",
          2666 => x"75",
          2667 => x"0c",
          2668 => x"04",
          2669 => x"7a",
          2670 => x"56",
          2671 => x"77",
          2672 => x"38",
          2673 => x"08",
          2674 => x"38",
          2675 => x"54",
          2676 => x"2e",
          2677 => x"72",
          2678 => x"38",
          2679 => x"8d",
          2680 => x"39",
          2681 => x"81",
          2682 => x"b6",
          2683 => x"2a",
          2684 => x"2a",
          2685 => x"05",
          2686 => x"55",
          2687 => x"82",
          2688 => x"81",
          2689 => x"83",
          2690 => x"b4",
          2691 => x"17",
          2692 => x"a4",
          2693 => x"55",
          2694 => x"57",
          2695 => x"3f",
          2696 => x"08",
          2697 => x"74",
          2698 => x"14",
          2699 => x"70",
          2700 => x"07",
          2701 => x"71",
          2702 => x"52",
          2703 => x"72",
          2704 => x"75",
          2705 => x"58",
          2706 => x"76",
          2707 => x"15",
          2708 => x"73",
          2709 => x"3f",
          2710 => x"08",
          2711 => x"76",
          2712 => x"06",
          2713 => x"05",
          2714 => x"3f",
          2715 => x"08",
          2716 => x"06",
          2717 => x"76",
          2718 => x"15",
          2719 => x"73",
          2720 => x"3f",
          2721 => x"08",
          2722 => x"82",
          2723 => x"06",
          2724 => x"05",
          2725 => x"3f",
          2726 => x"08",
          2727 => x"58",
          2728 => x"58",
          2729 => x"dc",
          2730 => x"0d",
          2731 => x"0d",
          2732 => x"5a",
          2733 => x"59",
          2734 => x"82",
          2735 => x"98",
          2736 => x"82",
          2737 => x"33",
          2738 => x"2e",
          2739 => x"72",
          2740 => x"38",
          2741 => x"8d",
          2742 => x"39",
          2743 => x"81",
          2744 => x"f7",
          2745 => x"2a",
          2746 => x"2a",
          2747 => x"05",
          2748 => x"55",
          2749 => x"82",
          2750 => x"59",
          2751 => x"08",
          2752 => x"74",
          2753 => x"16",
          2754 => x"16",
          2755 => x"59",
          2756 => x"53",
          2757 => x"8f",
          2758 => x"2b",
          2759 => x"74",
          2760 => x"71",
          2761 => x"72",
          2762 => x"0b",
          2763 => x"74",
          2764 => x"17",
          2765 => x"75",
          2766 => x"3f",
          2767 => x"08",
          2768 => x"dc",
          2769 => x"38",
          2770 => x"06",
          2771 => x"78",
          2772 => x"54",
          2773 => x"77",
          2774 => x"33",
          2775 => x"71",
          2776 => x"51",
          2777 => x"34",
          2778 => x"76",
          2779 => x"17",
          2780 => x"75",
          2781 => x"3f",
          2782 => x"08",
          2783 => x"dc",
          2784 => x"38",
          2785 => x"ff",
          2786 => x"10",
          2787 => x"76",
          2788 => x"51",
          2789 => x"be",
          2790 => x"2a",
          2791 => x"05",
          2792 => x"f9",
          2793 => x"8c",
          2794 => x"82",
          2795 => x"ab",
          2796 => x"0a",
          2797 => x"2b",
          2798 => x"70",
          2799 => x"70",
          2800 => x"54",
          2801 => x"82",
          2802 => x"8f",
          2803 => x"07",
          2804 => x"f7",
          2805 => x"0b",
          2806 => x"78",
          2807 => x"0c",
          2808 => x"04",
          2809 => x"7a",
          2810 => x"08",
          2811 => x"59",
          2812 => x"a4",
          2813 => x"17",
          2814 => x"38",
          2815 => x"aa",
          2816 => x"73",
          2817 => x"fd",
          2818 => x"8c",
          2819 => x"82",
          2820 => x"80",
          2821 => x"39",
          2822 => x"eb",
          2823 => x"80",
          2824 => x"8c",
          2825 => x"80",
          2826 => x"52",
          2827 => x"84",
          2828 => x"dc",
          2829 => x"8c",
          2830 => x"2e",
          2831 => x"82",
          2832 => x"81",
          2833 => x"82",
          2834 => x"ff",
          2835 => x"80",
          2836 => x"75",
          2837 => x"3f",
          2838 => x"08",
          2839 => x"16",
          2840 => x"90",
          2841 => x"55",
          2842 => x"27",
          2843 => x"15",
          2844 => x"84",
          2845 => x"07",
          2846 => x"17",
          2847 => x"76",
          2848 => x"a6",
          2849 => x"73",
          2850 => x"0c",
          2851 => x"04",
          2852 => x"7c",
          2853 => x"59",
          2854 => x"95",
          2855 => x"08",
          2856 => x"2e",
          2857 => x"17",
          2858 => x"b2",
          2859 => x"ae",
          2860 => x"7a",
          2861 => x"3f",
          2862 => x"82",
          2863 => x"27",
          2864 => x"82",
          2865 => x"55",
          2866 => x"08",
          2867 => x"d2",
          2868 => x"08",
          2869 => x"08",
          2870 => x"38",
          2871 => x"17",
          2872 => x"54",
          2873 => x"82",
          2874 => x"7a",
          2875 => x"06",
          2876 => x"81",
          2877 => x"17",
          2878 => x"83",
          2879 => x"75",
          2880 => x"f9",
          2881 => x"59",
          2882 => x"08",
          2883 => x"81",
          2884 => x"82",
          2885 => x"59",
          2886 => x"08",
          2887 => x"70",
          2888 => x"25",
          2889 => x"82",
          2890 => x"54",
          2891 => x"55",
          2892 => x"38",
          2893 => x"08",
          2894 => x"38",
          2895 => x"54",
          2896 => x"90",
          2897 => x"18",
          2898 => x"38",
          2899 => x"39",
          2900 => x"38",
          2901 => x"16",
          2902 => x"08",
          2903 => x"38",
          2904 => x"78",
          2905 => x"38",
          2906 => x"51",
          2907 => x"82",
          2908 => x"80",
          2909 => x"80",
          2910 => x"dc",
          2911 => x"09",
          2912 => x"38",
          2913 => x"08",
          2914 => x"dc",
          2915 => x"30",
          2916 => x"80",
          2917 => x"07",
          2918 => x"55",
          2919 => x"38",
          2920 => x"09",
          2921 => x"ae",
          2922 => x"80",
          2923 => x"53",
          2924 => x"51",
          2925 => x"82",
          2926 => x"82",
          2927 => x"30",
          2928 => x"dc",
          2929 => x"25",
          2930 => x"79",
          2931 => x"38",
          2932 => x"8f",
          2933 => x"79",
          2934 => x"f9",
          2935 => x"8c",
          2936 => x"74",
          2937 => x"8c",
          2938 => x"17",
          2939 => x"90",
          2940 => x"54",
          2941 => x"86",
          2942 => x"90",
          2943 => x"17",
          2944 => x"54",
          2945 => x"34",
          2946 => x"56",
          2947 => x"90",
          2948 => x"80",
          2949 => x"82",
          2950 => x"55",
          2951 => x"56",
          2952 => x"82",
          2953 => x"8c",
          2954 => x"f8",
          2955 => x"70",
          2956 => x"f0",
          2957 => x"dc",
          2958 => x"56",
          2959 => x"08",
          2960 => x"7b",
          2961 => x"f6",
          2962 => x"8c",
          2963 => x"8c",
          2964 => x"17",
          2965 => x"80",
          2966 => x"b4",
          2967 => x"57",
          2968 => x"77",
          2969 => x"81",
          2970 => x"15",
          2971 => x"78",
          2972 => x"81",
          2973 => x"53",
          2974 => x"15",
          2975 => x"e9",
          2976 => x"dc",
          2977 => x"df",
          2978 => x"22",
          2979 => x"30",
          2980 => x"70",
          2981 => x"51",
          2982 => x"82",
          2983 => x"8a",
          2984 => x"f8",
          2985 => x"7c",
          2986 => x"56",
          2987 => x"80",
          2988 => x"f1",
          2989 => x"06",
          2990 => x"e9",
          2991 => x"18",
          2992 => x"08",
          2993 => x"38",
          2994 => x"82",
          2995 => x"38",
          2996 => x"54",
          2997 => x"74",
          2998 => x"82",
          2999 => x"22",
          3000 => x"79",
          3001 => x"38",
          3002 => x"98",
          3003 => x"cd",
          3004 => x"22",
          3005 => x"54",
          3006 => x"26",
          3007 => x"52",
          3008 => x"b0",
          3009 => x"dc",
          3010 => x"8c",
          3011 => x"2e",
          3012 => x"0b",
          3013 => x"08",
          3014 => x"98",
          3015 => x"8c",
          3016 => x"85",
          3017 => x"bd",
          3018 => x"31",
          3019 => x"73",
          3020 => x"f4",
          3021 => x"8c",
          3022 => x"18",
          3023 => x"18",
          3024 => x"08",
          3025 => x"72",
          3026 => x"38",
          3027 => x"58",
          3028 => x"89",
          3029 => x"18",
          3030 => x"ff",
          3031 => x"05",
          3032 => x"80",
          3033 => x"8c",
          3034 => x"3d",
          3035 => x"3d",
          3036 => x"08",
          3037 => x"a0",
          3038 => x"54",
          3039 => x"77",
          3040 => x"80",
          3041 => x"0c",
          3042 => x"53",
          3043 => x"80",
          3044 => x"38",
          3045 => x"06",
          3046 => x"b5",
          3047 => x"98",
          3048 => x"14",
          3049 => x"92",
          3050 => x"2a",
          3051 => x"56",
          3052 => x"26",
          3053 => x"80",
          3054 => x"16",
          3055 => x"77",
          3056 => x"53",
          3057 => x"38",
          3058 => x"51",
          3059 => x"82",
          3060 => x"53",
          3061 => x"0b",
          3062 => x"08",
          3063 => x"38",
          3064 => x"8c",
          3065 => x"2e",
          3066 => x"98",
          3067 => x"8c",
          3068 => x"80",
          3069 => x"8a",
          3070 => x"15",
          3071 => x"80",
          3072 => x"14",
          3073 => x"51",
          3074 => x"82",
          3075 => x"53",
          3076 => x"8c",
          3077 => x"2e",
          3078 => x"82",
          3079 => x"dc",
          3080 => x"ba",
          3081 => x"82",
          3082 => x"ff",
          3083 => x"82",
          3084 => x"52",
          3085 => x"f3",
          3086 => x"dc",
          3087 => x"72",
          3088 => x"72",
          3089 => x"f2",
          3090 => x"8c",
          3091 => x"15",
          3092 => x"15",
          3093 => x"b4",
          3094 => x"0c",
          3095 => x"82",
          3096 => x"8a",
          3097 => x"f7",
          3098 => x"7d",
          3099 => x"5b",
          3100 => x"76",
          3101 => x"3f",
          3102 => x"08",
          3103 => x"dc",
          3104 => x"38",
          3105 => x"08",
          3106 => x"08",
          3107 => x"f0",
          3108 => x"8c",
          3109 => x"82",
          3110 => x"80",
          3111 => x"8c",
          3112 => x"18",
          3113 => x"51",
          3114 => x"81",
          3115 => x"81",
          3116 => x"81",
          3117 => x"dc",
          3118 => x"83",
          3119 => x"77",
          3120 => x"72",
          3121 => x"38",
          3122 => x"75",
          3123 => x"81",
          3124 => x"a5",
          3125 => x"dc",
          3126 => x"52",
          3127 => x"8e",
          3128 => x"dc",
          3129 => x"8c",
          3130 => x"2e",
          3131 => x"73",
          3132 => x"81",
          3133 => x"87",
          3134 => x"8c",
          3135 => x"3d",
          3136 => x"3d",
          3137 => x"11",
          3138 => x"ec",
          3139 => x"dc",
          3140 => x"ff",
          3141 => x"33",
          3142 => x"71",
          3143 => x"81",
          3144 => x"94",
          3145 => x"d0",
          3146 => x"dc",
          3147 => x"73",
          3148 => x"82",
          3149 => x"85",
          3150 => x"fc",
          3151 => x"79",
          3152 => x"ff",
          3153 => x"12",
          3154 => x"eb",
          3155 => x"70",
          3156 => x"72",
          3157 => x"81",
          3158 => x"73",
          3159 => x"94",
          3160 => x"d6",
          3161 => x"0d",
          3162 => x"0d",
          3163 => x"55",
          3164 => x"5a",
          3165 => x"08",
          3166 => x"8a",
          3167 => x"08",
          3168 => x"ee",
          3169 => x"8c",
          3170 => x"82",
          3171 => x"80",
          3172 => x"15",
          3173 => x"55",
          3174 => x"38",
          3175 => x"e6",
          3176 => x"33",
          3177 => x"70",
          3178 => x"58",
          3179 => x"86",
          3180 => x"8c",
          3181 => x"73",
          3182 => x"83",
          3183 => x"73",
          3184 => x"38",
          3185 => x"06",
          3186 => x"80",
          3187 => x"75",
          3188 => x"38",
          3189 => x"08",
          3190 => x"54",
          3191 => x"2e",
          3192 => x"83",
          3193 => x"73",
          3194 => x"38",
          3195 => x"51",
          3196 => x"82",
          3197 => x"58",
          3198 => x"08",
          3199 => x"15",
          3200 => x"38",
          3201 => x"0b",
          3202 => x"77",
          3203 => x"0c",
          3204 => x"04",
          3205 => x"77",
          3206 => x"54",
          3207 => x"51",
          3208 => x"82",
          3209 => x"55",
          3210 => x"08",
          3211 => x"14",
          3212 => x"51",
          3213 => x"82",
          3214 => x"55",
          3215 => x"08",
          3216 => x"53",
          3217 => x"08",
          3218 => x"08",
          3219 => x"3f",
          3220 => x"14",
          3221 => x"08",
          3222 => x"3f",
          3223 => x"17",
          3224 => x"8c",
          3225 => x"3d",
          3226 => x"3d",
          3227 => x"08",
          3228 => x"54",
          3229 => x"53",
          3230 => x"82",
          3231 => x"8d",
          3232 => x"08",
          3233 => x"34",
          3234 => x"15",
          3235 => x"0d",
          3236 => x"0d",
          3237 => x"57",
          3238 => x"17",
          3239 => x"08",
          3240 => x"82",
          3241 => x"89",
          3242 => x"55",
          3243 => x"14",
          3244 => x"16",
          3245 => x"71",
          3246 => x"38",
          3247 => x"09",
          3248 => x"38",
          3249 => x"73",
          3250 => x"81",
          3251 => x"ae",
          3252 => x"05",
          3253 => x"15",
          3254 => x"70",
          3255 => x"34",
          3256 => x"8a",
          3257 => x"38",
          3258 => x"05",
          3259 => x"81",
          3260 => x"17",
          3261 => x"12",
          3262 => x"34",
          3263 => x"9c",
          3264 => x"e8",
          3265 => x"8c",
          3266 => x"0c",
          3267 => x"e7",
          3268 => x"8c",
          3269 => x"17",
          3270 => x"51",
          3271 => x"82",
          3272 => x"84",
          3273 => x"3d",
          3274 => x"3d",
          3275 => x"08",
          3276 => x"61",
          3277 => x"55",
          3278 => x"2e",
          3279 => x"55",
          3280 => x"2e",
          3281 => x"80",
          3282 => x"94",
          3283 => x"1c",
          3284 => x"81",
          3285 => x"61",
          3286 => x"56",
          3287 => x"2e",
          3288 => x"83",
          3289 => x"73",
          3290 => x"70",
          3291 => x"25",
          3292 => x"51",
          3293 => x"38",
          3294 => x"0c",
          3295 => x"51",
          3296 => x"26",
          3297 => x"80",
          3298 => x"34",
          3299 => x"51",
          3300 => x"82",
          3301 => x"55",
          3302 => x"91",
          3303 => x"1d",
          3304 => x"8b",
          3305 => x"79",
          3306 => x"3f",
          3307 => x"57",
          3308 => x"55",
          3309 => x"2e",
          3310 => x"80",
          3311 => x"18",
          3312 => x"1a",
          3313 => x"70",
          3314 => x"2a",
          3315 => x"07",
          3316 => x"5a",
          3317 => x"8c",
          3318 => x"54",
          3319 => x"81",
          3320 => x"39",
          3321 => x"70",
          3322 => x"2a",
          3323 => x"75",
          3324 => x"8c",
          3325 => x"2e",
          3326 => x"a0",
          3327 => x"38",
          3328 => x"0c",
          3329 => x"76",
          3330 => x"38",
          3331 => x"b8",
          3332 => x"70",
          3333 => x"5a",
          3334 => x"76",
          3335 => x"38",
          3336 => x"70",
          3337 => x"dc",
          3338 => x"72",
          3339 => x"80",
          3340 => x"51",
          3341 => x"73",
          3342 => x"38",
          3343 => x"18",
          3344 => x"1a",
          3345 => x"55",
          3346 => x"2e",
          3347 => x"83",
          3348 => x"73",
          3349 => x"70",
          3350 => x"25",
          3351 => x"51",
          3352 => x"38",
          3353 => x"75",
          3354 => x"81",
          3355 => x"81",
          3356 => x"27",
          3357 => x"73",
          3358 => x"38",
          3359 => x"70",
          3360 => x"32",
          3361 => x"80",
          3362 => x"2a",
          3363 => x"56",
          3364 => x"81",
          3365 => x"57",
          3366 => x"f5",
          3367 => x"2b",
          3368 => x"25",
          3369 => x"80",
          3370 => x"fa",
          3371 => x"57",
          3372 => x"e6",
          3373 => x"8c",
          3374 => x"2e",
          3375 => x"18",
          3376 => x"1a",
          3377 => x"56",
          3378 => x"3f",
          3379 => x"08",
          3380 => x"e8",
          3381 => x"54",
          3382 => x"80",
          3383 => x"17",
          3384 => x"34",
          3385 => x"11",
          3386 => x"74",
          3387 => x"75",
          3388 => x"8c",
          3389 => x"3f",
          3390 => x"08",
          3391 => x"9f",
          3392 => x"99",
          3393 => x"e0",
          3394 => x"ff",
          3395 => x"79",
          3396 => x"74",
          3397 => x"57",
          3398 => x"77",
          3399 => x"76",
          3400 => x"38",
          3401 => x"73",
          3402 => x"09",
          3403 => x"38",
          3404 => x"84",
          3405 => x"27",
          3406 => x"39",
          3407 => x"f2",
          3408 => x"80",
          3409 => x"54",
          3410 => x"34",
          3411 => x"58",
          3412 => x"f2",
          3413 => x"8c",
          3414 => x"82",
          3415 => x"80",
          3416 => x"1b",
          3417 => x"51",
          3418 => x"82",
          3419 => x"56",
          3420 => x"08",
          3421 => x"9c",
          3422 => x"33",
          3423 => x"80",
          3424 => x"38",
          3425 => x"bf",
          3426 => x"86",
          3427 => x"15",
          3428 => x"2a",
          3429 => x"51",
          3430 => x"92",
          3431 => x"79",
          3432 => x"e4",
          3433 => x"8c",
          3434 => x"2e",
          3435 => x"52",
          3436 => x"ba",
          3437 => x"39",
          3438 => x"33",
          3439 => x"80",
          3440 => x"74",
          3441 => x"81",
          3442 => x"38",
          3443 => x"70",
          3444 => x"82",
          3445 => x"54",
          3446 => x"96",
          3447 => x"06",
          3448 => x"2e",
          3449 => x"ff",
          3450 => x"1c",
          3451 => x"80",
          3452 => x"81",
          3453 => x"ba",
          3454 => x"b6",
          3455 => x"2a",
          3456 => x"51",
          3457 => x"38",
          3458 => x"70",
          3459 => x"81",
          3460 => x"55",
          3461 => x"e1",
          3462 => x"08",
          3463 => x"1d",
          3464 => x"7c",
          3465 => x"3f",
          3466 => x"08",
          3467 => x"fa",
          3468 => x"82",
          3469 => x"8f",
          3470 => x"f6",
          3471 => x"5b",
          3472 => x"70",
          3473 => x"59",
          3474 => x"73",
          3475 => x"c6",
          3476 => x"81",
          3477 => x"70",
          3478 => x"52",
          3479 => x"8d",
          3480 => x"38",
          3481 => x"09",
          3482 => x"a5",
          3483 => x"d0",
          3484 => x"ff",
          3485 => x"53",
          3486 => x"91",
          3487 => x"73",
          3488 => x"d0",
          3489 => x"71",
          3490 => x"f7",
          3491 => x"81",
          3492 => x"55",
          3493 => x"55",
          3494 => x"81",
          3495 => x"74",
          3496 => x"56",
          3497 => x"12",
          3498 => x"70",
          3499 => x"38",
          3500 => x"81",
          3501 => x"51",
          3502 => x"51",
          3503 => x"89",
          3504 => x"70",
          3505 => x"53",
          3506 => x"70",
          3507 => x"51",
          3508 => x"09",
          3509 => x"38",
          3510 => x"38",
          3511 => x"77",
          3512 => x"70",
          3513 => x"2a",
          3514 => x"07",
          3515 => x"51",
          3516 => x"8f",
          3517 => x"84",
          3518 => x"83",
          3519 => x"94",
          3520 => x"74",
          3521 => x"38",
          3522 => x"0c",
          3523 => x"86",
          3524 => x"a0",
          3525 => x"82",
          3526 => x"8c",
          3527 => x"fa",
          3528 => x"56",
          3529 => x"17",
          3530 => x"b0",
          3531 => x"52",
          3532 => x"e0",
          3533 => x"82",
          3534 => x"81",
          3535 => x"b2",
          3536 => x"b4",
          3537 => x"dc",
          3538 => x"ff",
          3539 => x"55",
          3540 => x"d5",
          3541 => x"06",
          3542 => x"80",
          3543 => x"33",
          3544 => x"81",
          3545 => x"81",
          3546 => x"81",
          3547 => x"eb",
          3548 => x"70",
          3549 => x"07",
          3550 => x"73",
          3551 => x"81",
          3552 => x"81",
          3553 => x"83",
          3554 => x"9c",
          3555 => x"16",
          3556 => x"3f",
          3557 => x"08",
          3558 => x"dc",
          3559 => x"9d",
          3560 => x"81",
          3561 => x"81",
          3562 => x"e0",
          3563 => x"8c",
          3564 => x"82",
          3565 => x"80",
          3566 => x"82",
          3567 => x"8c",
          3568 => x"3d",
          3569 => x"3d",
          3570 => x"84",
          3571 => x"05",
          3572 => x"80",
          3573 => x"51",
          3574 => x"82",
          3575 => x"58",
          3576 => x"0b",
          3577 => x"08",
          3578 => x"38",
          3579 => x"08",
          3580 => x"8d",
          3581 => x"08",
          3582 => x"56",
          3583 => x"86",
          3584 => x"75",
          3585 => x"fe",
          3586 => x"54",
          3587 => x"2e",
          3588 => x"14",
          3589 => x"ca",
          3590 => x"dc",
          3591 => x"06",
          3592 => x"54",
          3593 => x"38",
          3594 => x"86",
          3595 => x"82",
          3596 => x"06",
          3597 => x"56",
          3598 => x"38",
          3599 => x"80",
          3600 => x"81",
          3601 => x"52",
          3602 => x"51",
          3603 => x"82",
          3604 => x"81",
          3605 => x"81",
          3606 => x"83",
          3607 => x"87",
          3608 => x"2e",
          3609 => x"82",
          3610 => x"06",
          3611 => x"56",
          3612 => x"38",
          3613 => x"74",
          3614 => x"a3",
          3615 => x"dc",
          3616 => x"06",
          3617 => x"2e",
          3618 => x"80",
          3619 => x"3d",
          3620 => x"83",
          3621 => x"15",
          3622 => x"53",
          3623 => x"8d",
          3624 => x"15",
          3625 => x"3f",
          3626 => x"08",
          3627 => x"70",
          3628 => x"0c",
          3629 => x"16",
          3630 => x"80",
          3631 => x"80",
          3632 => x"54",
          3633 => x"84",
          3634 => x"5b",
          3635 => x"80",
          3636 => x"7a",
          3637 => x"fc",
          3638 => x"8c",
          3639 => x"ff",
          3640 => x"77",
          3641 => x"81",
          3642 => x"76",
          3643 => x"81",
          3644 => x"2e",
          3645 => x"8d",
          3646 => x"26",
          3647 => x"bf",
          3648 => x"f4",
          3649 => x"dc",
          3650 => x"ff",
          3651 => x"84",
          3652 => x"81",
          3653 => x"38",
          3654 => x"51",
          3655 => x"82",
          3656 => x"83",
          3657 => x"58",
          3658 => x"80",
          3659 => x"db",
          3660 => x"8c",
          3661 => x"77",
          3662 => x"80",
          3663 => x"82",
          3664 => x"c4",
          3665 => x"11",
          3666 => x"06",
          3667 => x"8d",
          3668 => x"26",
          3669 => x"74",
          3670 => x"78",
          3671 => x"c1",
          3672 => x"59",
          3673 => x"15",
          3674 => x"2e",
          3675 => x"13",
          3676 => x"72",
          3677 => x"38",
          3678 => x"eb",
          3679 => x"14",
          3680 => x"3f",
          3681 => x"08",
          3682 => x"dc",
          3683 => x"23",
          3684 => x"57",
          3685 => x"83",
          3686 => x"c7",
          3687 => x"d8",
          3688 => x"dc",
          3689 => x"ff",
          3690 => x"8d",
          3691 => x"14",
          3692 => x"3f",
          3693 => x"08",
          3694 => x"14",
          3695 => x"3f",
          3696 => x"08",
          3697 => x"06",
          3698 => x"72",
          3699 => x"97",
          3700 => x"22",
          3701 => x"84",
          3702 => x"5a",
          3703 => x"83",
          3704 => x"14",
          3705 => x"79",
          3706 => x"96",
          3707 => x"8c",
          3708 => x"82",
          3709 => x"80",
          3710 => x"38",
          3711 => x"08",
          3712 => x"ff",
          3713 => x"38",
          3714 => x"83",
          3715 => x"83",
          3716 => x"74",
          3717 => x"85",
          3718 => x"89",
          3719 => x"76",
          3720 => x"c3",
          3721 => x"70",
          3722 => x"7b",
          3723 => x"73",
          3724 => x"17",
          3725 => x"ac",
          3726 => x"55",
          3727 => x"09",
          3728 => x"38",
          3729 => x"51",
          3730 => x"82",
          3731 => x"83",
          3732 => x"53",
          3733 => x"82",
          3734 => x"82",
          3735 => x"e0",
          3736 => x"ab",
          3737 => x"dc",
          3738 => x"0c",
          3739 => x"53",
          3740 => x"56",
          3741 => x"81",
          3742 => x"13",
          3743 => x"74",
          3744 => x"82",
          3745 => x"74",
          3746 => x"81",
          3747 => x"06",
          3748 => x"83",
          3749 => x"2a",
          3750 => x"72",
          3751 => x"26",
          3752 => x"ff",
          3753 => x"0c",
          3754 => x"15",
          3755 => x"0b",
          3756 => x"76",
          3757 => x"81",
          3758 => x"38",
          3759 => x"51",
          3760 => x"82",
          3761 => x"83",
          3762 => x"53",
          3763 => x"09",
          3764 => x"f9",
          3765 => x"52",
          3766 => x"b8",
          3767 => x"dc",
          3768 => x"38",
          3769 => x"08",
          3770 => x"84",
          3771 => x"d8",
          3772 => x"8c",
          3773 => x"ff",
          3774 => x"72",
          3775 => x"2e",
          3776 => x"80",
          3777 => x"14",
          3778 => x"3f",
          3779 => x"08",
          3780 => x"a4",
          3781 => x"81",
          3782 => x"84",
          3783 => x"d7",
          3784 => x"8c",
          3785 => x"8a",
          3786 => x"2e",
          3787 => x"9d",
          3788 => x"14",
          3789 => x"3f",
          3790 => x"08",
          3791 => x"84",
          3792 => x"d7",
          3793 => x"8c",
          3794 => x"15",
          3795 => x"34",
          3796 => x"22",
          3797 => x"72",
          3798 => x"23",
          3799 => x"23",
          3800 => x"15",
          3801 => x"75",
          3802 => x"0c",
          3803 => x"04",
          3804 => x"77",
          3805 => x"73",
          3806 => x"38",
          3807 => x"72",
          3808 => x"38",
          3809 => x"71",
          3810 => x"38",
          3811 => x"84",
          3812 => x"52",
          3813 => x"09",
          3814 => x"38",
          3815 => x"51",
          3816 => x"82",
          3817 => x"81",
          3818 => x"88",
          3819 => x"08",
          3820 => x"39",
          3821 => x"73",
          3822 => x"74",
          3823 => x"0c",
          3824 => x"04",
          3825 => x"02",
          3826 => x"7a",
          3827 => x"fc",
          3828 => x"f4",
          3829 => x"54",
          3830 => x"8c",
          3831 => x"bc",
          3832 => x"dc",
          3833 => x"82",
          3834 => x"70",
          3835 => x"73",
          3836 => x"38",
          3837 => x"78",
          3838 => x"2e",
          3839 => x"74",
          3840 => x"0c",
          3841 => x"80",
          3842 => x"80",
          3843 => x"70",
          3844 => x"51",
          3845 => x"82",
          3846 => x"54",
          3847 => x"dc",
          3848 => x"0d",
          3849 => x"0d",
          3850 => x"05",
          3851 => x"33",
          3852 => x"54",
          3853 => x"84",
          3854 => x"bf",
          3855 => x"98",
          3856 => x"53",
          3857 => x"05",
          3858 => x"fa",
          3859 => x"dc",
          3860 => x"8c",
          3861 => x"a4",
          3862 => x"68",
          3863 => x"70",
          3864 => x"c6",
          3865 => x"dc",
          3866 => x"8c",
          3867 => x"38",
          3868 => x"05",
          3869 => x"2b",
          3870 => x"80",
          3871 => x"86",
          3872 => x"06",
          3873 => x"2e",
          3874 => x"74",
          3875 => x"38",
          3876 => x"09",
          3877 => x"38",
          3878 => x"f8",
          3879 => x"dc",
          3880 => x"39",
          3881 => x"33",
          3882 => x"73",
          3883 => x"77",
          3884 => x"81",
          3885 => x"73",
          3886 => x"38",
          3887 => x"bc",
          3888 => x"07",
          3889 => x"b4",
          3890 => x"2a",
          3891 => x"51",
          3892 => x"2e",
          3893 => x"62",
          3894 => x"e8",
          3895 => x"8c",
          3896 => x"82",
          3897 => x"52",
          3898 => x"51",
          3899 => x"62",
          3900 => x"8b",
          3901 => x"53",
          3902 => x"51",
          3903 => x"80",
          3904 => x"05",
          3905 => x"3f",
          3906 => x"0b",
          3907 => x"75",
          3908 => x"f1",
          3909 => x"11",
          3910 => x"80",
          3911 => x"97",
          3912 => x"51",
          3913 => x"82",
          3914 => x"55",
          3915 => x"08",
          3916 => x"b7",
          3917 => x"c4",
          3918 => x"05",
          3919 => x"2a",
          3920 => x"51",
          3921 => x"80",
          3922 => x"84",
          3923 => x"39",
          3924 => x"70",
          3925 => x"54",
          3926 => x"a9",
          3927 => x"06",
          3928 => x"2e",
          3929 => x"55",
          3930 => x"73",
          3931 => x"d6",
          3932 => x"8c",
          3933 => x"ff",
          3934 => x"0c",
          3935 => x"8c",
          3936 => x"f8",
          3937 => x"2a",
          3938 => x"51",
          3939 => x"2e",
          3940 => x"80",
          3941 => x"7a",
          3942 => x"a0",
          3943 => x"a4",
          3944 => x"53",
          3945 => x"e6",
          3946 => x"8c",
          3947 => x"8c",
          3948 => x"1b",
          3949 => x"05",
          3950 => x"d3",
          3951 => x"dc",
          3952 => x"dc",
          3953 => x"0c",
          3954 => x"56",
          3955 => x"84",
          3956 => x"90",
          3957 => x"0b",
          3958 => x"80",
          3959 => x"0c",
          3960 => x"1a",
          3961 => x"2a",
          3962 => x"51",
          3963 => x"2e",
          3964 => x"82",
          3965 => x"80",
          3966 => x"38",
          3967 => x"08",
          3968 => x"8a",
          3969 => x"89",
          3970 => x"59",
          3971 => x"76",
          3972 => x"d7",
          3973 => x"8c",
          3974 => x"82",
          3975 => x"81",
          3976 => x"82",
          3977 => x"dc",
          3978 => x"09",
          3979 => x"38",
          3980 => x"78",
          3981 => x"30",
          3982 => x"80",
          3983 => x"77",
          3984 => x"38",
          3985 => x"06",
          3986 => x"c3",
          3987 => x"1a",
          3988 => x"38",
          3989 => x"06",
          3990 => x"2e",
          3991 => x"52",
          3992 => x"a6",
          3993 => x"dc",
          3994 => x"82",
          3995 => x"75",
          3996 => x"8c",
          3997 => x"9c",
          3998 => x"39",
          3999 => x"74",
          4000 => x"8c",
          4001 => x"3d",
          4002 => x"3d",
          4003 => x"65",
          4004 => x"5d",
          4005 => x"0c",
          4006 => x"05",
          4007 => x"f9",
          4008 => x"8c",
          4009 => x"82",
          4010 => x"8a",
          4011 => x"33",
          4012 => x"2e",
          4013 => x"56",
          4014 => x"90",
          4015 => x"06",
          4016 => x"74",
          4017 => x"b6",
          4018 => x"82",
          4019 => x"34",
          4020 => x"aa",
          4021 => x"91",
          4022 => x"56",
          4023 => x"8c",
          4024 => x"1a",
          4025 => x"74",
          4026 => x"38",
          4027 => x"80",
          4028 => x"38",
          4029 => x"70",
          4030 => x"56",
          4031 => x"b2",
          4032 => x"11",
          4033 => x"77",
          4034 => x"5b",
          4035 => x"38",
          4036 => x"88",
          4037 => x"8f",
          4038 => x"08",
          4039 => x"d5",
          4040 => x"8c",
          4041 => x"81",
          4042 => x"9f",
          4043 => x"2e",
          4044 => x"74",
          4045 => x"98",
          4046 => x"7e",
          4047 => x"3f",
          4048 => x"08",
          4049 => x"83",
          4050 => x"dc",
          4051 => x"89",
          4052 => x"77",
          4053 => x"d6",
          4054 => x"7f",
          4055 => x"58",
          4056 => x"75",
          4057 => x"75",
          4058 => x"77",
          4059 => x"7c",
          4060 => x"33",
          4061 => x"3f",
          4062 => x"08",
          4063 => x"7e",
          4064 => x"56",
          4065 => x"2e",
          4066 => x"16",
          4067 => x"55",
          4068 => x"94",
          4069 => x"53",
          4070 => x"b0",
          4071 => x"31",
          4072 => x"05",
          4073 => x"3f",
          4074 => x"56",
          4075 => x"9c",
          4076 => x"19",
          4077 => x"06",
          4078 => x"31",
          4079 => x"76",
          4080 => x"7b",
          4081 => x"08",
          4082 => x"d1",
          4083 => x"8c",
          4084 => x"81",
          4085 => x"94",
          4086 => x"ff",
          4087 => x"05",
          4088 => x"cf",
          4089 => x"76",
          4090 => x"17",
          4091 => x"1e",
          4092 => x"18",
          4093 => x"5e",
          4094 => x"39",
          4095 => x"82",
          4096 => x"90",
          4097 => x"f2",
          4098 => x"63",
          4099 => x"40",
          4100 => x"7e",
          4101 => x"fc",
          4102 => x"51",
          4103 => x"82",
          4104 => x"55",
          4105 => x"08",
          4106 => x"18",
          4107 => x"80",
          4108 => x"74",
          4109 => x"39",
          4110 => x"70",
          4111 => x"81",
          4112 => x"56",
          4113 => x"80",
          4114 => x"38",
          4115 => x"0b",
          4116 => x"82",
          4117 => x"39",
          4118 => x"19",
          4119 => x"83",
          4120 => x"18",
          4121 => x"56",
          4122 => x"27",
          4123 => x"09",
          4124 => x"2e",
          4125 => x"94",
          4126 => x"83",
          4127 => x"56",
          4128 => x"38",
          4129 => x"22",
          4130 => x"89",
          4131 => x"55",
          4132 => x"75",
          4133 => x"18",
          4134 => x"9c",
          4135 => x"85",
          4136 => x"08",
          4137 => x"d7",
          4138 => x"8c",
          4139 => x"82",
          4140 => x"80",
          4141 => x"38",
          4142 => x"ff",
          4143 => x"ff",
          4144 => x"38",
          4145 => x"0c",
          4146 => x"85",
          4147 => x"19",
          4148 => x"b0",
          4149 => x"19",
          4150 => x"81",
          4151 => x"74",
          4152 => x"3f",
          4153 => x"08",
          4154 => x"98",
          4155 => x"7e",
          4156 => x"3f",
          4157 => x"08",
          4158 => x"d2",
          4159 => x"dc",
          4160 => x"89",
          4161 => x"78",
          4162 => x"d5",
          4163 => x"7f",
          4164 => x"58",
          4165 => x"75",
          4166 => x"75",
          4167 => x"78",
          4168 => x"7c",
          4169 => x"33",
          4170 => x"3f",
          4171 => x"08",
          4172 => x"7e",
          4173 => x"78",
          4174 => x"74",
          4175 => x"38",
          4176 => x"b0",
          4177 => x"31",
          4178 => x"05",
          4179 => x"51",
          4180 => x"7e",
          4181 => x"83",
          4182 => x"89",
          4183 => x"db",
          4184 => x"08",
          4185 => x"26",
          4186 => x"51",
          4187 => x"82",
          4188 => x"fd",
          4189 => x"77",
          4190 => x"55",
          4191 => x"0c",
          4192 => x"83",
          4193 => x"80",
          4194 => x"55",
          4195 => x"83",
          4196 => x"9c",
          4197 => x"7e",
          4198 => x"3f",
          4199 => x"08",
          4200 => x"75",
          4201 => x"94",
          4202 => x"ff",
          4203 => x"05",
          4204 => x"3f",
          4205 => x"0b",
          4206 => x"7b",
          4207 => x"08",
          4208 => x"76",
          4209 => x"08",
          4210 => x"1c",
          4211 => x"08",
          4212 => x"5c",
          4213 => x"83",
          4214 => x"74",
          4215 => x"fd",
          4216 => x"18",
          4217 => x"07",
          4218 => x"19",
          4219 => x"75",
          4220 => x"0c",
          4221 => x"04",
          4222 => x"7a",
          4223 => x"05",
          4224 => x"56",
          4225 => x"82",
          4226 => x"57",
          4227 => x"08",
          4228 => x"90",
          4229 => x"86",
          4230 => x"06",
          4231 => x"73",
          4232 => x"e9",
          4233 => x"08",
          4234 => x"cc",
          4235 => x"8c",
          4236 => x"82",
          4237 => x"80",
          4238 => x"16",
          4239 => x"33",
          4240 => x"55",
          4241 => x"34",
          4242 => x"53",
          4243 => x"08",
          4244 => x"3f",
          4245 => x"52",
          4246 => x"c9",
          4247 => x"88",
          4248 => x"96",
          4249 => x"f0",
          4250 => x"92",
          4251 => x"ca",
          4252 => x"81",
          4253 => x"34",
          4254 => x"df",
          4255 => x"dc",
          4256 => x"33",
          4257 => x"55",
          4258 => x"17",
          4259 => x"8c",
          4260 => x"3d",
          4261 => x"3d",
          4262 => x"52",
          4263 => x"3f",
          4264 => x"08",
          4265 => x"dc",
          4266 => x"86",
          4267 => x"52",
          4268 => x"bc",
          4269 => x"dc",
          4270 => x"8c",
          4271 => x"38",
          4272 => x"08",
          4273 => x"82",
          4274 => x"86",
          4275 => x"ff",
          4276 => x"3d",
          4277 => x"3f",
          4278 => x"0b",
          4279 => x"08",
          4280 => x"82",
          4281 => x"82",
          4282 => x"80",
          4283 => x"8c",
          4284 => x"3d",
          4285 => x"3d",
          4286 => x"93",
          4287 => x"52",
          4288 => x"e9",
          4289 => x"8c",
          4290 => x"82",
          4291 => x"80",
          4292 => x"58",
          4293 => x"3d",
          4294 => x"e0",
          4295 => x"8c",
          4296 => x"82",
          4297 => x"bc",
          4298 => x"c7",
          4299 => x"98",
          4300 => x"73",
          4301 => x"38",
          4302 => x"12",
          4303 => x"39",
          4304 => x"33",
          4305 => x"70",
          4306 => x"55",
          4307 => x"2e",
          4308 => x"7f",
          4309 => x"54",
          4310 => x"82",
          4311 => x"94",
          4312 => x"39",
          4313 => x"08",
          4314 => x"81",
          4315 => x"85",
          4316 => x"8c",
          4317 => x"3d",
          4318 => x"3d",
          4319 => x"5b",
          4320 => x"34",
          4321 => x"3d",
          4322 => x"52",
          4323 => x"e8",
          4324 => x"8c",
          4325 => x"82",
          4326 => x"82",
          4327 => x"43",
          4328 => x"11",
          4329 => x"58",
          4330 => x"80",
          4331 => x"38",
          4332 => x"3d",
          4333 => x"d5",
          4334 => x"8c",
          4335 => x"82",
          4336 => x"82",
          4337 => x"52",
          4338 => x"c8",
          4339 => x"dc",
          4340 => x"8c",
          4341 => x"c1",
          4342 => x"7b",
          4343 => x"3f",
          4344 => x"08",
          4345 => x"74",
          4346 => x"3f",
          4347 => x"08",
          4348 => x"dc",
          4349 => x"38",
          4350 => x"51",
          4351 => x"82",
          4352 => x"57",
          4353 => x"08",
          4354 => x"52",
          4355 => x"f2",
          4356 => x"8c",
          4357 => x"a6",
          4358 => x"74",
          4359 => x"3f",
          4360 => x"08",
          4361 => x"dc",
          4362 => x"cc",
          4363 => x"2e",
          4364 => x"86",
          4365 => x"81",
          4366 => x"81",
          4367 => x"3d",
          4368 => x"52",
          4369 => x"c9",
          4370 => x"3d",
          4371 => x"11",
          4372 => x"5a",
          4373 => x"2e",
          4374 => x"b9",
          4375 => x"16",
          4376 => x"33",
          4377 => x"73",
          4378 => x"16",
          4379 => x"26",
          4380 => x"75",
          4381 => x"38",
          4382 => x"05",
          4383 => x"6f",
          4384 => x"ff",
          4385 => x"55",
          4386 => x"74",
          4387 => x"38",
          4388 => x"11",
          4389 => x"74",
          4390 => x"39",
          4391 => x"09",
          4392 => x"38",
          4393 => x"11",
          4394 => x"74",
          4395 => x"82",
          4396 => x"70",
          4397 => x"fa",
          4398 => x"08",
          4399 => x"5c",
          4400 => x"73",
          4401 => x"38",
          4402 => x"1a",
          4403 => x"55",
          4404 => x"38",
          4405 => x"73",
          4406 => x"38",
          4407 => x"76",
          4408 => x"74",
          4409 => x"33",
          4410 => x"05",
          4411 => x"15",
          4412 => x"ba",
          4413 => x"05",
          4414 => x"ff",
          4415 => x"06",
          4416 => x"57",
          4417 => x"18",
          4418 => x"54",
          4419 => x"70",
          4420 => x"34",
          4421 => x"ee",
          4422 => x"34",
          4423 => x"dc",
          4424 => x"0d",
          4425 => x"0d",
          4426 => x"3d",
          4427 => x"71",
          4428 => x"ec",
          4429 => x"8c",
          4430 => x"82",
          4431 => x"82",
          4432 => x"15",
          4433 => x"82",
          4434 => x"15",
          4435 => x"76",
          4436 => x"90",
          4437 => x"81",
          4438 => x"06",
          4439 => x"72",
          4440 => x"56",
          4441 => x"54",
          4442 => x"17",
          4443 => x"78",
          4444 => x"38",
          4445 => x"22",
          4446 => x"59",
          4447 => x"78",
          4448 => x"76",
          4449 => x"51",
          4450 => x"3f",
          4451 => x"08",
          4452 => x"54",
          4453 => x"53",
          4454 => x"3f",
          4455 => x"08",
          4456 => x"38",
          4457 => x"75",
          4458 => x"18",
          4459 => x"31",
          4460 => x"57",
          4461 => x"b1",
          4462 => x"08",
          4463 => x"38",
          4464 => x"51",
          4465 => x"82",
          4466 => x"54",
          4467 => x"08",
          4468 => x"9a",
          4469 => x"dc",
          4470 => x"81",
          4471 => x"8c",
          4472 => x"16",
          4473 => x"16",
          4474 => x"2e",
          4475 => x"76",
          4476 => x"dc",
          4477 => x"31",
          4478 => x"18",
          4479 => x"90",
          4480 => x"81",
          4481 => x"06",
          4482 => x"56",
          4483 => x"9a",
          4484 => x"74",
          4485 => x"3f",
          4486 => x"08",
          4487 => x"dc",
          4488 => x"82",
          4489 => x"56",
          4490 => x"52",
          4491 => x"84",
          4492 => x"dc",
          4493 => x"ff",
          4494 => x"81",
          4495 => x"38",
          4496 => x"98",
          4497 => x"a6",
          4498 => x"16",
          4499 => x"39",
          4500 => x"16",
          4501 => x"75",
          4502 => x"53",
          4503 => x"aa",
          4504 => x"79",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"0b",
          4508 => x"82",
          4509 => x"39",
          4510 => x"16",
          4511 => x"bb",
          4512 => x"2a",
          4513 => x"08",
          4514 => x"15",
          4515 => x"15",
          4516 => x"90",
          4517 => x"16",
          4518 => x"33",
          4519 => x"53",
          4520 => x"34",
          4521 => x"06",
          4522 => x"2e",
          4523 => x"9c",
          4524 => x"85",
          4525 => x"16",
          4526 => x"72",
          4527 => x"0c",
          4528 => x"04",
          4529 => x"79",
          4530 => x"75",
          4531 => x"8a",
          4532 => x"89",
          4533 => x"52",
          4534 => x"05",
          4535 => x"3f",
          4536 => x"08",
          4537 => x"dc",
          4538 => x"38",
          4539 => x"7a",
          4540 => x"d8",
          4541 => x"8c",
          4542 => x"82",
          4543 => x"80",
          4544 => x"16",
          4545 => x"2b",
          4546 => x"74",
          4547 => x"86",
          4548 => x"84",
          4549 => x"06",
          4550 => x"73",
          4551 => x"38",
          4552 => x"52",
          4553 => x"da",
          4554 => x"dc",
          4555 => x"0c",
          4556 => x"14",
          4557 => x"23",
          4558 => x"51",
          4559 => x"82",
          4560 => x"55",
          4561 => x"09",
          4562 => x"38",
          4563 => x"39",
          4564 => x"84",
          4565 => x"0c",
          4566 => x"82",
          4567 => x"89",
          4568 => x"fc",
          4569 => x"87",
          4570 => x"53",
          4571 => x"e7",
          4572 => x"8c",
          4573 => x"38",
          4574 => x"08",
          4575 => x"3d",
          4576 => x"3d",
          4577 => x"89",
          4578 => x"54",
          4579 => x"54",
          4580 => x"82",
          4581 => x"53",
          4582 => x"08",
          4583 => x"74",
          4584 => x"8c",
          4585 => x"73",
          4586 => x"3f",
          4587 => x"08",
          4588 => x"39",
          4589 => x"08",
          4590 => x"d3",
          4591 => x"8c",
          4592 => x"82",
          4593 => x"84",
          4594 => x"06",
          4595 => x"53",
          4596 => x"8c",
          4597 => x"38",
          4598 => x"51",
          4599 => x"72",
          4600 => x"cf",
          4601 => x"8c",
          4602 => x"32",
          4603 => x"72",
          4604 => x"70",
          4605 => x"08",
          4606 => x"54",
          4607 => x"8c",
          4608 => x"3d",
          4609 => x"3d",
          4610 => x"80",
          4611 => x"70",
          4612 => x"52",
          4613 => x"3f",
          4614 => x"08",
          4615 => x"dc",
          4616 => x"64",
          4617 => x"d6",
          4618 => x"8c",
          4619 => x"82",
          4620 => x"a0",
          4621 => x"cb",
          4622 => x"98",
          4623 => x"73",
          4624 => x"38",
          4625 => x"39",
          4626 => x"88",
          4627 => x"75",
          4628 => x"3f",
          4629 => x"dc",
          4630 => x"0d",
          4631 => x"0d",
          4632 => x"5c",
          4633 => x"3d",
          4634 => x"93",
          4635 => x"d6",
          4636 => x"dc",
          4637 => x"8c",
          4638 => x"80",
          4639 => x"0c",
          4640 => x"11",
          4641 => x"90",
          4642 => x"56",
          4643 => x"74",
          4644 => x"75",
          4645 => x"e4",
          4646 => x"81",
          4647 => x"5b",
          4648 => x"82",
          4649 => x"75",
          4650 => x"73",
          4651 => x"81",
          4652 => x"82",
          4653 => x"76",
          4654 => x"f0",
          4655 => x"f4",
          4656 => x"dc",
          4657 => x"d1",
          4658 => x"dc",
          4659 => x"ce",
          4660 => x"dc",
          4661 => x"82",
          4662 => x"07",
          4663 => x"05",
          4664 => x"53",
          4665 => x"98",
          4666 => x"26",
          4667 => x"f9",
          4668 => x"08",
          4669 => x"08",
          4670 => x"98",
          4671 => x"81",
          4672 => x"58",
          4673 => x"3f",
          4674 => x"08",
          4675 => x"dc",
          4676 => x"38",
          4677 => x"77",
          4678 => x"5d",
          4679 => x"74",
          4680 => x"81",
          4681 => x"b4",
          4682 => x"bb",
          4683 => x"8c",
          4684 => x"ff",
          4685 => x"30",
          4686 => x"1b",
          4687 => x"5b",
          4688 => x"39",
          4689 => x"ff",
          4690 => x"82",
          4691 => x"f0",
          4692 => x"30",
          4693 => x"1b",
          4694 => x"5b",
          4695 => x"83",
          4696 => x"58",
          4697 => x"92",
          4698 => x"0c",
          4699 => x"12",
          4700 => x"33",
          4701 => x"54",
          4702 => x"34",
          4703 => x"dc",
          4704 => x"0d",
          4705 => x"0d",
          4706 => x"fc",
          4707 => x"52",
          4708 => x"3f",
          4709 => x"08",
          4710 => x"dc",
          4711 => x"38",
          4712 => x"56",
          4713 => x"38",
          4714 => x"70",
          4715 => x"81",
          4716 => x"55",
          4717 => x"80",
          4718 => x"38",
          4719 => x"54",
          4720 => x"08",
          4721 => x"38",
          4722 => x"82",
          4723 => x"53",
          4724 => x"52",
          4725 => x"8c",
          4726 => x"dc",
          4727 => x"19",
          4728 => x"c9",
          4729 => x"08",
          4730 => x"ff",
          4731 => x"82",
          4732 => x"ff",
          4733 => x"06",
          4734 => x"56",
          4735 => x"08",
          4736 => x"81",
          4737 => x"82",
          4738 => x"75",
          4739 => x"54",
          4740 => x"08",
          4741 => x"27",
          4742 => x"17",
          4743 => x"8c",
          4744 => x"76",
          4745 => x"3f",
          4746 => x"08",
          4747 => x"08",
          4748 => x"90",
          4749 => x"c0",
          4750 => x"90",
          4751 => x"80",
          4752 => x"75",
          4753 => x"75",
          4754 => x"8c",
          4755 => x"3d",
          4756 => x"3d",
          4757 => x"a0",
          4758 => x"05",
          4759 => x"51",
          4760 => x"82",
          4761 => x"55",
          4762 => x"08",
          4763 => x"78",
          4764 => x"08",
          4765 => x"70",
          4766 => x"ae",
          4767 => x"dc",
          4768 => x"8c",
          4769 => x"db",
          4770 => x"fb",
          4771 => x"85",
          4772 => x"06",
          4773 => x"86",
          4774 => x"c7",
          4775 => x"2b",
          4776 => x"24",
          4777 => x"02",
          4778 => x"33",
          4779 => x"58",
          4780 => x"76",
          4781 => x"6b",
          4782 => x"cc",
          4783 => x"8c",
          4784 => x"84",
          4785 => x"06",
          4786 => x"73",
          4787 => x"d4",
          4788 => x"82",
          4789 => x"94",
          4790 => x"81",
          4791 => x"5a",
          4792 => x"08",
          4793 => x"8a",
          4794 => x"54",
          4795 => x"82",
          4796 => x"55",
          4797 => x"08",
          4798 => x"82",
          4799 => x"52",
          4800 => x"e5",
          4801 => x"dc",
          4802 => x"8c",
          4803 => x"38",
          4804 => x"cf",
          4805 => x"dc",
          4806 => x"88",
          4807 => x"dc",
          4808 => x"38",
          4809 => x"c2",
          4810 => x"dc",
          4811 => x"dc",
          4812 => x"82",
          4813 => x"07",
          4814 => x"55",
          4815 => x"2e",
          4816 => x"80",
          4817 => x"80",
          4818 => x"77",
          4819 => x"3f",
          4820 => x"08",
          4821 => x"38",
          4822 => x"ba",
          4823 => x"8c",
          4824 => x"74",
          4825 => x"0c",
          4826 => x"04",
          4827 => x"82",
          4828 => x"c0",
          4829 => x"3d",
          4830 => x"3f",
          4831 => x"08",
          4832 => x"dc",
          4833 => x"38",
          4834 => x"52",
          4835 => x"52",
          4836 => x"3f",
          4837 => x"08",
          4838 => x"dc",
          4839 => x"88",
          4840 => x"39",
          4841 => x"08",
          4842 => x"81",
          4843 => x"38",
          4844 => x"05",
          4845 => x"2a",
          4846 => x"55",
          4847 => x"81",
          4848 => x"5a",
          4849 => x"3d",
          4850 => x"c1",
          4851 => x"8c",
          4852 => x"55",
          4853 => x"dc",
          4854 => x"87",
          4855 => x"dc",
          4856 => x"09",
          4857 => x"38",
          4858 => x"8c",
          4859 => x"2e",
          4860 => x"86",
          4861 => x"81",
          4862 => x"81",
          4863 => x"8c",
          4864 => x"78",
          4865 => x"3f",
          4866 => x"08",
          4867 => x"dc",
          4868 => x"38",
          4869 => x"52",
          4870 => x"ff",
          4871 => x"78",
          4872 => x"b4",
          4873 => x"54",
          4874 => x"15",
          4875 => x"b2",
          4876 => x"ca",
          4877 => x"b6",
          4878 => x"53",
          4879 => x"53",
          4880 => x"3f",
          4881 => x"b4",
          4882 => x"d4",
          4883 => x"b6",
          4884 => x"54",
          4885 => x"d5",
          4886 => x"53",
          4887 => x"11",
          4888 => x"d7",
          4889 => x"81",
          4890 => x"34",
          4891 => x"a4",
          4892 => x"dc",
          4893 => x"8c",
          4894 => x"38",
          4895 => x"0a",
          4896 => x"05",
          4897 => x"d0",
          4898 => x"64",
          4899 => x"c9",
          4900 => x"54",
          4901 => x"15",
          4902 => x"81",
          4903 => x"34",
          4904 => x"b8",
          4905 => x"8c",
          4906 => x"8b",
          4907 => x"75",
          4908 => x"ff",
          4909 => x"73",
          4910 => x"0c",
          4911 => x"04",
          4912 => x"a9",
          4913 => x"51",
          4914 => x"82",
          4915 => x"ff",
          4916 => x"a9",
          4917 => x"ee",
          4918 => x"dc",
          4919 => x"8c",
          4920 => x"d3",
          4921 => x"a9",
          4922 => x"9d",
          4923 => x"58",
          4924 => x"82",
          4925 => x"55",
          4926 => x"08",
          4927 => x"02",
          4928 => x"33",
          4929 => x"54",
          4930 => x"82",
          4931 => x"53",
          4932 => x"52",
          4933 => x"88",
          4934 => x"b4",
          4935 => x"53",
          4936 => x"3d",
          4937 => x"ff",
          4938 => x"aa",
          4939 => x"73",
          4940 => x"3f",
          4941 => x"08",
          4942 => x"dc",
          4943 => x"63",
          4944 => x"81",
          4945 => x"65",
          4946 => x"2e",
          4947 => x"55",
          4948 => x"82",
          4949 => x"84",
          4950 => x"06",
          4951 => x"73",
          4952 => x"3f",
          4953 => x"08",
          4954 => x"dc",
          4955 => x"38",
          4956 => x"53",
          4957 => x"95",
          4958 => x"16",
          4959 => x"87",
          4960 => x"05",
          4961 => x"34",
          4962 => x"70",
          4963 => x"81",
          4964 => x"55",
          4965 => x"74",
          4966 => x"73",
          4967 => x"78",
          4968 => x"83",
          4969 => x"16",
          4970 => x"2a",
          4971 => x"51",
          4972 => x"80",
          4973 => x"38",
          4974 => x"80",
          4975 => x"52",
          4976 => x"be",
          4977 => x"dc",
          4978 => x"51",
          4979 => x"3f",
          4980 => x"8c",
          4981 => x"2e",
          4982 => x"82",
          4983 => x"52",
          4984 => x"b5",
          4985 => x"8c",
          4986 => x"80",
          4987 => x"58",
          4988 => x"dc",
          4989 => x"38",
          4990 => x"54",
          4991 => x"09",
          4992 => x"38",
          4993 => x"52",
          4994 => x"af",
          4995 => x"81",
          4996 => x"34",
          4997 => x"8c",
          4998 => x"38",
          4999 => x"ca",
          5000 => x"dc",
          5001 => x"8c",
          5002 => x"38",
          5003 => x"b5",
          5004 => x"8c",
          5005 => x"74",
          5006 => x"0c",
          5007 => x"04",
          5008 => x"02",
          5009 => x"33",
          5010 => x"80",
          5011 => x"57",
          5012 => x"95",
          5013 => x"52",
          5014 => x"d2",
          5015 => x"8c",
          5016 => x"82",
          5017 => x"80",
          5018 => x"5a",
          5019 => x"3d",
          5020 => x"c9",
          5021 => x"8c",
          5022 => x"82",
          5023 => x"b8",
          5024 => x"cf",
          5025 => x"a0",
          5026 => x"55",
          5027 => x"75",
          5028 => x"71",
          5029 => x"33",
          5030 => x"74",
          5031 => x"57",
          5032 => x"8b",
          5033 => x"54",
          5034 => x"15",
          5035 => x"ff",
          5036 => x"82",
          5037 => x"55",
          5038 => x"dc",
          5039 => x"0d",
          5040 => x"0d",
          5041 => x"53",
          5042 => x"05",
          5043 => x"51",
          5044 => x"82",
          5045 => x"55",
          5046 => x"08",
          5047 => x"76",
          5048 => x"93",
          5049 => x"51",
          5050 => x"82",
          5051 => x"55",
          5052 => x"08",
          5053 => x"80",
          5054 => x"81",
          5055 => x"86",
          5056 => x"38",
          5057 => x"86",
          5058 => x"90",
          5059 => x"54",
          5060 => x"ff",
          5061 => x"76",
          5062 => x"83",
          5063 => x"51",
          5064 => x"3f",
          5065 => x"08",
          5066 => x"8c",
          5067 => x"3d",
          5068 => x"3d",
          5069 => x"5c",
          5070 => x"98",
          5071 => x"52",
          5072 => x"d1",
          5073 => x"8c",
          5074 => x"8c",
          5075 => x"70",
          5076 => x"08",
          5077 => x"51",
          5078 => x"80",
          5079 => x"38",
          5080 => x"06",
          5081 => x"80",
          5082 => x"38",
          5083 => x"5f",
          5084 => x"3d",
          5085 => x"ff",
          5086 => x"82",
          5087 => x"57",
          5088 => x"08",
          5089 => x"74",
          5090 => x"c3",
          5091 => x"8c",
          5092 => x"82",
          5093 => x"bf",
          5094 => x"dc",
          5095 => x"dc",
          5096 => x"59",
          5097 => x"81",
          5098 => x"56",
          5099 => x"33",
          5100 => x"16",
          5101 => x"27",
          5102 => x"56",
          5103 => x"80",
          5104 => x"80",
          5105 => x"ff",
          5106 => x"70",
          5107 => x"56",
          5108 => x"e8",
          5109 => x"76",
          5110 => x"81",
          5111 => x"80",
          5112 => x"57",
          5113 => x"78",
          5114 => x"51",
          5115 => x"2e",
          5116 => x"73",
          5117 => x"38",
          5118 => x"08",
          5119 => x"b1",
          5120 => x"8c",
          5121 => x"82",
          5122 => x"a7",
          5123 => x"33",
          5124 => x"c3",
          5125 => x"2e",
          5126 => x"e4",
          5127 => x"2e",
          5128 => x"56",
          5129 => x"05",
          5130 => x"e3",
          5131 => x"dc",
          5132 => x"76",
          5133 => x"0c",
          5134 => x"04",
          5135 => x"82",
          5136 => x"ff",
          5137 => x"9d",
          5138 => x"fa",
          5139 => x"dc",
          5140 => x"dc",
          5141 => x"82",
          5142 => x"83",
          5143 => x"53",
          5144 => x"3d",
          5145 => x"ff",
          5146 => x"73",
          5147 => x"70",
          5148 => x"52",
          5149 => x"9f",
          5150 => x"bc",
          5151 => x"74",
          5152 => x"6d",
          5153 => x"70",
          5154 => x"af",
          5155 => x"8c",
          5156 => x"2e",
          5157 => x"70",
          5158 => x"57",
          5159 => x"fd",
          5160 => x"dc",
          5161 => x"8d",
          5162 => x"2b",
          5163 => x"81",
          5164 => x"86",
          5165 => x"dc",
          5166 => x"9f",
          5167 => x"ff",
          5168 => x"54",
          5169 => x"8a",
          5170 => x"70",
          5171 => x"06",
          5172 => x"ff",
          5173 => x"38",
          5174 => x"15",
          5175 => x"80",
          5176 => x"74",
          5177 => x"ec",
          5178 => x"89",
          5179 => x"dc",
          5180 => x"81",
          5181 => x"88",
          5182 => x"26",
          5183 => x"39",
          5184 => x"86",
          5185 => x"81",
          5186 => x"ff",
          5187 => x"38",
          5188 => x"54",
          5189 => x"81",
          5190 => x"81",
          5191 => x"78",
          5192 => x"5a",
          5193 => x"6d",
          5194 => x"81",
          5195 => x"57",
          5196 => x"9f",
          5197 => x"38",
          5198 => x"54",
          5199 => x"81",
          5200 => x"b1",
          5201 => x"2e",
          5202 => x"a7",
          5203 => x"15",
          5204 => x"54",
          5205 => x"09",
          5206 => x"38",
          5207 => x"76",
          5208 => x"41",
          5209 => x"52",
          5210 => x"52",
          5211 => x"b3",
          5212 => x"dc",
          5213 => x"8c",
          5214 => x"f7",
          5215 => x"74",
          5216 => x"e5",
          5217 => x"dc",
          5218 => x"8c",
          5219 => x"38",
          5220 => x"38",
          5221 => x"74",
          5222 => x"39",
          5223 => x"08",
          5224 => x"81",
          5225 => x"38",
          5226 => x"74",
          5227 => x"38",
          5228 => x"51",
          5229 => x"3f",
          5230 => x"08",
          5231 => x"dc",
          5232 => x"a0",
          5233 => x"dc",
          5234 => x"51",
          5235 => x"3f",
          5236 => x"0b",
          5237 => x"8b",
          5238 => x"67",
          5239 => x"a7",
          5240 => x"81",
          5241 => x"34",
          5242 => x"ad",
          5243 => x"8c",
          5244 => x"73",
          5245 => x"8c",
          5246 => x"3d",
          5247 => x"3d",
          5248 => x"02",
          5249 => x"cb",
          5250 => x"3d",
          5251 => x"72",
          5252 => x"5a",
          5253 => x"82",
          5254 => x"58",
          5255 => x"08",
          5256 => x"91",
          5257 => x"77",
          5258 => x"7c",
          5259 => x"38",
          5260 => x"59",
          5261 => x"90",
          5262 => x"81",
          5263 => x"06",
          5264 => x"73",
          5265 => x"54",
          5266 => x"82",
          5267 => x"39",
          5268 => x"8b",
          5269 => x"11",
          5270 => x"2b",
          5271 => x"54",
          5272 => x"fe",
          5273 => x"ff",
          5274 => x"70",
          5275 => x"07",
          5276 => x"8c",
          5277 => x"8c",
          5278 => x"40",
          5279 => x"55",
          5280 => x"88",
          5281 => x"08",
          5282 => x"38",
          5283 => x"77",
          5284 => x"56",
          5285 => x"51",
          5286 => x"3f",
          5287 => x"55",
          5288 => x"08",
          5289 => x"38",
          5290 => x"8c",
          5291 => x"2e",
          5292 => x"82",
          5293 => x"ff",
          5294 => x"38",
          5295 => x"08",
          5296 => x"16",
          5297 => x"2e",
          5298 => x"87",
          5299 => x"74",
          5300 => x"74",
          5301 => x"81",
          5302 => x"38",
          5303 => x"ff",
          5304 => x"2e",
          5305 => x"7b",
          5306 => x"80",
          5307 => x"81",
          5308 => x"81",
          5309 => x"06",
          5310 => x"56",
          5311 => x"52",
          5312 => x"af",
          5313 => x"8c",
          5314 => x"82",
          5315 => x"80",
          5316 => x"81",
          5317 => x"56",
          5318 => x"d3",
          5319 => x"ff",
          5320 => x"7c",
          5321 => x"55",
          5322 => x"b3",
          5323 => x"1b",
          5324 => x"1b",
          5325 => x"33",
          5326 => x"54",
          5327 => x"34",
          5328 => x"fe",
          5329 => x"08",
          5330 => x"74",
          5331 => x"75",
          5332 => x"16",
          5333 => x"33",
          5334 => x"73",
          5335 => x"77",
          5336 => x"8c",
          5337 => x"3d",
          5338 => x"3d",
          5339 => x"02",
          5340 => x"eb",
          5341 => x"3d",
          5342 => x"59",
          5343 => x"8b",
          5344 => x"82",
          5345 => x"24",
          5346 => x"82",
          5347 => x"84",
          5348 => x"8c",
          5349 => x"51",
          5350 => x"2e",
          5351 => x"75",
          5352 => x"dc",
          5353 => x"06",
          5354 => x"7e",
          5355 => x"d0",
          5356 => x"dc",
          5357 => x"06",
          5358 => x"56",
          5359 => x"74",
          5360 => x"76",
          5361 => x"81",
          5362 => x"8a",
          5363 => x"b2",
          5364 => x"fc",
          5365 => x"52",
          5366 => x"a4",
          5367 => x"8c",
          5368 => x"38",
          5369 => x"80",
          5370 => x"74",
          5371 => x"26",
          5372 => x"15",
          5373 => x"74",
          5374 => x"38",
          5375 => x"80",
          5376 => x"84",
          5377 => x"92",
          5378 => x"80",
          5379 => x"38",
          5380 => x"06",
          5381 => x"2e",
          5382 => x"56",
          5383 => x"78",
          5384 => x"89",
          5385 => x"2b",
          5386 => x"43",
          5387 => x"38",
          5388 => x"30",
          5389 => x"77",
          5390 => x"91",
          5391 => x"c2",
          5392 => x"f8",
          5393 => x"52",
          5394 => x"a4",
          5395 => x"56",
          5396 => x"08",
          5397 => x"77",
          5398 => x"77",
          5399 => x"dc",
          5400 => x"45",
          5401 => x"bf",
          5402 => x"8e",
          5403 => x"26",
          5404 => x"74",
          5405 => x"48",
          5406 => x"75",
          5407 => x"38",
          5408 => x"81",
          5409 => x"fa",
          5410 => x"2a",
          5411 => x"56",
          5412 => x"2e",
          5413 => x"87",
          5414 => x"82",
          5415 => x"38",
          5416 => x"55",
          5417 => x"83",
          5418 => x"81",
          5419 => x"56",
          5420 => x"80",
          5421 => x"38",
          5422 => x"83",
          5423 => x"06",
          5424 => x"78",
          5425 => x"91",
          5426 => x"0b",
          5427 => x"22",
          5428 => x"80",
          5429 => x"74",
          5430 => x"38",
          5431 => x"56",
          5432 => x"17",
          5433 => x"57",
          5434 => x"2e",
          5435 => x"75",
          5436 => x"79",
          5437 => x"fe",
          5438 => x"82",
          5439 => x"84",
          5440 => x"05",
          5441 => x"5e",
          5442 => x"80",
          5443 => x"dc",
          5444 => x"8a",
          5445 => x"fd",
          5446 => x"75",
          5447 => x"38",
          5448 => x"78",
          5449 => x"8c",
          5450 => x"0b",
          5451 => x"22",
          5452 => x"80",
          5453 => x"74",
          5454 => x"38",
          5455 => x"56",
          5456 => x"17",
          5457 => x"57",
          5458 => x"2e",
          5459 => x"75",
          5460 => x"79",
          5461 => x"fe",
          5462 => x"82",
          5463 => x"10",
          5464 => x"82",
          5465 => x"9f",
          5466 => x"38",
          5467 => x"8c",
          5468 => x"82",
          5469 => x"05",
          5470 => x"2a",
          5471 => x"56",
          5472 => x"17",
          5473 => x"81",
          5474 => x"60",
          5475 => x"65",
          5476 => x"12",
          5477 => x"30",
          5478 => x"74",
          5479 => x"59",
          5480 => x"7d",
          5481 => x"81",
          5482 => x"76",
          5483 => x"41",
          5484 => x"76",
          5485 => x"90",
          5486 => x"62",
          5487 => x"51",
          5488 => x"26",
          5489 => x"75",
          5490 => x"31",
          5491 => x"65",
          5492 => x"fe",
          5493 => x"82",
          5494 => x"58",
          5495 => x"09",
          5496 => x"38",
          5497 => x"08",
          5498 => x"26",
          5499 => x"78",
          5500 => x"79",
          5501 => x"78",
          5502 => x"86",
          5503 => x"82",
          5504 => x"06",
          5505 => x"83",
          5506 => x"82",
          5507 => x"27",
          5508 => x"8f",
          5509 => x"55",
          5510 => x"26",
          5511 => x"59",
          5512 => x"62",
          5513 => x"74",
          5514 => x"38",
          5515 => x"88",
          5516 => x"dc",
          5517 => x"26",
          5518 => x"86",
          5519 => x"1a",
          5520 => x"79",
          5521 => x"38",
          5522 => x"80",
          5523 => x"2e",
          5524 => x"83",
          5525 => x"9f",
          5526 => x"8b",
          5527 => x"06",
          5528 => x"74",
          5529 => x"84",
          5530 => x"52",
          5531 => x"a2",
          5532 => x"53",
          5533 => x"52",
          5534 => x"a2",
          5535 => x"80",
          5536 => x"51",
          5537 => x"3f",
          5538 => x"34",
          5539 => x"ff",
          5540 => x"1b",
          5541 => x"a2",
          5542 => x"90",
          5543 => x"83",
          5544 => x"70",
          5545 => x"80",
          5546 => x"55",
          5547 => x"ff",
          5548 => x"66",
          5549 => x"ff",
          5550 => x"38",
          5551 => x"ff",
          5552 => x"1b",
          5553 => x"f2",
          5554 => x"74",
          5555 => x"51",
          5556 => x"3f",
          5557 => x"1c",
          5558 => x"98",
          5559 => x"a0",
          5560 => x"ff",
          5561 => x"51",
          5562 => x"3f",
          5563 => x"1b",
          5564 => x"e4",
          5565 => x"2e",
          5566 => x"80",
          5567 => x"88",
          5568 => x"80",
          5569 => x"ff",
          5570 => x"7c",
          5571 => x"51",
          5572 => x"3f",
          5573 => x"1b",
          5574 => x"bc",
          5575 => x"b0",
          5576 => x"a0",
          5577 => x"52",
          5578 => x"ff",
          5579 => x"ff",
          5580 => x"c0",
          5581 => x"0b",
          5582 => x"34",
          5583 => x"fa",
          5584 => x"c7",
          5585 => x"39",
          5586 => x"0a",
          5587 => x"51",
          5588 => x"3f",
          5589 => x"ff",
          5590 => x"1b",
          5591 => x"da",
          5592 => x"0b",
          5593 => x"a9",
          5594 => x"34",
          5595 => x"fa",
          5596 => x"1b",
          5597 => x"8f",
          5598 => x"d5",
          5599 => x"1b",
          5600 => x"ff",
          5601 => x"81",
          5602 => x"7a",
          5603 => x"ff",
          5604 => x"81",
          5605 => x"dc",
          5606 => x"38",
          5607 => x"09",
          5608 => x"ee",
          5609 => x"60",
          5610 => x"7a",
          5611 => x"ff",
          5612 => x"84",
          5613 => x"52",
          5614 => x"9f",
          5615 => x"8b",
          5616 => x"52",
          5617 => x"9f",
          5618 => x"8a",
          5619 => x"52",
          5620 => x"51",
          5621 => x"3f",
          5622 => x"83",
          5623 => x"ff",
          5624 => x"82",
          5625 => x"1b",
          5626 => x"ec",
          5627 => x"d5",
          5628 => x"ff",
          5629 => x"75",
          5630 => x"05",
          5631 => x"7e",
          5632 => x"e5",
          5633 => x"60",
          5634 => x"52",
          5635 => x"9a",
          5636 => x"53",
          5637 => x"51",
          5638 => x"3f",
          5639 => x"58",
          5640 => x"09",
          5641 => x"38",
          5642 => x"51",
          5643 => x"3f",
          5644 => x"1b",
          5645 => x"a0",
          5646 => x"52",
          5647 => x"91",
          5648 => x"ff",
          5649 => x"81",
          5650 => x"f8",
          5651 => x"7a",
          5652 => x"84",
          5653 => x"61",
          5654 => x"26",
          5655 => x"57",
          5656 => x"53",
          5657 => x"51",
          5658 => x"3f",
          5659 => x"08",
          5660 => x"84",
          5661 => x"8c",
          5662 => x"7a",
          5663 => x"aa",
          5664 => x"75",
          5665 => x"56",
          5666 => x"81",
          5667 => x"80",
          5668 => x"38",
          5669 => x"83",
          5670 => x"63",
          5671 => x"74",
          5672 => x"38",
          5673 => x"54",
          5674 => x"52",
          5675 => x"99",
          5676 => x"8c",
          5677 => x"c1",
          5678 => x"75",
          5679 => x"56",
          5680 => x"8c",
          5681 => x"2e",
          5682 => x"56",
          5683 => x"ff",
          5684 => x"84",
          5685 => x"2e",
          5686 => x"56",
          5687 => x"58",
          5688 => x"38",
          5689 => x"77",
          5690 => x"ff",
          5691 => x"82",
          5692 => x"78",
          5693 => x"c2",
          5694 => x"1b",
          5695 => x"34",
          5696 => x"16",
          5697 => x"82",
          5698 => x"83",
          5699 => x"84",
          5700 => x"67",
          5701 => x"fd",
          5702 => x"51",
          5703 => x"3f",
          5704 => x"16",
          5705 => x"dc",
          5706 => x"bf",
          5707 => x"86",
          5708 => x"8c",
          5709 => x"16",
          5710 => x"83",
          5711 => x"ff",
          5712 => x"66",
          5713 => x"1b",
          5714 => x"8c",
          5715 => x"77",
          5716 => x"7e",
          5717 => x"91",
          5718 => x"82",
          5719 => x"a2",
          5720 => x"80",
          5721 => x"ff",
          5722 => x"81",
          5723 => x"dc",
          5724 => x"89",
          5725 => x"8a",
          5726 => x"86",
          5727 => x"dc",
          5728 => x"82",
          5729 => x"99",
          5730 => x"f5",
          5731 => x"60",
          5732 => x"79",
          5733 => x"5a",
          5734 => x"78",
          5735 => x"8d",
          5736 => x"55",
          5737 => x"fc",
          5738 => x"51",
          5739 => x"7a",
          5740 => x"81",
          5741 => x"8c",
          5742 => x"74",
          5743 => x"38",
          5744 => x"81",
          5745 => x"81",
          5746 => x"8a",
          5747 => x"06",
          5748 => x"76",
          5749 => x"76",
          5750 => x"55",
          5751 => x"dc",
          5752 => x"0d",
          5753 => x"0d",
          5754 => x"05",
          5755 => x"59",
          5756 => x"2e",
          5757 => x"87",
          5758 => x"76",
          5759 => x"84",
          5760 => x"80",
          5761 => x"38",
          5762 => x"77",
          5763 => x"56",
          5764 => x"34",
          5765 => x"bb",
          5766 => x"38",
          5767 => x"05",
          5768 => x"8c",
          5769 => x"08",
          5770 => x"3f",
          5771 => x"70",
          5772 => x"07",
          5773 => x"30",
          5774 => x"56",
          5775 => x"0c",
          5776 => x"18",
          5777 => x"0d",
          5778 => x"0d",
          5779 => x"08",
          5780 => x"75",
          5781 => x"89",
          5782 => x"54",
          5783 => x"16",
          5784 => x"51",
          5785 => x"82",
          5786 => x"91",
          5787 => x"08",
          5788 => x"81",
          5789 => x"88",
          5790 => x"83",
          5791 => x"74",
          5792 => x"0c",
          5793 => x"04",
          5794 => x"75",
          5795 => x"53",
          5796 => x"51",
          5797 => x"3f",
          5798 => x"85",
          5799 => x"ea",
          5800 => x"80",
          5801 => x"6a",
          5802 => x"70",
          5803 => x"d8",
          5804 => x"72",
          5805 => x"3f",
          5806 => x"8d",
          5807 => x"0d",
          5808 => x"0d",
          5809 => x"70",
          5810 => x"74",
          5811 => x"e1",
          5812 => x"77",
          5813 => x"85",
          5814 => x"80",
          5815 => x"33",
          5816 => x"2e",
          5817 => x"86",
          5818 => x"55",
          5819 => x"57",
          5820 => x"82",
          5821 => x"70",
          5822 => x"fe",
          5823 => x"82",
          5824 => x"82",
          5825 => x"54",
          5826 => x"08",
          5827 => x"db",
          5828 => x"8c",
          5829 => x"38",
          5830 => x"54",
          5831 => x"ff",
          5832 => x"17",
          5833 => x"06",
          5834 => x"77",
          5835 => x"ff",
          5836 => x"8c",
          5837 => x"3d",
          5838 => x"3d",
          5839 => x"71",
          5840 => x"8e",
          5841 => x"29",
          5842 => x"05",
          5843 => x"04",
          5844 => x"51",
          5845 => x"81",
          5846 => x"80",
          5847 => x"fd",
          5848 => x"f2",
          5849 => x"fc",
          5850 => x"39",
          5851 => x"51",
          5852 => x"81",
          5853 => x"80",
          5854 => x"fe",
          5855 => x"d6",
          5856 => x"c0",
          5857 => x"39",
          5858 => x"51",
          5859 => x"81",
          5860 => x"80",
          5861 => x"ff",
          5862 => x"39",
          5863 => x"51",
          5864 => x"ff",
          5865 => x"39",
          5866 => x"51",
          5867 => x"ff",
          5868 => x"39",
          5869 => x"51",
          5870 => x"80",
          5871 => x"39",
          5872 => x"51",
          5873 => x"80",
          5874 => x"39",
          5875 => x"51",
          5876 => x"81",
          5877 => x"f2",
          5878 => x"3d",
          5879 => x"3d",
          5880 => x"56",
          5881 => x"e7",
          5882 => x"74",
          5883 => x"e8",
          5884 => x"39",
          5885 => x"74",
          5886 => x"df",
          5887 => x"dc",
          5888 => x"51",
          5889 => x"3f",
          5890 => x"08",
          5891 => x"75",
          5892 => x"90",
          5893 => x"d3",
          5894 => x"0d",
          5895 => x"0d",
          5896 => x"05",
          5897 => x"33",
          5898 => x"68",
          5899 => x"7a",
          5900 => x"51",
          5901 => x"78",
          5902 => x"ff",
          5903 => x"81",
          5904 => x"07",
          5905 => x"06",
          5906 => x"56",
          5907 => x"38",
          5908 => x"52",
          5909 => x"52",
          5910 => x"c9",
          5911 => x"dc",
          5912 => x"8c",
          5913 => x"38",
          5914 => x"08",
          5915 => x"88",
          5916 => x"dc",
          5917 => x"3d",
          5918 => x"84",
          5919 => x"52",
          5920 => x"86",
          5921 => x"dc",
          5922 => x"8c",
          5923 => x"38",
          5924 => x"80",
          5925 => x"74",
          5926 => x"59",
          5927 => x"96",
          5928 => x"51",
          5929 => x"76",
          5930 => x"07",
          5931 => x"30",
          5932 => x"72",
          5933 => x"51",
          5934 => x"2e",
          5935 => x"81",
          5936 => x"c0",
          5937 => x"52",
          5938 => x"92",
          5939 => x"75",
          5940 => x"0c",
          5941 => x"04",
          5942 => x"7b",
          5943 => x"b3",
          5944 => x"58",
          5945 => x"53",
          5946 => x"51",
          5947 => x"82",
          5948 => x"a4",
          5949 => x"2e",
          5950 => x"81",
          5951 => x"98",
          5952 => x"7f",
          5953 => x"dc",
          5954 => x"7d",
          5955 => x"82",
          5956 => x"57",
          5957 => x"04",
          5958 => x"dc",
          5959 => x"0d",
          5960 => x"0d",
          5961 => x"02",
          5962 => x"cf",
          5963 => x"73",
          5964 => x"5f",
          5965 => x"5e",
          5966 => x"82",
          5967 => x"fe",
          5968 => x"82",
          5969 => x"fe",
          5970 => x"80",
          5971 => x"27",
          5972 => x"7b",
          5973 => x"38",
          5974 => x"a7",
          5975 => x"39",
          5976 => x"72",
          5977 => x"38",
          5978 => x"82",
          5979 => x"fe",
          5980 => x"89",
          5981 => x"d4",
          5982 => x"8b",
          5983 => x"55",
          5984 => x"74",
          5985 => x"7a",
          5986 => x"72",
          5987 => x"81",
          5988 => x"f4",
          5989 => x"39",
          5990 => x"51",
          5991 => x"3f",
          5992 => x"a1",
          5993 => x"53",
          5994 => x"8e",
          5995 => x"52",
          5996 => x"51",
          5997 => x"3f",
          5998 => x"81",
          5999 => x"ee",
          6000 => x"15",
          6001 => x"fe",
          6002 => x"ff",
          6003 => x"81",
          6004 => x"ee",
          6005 => x"55",
          6006 => x"bc",
          6007 => x"70",
          6008 => x"80",
          6009 => x"27",
          6010 => x"56",
          6011 => x"74",
          6012 => x"81",
          6013 => x"06",
          6014 => x"06",
          6015 => x"80",
          6016 => x"73",
          6017 => x"85",
          6018 => x"83",
          6019 => x"fe",
          6020 => x"81",
          6021 => x"39",
          6022 => x"51",
          6023 => x"3f",
          6024 => x"1c",
          6025 => x"de",
          6026 => x"8c",
          6027 => x"2b",
          6028 => x"51",
          6029 => x"2e",
          6030 => x"ab",
          6031 => x"be",
          6032 => x"dc",
          6033 => x"70",
          6034 => x"a0",
          6035 => x"72",
          6036 => x"30",
          6037 => x"73",
          6038 => x"51",
          6039 => x"57",
          6040 => x"73",
          6041 => x"76",
          6042 => x"81",
          6043 => x"80",
          6044 => x"7c",
          6045 => x"78",
          6046 => x"38",
          6047 => x"82",
          6048 => x"8f",
          6049 => x"fc",
          6050 => x"9b",
          6051 => x"81",
          6052 => x"81",
          6053 => x"fe",
          6054 => x"82",
          6055 => x"51",
          6056 => x"3f",
          6057 => x"54",
          6058 => x"53",
          6059 => x"33",
          6060 => x"94",
          6061 => x"b3",
          6062 => x"2e",
          6063 => x"e2",
          6064 => x"3d",
          6065 => x"3d",
          6066 => x"96",
          6067 => x"fe",
          6068 => x"81",
          6069 => x"ba",
          6070 => x"b0",
          6071 => x"b2",
          6072 => x"fe",
          6073 => x"72",
          6074 => x"81",
          6075 => x"71",
          6076 => x"38",
          6077 => x"d9",
          6078 => x"82",
          6079 => x"db",
          6080 => x"51",
          6081 => x"3f",
          6082 => x"70",
          6083 => x"52",
          6084 => x"95",
          6085 => x"fe",
          6086 => x"82",
          6087 => x"fe",
          6088 => x"80",
          6089 => x"ea",
          6090 => x"2a",
          6091 => x"51",
          6092 => x"2e",
          6093 => x"51",
          6094 => x"3f",
          6095 => x"51",
          6096 => x"3f",
          6097 => x"d8",
          6098 => x"84",
          6099 => x"06",
          6100 => x"80",
          6101 => x"81",
          6102 => x"b6",
          6103 => x"80",
          6104 => x"ae",
          6105 => x"fe",
          6106 => x"72",
          6107 => x"81",
          6108 => x"71",
          6109 => x"38",
          6110 => x"d8",
          6111 => x"83",
          6112 => x"da",
          6113 => x"51",
          6114 => x"3f",
          6115 => x"70",
          6116 => x"52",
          6117 => x"95",
          6118 => x"fe",
          6119 => x"82",
          6120 => x"fe",
          6121 => x"80",
          6122 => x"e6",
          6123 => x"2a",
          6124 => x"51",
          6125 => x"2e",
          6126 => x"51",
          6127 => x"3f",
          6128 => x"51",
          6129 => x"3f",
          6130 => x"d7",
          6131 => x"88",
          6132 => x"06",
          6133 => x"80",
          6134 => x"81",
          6135 => x"b2",
          6136 => x"d0",
          6137 => x"aa",
          6138 => x"fe",
          6139 => x"fe",
          6140 => x"84",
          6141 => x"fb",
          6142 => x"02",
          6143 => x"05",
          6144 => x"56",
          6145 => x"75",
          6146 => x"e2",
          6147 => x"c8",
          6148 => x"a7",
          6149 => x"82",
          6150 => x"82",
          6151 => x"ff",
          6152 => x"82",
          6153 => x"30",
          6154 => x"dc",
          6155 => x"25",
          6156 => x"51",
          6157 => x"82",
          6158 => x"82",
          6159 => x"54",
          6160 => x"09",
          6161 => x"38",
          6162 => x"53",
          6163 => x"51",
          6164 => x"82",
          6165 => x"80",
          6166 => x"82",
          6167 => x"51",
          6168 => x"3f",
          6169 => x"a3",
          6170 => x"aa",
          6171 => x"82",
          6172 => x"82",
          6173 => x"54",
          6174 => x"09",
          6175 => x"38",
          6176 => x"51",
          6177 => x"3f",
          6178 => x"8c",
          6179 => x"3d",
          6180 => x"3d",
          6181 => x"71",
          6182 => x"0c",
          6183 => x"52",
          6184 => x"86",
          6185 => x"8c",
          6186 => x"ff",
          6187 => x"7d",
          6188 => x"06",
          6189 => x"84",
          6190 => x"3d",
          6191 => x"fe",
          6192 => x"7c",
          6193 => x"82",
          6194 => x"ff",
          6195 => x"82",
          6196 => x"7d",
          6197 => x"82",
          6198 => x"8d",
          6199 => x"70",
          6200 => x"84",
          6201 => x"e8",
          6202 => x"3d",
          6203 => x"80",
          6204 => x"51",
          6205 => x"b4",
          6206 => x"05",
          6207 => x"3f",
          6208 => x"08",
          6209 => x"90",
          6210 => x"78",
          6211 => x"87",
          6212 => x"80",
          6213 => x"38",
          6214 => x"81",
          6215 => x"bd",
          6216 => x"78",
          6217 => x"ba",
          6218 => x"2e",
          6219 => x"8a",
          6220 => x"80",
          6221 => x"a1",
          6222 => x"c0",
          6223 => x"38",
          6224 => x"82",
          6225 => x"d2",
          6226 => x"f9",
          6227 => x"38",
          6228 => x"24",
          6229 => x"80",
          6230 => x"98",
          6231 => x"f8",
          6232 => x"38",
          6233 => x"78",
          6234 => x"8a",
          6235 => x"81",
          6236 => x"38",
          6237 => x"2e",
          6238 => x"8a",
          6239 => x"81",
          6240 => x"8f",
          6241 => x"39",
          6242 => x"80",
          6243 => x"84",
          6244 => x"ee",
          6245 => x"8c",
          6246 => x"2e",
          6247 => x"b4",
          6248 => x"11",
          6249 => x"05",
          6250 => x"b4",
          6251 => x"dc",
          6252 => x"fe",
          6253 => x"3d",
          6254 => x"53",
          6255 => x"51",
          6256 => x"3f",
          6257 => x"08",
          6258 => x"8c",
          6259 => x"82",
          6260 => x"fe",
          6261 => x"63",
          6262 => x"79",
          6263 => x"f2",
          6264 => x"78",
          6265 => x"05",
          6266 => x"7a",
          6267 => x"81",
          6268 => x"3d",
          6269 => x"53",
          6270 => x"51",
          6271 => x"3f",
          6272 => x"08",
          6273 => x"da",
          6274 => x"fe",
          6275 => x"ff",
          6276 => x"fe",
          6277 => x"82",
          6278 => x"80",
          6279 => x"38",
          6280 => x"f8",
          6281 => x"84",
          6282 => x"ed",
          6283 => x"8c",
          6284 => x"2e",
          6285 => x"82",
          6286 => x"fe",
          6287 => x"63",
          6288 => x"27",
          6289 => x"61",
          6290 => x"81",
          6291 => x"79",
          6292 => x"05",
          6293 => x"b4",
          6294 => x"11",
          6295 => x"05",
          6296 => x"fc",
          6297 => x"dc",
          6298 => x"fc",
          6299 => x"3d",
          6300 => x"53",
          6301 => x"51",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"de",
          6305 => x"fe",
          6306 => x"ff",
          6307 => x"fe",
          6308 => x"82",
          6309 => x"80",
          6310 => x"38",
          6311 => x"51",
          6312 => x"3f",
          6313 => x"63",
          6314 => x"61",
          6315 => x"33",
          6316 => x"78",
          6317 => x"38",
          6318 => x"54",
          6319 => x"79",
          6320 => x"8c",
          6321 => x"a3",
          6322 => x"62",
          6323 => x"5a",
          6324 => x"85",
          6325 => x"bd",
          6326 => x"ff",
          6327 => x"ff",
          6328 => x"fe",
          6329 => x"82",
          6330 => x"80",
          6331 => x"88",
          6332 => x"78",
          6333 => x"38",
          6334 => x"08",
          6335 => x"39",
          6336 => x"33",
          6337 => x"2e",
          6338 => x"87",
          6339 => x"bc",
          6340 => x"a2",
          6341 => x"80",
          6342 => x"82",
          6343 => x"44",
          6344 => x"88",
          6345 => x"78",
          6346 => x"38",
          6347 => x"08",
          6348 => x"82",
          6349 => x"59",
          6350 => x"88",
          6351 => x"f8",
          6352 => x"39",
          6353 => x"08",
          6354 => x"44",
          6355 => x"fc",
          6356 => x"84",
          6357 => x"eb",
          6358 => x"8c",
          6359 => x"de",
          6360 => x"a0",
          6361 => x"80",
          6362 => x"82",
          6363 => x"43",
          6364 => x"82",
          6365 => x"59",
          6366 => x"88",
          6367 => x"e4",
          6368 => x"39",
          6369 => x"33",
          6370 => x"2e",
          6371 => x"87",
          6372 => x"aa",
          6373 => x"a3",
          6374 => x"80",
          6375 => x"82",
          6376 => x"43",
          6377 => x"88",
          6378 => x"78",
          6379 => x"38",
          6380 => x"08",
          6381 => x"82",
          6382 => x"88",
          6383 => x"3d",
          6384 => x"53",
          6385 => x"51",
          6386 => x"3f",
          6387 => x"08",
          6388 => x"38",
          6389 => x"5c",
          6390 => x"83",
          6391 => x"7a",
          6392 => x"30",
          6393 => x"9f",
          6394 => x"06",
          6395 => x"5a",
          6396 => x"88",
          6397 => x"2e",
          6398 => x"42",
          6399 => x"51",
          6400 => x"3f",
          6401 => x"54",
          6402 => x"52",
          6403 => x"91",
          6404 => x"b8",
          6405 => x"ef",
          6406 => x"39",
          6407 => x"80",
          6408 => x"84",
          6409 => x"e9",
          6410 => x"8c",
          6411 => x"2e",
          6412 => x"b4",
          6413 => x"11",
          6414 => x"05",
          6415 => x"a0",
          6416 => x"dc",
          6417 => x"a5",
          6418 => x"02",
          6419 => x"33",
          6420 => x"81",
          6421 => x"3d",
          6422 => x"53",
          6423 => x"51",
          6424 => x"3f",
          6425 => x"08",
          6426 => x"f6",
          6427 => x"33",
          6428 => x"85",
          6429 => x"e6",
          6430 => x"f8",
          6431 => x"fe",
          6432 => x"79",
          6433 => x"59",
          6434 => x"f8",
          6435 => x"79",
          6436 => x"b4",
          6437 => x"11",
          6438 => x"05",
          6439 => x"c0",
          6440 => x"dc",
          6441 => x"91",
          6442 => x"02",
          6443 => x"33",
          6444 => x"81",
          6445 => x"b5",
          6446 => x"d0",
          6447 => x"c7",
          6448 => x"39",
          6449 => x"f4",
          6450 => x"84",
          6451 => x"ea",
          6452 => x"8c",
          6453 => x"2e",
          6454 => x"b4",
          6455 => x"11",
          6456 => x"05",
          6457 => x"ea",
          6458 => x"dc",
          6459 => x"a6",
          6460 => x"02",
          6461 => x"79",
          6462 => x"5b",
          6463 => x"b4",
          6464 => x"11",
          6465 => x"05",
          6466 => x"c6",
          6467 => x"dc",
          6468 => x"f7",
          6469 => x"70",
          6470 => x"82",
          6471 => x"fe",
          6472 => x"80",
          6473 => x"51",
          6474 => x"3f",
          6475 => x"33",
          6476 => x"2e",
          6477 => x"78",
          6478 => x"38",
          6479 => x"41",
          6480 => x"3d",
          6481 => x"53",
          6482 => x"51",
          6483 => x"3f",
          6484 => x"08",
          6485 => x"38",
          6486 => x"be",
          6487 => x"70",
          6488 => x"23",
          6489 => x"ae",
          6490 => x"d0",
          6491 => x"97",
          6492 => x"39",
          6493 => x"f4",
          6494 => x"84",
          6495 => x"e8",
          6496 => x"8c",
          6497 => x"2e",
          6498 => x"b4",
          6499 => x"11",
          6500 => x"05",
          6501 => x"ba",
          6502 => x"dc",
          6503 => x"a1",
          6504 => x"71",
          6505 => x"84",
          6506 => x"3d",
          6507 => x"53",
          6508 => x"51",
          6509 => x"3f",
          6510 => x"08",
          6511 => x"a2",
          6512 => x"08",
          6513 => x"85",
          6514 => x"e4",
          6515 => x"f8",
          6516 => x"fe",
          6517 => x"79",
          6518 => x"59",
          6519 => x"f6",
          6520 => x"79",
          6521 => x"b4",
          6522 => x"11",
          6523 => x"05",
          6524 => x"de",
          6525 => x"dc",
          6526 => x"8d",
          6527 => x"71",
          6528 => x"84",
          6529 => x"b9",
          6530 => x"d0",
          6531 => x"f7",
          6532 => x"39",
          6533 => x"80",
          6534 => x"84",
          6535 => x"e5",
          6536 => x"8c",
          6537 => x"2e",
          6538 => x"63",
          6539 => x"f0",
          6540 => x"b7",
          6541 => x"78",
          6542 => x"ff",
          6543 => x"ff",
          6544 => x"fe",
          6545 => x"82",
          6546 => x"80",
          6547 => x"38",
          6548 => x"86",
          6549 => x"e3",
          6550 => x"59",
          6551 => x"8c",
          6552 => x"2e",
          6553 => x"82",
          6554 => x"52",
          6555 => x"51",
          6556 => x"3f",
          6557 => x"82",
          6558 => x"fe",
          6559 => x"fe",
          6560 => x"f4",
          6561 => x"86",
          6562 => x"dc",
          6563 => x"59",
          6564 => x"fe",
          6565 => x"f4",
          6566 => x"45",
          6567 => x"78",
          6568 => x"be",
          6569 => x"06",
          6570 => x"2e",
          6571 => x"b4",
          6572 => x"05",
          6573 => x"8b",
          6574 => x"dc",
          6575 => x"5b",
          6576 => x"b2",
          6577 => x"24",
          6578 => x"81",
          6579 => x"80",
          6580 => x"83",
          6581 => x"80",
          6582 => x"86",
          6583 => x"55",
          6584 => x"54",
          6585 => x"86",
          6586 => x"3d",
          6587 => x"51",
          6588 => x"3f",
          6589 => x"87",
          6590 => x"3d",
          6591 => x"51",
          6592 => x"3f",
          6593 => x"55",
          6594 => x"54",
          6595 => x"87",
          6596 => x"3d",
          6597 => x"51",
          6598 => x"3f",
          6599 => x"54",
          6600 => x"87",
          6601 => x"3d",
          6602 => x"51",
          6603 => x"3f",
          6604 => x"58",
          6605 => x"57",
          6606 => x"55",
          6607 => x"80",
          6608 => x"80",
          6609 => x"3d",
          6610 => x"51",
          6611 => x"82",
          6612 => x"82",
          6613 => x"09",
          6614 => x"72",
          6615 => x"51",
          6616 => x"80",
          6617 => x"26",
          6618 => x"5a",
          6619 => x"59",
          6620 => x"8d",
          6621 => x"70",
          6622 => x"5c",
          6623 => x"c0",
          6624 => x"32",
          6625 => x"07",
          6626 => x"38",
          6627 => x"09",
          6628 => x"ce",
          6629 => x"a0",
          6630 => x"cf",
          6631 => x"39",
          6632 => x"80",
          6633 => x"a4",
          6634 => x"94",
          6635 => x"54",
          6636 => x"80",
          6637 => x"fe",
          6638 => x"82",
          6639 => x"90",
          6640 => x"55",
          6641 => x"80",
          6642 => x"fe",
          6643 => x"72",
          6644 => x"08",
          6645 => x"87",
          6646 => x"70",
          6647 => x"87",
          6648 => x"72",
          6649 => x"f3",
          6650 => x"dc",
          6651 => x"75",
          6652 => x"87",
          6653 => x"73",
          6654 => x"df",
          6655 => x"8c",
          6656 => x"75",
          6657 => x"83",
          6658 => x"94",
          6659 => x"80",
          6660 => x"c0",
          6661 => x"b7",
          6662 => x"8c",
          6663 => x"ad",
          6664 => x"f4",
          6665 => x"ae",
          6666 => x"d7",
          6667 => x"b0",
          6668 => x"d3",
          6669 => x"bc",
          6670 => x"cb",
          6671 => x"c6",
          6672 => x"ba",
          6673 => x"ec",
          6674 => x"c6",
          6675 => x"00",
          6676 => x"55",
          6677 => x"5b",
          6678 => x"61",
          6679 => x"67",
          6680 => x"6d",
          6681 => x"d8",
          6682 => x"b4",
          6683 => x"57",
          6684 => x"97",
          6685 => x"ba",
          6686 => x"47",
          6687 => x"ad",
          6688 => x"ad",
          6689 => x"84",
          6690 => x"fa",
          6691 => x"85",
          6692 => x"ae",
          6693 => x"cc",
          6694 => x"50",
          6695 => x"57",
          6696 => x"5e",
          6697 => x"65",
          6698 => x"6c",
          6699 => x"73",
          6700 => x"7a",
          6701 => x"81",
          6702 => x"88",
          6703 => x"8f",
          6704 => x"96",
          6705 => x"9c",
          6706 => x"a2",
          6707 => x"a8",
          6708 => x"ae",
          6709 => x"b4",
          6710 => x"ba",
          6711 => x"c0",
          6712 => x"c6",
          6713 => x"25",
          6714 => x"64",
          6715 => x"3a",
          6716 => x"25",
          6717 => x"64",
          6718 => x"00",
          6719 => x"20",
          6720 => x"66",
          6721 => x"72",
          6722 => x"6f",
          6723 => x"00",
          6724 => x"72",
          6725 => x"53",
          6726 => x"63",
          6727 => x"69",
          6728 => x"00",
          6729 => x"65",
          6730 => x"65",
          6731 => x"6d",
          6732 => x"6d",
          6733 => x"65",
          6734 => x"00",
          6735 => x"20",
          6736 => x"53",
          6737 => x"4d",
          6738 => x"25",
          6739 => x"3a",
          6740 => x"58",
          6741 => x"00",
          6742 => x"20",
          6743 => x"41",
          6744 => x"20",
          6745 => x"25",
          6746 => x"3a",
          6747 => x"58",
          6748 => x"00",
          6749 => x"20",
          6750 => x"4e",
          6751 => x"41",
          6752 => x"25",
          6753 => x"3a",
          6754 => x"58",
          6755 => x"00",
          6756 => x"20",
          6757 => x"4d",
          6758 => x"20",
          6759 => x"25",
          6760 => x"3a",
          6761 => x"58",
          6762 => x"00",
          6763 => x"20",
          6764 => x"20",
          6765 => x"20",
          6766 => x"25",
          6767 => x"3a",
          6768 => x"58",
          6769 => x"00",
          6770 => x"20",
          6771 => x"43",
          6772 => x"20",
          6773 => x"44",
          6774 => x"63",
          6775 => x"3d",
          6776 => x"64",
          6777 => x"00",
          6778 => x"20",
          6779 => x"45",
          6780 => x"20",
          6781 => x"54",
          6782 => x"72",
          6783 => x"3d",
          6784 => x"64",
          6785 => x"00",
          6786 => x"20",
          6787 => x"52",
          6788 => x"52",
          6789 => x"43",
          6790 => x"6e",
          6791 => x"3d",
          6792 => x"64",
          6793 => x"00",
          6794 => x"20",
          6795 => x"48",
          6796 => x"45",
          6797 => x"53",
          6798 => x"00",
          6799 => x"20",
          6800 => x"49",
          6801 => x"00",
          6802 => x"20",
          6803 => x"54",
          6804 => x"00",
          6805 => x"20",
          6806 => x"0a",
          6807 => x"00",
          6808 => x"20",
          6809 => x"0a",
          6810 => x"00",
          6811 => x"72",
          6812 => x"65",
          6813 => x"00",
          6814 => x"20",
          6815 => x"20",
          6816 => x"65",
          6817 => x"65",
          6818 => x"72",
          6819 => x"64",
          6820 => x"73",
          6821 => x"25",
          6822 => x"0a",
          6823 => x"00",
          6824 => x"20",
          6825 => x"20",
          6826 => x"6f",
          6827 => x"53",
          6828 => x"74",
          6829 => x"64",
          6830 => x"73",
          6831 => x"25",
          6832 => x"0a",
          6833 => x"00",
          6834 => x"20",
          6835 => x"63",
          6836 => x"74",
          6837 => x"20",
          6838 => x"72",
          6839 => x"20",
          6840 => x"20",
          6841 => x"25",
          6842 => x"0a",
          6843 => x"00",
          6844 => x"63",
          6845 => x"00",
          6846 => x"20",
          6847 => x"20",
          6848 => x"20",
          6849 => x"20",
          6850 => x"20",
          6851 => x"20",
          6852 => x"20",
          6853 => x"25",
          6854 => x"0a",
          6855 => x"00",
          6856 => x"20",
          6857 => x"74",
          6858 => x"43",
          6859 => x"6b",
          6860 => x"65",
          6861 => x"20",
          6862 => x"20",
          6863 => x"25",
          6864 => x"30",
          6865 => x"48",
          6866 => x"00",
          6867 => x"20",
          6868 => x"41",
          6869 => x"6c",
          6870 => x"20",
          6871 => x"71",
          6872 => x"20",
          6873 => x"20",
          6874 => x"25",
          6875 => x"30",
          6876 => x"48",
          6877 => x"00",
          6878 => x"20",
          6879 => x"68",
          6880 => x"65",
          6881 => x"52",
          6882 => x"43",
          6883 => x"6b",
          6884 => x"65",
          6885 => x"25",
          6886 => x"30",
          6887 => x"48",
          6888 => x"00",
          6889 => x"6c",
          6890 => x"00",
          6891 => x"69",
          6892 => x"00",
          6893 => x"78",
          6894 => x"00",
          6895 => x"00",
          6896 => x"6d",
          6897 => x"00",
          6898 => x"6e",
          6899 => x"00",
          6900 => x"74",
          6901 => x"2e",
          6902 => x"00",
          6903 => x"74",
          6904 => x"00",
          6905 => x"74",
          6906 => x"00",
          6907 => x"00",
          6908 => x"64",
          6909 => x"73",
          6910 => x"00",
          6911 => x"6c",
          6912 => x"74",
          6913 => x"65",
          6914 => x"20",
          6915 => x"20",
          6916 => x"74",
          6917 => x"20",
          6918 => x"65",
          6919 => x"20",
          6920 => x"2e",
          6921 => x"00",
          6922 => x"6e",
          6923 => x"6f",
          6924 => x"2f",
          6925 => x"61",
          6926 => x"68",
          6927 => x"6f",
          6928 => x"66",
          6929 => x"2c",
          6930 => x"73",
          6931 => x"69",
          6932 => x"0a",
          6933 => x"00",
          6934 => x"04",
          6935 => x"00",
          6936 => x"01",
          6937 => x"00",
          6938 => x"00",
          6939 => x"02",
          6940 => x"fc",
          6941 => x"00",
          6942 => x"03",
          6943 => x"f8",
          6944 => x"00",
          6945 => x"04",
          6946 => x"f4",
          6947 => x"00",
          6948 => x"05",
          6949 => x"f0",
          6950 => x"00",
          6951 => x"06",
          6952 => x"ec",
          6953 => x"00",
          6954 => x"07",
          6955 => x"e8",
          6956 => x"00",
          6957 => x"08",
          6958 => x"e4",
          6959 => x"00",
          6960 => x"09",
          6961 => x"e0",
          6962 => x"00",
          6963 => x"0a",
          6964 => x"dc",
          6965 => x"00",
          6966 => x"0b",
          6967 => x"00",
          6968 => x"00",
          6969 => x"00",
          6970 => x"00",
          6971 => x"7e",
          6972 => x"7e",
          6973 => x"7e",
          6974 => x"7e",
          6975 => x"7e",
          6976 => x"00",
          6977 => x"00",
          6978 => x"00",
          6979 => x"2c",
          6980 => x"3d",
          6981 => x"5d",
          6982 => x"00",
          6983 => x"00",
          6984 => x"33",
          6985 => x"00",
          6986 => x"4d",
          6987 => x"53",
          6988 => x"00",
          6989 => x"4e",
          6990 => x"20",
          6991 => x"46",
          6992 => x"32",
          6993 => x"00",
          6994 => x"4e",
          6995 => x"20",
          6996 => x"46",
          6997 => x"20",
          6998 => x"00",
          6999 => x"08",
          7000 => x"00",
          7001 => x"00",
          7002 => x"00",
          7003 => x"41",
          7004 => x"80",
          7005 => x"49",
          7006 => x"8f",
          7007 => x"4f",
          7008 => x"55",
          7009 => x"9b",
          7010 => x"9f",
          7011 => x"55",
          7012 => x"a7",
          7013 => x"ab",
          7014 => x"af",
          7015 => x"b3",
          7016 => x"b7",
          7017 => x"bb",
          7018 => x"bf",
          7019 => x"c3",
          7020 => x"c7",
          7021 => x"cb",
          7022 => x"cf",
          7023 => x"d3",
          7024 => x"d7",
          7025 => x"db",
          7026 => x"df",
          7027 => x"e3",
          7028 => x"e7",
          7029 => x"eb",
          7030 => x"ef",
          7031 => x"f3",
          7032 => x"f7",
          7033 => x"fb",
          7034 => x"ff",
          7035 => x"3b",
          7036 => x"2f",
          7037 => x"3a",
          7038 => x"7c",
          7039 => x"00",
          7040 => x"04",
          7041 => x"40",
          7042 => x"00",
          7043 => x"00",
          7044 => x"02",
          7045 => x"08",
          7046 => x"20",
          7047 => x"00",
          7048 => x"69",
          7049 => x"00",
          7050 => x"63",
          7051 => x"00",
          7052 => x"69",
          7053 => x"00",
          7054 => x"61",
          7055 => x"00",
          7056 => x"65",
          7057 => x"00",
          7058 => x"65",
          7059 => x"00",
          7060 => x"70",
          7061 => x"00",
          7062 => x"66",
          7063 => x"00",
          7064 => x"6d",
          7065 => x"00",
          7066 => x"00",
          7067 => x"00",
          7068 => x"00",
          7069 => x"00",
          7070 => x"00",
          7071 => x"00",
          7072 => x"00",
          7073 => x"6c",
          7074 => x"00",
          7075 => x"00",
          7076 => x"74",
          7077 => x"00",
          7078 => x"65",
          7079 => x"00",
          7080 => x"6f",
          7081 => x"00",
          7082 => x"74",
          7083 => x"00",
          7084 => x"73",
          7085 => x"00",
          7086 => x"73",
          7087 => x"00",
          7088 => x"6f",
          7089 => x"00",
          7090 => x"6b",
          7091 => x"72",
          7092 => x"00",
          7093 => x"65",
          7094 => x"6c",
          7095 => x"72",
          7096 => x"0a",
          7097 => x"00",
          7098 => x"6b",
          7099 => x"74",
          7100 => x"61",
          7101 => x"0a",
          7102 => x"00",
          7103 => x"66",
          7104 => x"20",
          7105 => x"6e",
          7106 => x"00",
          7107 => x"70",
          7108 => x"20",
          7109 => x"6e",
          7110 => x"00",
          7111 => x"61",
          7112 => x"20",
          7113 => x"65",
          7114 => x"65",
          7115 => x"00",
          7116 => x"65",
          7117 => x"64",
          7118 => x"65",
          7119 => x"00",
          7120 => x"65",
          7121 => x"72",
          7122 => x"79",
          7123 => x"69",
          7124 => x"2e",
          7125 => x"00",
          7126 => x"65",
          7127 => x"6e",
          7128 => x"20",
          7129 => x"61",
          7130 => x"2e",
          7131 => x"00",
          7132 => x"69",
          7133 => x"72",
          7134 => x"20",
          7135 => x"74",
          7136 => x"65",
          7137 => x"00",
          7138 => x"76",
          7139 => x"75",
          7140 => x"72",
          7141 => x"20",
          7142 => x"61",
          7143 => x"2e",
          7144 => x"00",
          7145 => x"6b",
          7146 => x"74",
          7147 => x"61",
          7148 => x"64",
          7149 => x"00",
          7150 => x"63",
          7151 => x"61",
          7152 => x"6c",
          7153 => x"69",
          7154 => x"79",
          7155 => x"6d",
          7156 => x"75",
          7157 => x"6f",
          7158 => x"69",
          7159 => x"0a",
          7160 => x"00",
          7161 => x"6d",
          7162 => x"61",
          7163 => x"74",
          7164 => x"0a",
          7165 => x"00",
          7166 => x"65",
          7167 => x"2c",
          7168 => x"65",
          7169 => x"69",
          7170 => x"63",
          7171 => x"65",
          7172 => x"64",
          7173 => x"00",
          7174 => x"65",
          7175 => x"20",
          7176 => x"6b",
          7177 => x"0a",
          7178 => x"00",
          7179 => x"75",
          7180 => x"63",
          7181 => x"74",
          7182 => x"6d",
          7183 => x"2e",
          7184 => x"00",
          7185 => x"20",
          7186 => x"79",
          7187 => x"65",
          7188 => x"69",
          7189 => x"2e",
          7190 => x"00",
          7191 => x"61",
          7192 => x"65",
          7193 => x"69",
          7194 => x"72",
          7195 => x"74",
          7196 => x"00",
          7197 => x"63",
          7198 => x"2e",
          7199 => x"00",
          7200 => x"6e",
          7201 => x"20",
          7202 => x"6f",
          7203 => x"00",
          7204 => x"75",
          7205 => x"74",
          7206 => x"25",
          7207 => x"74",
          7208 => x"75",
          7209 => x"74",
          7210 => x"73",
          7211 => x"0a",
          7212 => x"00",
          7213 => x"64",
          7214 => x"00",
          7215 => x"58",
          7216 => x"00",
          7217 => x"00",
          7218 => x"58",
          7219 => x"00",
          7220 => x"20",
          7221 => x"20",
          7222 => x"00",
          7223 => x"58",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"00",
          7228 => x"00",
          7229 => x"20",
          7230 => x"28",
          7231 => x"00",
          7232 => x"30",
          7233 => x"30",
          7234 => x"00",
          7235 => x"30",
          7236 => x"00",
          7237 => x"55",
          7238 => x"65",
          7239 => x"30",
          7240 => x"20",
          7241 => x"25",
          7242 => x"2a",
          7243 => x"00",
          7244 => x"20",
          7245 => x"65",
          7246 => x"70",
          7247 => x"61",
          7248 => x"65",
          7249 => x"00",
          7250 => x"65",
          7251 => x"6e",
          7252 => x"72",
          7253 => x"0a",
          7254 => x"00",
          7255 => x"20",
          7256 => x"65",
          7257 => x"70",
          7258 => x"00",
          7259 => x"54",
          7260 => x"44",
          7261 => x"74",
          7262 => x"75",
          7263 => x"00",
          7264 => x"54",
          7265 => x"52",
          7266 => x"74",
          7267 => x"75",
          7268 => x"00",
          7269 => x"54",
          7270 => x"58",
          7271 => x"74",
          7272 => x"75",
          7273 => x"00",
          7274 => x"54",
          7275 => x"58",
          7276 => x"74",
          7277 => x"75",
          7278 => x"00",
          7279 => x"54",
          7280 => x"58",
          7281 => x"74",
          7282 => x"75",
          7283 => x"00",
          7284 => x"54",
          7285 => x"58",
          7286 => x"74",
          7287 => x"75",
          7288 => x"00",
          7289 => x"74",
          7290 => x"20",
          7291 => x"74",
          7292 => x"72",
          7293 => x"0a",
          7294 => x"00",
          7295 => x"62",
          7296 => x"67",
          7297 => x"6d",
          7298 => x"2e",
          7299 => x"00",
          7300 => x"6f",
          7301 => x"63",
          7302 => x"74",
          7303 => x"00",
          7304 => x"00",
          7305 => x"6c",
          7306 => x"74",
          7307 => x"6e",
          7308 => x"61",
          7309 => x"65",
          7310 => x"20",
          7311 => x"64",
          7312 => x"20",
          7313 => x"61",
          7314 => x"69",
          7315 => x"20",
          7316 => x"75",
          7317 => x"79",
          7318 => x"00",
          7319 => x"00",
          7320 => x"61",
          7321 => x"67",
          7322 => x"2e",
          7323 => x"00",
          7324 => x"79",
          7325 => x"2e",
          7326 => x"00",
          7327 => x"70",
          7328 => x"6e",
          7329 => x"2e",
          7330 => x"00",
          7331 => x"6c",
          7332 => x"30",
          7333 => x"2d",
          7334 => x"38",
          7335 => x"25",
          7336 => x"29",
          7337 => x"00",
          7338 => x"70",
          7339 => x"6d",
          7340 => x"0a",
          7341 => x"00",
          7342 => x"6d",
          7343 => x"74",
          7344 => x"00",
          7345 => x"58",
          7346 => x"32",
          7347 => x"00",
          7348 => x"0a",
          7349 => x"00",
          7350 => x"58",
          7351 => x"34",
          7352 => x"00",
          7353 => x"58",
          7354 => x"38",
          7355 => x"00",
          7356 => x"63",
          7357 => x"6e",
          7358 => x"6f",
          7359 => x"40",
          7360 => x"38",
          7361 => x"2e",
          7362 => x"00",
          7363 => x"6c",
          7364 => x"20",
          7365 => x"65",
          7366 => x"25",
          7367 => x"20",
          7368 => x"0a",
          7369 => x"00",
          7370 => x"6c",
          7371 => x"74",
          7372 => x"65",
          7373 => x"6f",
          7374 => x"28",
          7375 => x"2e",
          7376 => x"00",
          7377 => x"74",
          7378 => x"69",
          7379 => x"61",
          7380 => x"69",
          7381 => x"69",
          7382 => x"2e",
          7383 => x"00",
          7384 => x"64",
          7385 => x"62",
          7386 => x"69",
          7387 => x"2e",
          7388 => x"00",
          7389 => x"00",
          7390 => x"00",
          7391 => x"5c",
          7392 => x"25",
          7393 => x"73",
          7394 => x"00",
          7395 => x"5c",
          7396 => x"25",
          7397 => x"00",
          7398 => x"5c",
          7399 => x"00",
          7400 => x"20",
          7401 => x"6d",
          7402 => x"2e",
          7403 => x"00",
          7404 => x"6e",
          7405 => x"2e",
          7406 => x"00",
          7407 => x"62",
          7408 => x"67",
          7409 => x"74",
          7410 => x"75",
          7411 => x"2e",
          7412 => x"00",
          7413 => x"00",
          7414 => x"00",
          7415 => x"ff",
          7416 => x"00",
          7417 => x"ff",
          7418 => x"00",
          7419 => x"ff",
          7420 => x"00",
          7421 => x"00",
          7422 => x"00",
          7423 => x"ff",
          7424 => x"00",
          7425 => x"00",
          7426 => x"00",
          7427 => x"00",
          7428 => x"00",
          7429 => x"00",
          7430 => x"00",
          7431 => x"00",
          7432 => x"01",
          7433 => x"01",
          7434 => x"01",
          7435 => x"00",
          7436 => x"00",
          7437 => x"02",
          7438 => x"00",
          7439 => x"34",
          7440 => x"34",
          7441 => x"34",
          7442 => x"34",
          7443 => x"d0",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"dc",
          7468 => x"00",
          7469 => x"e4",
          7470 => x"00",
          7471 => x"ec",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"20",
          7476 => x"00",
          7477 => x"00",
          7478 => x"00",
          7479 => x"28",
          7480 => x"00",
          7481 => x"00",
          7482 => x"00",
          7483 => x"30",
          7484 => x"00",
          7485 => x"00",
          7486 => x"00",
          7487 => x"38",
          7488 => x"00",
          7489 => x"00",
          7490 => x"00",
          7491 => x"40",
          7492 => x"00",
          7493 => x"00",
          7494 => x"00",
          7495 => x"48",
          7496 => x"00",
          7497 => x"00",
          7498 => x"00",
          7499 => x"50",
          7500 => x"00",
          7501 => x"00",
          7502 => x"00",
          7503 => x"58",
          7504 => x"00",
          7505 => x"00",
          7506 => x"00",
          7507 => x"60",
          7508 => x"00",
          7509 => x"00",
          7510 => x"00",
          7511 => x"68",
          7512 => x"00",
          7513 => x"00",
          7514 => x"00",
          7515 => x"6c",
          7516 => x"00",
          7517 => x"00",
          7518 => x"00",
          7519 => x"70",
          7520 => x"00",
          7521 => x"00",
          7522 => x"00",
          7523 => x"74",
          7524 => x"00",
          7525 => x"00",
          7526 => x"00",
          7527 => x"78",
          7528 => x"00",
          7529 => x"00",
          7530 => x"00",
          7531 => x"7c",
          7532 => x"00",
          7533 => x"00",
          7534 => x"00",
          7535 => x"80",
          7536 => x"00",
          7537 => x"00",
          7538 => x"00",
          7539 => x"84",
          7540 => x"00",
          7541 => x"00",
          7542 => x"00",
          7543 => x"8c",
          7544 => x"00",
          7545 => x"00",
          7546 => x"00",
          7547 => x"90",
          7548 => x"00",
          7549 => x"00",
          7550 => x"00",
          7551 => x"98",
          7552 => x"00",
          7553 => x"00",
          7554 => x"00",
          7555 => x"a0",
          7556 => x"00",
          7557 => x"00",
          7558 => x"00",
          7559 => x"a8",
          7560 => x"00",
          7561 => x"00",
          7562 => x"00",
          7563 => x"b0",
          7564 => x"00",
          7565 => x"00",
          7566 => x"00",
          7567 => x"b8",
          7568 => x"00",
          7569 => x"00",
          7570 => x"00",
          7571 => x"c0",
          7572 => x"00",
          7573 => x"00",
          7574 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"bb",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"0b",
            10 => x"84",
            11 => x"0b",
            12 => x"0b",
            13 => x"a3",
            14 => x"0b",
            15 => x"0b",
            16 => x"c3",
            17 => x"0b",
            18 => x"0b",
            19 => x"e3",
            20 => x"0b",
            21 => x"0b",
            22 => x"83",
            23 => x"0b",
            24 => x"0b",
            25 => x"a3",
            26 => x"0b",
            27 => x"0b",
            28 => x"c3",
            29 => x"0b",
            30 => x"0b",
            31 => x"e2",
            32 => x"0b",
            33 => x"0b",
            34 => x"80",
            35 => x"0b",
            36 => x"0b",
            37 => x"9e",
            38 => x"0b",
            39 => x"0b",
            40 => x"be",
            41 => x"0b",
            42 => x"0b",
            43 => x"de",
            44 => x"0b",
            45 => x"0b",
            46 => x"fe",
            47 => x"0b",
            48 => x"0b",
            49 => x"9e",
            50 => x"0b",
            51 => x"0b",
            52 => x"be",
            53 => x"0b",
            54 => x"0b",
            55 => x"de",
            56 => x"0b",
            57 => x"0b",
            58 => x"fe",
            59 => x"0b",
            60 => x"0b",
            61 => x"9e",
            62 => x"0b",
            63 => x"0b",
            64 => x"be",
            65 => x"0b",
            66 => x"0b",
            67 => x"de",
            68 => x"0b",
            69 => x"0b",
            70 => x"fe",
            71 => x"0b",
            72 => x"0b",
            73 => x"9e",
            74 => x"0b",
            75 => x"0b",
            76 => x"be",
            77 => x"0b",
            78 => x"0b",
            79 => x"de",
            80 => x"0b",
            81 => x"0b",
            82 => x"fe",
            83 => x"0b",
            84 => x"0b",
            85 => x"9c",
            86 => x"0b",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"80",
           129 => x"e8",
           130 => x"2d",
           131 => x"08",
           132 => x"04",
           133 => x"0c",
           134 => x"2d",
           135 => x"08",
           136 => x"04",
           137 => x"0c",
           138 => x"2d",
           139 => x"08",
           140 => x"04",
           141 => x"0c",
           142 => x"2d",
           143 => x"08",
           144 => x"04",
           145 => x"0c",
           146 => x"2d",
           147 => x"08",
           148 => x"04",
           149 => x"0c",
           150 => x"2d",
           151 => x"08",
           152 => x"04",
           153 => x"0c",
           154 => x"2d",
           155 => x"08",
           156 => x"04",
           157 => x"0c",
           158 => x"2d",
           159 => x"08",
           160 => x"04",
           161 => x"0c",
           162 => x"2d",
           163 => x"08",
           164 => x"04",
           165 => x"0c",
           166 => x"2d",
           167 => x"08",
           168 => x"04",
           169 => x"0c",
           170 => x"2d",
           171 => x"08",
           172 => x"04",
           173 => x"0c",
           174 => x"2d",
           175 => x"08",
           176 => x"04",
           177 => x"0c",
           178 => x"2d",
           179 => x"08",
           180 => x"04",
           181 => x"0c",
           182 => x"82",
           183 => x"83",
           184 => x"82",
           185 => x"ba",
           186 => x"8c",
           187 => x"80",
           188 => x"8c",
           189 => x"9a",
           190 => x"e8",
           191 => x"90",
           192 => x"e8",
           193 => x"2d",
           194 => x"08",
           195 => x"04",
           196 => x"0c",
           197 => x"82",
           198 => x"83",
           199 => x"82",
           200 => x"81",
           201 => x"82",
           202 => x"83",
           203 => x"82",
           204 => x"81",
           205 => x"82",
           206 => x"83",
           207 => x"82",
           208 => x"81",
           209 => x"82",
           210 => x"83",
           211 => x"82",
           212 => x"81",
           213 => x"82",
           214 => x"83",
           215 => x"82",
           216 => x"81",
           217 => x"82",
           218 => x"83",
           219 => x"82",
           220 => x"81",
           221 => x"82",
           222 => x"83",
           223 => x"82",
           224 => x"81",
           225 => x"82",
           226 => x"83",
           227 => x"82",
           228 => x"81",
           229 => x"82",
           230 => x"83",
           231 => x"82",
           232 => x"81",
           233 => x"82",
           234 => x"83",
           235 => x"82",
           236 => x"81",
           237 => x"82",
           238 => x"83",
           239 => x"82",
           240 => x"81",
           241 => x"82",
           242 => x"83",
           243 => x"82",
           244 => x"81",
           245 => x"82",
           246 => x"83",
           247 => x"82",
           248 => x"81",
           249 => x"82",
           250 => x"83",
           251 => x"82",
           252 => x"81",
           253 => x"82",
           254 => x"83",
           255 => x"82",
           256 => x"81",
           257 => x"82",
           258 => x"83",
           259 => x"82",
           260 => x"81",
           261 => x"82",
           262 => x"83",
           263 => x"82",
           264 => x"81",
           265 => x"82",
           266 => x"83",
           267 => x"82",
           268 => x"81",
           269 => x"82",
           270 => x"83",
           271 => x"82",
           272 => x"81",
           273 => x"82",
           274 => x"83",
           275 => x"82",
           276 => x"81",
           277 => x"82",
           278 => x"83",
           279 => x"82",
           280 => x"81",
           281 => x"82",
           282 => x"83",
           283 => x"82",
           284 => x"81",
           285 => x"82",
           286 => x"83",
           287 => x"82",
           288 => x"81",
           289 => x"82",
           290 => x"83",
           291 => x"82",
           292 => x"81",
           293 => x"82",
           294 => x"83",
           295 => x"82",
           296 => x"81",
           297 => x"82",
           298 => x"83",
           299 => x"82",
           300 => x"81",
           301 => x"82",
           302 => x"83",
           303 => x"82",
           304 => x"81",
           305 => x"82",
           306 => x"83",
           307 => x"82",
           308 => x"80",
           309 => x"82",
           310 => x"83",
           311 => x"82",
           312 => x"80",
           313 => x"82",
           314 => x"83",
           315 => x"82",
           316 => x"80",
           317 => x"82",
           318 => x"83",
           319 => x"82",
           320 => x"b3",
           321 => x"8c",
           322 => x"80",
           323 => x"8c",
           324 => x"a5",
           325 => x"e8",
           326 => x"90",
           327 => x"e8",
           328 => x"2d",
           329 => x"08",
           330 => x"04",
           331 => x"0c",
           332 => x"2d",
           333 => x"08",
           334 => x"04",
           335 => x"70",
           336 => x"27",
           337 => x"71",
           338 => x"53",
           339 => x"0b",
           340 => x"a4",
           341 => x"ef",
           342 => x"04",
           343 => x"08",
           344 => x"e8",
           345 => x"0d",
           346 => x"8c",
           347 => x"05",
           348 => x"8c",
           349 => x"05",
           350 => x"c5",
           351 => x"dc",
           352 => x"8c",
           353 => x"85",
           354 => x"8c",
           355 => x"82",
           356 => x"02",
           357 => x"0c",
           358 => x"81",
           359 => x"e8",
           360 => x"08",
           361 => x"e8",
           362 => x"08",
           363 => x"82",
           364 => x"70",
           365 => x"0c",
           366 => x"0d",
           367 => x"0c",
           368 => x"e8",
           369 => x"8c",
           370 => x"3d",
           371 => x"82",
           372 => x"fc",
           373 => x"0b",
           374 => x"08",
           375 => x"82",
           376 => x"8c",
           377 => x"8c",
           378 => x"05",
           379 => x"38",
           380 => x"08",
           381 => x"80",
           382 => x"80",
           383 => x"e8",
           384 => x"08",
           385 => x"82",
           386 => x"8c",
           387 => x"82",
           388 => x"8c",
           389 => x"8c",
           390 => x"05",
           391 => x"8c",
           392 => x"05",
           393 => x"39",
           394 => x"08",
           395 => x"80",
           396 => x"38",
           397 => x"08",
           398 => x"82",
           399 => x"88",
           400 => x"ad",
           401 => x"e8",
           402 => x"08",
           403 => x"08",
           404 => x"31",
           405 => x"08",
           406 => x"82",
           407 => x"f8",
           408 => x"8c",
           409 => x"05",
           410 => x"8c",
           411 => x"05",
           412 => x"e8",
           413 => x"08",
           414 => x"8c",
           415 => x"05",
           416 => x"e8",
           417 => x"08",
           418 => x"8c",
           419 => x"05",
           420 => x"39",
           421 => x"08",
           422 => x"80",
           423 => x"82",
           424 => x"88",
           425 => x"82",
           426 => x"f4",
           427 => x"91",
           428 => x"e8",
           429 => x"08",
           430 => x"e8",
           431 => x"0c",
           432 => x"e8",
           433 => x"08",
           434 => x"0c",
           435 => x"82",
           436 => x"04",
           437 => x"76",
           438 => x"55",
           439 => x"8f",
           440 => x"38",
           441 => x"83",
           442 => x"80",
           443 => x"ff",
           444 => x"ff",
           445 => x"72",
           446 => x"54",
           447 => x"81",
           448 => x"ff",
           449 => x"ff",
           450 => x"06",
           451 => x"82",
           452 => x"86",
           453 => x"74",
           454 => x"84",
           455 => x"71",
           456 => x"53",
           457 => x"84",
           458 => x"71",
           459 => x"53",
           460 => x"84",
           461 => x"71",
           462 => x"53",
           463 => x"84",
           464 => x"71",
           465 => x"53",
           466 => x"52",
           467 => x"c9",
           468 => x"27",
           469 => x"70",
           470 => x"08",
           471 => x"05",
           472 => x"12",
           473 => x"26",
           474 => x"54",
           475 => x"fc",
           476 => x"79",
           477 => x"05",
           478 => x"57",
           479 => x"83",
           480 => x"38",
           481 => x"51",
           482 => x"a4",
           483 => x"52",
           484 => x"93",
           485 => x"70",
           486 => x"34",
           487 => x"71",
           488 => x"81",
           489 => x"74",
           490 => x"0c",
           491 => x"04",
           492 => x"2b",
           493 => x"71",
           494 => x"51",
           495 => x"72",
           496 => x"72",
           497 => x"05",
           498 => x"71",
           499 => x"53",
           500 => x"70",
           501 => x"0c",
           502 => x"84",
           503 => x"f0",
           504 => x"8f",
           505 => x"83",
           506 => x"38",
           507 => x"84",
           508 => x"fc",
           509 => x"83",
           510 => x"70",
           511 => x"39",
           512 => x"76",
           513 => x"73",
           514 => x"54",
           515 => x"70",
           516 => x"71",
           517 => x"09",
           518 => x"fd",
           519 => x"70",
           520 => x"81",
           521 => x"51",
           522 => x"70",
           523 => x"14",
           524 => x"84",
           525 => x"70",
           526 => x"70",
           527 => x"ff",
           528 => x"f8",
           529 => x"80",
           530 => x"53",
           531 => x"80",
           532 => x"73",
           533 => x"81",
           534 => x"51",
           535 => x"81",
           536 => x"70",
           537 => x"82",
           538 => x"86",
           539 => x"fd",
           540 => x"70",
           541 => x"53",
           542 => x"b8",
           543 => x"08",
           544 => x"fb",
           545 => x"06",
           546 => x"82",
           547 => x"51",
           548 => x"70",
           549 => x"13",
           550 => x"09",
           551 => x"ff",
           552 => x"f8",
           553 => x"80",
           554 => x"52",
           555 => x"2e",
           556 => x"52",
           557 => x"70",
           558 => x"38",
           559 => x"33",
           560 => x"f8",
           561 => x"31",
           562 => x"0c",
           563 => x"04",
           564 => x"78",
           565 => x"54",
           566 => x"72",
           567 => x"d9",
           568 => x"07",
           569 => x"70",
           570 => x"d6",
           571 => x"53",
           572 => x"b1",
           573 => x"74",
           574 => x"74",
           575 => x"81",
           576 => x"72",
           577 => x"89",
           578 => x"ff",
           579 => x"80",
           580 => x"38",
           581 => x"15",
           582 => x"55",
           583 => x"2e",
           584 => x"d1",
           585 => x"74",
           586 => x"70",
           587 => x"75",
           588 => x"71",
           589 => x"52",
           590 => x"8c",
           591 => x"3d",
           592 => x"74",
           593 => x"73",
           594 => x"71",
           595 => x"2e",
           596 => x"76",
           597 => x"95",
           598 => x"53",
           599 => x"b1",
           600 => x"70",
           601 => x"fd",
           602 => x"70",
           603 => x"81",
           604 => x"51",
           605 => x"38",
           606 => x"17",
           607 => x"73",
           608 => x"74",
           609 => x"2e",
           610 => x"76",
           611 => x"dd",
           612 => x"82",
           613 => x"88",
           614 => x"fe",
           615 => x"52",
           616 => x"88",
           617 => x"86",
           618 => x"dc",
           619 => x"06",
           620 => x"14",
           621 => x"80",
           622 => x"71",
           623 => x"0c",
           624 => x"04",
           625 => x"77",
           626 => x"53",
           627 => x"80",
           628 => x"38",
           629 => x"70",
           630 => x"81",
           631 => x"81",
           632 => x"39",
           633 => x"39",
           634 => x"80",
           635 => x"81",
           636 => x"55",
           637 => x"2e",
           638 => x"55",
           639 => x"84",
           640 => x"38",
           641 => x"06",
           642 => x"2e",
           643 => x"88",
           644 => x"70",
           645 => x"34",
           646 => x"71",
           647 => x"8c",
           648 => x"3d",
           649 => x"3d",
           650 => x"72",
           651 => x"91",
           652 => x"fc",
           653 => x"51",
           654 => x"82",
           655 => x"85",
           656 => x"83",
           657 => x"72",
           658 => x"0c",
           659 => x"04",
           660 => x"76",
           661 => x"ff",
           662 => x"81",
           663 => x"26",
           664 => x"83",
           665 => x"05",
           666 => x"70",
           667 => x"8a",
           668 => x"33",
           669 => x"70",
           670 => x"fe",
           671 => x"33",
           672 => x"70",
           673 => x"f2",
           674 => x"33",
           675 => x"70",
           676 => x"e6",
           677 => x"22",
           678 => x"74",
           679 => x"80",
           680 => x"13",
           681 => x"52",
           682 => x"26",
           683 => x"81",
           684 => x"98",
           685 => x"22",
           686 => x"bc",
           687 => x"33",
           688 => x"b8",
           689 => x"33",
           690 => x"b4",
           691 => x"33",
           692 => x"b0",
           693 => x"33",
           694 => x"ac",
           695 => x"33",
           696 => x"a8",
           697 => x"c0",
           698 => x"73",
           699 => x"a0",
           700 => x"87",
           701 => x"0c",
           702 => x"82",
           703 => x"86",
           704 => x"f3",
           705 => x"5b",
           706 => x"9c",
           707 => x"0c",
           708 => x"bc",
           709 => x"7b",
           710 => x"98",
           711 => x"79",
           712 => x"87",
           713 => x"08",
           714 => x"1c",
           715 => x"98",
           716 => x"79",
           717 => x"87",
           718 => x"08",
           719 => x"1c",
           720 => x"98",
           721 => x"79",
           722 => x"87",
           723 => x"08",
           724 => x"1c",
           725 => x"98",
           726 => x"79",
           727 => x"80",
           728 => x"83",
           729 => x"59",
           730 => x"ff",
           731 => x"1b",
           732 => x"1b",
           733 => x"1b",
           734 => x"1b",
           735 => x"1b",
           736 => x"83",
           737 => x"52",
           738 => x"51",
           739 => x"8f",
           740 => x"ff",
           741 => x"8f",
           742 => x"30",
           743 => x"51",
           744 => x"0b",
           745 => x"d4",
           746 => x"0d",
           747 => x"0d",
           748 => x"82",
           749 => x"70",
           750 => x"57",
           751 => x"c0",
           752 => x"74",
           753 => x"38",
           754 => x"94",
           755 => x"70",
           756 => x"81",
           757 => x"52",
           758 => x"8c",
           759 => x"2a",
           760 => x"51",
           761 => x"38",
           762 => x"70",
           763 => x"51",
           764 => x"8d",
           765 => x"2a",
           766 => x"51",
           767 => x"be",
           768 => x"ff",
           769 => x"c0",
           770 => x"70",
           771 => x"38",
           772 => x"90",
           773 => x"0c",
           774 => x"dc",
           775 => x"0d",
           776 => x"0d",
           777 => x"33",
           778 => x"87",
           779 => x"81",
           780 => x"55",
           781 => x"94",
           782 => x"80",
           783 => x"87",
           784 => x"51",
           785 => x"96",
           786 => x"06",
           787 => x"70",
           788 => x"38",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"81",
           793 => x"70",
           794 => x"38",
           795 => x"70",
           796 => x"51",
           797 => x"38",
           798 => x"06",
           799 => x"94",
           800 => x"80",
           801 => x"87",
           802 => x"52",
           803 => x"87",
           804 => x"f9",
           805 => x"54",
           806 => x"70",
           807 => x"53",
           808 => x"77",
           809 => x"38",
           810 => x"06",
           811 => x"0b",
           812 => x"33",
           813 => x"06",
           814 => x"58",
           815 => x"84",
           816 => x"2e",
           817 => x"c0",
           818 => x"70",
           819 => x"2a",
           820 => x"53",
           821 => x"80",
           822 => x"71",
           823 => x"81",
           824 => x"70",
           825 => x"81",
           826 => x"06",
           827 => x"80",
           828 => x"71",
           829 => x"81",
           830 => x"70",
           831 => x"74",
           832 => x"51",
           833 => x"80",
           834 => x"2e",
           835 => x"c0",
           836 => x"77",
           837 => x"17",
           838 => x"81",
           839 => x"53",
           840 => x"84",
           841 => x"8c",
           842 => x"3d",
           843 => x"3d",
           844 => x"82",
           845 => x"70",
           846 => x"54",
           847 => x"94",
           848 => x"80",
           849 => x"87",
           850 => x"51",
           851 => x"82",
           852 => x"06",
           853 => x"70",
           854 => x"38",
           855 => x"06",
           856 => x"94",
           857 => x"80",
           858 => x"87",
           859 => x"52",
           860 => x"81",
           861 => x"8c",
           862 => x"84",
           863 => x"fe",
           864 => x"0b",
           865 => x"33",
           866 => x"06",
           867 => x"c0",
           868 => x"70",
           869 => x"38",
           870 => x"94",
           871 => x"70",
           872 => x"81",
           873 => x"51",
           874 => x"80",
           875 => x"72",
           876 => x"51",
           877 => x"80",
           878 => x"2e",
           879 => x"c0",
           880 => x"71",
           881 => x"2b",
           882 => x"51",
           883 => x"82",
           884 => x"84",
           885 => x"ff",
           886 => x"c0",
           887 => x"70",
           888 => x"06",
           889 => x"80",
           890 => x"38",
           891 => x"a4",
           892 => x"d8",
           893 => x"9e",
           894 => x"87",
           895 => x"c0",
           896 => x"82",
           897 => x"87",
           898 => x"08",
           899 => x"0c",
           900 => x"9c",
           901 => x"e8",
           902 => x"9e",
           903 => x"87",
           904 => x"c0",
           905 => x"82",
           906 => x"87",
           907 => x"08",
           908 => x"0c",
           909 => x"b4",
           910 => x"f8",
           911 => x"9e",
           912 => x"87",
           913 => x"c0",
           914 => x"82",
           915 => x"87",
           916 => x"08",
           917 => x"0c",
           918 => x"c4",
           919 => x"88",
           920 => x"9e",
           921 => x"70",
           922 => x"23",
           923 => x"84",
           924 => x"90",
           925 => x"9e",
           926 => x"88",
           927 => x"c0",
           928 => x"82",
           929 => x"81",
           930 => x"9c",
           931 => x"87",
           932 => x"08",
           933 => x"0a",
           934 => x"52",
           935 => x"83",
           936 => x"71",
           937 => x"34",
           938 => x"c0",
           939 => x"70",
           940 => x"06",
           941 => x"70",
           942 => x"38",
           943 => x"82",
           944 => x"80",
           945 => x"9e",
           946 => x"90",
           947 => x"51",
           948 => x"80",
           949 => x"81",
           950 => x"88",
           951 => x"0b",
           952 => x"90",
           953 => x"80",
           954 => x"52",
           955 => x"2e",
           956 => x"52",
           957 => x"a0",
           958 => x"87",
           959 => x"08",
           960 => x"80",
           961 => x"52",
           962 => x"83",
           963 => x"71",
           964 => x"34",
           965 => x"c0",
           966 => x"70",
           967 => x"06",
           968 => x"70",
           969 => x"38",
           970 => x"82",
           971 => x"80",
           972 => x"9e",
           973 => x"84",
           974 => x"51",
           975 => x"80",
           976 => x"81",
           977 => x"88",
           978 => x"0b",
           979 => x"90",
           980 => x"80",
           981 => x"52",
           982 => x"2e",
           983 => x"52",
           984 => x"a4",
           985 => x"87",
           986 => x"08",
           987 => x"80",
           988 => x"52",
           989 => x"83",
           990 => x"71",
           991 => x"34",
           992 => x"c0",
           993 => x"70",
           994 => x"06",
           995 => x"70",
           996 => x"38",
           997 => x"82",
           998 => x"80",
           999 => x"9e",
          1000 => x"a0",
          1001 => x"52",
          1002 => x"2e",
          1003 => x"52",
          1004 => x"a7",
          1005 => x"9e",
          1006 => x"98",
          1007 => x"8a",
          1008 => x"51",
          1009 => x"a8",
          1010 => x"87",
          1011 => x"08",
          1012 => x"06",
          1013 => x"70",
          1014 => x"38",
          1015 => x"82",
          1016 => x"87",
          1017 => x"08",
          1018 => x"06",
          1019 => x"51",
          1020 => x"82",
          1021 => x"80",
          1022 => x"9e",
          1023 => x"88",
          1024 => x"52",
          1025 => x"83",
          1026 => x"71",
          1027 => x"34",
          1028 => x"90",
          1029 => x"06",
          1030 => x"82",
          1031 => x"83",
          1032 => x"fb",
          1033 => x"f1",
          1034 => x"dc",
          1035 => x"9c",
          1036 => x"80",
          1037 => x"81",
          1038 => x"89",
          1039 => x"f2",
          1040 => x"c4",
          1041 => x"9e",
          1042 => x"80",
          1043 => x"82",
          1044 => x"82",
          1045 => x"11",
          1046 => x"f2",
          1047 => x"8c",
          1048 => x"a3",
          1049 => x"80",
          1050 => x"82",
          1051 => x"82",
          1052 => x"11",
          1053 => x"f2",
          1054 => x"f0",
          1055 => x"a0",
          1056 => x"80",
          1057 => x"82",
          1058 => x"82",
          1059 => x"11",
          1060 => x"f2",
          1061 => x"d4",
          1062 => x"a1",
          1063 => x"80",
          1064 => x"82",
          1065 => x"82",
          1066 => x"11",
          1067 => x"f3",
          1068 => x"b8",
          1069 => x"a2",
          1070 => x"80",
          1071 => x"82",
          1072 => x"82",
          1073 => x"11",
          1074 => x"f3",
          1075 => x"9c",
          1076 => x"a7",
          1077 => x"80",
          1078 => x"82",
          1079 => x"52",
          1080 => x"51",
          1081 => x"82",
          1082 => x"54",
          1083 => x"8d",
          1084 => x"ac",
          1085 => x"f3",
          1086 => x"f0",
          1087 => x"a9",
          1088 => x"80",
          1089 => x"82",
          1090 => x"52",
          1091 => x"51",
          1092 => x"82",
          1093 => x"54",
          1094 => x"88",
          1095 => x"a8",
          1096 => x"3f",
          1097 => x"33",
          1098 => x"2e",
          1099 => x"f4",
          1100 => x"d4",
          1101 => x"a4",
          1102 => x"80",
          1103 => x"81",
          1104 => x"87",
          1105 => x"88",
          1106 => x"73",
          1107 => x"38",
          1108 => x"51",
          1109 => x"82",
          1110 => x"54",
          1111 => x"88",
          1112 => x"e0",
          1113 => x"3f",
          1114 => x"51",
          1115 => x"82",
          1116 => x"52",
          1117 => x"51",
          1118 => x"82",
          1119 => x"52",
          1120 => x"51",
          1121 => x"82",
          1122 => x"52",
          1123 => x"51",
          1124 => x"81",
          1125 => x"86",
          1126 => x"88",
          1127 => x"81",
          1128 => x"8c",
          1129 => x"88",
          1130 => x"bd",
          1131 => x"75",
          1132 => x"3f",
          1133 => x"08",
          1134 => x"29",
          1135 => x"54",
          1136 => x"dc",
          1137 => x"f6",
          1138 => x"a0",
          1139 => x"a3",
          1140 => x"80",
          1141 => x"82",
          1142 => x"56",
          1143 => x"52",
          1144 => x"f8",
          1145 => x"dc",
          1146 => x"c0",
          1147 => x"31",
          1148 => x"8c",
          1149 => x"81",
          1150 => x"8b",
          1151 => x"88",
          1152 => x"73",
          1153 => x"38",
          1154 => x"08",
          1155 => x"c0",
          1156 => x"e6",
          1157 => x"8c",
          1158 => x"84",
          1159 => x"71",
          1160 => x"82",
          1161 => x"52",
          1162 => x"51",
          1163 => x"82",
          1164 => x"85",
          1165 => x"3d",
          1166 => x"3d",
          1167 => x"05",
          1168 => x"52",
          1169 => x"ac",
          1170 => x"29",
          1171 => x"f0",
          1172 => x"71",
          1173 => x"f7",
          1174 => x"39",
          1175 => x"51",
          1176 => x"f7",
          1177 => x"39",
          1178 => x"51",
          1179 => x"f7",
          1180 => x"39",
          1181 => x"51",
          1182 => x"84",
          1183 => x"71",
          1184 => x"04",
          1185 => x"c0",
          1186 => x"04",
          1187 => x"08",
          1188 => x"84",
          1189 => x"3d",
          1190 => x"ec",
          1191 => x"82",
          1192 => x"82",
          1193 => x"82",
          1194 => x"75",
          1195 => x"ff",
          1196 => x"b7",
          1197 => x"38",
          1198 => x"ec",
          1199 => x"72",
          1200 => x"0c",
          1201 => x"04",
          1202 => x"79",
          1203 => x"08",
          1204 => x"14",
          1205 => x"08",
          1206 => x"5a",
          1207 => x"57",
          1208 => x"26",
          1209 => x"13",
          1210 => x"53",
          1211 => x"0c",
          1212 => x"84",
          1213 => x"73",
          1214 => x"14",
          1215 => x"12",
          1216 => x"12",
          1217 => x"13",
          1218 => x"14",
          1219 => x"12",
          1220 => x"12",
          1221 => x"15",
          1222 => x"16",
          1223 => x"80",
          1224 => x"90",
          1225 => x"94",
          1226 => x"82",
          1227 => x"89",
          1228 => x"fc",
          1229 => x"8c",
          1230 => x"12",
          1231 => x"53",
          1232 => x"2e",
          1233 => x"a3",
          1234 => x"08",
          1235 => x"55",
          1236 => x"09",
          1237 => x"38",
          1238 => x"15",
          1239 => x"73",
          1240 => x"71",
          1241 => x"71",
          1242 => x"81",
          1243 => x"88",
          1244 => x"14",
          1245 => x"b4",
          1246 => x"0c",
          1247 => x"c4",
          1248 => x"08",
          1249 => x"0c",
          1250 => x"81",
          1251 => x"06",
          1252 => x"13",
          1253 => x"52",
          1254 => x"2e",
          1255 => x"a4",
          1256 => x"08",
          1257 => x"0c",
          1258 => x"90",
          1259 => x"90",
          1260 => x"94",
          1261 => x"14",
          1262 => x"08",
          1263 => x"0c",
          1264 => x"0c",
          1265 => x"dc",
          1266 => x"0d",
          1267 => x"0d",
          1268 => x"57",
          1269 => x"81",
          1270 => x"17",
          1271 => x"88",
          1272 => x"57",
          1273 => x"2e",
          1274 => x"16",
          1275 => x"80",
          1276 => x"16",
          1277 => x"39",
          1278 => x"17",
          1279 => x"06",
          1280 => x"fd",
          1281 => x"8c",
          1282 => x"8c",
          1283 => x"70",
          1284 => x"08",
          1285 => x"82",
          1286 => x"09",
          1287 => x"72",
          1288 => x"73",
          1289 => x"58",
          1290 => x"80",
          1291 => x"2e",
          1292 => x"80",
          1293 => x"39",
          1294 => x"51",
          1295 => x"81",
          1296 => x"dc",
          1297 => x"82",
          1298 => x"84",
          1299 => x"88",
          1300 => x"72",
          1301 => x"8c",
          1302 => x"26",
          1303 => x"13",
          1304 => x"39",
          1305 => x"88",
          1306 => x"8c",
          1307 => x"88",
          1308 => x"16",
          1309 => x"12",
          1310 => x"51",
          1311 => x"76",
          1312 => x"dc",
          1313 => x"c0",
          1314 => x"dc",
          1315 => x"82",
          1316 => x"89",
          1317 => x"ff",
          1318 => x"52",
          1319 => x"87",
          1320 => x"51",
          1321 => x"83",
          1322 => x"fe",
          1323 => x"93",
          1324 => x"72",
          1325 => x"81",
          1326 => x"8d",
          1327 => x"82",
          1328 => x"52",
          1329 => x"90",
          1330 => x"34",
          1331 => x"08",
          1332 => x"8c",
          1333 => x"39",
          1334 => x"08",
          1335 => x"2e",
          1336 => x"51",
          1337 => x"3d",
          1338 => x"3d",
          1339 => x"05",
          1340 => x"f0",
          1341 => x"8c",
          1342 => x"51",
          1343 => x"72",
          1344 => x"0c",
          1345 => x"04",
          1346 => x"75",
          1347 => x"70",
          1348 => x"53",
          1349 => x"2e",
          1350 => x"81",
          1351 => x"81",
          1352 => x"87",
          1353 => x"85",
          1354 => x"fc",
          1355 => x"82",
          1356 => x"78",
          1357 => x"0c",
          1358 => x"33",
          1359 => x"06",
          1360 => x"80",
          1361 => x"72",
          1362 => x"51",
          1363 => x"fe",
          1364 => x"39",
          1365 => x"f0",
          1366 => x"0d",
          1367 => x"0d",
          1368 => x"59",
          1369 => x"05",
          1370 => x"75",
          1371 => x"f8",
          1372 => x"2e",
          1373 => x"82",
          1374 => x"70",
          1375 => x"05",
          1376 => x"5b",
          1377 => x"2e",
          1378 => x"85",
          1379 => x"8b",
          1380 => x"2e",
          1381 => x"8a",
          1382 => x"78",
          1383 => x"5a",
          1384 => x"aa",
          1385 => x"06",
          1386 => x"84",
          1387 => x"7b",
          1388 => x"5d",
          1389 => x"59",
          1390 => x"d0",
          1391 => x"89",
          1392 => x"7a",
          1393 => x"10",
          1394 => x"d0",
          1395 => x"81",
          1396 => x"57",
          1397 => x"75",
          1398 => x"70",
          1399 => x"07",
          1400 => x"80",
          1401 => x"30",
          1402 => x"80",
          1403 => x"53",
          1404 => x"55",
          1405 => x"2e",
          1406 => x"84",
          1407 => x"81",
          1408 => x"57",
          1409 => x"2e",
          1410 => x"75",
          1411 => x"76",
          1412 => x"e0",
          1413 => x"ff",
          1414 => x"73",
          1415 => x"81",
          1416 => x"80",
          1417 => x"38",
          1418 => x"2e",
          1419 => x"73",
          1420 => x"8b",
          1421 => x"c2",
          1422 => x"38",
          1423 => x"73",
          1424 => x"81",
          1425 => x"8f",
          1426 => x"d5",
          1427 => x"38",
          1428 => x"24",
          1429 => x"80",
          1430 => x"38",
          1431 => x"73",
          1432 => x"80",
          1433 => x"ef",
          1434 => x"19",
          1435 => x"59",
          1436 => x"33",
          1437 => x"75",
          1438 => x"81",
          1439 => x"70",
          1440 => x"55",
          1441 => x"79",
          1442 => x"90",
          1443 => x"16",
          1444 => x"7b",
          1445 => x"a0",
          1446 => x"3f",
          1447 => x"53",
          1448 => x"e9",
          1449 => x"fc",
          1450 => x"81",
          1451 => x"72",
          1452 => x"b0",
          1453 => x"fb",
          1454 => x"39",
          1455 => x"83",
          1456 => x"59",
          1457 => x"82",
          1458 => x"88",
          1459 => x"8a",
          1460 => x"90",
          1461 => x"75",
          1462 => x"3f",
          1463 => x"79",
          1464 => x"81",
          1465 => x"72",
          1466 => x"38",
          1467 => x"59",
          1468 => x"84",
          1469 => x"58",
          1470 => x"80",
          1471 => x"30",
          1472 => x"80",
          1473 => x"55",
          1474 => x"25",
          1475 => x"80",
          1476 => x"74",
          1477 => x"07",
          1478 => x"0b",
          1479 => x"57",
          1480 => x"51",
          1481 => x"82",
          1482 => x"81",
          1483 => x"53",
          1484 => x"dc",
          1485 => x"8c",
          1486 => x"89",
          1487 => x"38",
          1488 => x"75",
          1489 => x"84",
          1490 => x"53",
          1491 => x"06",
          1492 => x"53",
          1493 => x"81",
          1494 => x"81",
          1495 => x"70",
          1496 => x"2a",
          1497 => x"76",
          1498 => x"38",
          1499 => x"38",
          1500 => x"70",
          1501 => x"53",
          1502 => x"8e",
          1503 => x"77",
          1504 => x"53",
          1505 => x"81",
          1506 => x"7a",
          1507 => x"55",
          1508 => x"83",
          1509 => x"79",
          1510 => x"81",
          1511 => x"72",
          1512 => x"17",
          1513 => x"27",
          1514 => x"51",
          1515 => x"75",
          1516 => x"72",
          1517 => x"81",
          1518 => x"7a",
          1519 => x"38",
          1520 => x"05",
          1521 => x"ff",
          1522 => x"70",
          1523 => x"57",
          1524 => x"76",
          1525 => x"81",
          1526 => x"72",
          1527 => x"84",
          1528 => x"f9",
          1529 => x"39",
          1530 => x"04",
          1531 => x"86",
          1532 => x"84",
          1533 => x"55",
          1534 => x"fa",
          1535 => x"3d",
          1536 => x"3d",
          1537 => x"8c",
          1538 => x"3d",
          1539 => x"75",
          1540 => x"3f",
          1541 => x"08",
          1542 => x"34",
          1543 => x"8c",
          1544 => x"3d",
          1545 => x"3d",
          1546 => x"f0",
          1547 => x"8c",
          1548 => x"3d",
          1549 => x"77",
          1550 => x"a1",
          1551 => x"8c",
          1552 => x"3d",
          1553 => x"3d",
          1554 => x"82",
          1555 => x"70",
          1556 => x"55",
          1557 => x"80",
          1558 => x"38",
          1559 => x"08",
          1560 => x"82",
          1561 => x"81",
          1562 => x"72",
          1563 => x"cb",
          1564 => x"2e",
          1565 => x"88",
          1566 => x"70",
          1567 => x"51",
          1568 => x"2e",
          1569 => x"80",
          1570 => x"ff",
          1571 => x"39",
          1572 => x"c8",
          1573 => x"52",
          1574 => x"c0",
          1575 => x"52",
          1576 => x"81",
          1577 => x"51",
          1578 => x"ff",
          1579 => x"15",
          1580 => x"34",
          1581 => x"f3",
          1582 => x"72",
          1583 => x"0c",
          1584 => x"04",
          1585 => x"82",
          1586 => x"75",
          1587 => x"0c",
          1588 => x"52",
          1589 => x"3f",
          1590 => x"f4",
          1591 => x"0d",
          1592 => x"0d",
          1593 => x"56",
          1594 => x"0c",
          1595 => x"70",
          1596 => x"73",
          1597 => x"81",
          1598 => x"81",
          1599 => x"ed",
          1600 => x"2e",
          1601 => x"8e",
          1602 => x"08",
          1603 => x"76",
          1604 => x"56",
          1605 => x"b0",
          1606 => x"06",
          1607 => x"75",
          1608 => x"76",
          1609 => x"70",
          1610 => x"73",
          1611 => x"8b",
          1612 => x"73",
          1613 => x"85",
          1614 => x"82",
          1615 => x"76",
          1616 => x"70",
          1617 => x"ac",
          1618 => x"a0",
          1619 => x"fa",
          1620 => x"53",
          1621 => x"57",
          1622 => x"98",
          1623 => x"39",
          1624 => x"80",
          1625 => x"26",
          1626 => x"86",
          1627 => x"80",
          1628 => x"57",
          1629 => x"74",
          1630 => x"38",
          1631 => x"27",
          1632 => x"14",
          1633 => x"06",
          1634 => x"14",
          1635 => x"06",
          1636 => x"74",
          1637 => x"f9",
          1638 => x"ff",
          1639 => x"89",
          1640 => x"38",
          1641 => x"c5",
          1642 => x"29",
          1643 => x"81",
          1644 => x"76",
          1645 => x"56",
          1646 => x"ba",
          1647 => x"2e",
          1648 => x"30",
          1649 => x"0c",
          1650 => x"82",
          1651 => x"8a",
          1652 => x"f8",
          1653 => x"7c",
          1654 => x"70",
          1655 => x"75",
          1656 => x"55",
          1657 => x"2e",
          1658 => x"87",
          1659 => x"76",
          1660 => x"73",
          1661 => x"81",
          1662 => x"81",
          1663 => x"77",
          1664 => x"70",
          1665 => x"58",
          1666 => x"09",
          1667 => x"c2",
          1668 => x"81",
          1669 => x"75",
          1670 => x"55",
          1671 => x"e2",
          1672 => x"90",
          1673 => x"f8",
          1674 => x"8f",
          1675 => x"81",
          1676 => x"75",
          1677 => x"55",
          1678 => x"81",
          1679 => x"27",
          1680 => x"d0",
          1681 => x"55",
          1682 => x"73",
          1683 => x"80",
          1684 => x"14",
          1685 => x"72",
          1686 => x"e0",
          1687 => x"80",
          1688 => x"39",
          1689 => x"55",
          1690 => x"80",
          1691 => x"e0",
          1692 => x"38",
          1693 => x"81",
          1694 => x"53",
          1695 => x"81",
          1696 => x"53",
          1697 => x"8e",
          1698 => x"70",
          1699 => x"55",
          1700 => x"27",
          1701 => x"77",
          1702 => x"74",
          1703 => x"76",
          1704 => x"77",
          1705 => x"70",
          1706 => x"55",
          1707 => x"77",
          1708 => x"38",
          1709 => x"74",
          1710 => x"55",
          1711 => x"dc",
          1712 => x"0d",
          1713 => x"0d",
          1714 => x"70",
          1715 => x"98",
          1716 => x"2c",
          1717 => x"70",
          1718 => x"53",
          1719 => x"51",
          1720 => x"f8",
          1721 => x"55",
          1722 => x"25",
          1723 => x"f8",
          1724 => x"12",
          1725 => x"97",
          1726 => x"33",
          1727 => x"70",
          1728 => x"81",
          1729 => x"81",
          1730 => x"8c",
          1731 => x"3d",
          1732 => x"3d",
          1733 => x"84",
          1734 => x"33",
          1735 => x"55",
          1736 => x"2e",
          1737 => x"51",
          1738 => x"a0",
          1739 => x"3f",
          1740 => x"f7",
          1741 => x"ff",
          1742 => x"73",
          1743 => x"ff",
          1744 => x"39",
          1745 => x"c0",
          1746 => x"34",
          1747 => x"04",
          1748 => x"7c",
          1749 => x"b7",
          1750 => x"88",
          1751 => x"33",
          1752 => x"33",
          1753 => x"82",
          1754 => x"70",
          1755 => x"59",
          1756 => x"74",
          1757 => x"38",
          1758 => x"9b",
          1759 => x"a8",
          1760 => x"29",
          1761 => x"05",
          1762 => x"54",
          1763 => x"f0",
          1764 => x"8c",
          1765 => x"0c",
          1766 => x"33",
          1767 => x"82",
          1768 => x"70",
          1769 => x"5a",
          1770 => x"a6",
          1771 => x"78",
          1772 => x"d6",
          1773 => x"89",
          1774 => x"05",
          1775 => x"89",
          1776 => x"81",
          1777 => x"93",
          1778 => x"38",
          1779 => x"89",
          1780 => x"80",
          1781 => x"82",
          1782 => x"56",
          1783 => x"ac",
          1784 => x"a0",
          1785 => x"a4",
          1786 => x"fc",
          1787 => x"53",
          1788 => x"51",
          1789 => x"3f",
          1790 => x"08",
          1791 => x"80",
          1792 => x"82",
          1793 => x"51",
          1794 => x"3f",
          1795 => x"04",
          1796 => x"81",
          1797 => x"82",
          1798 => x"51",
          1799 => x"3f",
          1800 => x"08",
          1801 => x"82",
          1802 => x"53",
          1803 => x"88",
          1804 => x"56",
          1805 => x"3f",
          1806 => x"08",
          1807 => x"38",
          1808 => x"ab",
          1809 => x"dc",
          1810 => x"0b",
          1811 => x"08",
          1812 => x"82",
          1813 => x"ff",
          1814 => x"55",
          1815 => x"34",
          1816 => x"52",
          1817 => x"f7",
          1818 => x"f6",
          1819 => x"ff",
          1820 => x"06",
          1821 => x"a6",
          1822 => x"d9",
          1823 => x"3d",
          1824 => x"08",
          1825 => x"70",
          1826 => x"52",
          1827 => x"08",
          1828 => x"92",
          1829 => x"dc",
          1830 => x"38",
          1831 => x"89",
          1832 => x"55",
          1833 => x"8b",
          1834 => x"56",
          1835 => x"3f",
          1836 => x"08",
          1837 => x"38",
          1838 => x"b3",
          1839 => x"dc",
          1840 => x"58",
          1841 => x"82",
          1842 => x"25",
          1843 => x"8c",
          1844 => x"05",
          1845 => x"55",
          1846 => x"74",
          1847 => x"70",
          1848 => x"2a",
          1849 => x"78",
          1850 => x"38",
          1851 => x"38",
          1852 => x"08",
          1853 => x"53",
          1854 => x"aa",
          1855 => x"dc",
          1856 => x"88",
          1857 => x"fc",
          1858 => x"3f",
          1859 => x"09",
          1860 => x"38",
          1861 => x"51",
          1862 => x"79",
          1863 => x"3f",
          1864 => x"54",
          1865 => x"08",
          1866 => x"58",
          1867 => x"dc",
          1868 => x"0d",
          1869 => x"0d",
          1870 => x"5c",
          1871 => x"57",
          1872 => x"73",
          1873 => x"81",
          1874 => x"78",
          1875 => x"56",
          1876 => x"98",
          1877 => x"70",
          1878 => x"33",
          1879 => x"73",
          1880 => x"81",
          1881 => x"75",
          1882 => x"38",
          1883 => x"88",
          1884 => x"ac",
          1885 => x"52",
          1886 => x"3f",
          1887 => x"08",
          1888 => x"74",
          1889 => x"c8",
          1890 => x"dc",
          1891 => x"38",
          1892 => x"55",
          1893 => x"88",
          1894 => x"2e",
          1895 => x"39",
          1896 => x"ab",
          1897 => x"5a",
          1898 => x"11",
          1899 => x"51",
          1900 => x"82",
          1901 => x"80",
          1902 => x"7a",
          1903 => x"77",
          1904 => x"3f",
          1905 => x"08",
          1906 => x"55",
          1907 => x"74",
          1908 => x"81",
          1909 => x"ff",
          1910 => x"82",
          1911 => x"8e",
          1912 => x"73",
          1913 => x"0c",
          1914 => x"04",
          1915 => x"b0",
          1916 => x"84",
          1917 => x"05",
          1918 => x"80",
          1919 => x"34",
          1920 => x"33",
          1921 => x"a4",
          1922 => x"38",
          1923 => x"33",
          1924 => x"9a",
          1925 => x"eb",
          1926 => x"8c",
          1927 => x"89",
          1928 => x"8c",
          1929 => x"2e",
          1930 => x"93",
          1931 => x"cc",
          1932 => x"8c",
          1933 => x"bb",
          1934 => x"8c",
          1935 => x"2e",
          1936 => x"f8",
          1937 => x"a4",
          1938 => x"39",
          1939 => x"08",
          1940 => x"52",
          1941 => x"52",
          1942 => x"b0",
          1943 => x"dc",
          1944 => x"8c",
          1945 => x"2e",
          1946 => x"80",
          1947 => x"8c",
          1948 => x"d3",
          1949 => x"8c",
          1950 => x"80",
          1951 => x"dc",
          1952 => x"38",
          1953 => x"08",
          1954 => x"17",
          1955 => x"74",
          1956 => x"74",
          1957 => x"52",
          1958 => x"b4",
          1959 => x"2e",
          1960 => x"ff",
          1961 => x"39",
          1962 => x"89",
          1963 => x"3d",
          1964 => x"3f",
          1965 => x"08",
          1966 => x"98",
          1967 => x"78",
          1968 => x"38",
          1969 => x"06",
          1970 => x"33",
          1971 => x"70",
          1972 => x"8c",
          1973 => x"98",
          1974 => x"2c",
          1975 => x"05",
          1976 => x"81",
          1977 => x"70",
          1978 => x"33",
          1979 => x"51",
          1980 => x"59",
          1981 => x"56",
          1982 => x"80",
          1983 => x"74",
          1984 => x"74",
          1985 => x"29",
          1986 => x"05",
          1987 => x"51",
          1988 => x"24",
          1989 => x"76",
          1990 => x"77",
          1991 => x"3f",
          1992 => x"08",
          1993 => x"54",
          1994 => x"d7",
          1995 => x"8c",
          1996 => x"56",
          1997 => x"81",
          1998 => x"81",
          1999 => x"70",
          2000 => x"81",
          2001 => x"51",
          2002 => x"26",
          2003 => x"53",
          2004 => x"51",
          2005 => x"82",
          2006 => x"81",
          2007 => x"73",
          2008 => x"39",
          2009 => x"80",
          2010 => x"38",
          2011 => x"74",
          2012 => x"34",
          2013 => x"70",
          2014 => x"8c",
          2015 => x"98",
          2016 => x"2c",
          2017 => x"70",
          2018 => x"f8",
          2019 => x"5e",
          2020 => x"57",
          2021 => x"74",
          2022 => x"81",
          2023 => x"38",
          2024 => x"14",
          2025 => x"80",
          2026 => x"80",
          2027 => x"82",
          2028 => x"92",
          2029 => x"8d",
          2030 => x"82",
          2031 => x"78",
          2032 => x"75",
          2033 => x"54",
          2034 => x"fd",
          2035 => x"84",
          2036 => x"e4",
          2037 => x"08",
          2038 => x"88",
          2039 => x"7e",
          2040 => x"38",
          2041 => x"33",
          2042 => x"27",
          2043 => x"98",
          2044 => x"2c",
          2045 => x"75",
          2046 => x"74",
          2047 => x"33",
          2048 => x"74",
          2049 => x"29",
          2050 => x"05",
          2051 => x"82",
          2052 => x"56",
          2053 => x"39",
          2054 => x"33",
          2055 => x"54",
          2056 => x"88",
          2057 => x"54",
          2058 => x"74",
          2059 => x"84",
          2060 => x"7e",
          2061 => x"81",
          2062 => x"82",
          2063 => x"82",
          2064 => x"70",
          2065 => x"29",
          2066 => x"05",
          2067 => x"82",
          2068 => x"5a",
          2069 => x"74",
          2070 => x"38",
          2071 => x"33",
          2072 => x"c7",
          2073 => x"80",
          2074 => x"80",
          2075 => x"98",
          2076 => x"84",
          2077 => x"55",
          2078 => x"e0",
          2079 => x"88",
          2080 => x"2b",
          2081 => x"82",
          2082 => x"5a",
          2083 => x"74",
          2084 => x"9a",
          2085 => x"e8",
          2086 => x"81",
          2087 => x"81",
          2088 => x"70",
          2089 => x"8d",
          2090 => x"51",
          2091 => x"24",
          2092 => x"fa",
          2093 => x"88",
          2094 => x"ff",
          2095 => x"73",
          2096 => x"ea",
          2097 => x"84",
          2098 => x"54",
          2099 => x"84",
          2100 => x"54",
          2101 => x"88",
          2102 => x"e7",
          2103 => x"8d",
          2104 => x"98",
          2105 => x"2c",
          2106 => x"33",
          2107 => x"57",
          2108 => x"a7",
          2109 => x"54",
          2110 => x"74",
          2111 => x"51",
          2112 => x"74",
          2113 => x"29",
          2114 => x"05",
          2115 => x"82",
          2116 => x"58",
          2117 => x"75",
          2118 => x"a0",
          2119 => x"3f",
          2120 => x"33",
          2121 => x"70",
          2122 => x"8d",
          2123 => x"51",
          2124 => x"74",
          2125 => x"38",
          2126 => x"ef",
          2127 => x"80",
          2128 => x"80",
          2129 => x"98",
          2130 => x"84",
          2131 => x"55",
          2132 => x"e4",
          2133 => x"39",
          2134 => x"33",
          2135 => x"80",
          2136 => x"51",
          2137 => x"82",
          2138 => x"79",
          2139 => x"3f",
          2140 => x"08",
          2141 => x"54",
          2142 => x"82",
          2143 => x"54",
          2144 => x"84",
          2145 => x"53",
          2146 => x"51",
          2147 => x"84",
          2148 => x"7a",
          2149 => x"39",
          2150 => x"33",
          2151 => x"2e",
          2152 => x"88",
          2153 => x"3f",
          2154 => x"33",
          2155 => x"73",
          2156 => x"34",
          2157 => x"06",
          2158 => x"82",
          2159 => x"82",
          2160 => x"55",
          2161 => x"2e",
          2162 => x"ff",
          2163 => x"82",
          2164 => x"74",
          2165 => x"98",
          2166 => x"ff",
          2167 => x"55",
          2168 => x"a7",
          2169 => x"54",
          2170 => x"74",
          2171 => x"51",
          2172 => x"74",
          2173 => x"29",
          2174 => x"05",
          2175 => x"82",
          2176 => x"58",
          2177 => x"75",
          2178 => x"a0",
          2179 => x"3f",
          2180 => x"33",
          2181 => x"70",
          2182 => x"8d",
          2183 => x"51",
          2184 => x"74",
          2185 => x"38",
          2186 => x"ff",
          2187 => x"80",
          2188 => x"80",
          2189 => x"98",
          2190 => x"84",
          2191 => x"55",
          2192 => x"e4",
          2193 => x"39",
          2194 => x"33",
          2195 => x"06",
          2196 => x"33",
          2197 => x"74",
          2198 => x"d2",
          2199 => x"54",
          2200 => x"88",
          2201 => x"70",
          2202 => x"e4",
          2203 => x"8d",
          2204 => x"81",
          2205 => x"8d",
          2206 => x"56",
          2207 => x"26",
          2208 => x"aa",
          2209 => x"38",
          2210 => x"08",
          2211 => x"2e",
          2212 => x"51",
          2213 => x"82",
          2214 => x"82",
          2215 => x"82",
          2216 => x"81",
          2217 => x"05",
          2218 => x"79",
          2219 => x"3f",
          2220 => x"c1",
          2221 => x"29",
          2222 => x"05",
          2223 => x"56",
          2224 => x"2e",
          2225 => x"51",
          2226 => x"82",
          2227 => x"82",
          2228 => x"82",
          2229 => x"81",
          2230 => x"05",
          2231 => x"79",
          2232 => x"3f",
          2233 => x"80",
          2234 => x"08",
          2235 => x"2e",
          2236 => x"74",
          2237 => x"3f",
          2238 => x"7a",
          2239 => x"81",
          2240 => x"82",
          2241 => x"55",
          2242 => x"89",
          2243 => x"ca",
          2244 => x"c8",
          2245 => x"29",
          2246 => x"05",
          2247 => x"56",
          2248 => x"2e",
          2249 => x"51",
          2250 => x"82",
          2251 => x"82",
          2252 => x"82",
          2253 => x"81",
          2254 => x"05",
          2255 => x"79",
          2256 => x"3f",
          2257 => x"73",
          2258 => x"5b",
          2259 => x"08",
          2260 => x"2e",
          2261 => x"74",
          2262 => x"3f",
          2263 => x"08",
          2264 => x"34",
          2265 => x"08",
          2266 => x"81",
          2267 => x"52",
          2268 => x"e0",
          2269 => x"88",
          2270 => x"84",
          2271 => x"51",
          2272 => x"f6",
          2273 => x"8d",
          2274 => x"81",
          2275 => x"8d",
          2276 => x"56",
          2277 => x"27",
          2278 => x"81",
          2279 => x"82",
          2280 => x"74",
          2281 => x"52",
          2282 => x"3f",
          2283 => x"82",
          2284 => x"54",
          2285 => x"f5",
          2286 => x"51",
          2287 => x"82",
          2288 => x"ff",
          2289 => x"82",
          2290 => x"f5",
          2291 => x"0b",
          2292 => x"34",
          2293 => x"8d",
          2294 => x"82",
          2295 => x"af",
          2296 => x"ff",
          2297 => x"8f",
          2298 => x"81",
          2299 => x"26",
          2300 => x"89",
          2301 => x"52",
          2302 => x"dc",
          2303 => x"0d",
          2304 => x"0d",
          2305 => x"33",
          2306 => x"9f",
          2307 => x"53",
          2308 => x"81",
          2309 => x"38",
          2310 => x"87",
          2311 => x"11",
          2312 => x"54",
          2313 => x"84",
          2314 => x"54",
          2315 => x"87",
          2316 => x"11",
          2317 => x"0c",
          2318 => x"c0",
          2319 => x"70",
          2320 => x"70",
          2321 => x"51",
          2322 => x"8a",
          2323 => x"98",
          2324 => x"70",
          2325 => x"08",
          2326 => x"06",
          2327 => x"38",
          2328 => x"8c",
          2329 => x"80",
          2330 => x"71",
          2331 => x"14",
          2332 => x"c4",
          2333 => x"70",
          2334 => x"0c",
          2335 => x"04",
          2336 => x"60",
          2337 => x"8c",
          2338 => x"33",
          2339 => x"5b",
          2340 => x"5a",
          2341 => x"82",
          2342 => x"81",
          2343 => x"52",
          2344 => x"38",
          2345 => x"84",
          2346 => x"92",
          2347 => x"c0",
          2348 => x"87",
          2349 => x"13",
          2350 => x"57",
          2351 => x"0b",
          2352 => x"8c",
          2353 => x"0c",
          2354 => x"75",
          2355 => x"2a",
          2356 => x"51",
          2357 => x"80",
          2358 => x"7b",
          2359 => x"7b",
          2360 => x"5d",
          2361 => x"59",
          2362 => x"06",
          2363 => x"73",
          2364 => x"81",
          2365 => x"ff",
          2366 => x"72",
          2367 => x"38",
          2368 => x"8c",
          2369 => x"c3",
          2370 => x"98",
          2371 => x"71",
          2372 => x"38",
          2373 => x"2e",
          2374 => x"76",
          2375 => x"92",
          2376 => x"72",
          2377 => x"06",
          2378 => x"f7",
          2379 => x"5a",
          2380 => x"80",
          2381 => x"70",
          2382 => x"5a",
          2383 => x"80",
          2384 => x"73",
          2385 => x"06",
          2386 => x"38",
          2387 => x"fe",
          2388 => x"fc",
          2389 => x"52",
          2390 => x"83",
          2391 => x"71",
          2392 => x"8c",
          2393 => x"3d",
          2394 => x"3d",
          2395 => x"64",
          2396 => x"bf",
          2397 => x"40",
          2398 => x"59",
          2399 => x"58",
          2400 => x"82",
          2401 => x"81",
          2402 => x"52",
          2403 => x"09",
          2404 => x"b1",
          2405 => x"84",
          2406 => x"92",
          2407 => x"c0",
          2408 => x"87",
          2409 => x"13",
          2410 => x"56",
          2411 => x"87",
          2412 => x"0c",
          2413 => x"82",
          2414 => x"58",
          2415 => x"84",
          2416 => x"06",
          2417 => x"71",
          2418 => x"38",
          2419 => x"05",
          2420 => x"0c",
          2421 => x"73",
          2422 => x"81",
          2423 => x"71",
          2424 => x"38",
          2425 => x"8c",
          2426 => x"d0",
          2427 => x"98",
          2428 => x"71",
          2429 => x"38",
          2430 => x"2e",
          2431 => x"76",
          2432 => x"92",
          2433 => x"72",
          2434 => x"06",
          2435 => x"f7",
          2436 => x"59",
          2437 => x"1a",
          2438 => x"06",
          2439 => x"59",
          2440 => x"80",
          2441 => x"73",
          2442 => x"06",
          2443 => x"38",
          2444 => x"fe",
          2445 => x"fc",
          2446 => x"52",
          2447 => x"83",
          2448 => x"71",
          2449 => x"8c",
          2450 => x"3d",
          2451 => x"3d",
          2452 => x"84",
          2453 => x"33",
          2454 => x"a7",
          2455 => x"54",
          2456 => x"fa",
          2457 => x"8c",
          2458 => x"06",
          2459 => x"72",
          2460 => x"85",
          2461 => x"98",
          2462 => x"56",
          2463 => x"80",
          2464 => x"76",
          2465 => x"74",
          2466 => x"c0",
          2467 => x"54",
          2468 => x"2e",
          2469 => x"d4",
          2470 => x"2e",
          2471 => x"80",
          2472 => x"08",
          2473 => x"70",
          2474 => x"51",
          2475 => x"2e",
          2476 => x"c0",
          2477 => x"52",
          2478 => x"87",
          2479 => x"08",
          2480 => x"38",
          2481 => x"87",
          2482 => x"14",
          2483 => x"70",
          2484 => x"52",
          2485 => x"96",
          2486 => x"92",
          2487 => x"0a",
          2488 => x"39",
          2489 => x"0c",
          2490 => x"39",
          2491 => x"54",
          2492 => x"dc",
          2493 => x"0d",
          2494 => x"0d",
          2495 => x"33",
          2496 => x"88",
          2497 => x"8c",
          2498 => x"51",
          2499 => x"04",
          2500 => x"75",
          2501 => x"82",
          2502 => x"90",
          2503 => x"2b",
          2504 => x"33",
          2505 => x"88",
          2506 => x"71",
          2507 => x"dc",
          2508 => x"54",
          2509 => x"85",
          2510 => x"ff",
          2511 => x"02",
          2512 => x"05",
          2513 => x"70",
          2514 => x"05",
          2515 => x"88",
          2516 => x"72",
          2517 => x"0d",
          2518 => x"0d",
          2519 => x"52",
          2520 => x"81",
          2521 => x"70",
          2522 => x"70",
          2523 => x"05",
          2524 => x"88",
          2525 => x"72",
          2526 => x"54",
          2527 => x"2a",
          2528 => x"34",
          2529 => x"04",
          2530 => x"76",
          2531 => x"54",
          2532 => x"2e",
          2533 => x"70",
          2534 => x"33",
          2535 => x"05",
          2536 => x"11",
          2537 => x"84",
          2538 => x"fe",
          2539 => x"77",
          2540 => x"53",
          2541 => x"81",
          2542 => x"ff",
          2543 => x"f4",
          2544 => x"0d",
          2545 => x"0d",
          2546 => x"56",
          2547 => x"70",
          2548 => x"33",
          2549 => x"05",
          2550 => x"71",
          2551 => x"56",
          2552 => x"72",
          2553 => x"38",
          2554 => x"e2",
          2555 => x"8c",
          2556 => x"3d",
          2557 => x"3d",
          2558 => x"54",
          2559 => x"71",
          2560 => x"38",
          2561 => x"70",
          2562 => x"f3",
          2563 => x"82",
          2564 => x"84",
          2565 => x"80",
          2566 => x"dc",
          2567 => x"0b",
          2568 => x"0c",
          2569 => x"0d",
          2570 => x"0b",
          2571 => x"56",
          2572 => x"2e",
          2573 => x"81",
          2574 => x"08",
          2575 => x"70",
          2576 => x"33",
          2577 => x"a2",
          2578 => x"dc",
          2579 => x"09",
          2580 => x"38",
          2581 => x"08",
          2582 => x"b0",
          2583 => x"a4",
          2584 => x"9c",
          2585 => x"56",
          2586 => x"27",
          2587 => x"16",
          2588 => x"82",
          2589 => x"06",
          2590 => x"54",
          2591 => x"78",
          2592 => x"33",
          2593 => x"3f",
          2594 => x"5a",
          2595 => x"dc",
          2596 => x"0d",
          2597 => x"0d",
          2598 => x"56",
          2599 => x"b0",
          2600 => x"af",
          2601 => x"fe",
          2602 => x"8c",
          2603 => x"82",
          2604 => x"9f",
          2605 => x"74",
          2606 => x"52",
          2607 => x"51",
          2608 => x"82",
          2609 => x"80",
          2610 => x"ff",
          2611 => x"74",
          2612 => x"76",
          2613 => x"0c",
          2614 => x"04",
          2615 => x"7a",
          2616 => x"fe",
          2617 => x"8c",
          2618 => x"82",
          2619 => x"81",
          2620 => x"33",
          2621 => x"2e",
          2622 => x"80",
          2623 => x"17",
          2624 => x"81",
          2625 => x"06",
          2626 => x"84",
          2627 => x"8c",
          2628 => x"b4",
          2629 => x"56",
          2630 => x"82",
          2631 => x"84",
          2632 => x"fc",
          2633 => x"8b",
          2634 => x"52",
          2635 => x"a9",
          2636 => x"85",
          2637 => x"84",
          2638 => x"fc",
          2639 => x"17",
          2640 => x"9c",
          2641 => x"91",
          2642 => x"08",
          2643 => x"17",
          2644 => x"3f",
          2645 => x"81",
          2646 => x"19",
          2647 => x"53",
          2648 => x"17",
          2649 => x"82",
          2650 => x"18",
          2651 => x"80",
          2652 => x"33",
          2653 => x"3f",
          2654 => x"08",
          2655 => x"38",
          2656 => x"82",
          2657 => x"8a",
          2658 => x"fb",
          2659 => x"fe",
          2660 => x"08",
          2661 => x"56",
          2662 => x"74",
          2663 => x"38",
          2664 => x"75",
          2665 => x"16",
          2666 => x"53",
          2667 => x"dc",
          2668 => x"0d",
          2669 => x"0d",
          2670 => x"08",
          2671 => x"81",
          2672 => x"df",
          2673 => x"15",
          2674 => x"d7",
          2675 => x"33",
          2676 => x"82",
          2677 => x"38",
          2678 => x"89",
          2679 => x"2e",
          2680 => x"bf",
          2681 => x"2e",
          2682 => x"81",
          2683 => x"81",
          2684 => x"89",
          2685 => x"08",
          2686 => x"52",
          2687 => x"3f",
          2688 => x"08",
          2689 => x"74",
          2690 => x"14",
          2691 => x"81",
          2692 => x"2a",
          2693 => x"05",
          2694 => x"57",
          2695 => x"f5",
          2696 => x"dc",
          2697 => x"38",
          2698 => x"06",
          2699 => x"33",
          2700 => x"78",
          2701 => x"06",
          2702 => x"5c",
          2703 => x"53",
          2704 => x"38",
          2705 => x"06",
          2706 => x"39",
          2707 => x"a4",
          2708 => x"52",
          2709 => x"bd",
          2710 => x"dc",
          2711 => x"38",
          2712 => x"fe",
          2713 => x"b4",
          2714 => x"8d",
          2715 => x"dc",
          2716 => x"ff",
          2717 => x"39",
          2718 => x"a4",
          2719 => x"52",
          2720 => x"91",
          2721 => x"dc",
          2722 => x"76",
          2723 => x"fc",
          2724 => x"b4",
          2725 => x"f8",
          2726 => x"dc",
          2727 => x"06",
          2728 => x"81",
          2729 => x"8c",
          2730 => x"3d",
          2731 => x"3d",
          2732 => x"7e",
          2733 => x"82",
          2734 => x"27",
          2735 => x"76",
          2736 => x"27",
          2737 => x"75",
          2738 => x"79",
          2739 => x"38",
          2740 => x"89",
          2741 => x"2e",
          2742 => x"80",
          2743 => x"2e",
          2744 => x"81",
          2745 => x"81",
          2746 => x"89",
          2747 => x"08",
          2748 => x"52",
          2749 => x"3f",
          2750 => x"08",
          2751 => x"dc",
          2752 => x"38",
          2753 => x"06",
          2754 => x"81",
          2755 => x"06",
          2756 => x"77",
          2757 => x"2e",
          2758 => x"84",
          2759 => x"06",
          2760 => x"06",
          2761 => x"53",
          2762 => x"81",
          2763 => x"34",
          2764 => x"a4",
          2765 => x"52",
          2766 => x"d9",
          2767 => x"dc",
          2768 => x"8c",
          2769 => x"94",
          2770 => x"ff",
          2771 => x"05",
          2772 => x"54",
          2773 => x"38",
          2774 => x"74",
          2775 => x"06",
          2776 => x"07",
          2777 => x"74",
          2778 => x"39",
          2779 => x"a4",
          2780 => x"52",
          2781 => x"9d",
          2782 => x"dc",
          2783 => x"8c",
          2784 => x"d8",
          2785 => x"ff",
          2786 => x"76",
          2787 => x"06",
          2788 => x"05",
          2789 => x"3f",
          2790 => x"87",
          2791 => x"08",
          2792 => x"51",
          2793 => x"82",
          2794 => x"59",
          2795 => x"08",
          2796 => x"f0",
          2797 => x"82",
          2798 => x"06",
          2799 => x"05",
          2800 => x"54",
          2801 => x"3f",
          2802 => x"08",
          2803 => x"74",
          2804 => x"51",
          2805 => x"81",
          2806 => x"34",
          2807 => x"dc",
          2808 => x"0d",
          2809 => x"0d",
          2810 => x"72",
          2811 => x"56",
          2812 => x"27",
          2813 => x"98",
          2814 => x"9d",
          2815 => x"2e",
          2816 => x"53",
          2817 => x"51",
          2818 => x"82",
          2819 => x"54",
          2820 => x"08",
          2821 => x"93",
          2822 => x"80",
          2823 => x"54",
          2824 => x"82",
          2825 => x"54",
          2826 => x"74",
          2827 => x"fb",
          2828 => x"8c",
          2829 => x"82",
          2830 => x"80",
          2831 => x"38",
          2832 => x"08",
          2833 => x"38",
          2834 => x"08",
          2835 => x"38",
          2836 => x"52",
          2837 => x"d6",
          2838 => x"dc",
          2839 => x"98",
          2840 => x"11",
          2841 => x"57",
          2842 => x"74",
          2843 => x"81",
          2844 => x"0c",
          2845 => x"81",
          2846 => x"84",
          2847 => x"55",
          2848 => x"ff",
          2849 => x"54",
          2850 => x"dc",
          2851 => x"0d",
          2852 => x"0d",
          2853 => x"08",
          2854 => x"79",
          2855 => x"17",
          2856 => x"80",
          2857 => x"98",
          2858 => x"26",
          2859 => x"58",
          2860 => x"52",
          2861 => x"fd",
          2862 => x"74",
          2863 => x"08",
          2864 => x"38",
          2865 => x"08",
          2866 => x"dc",
          2867 => x"82",
          2868 => x"17",
          2869 => x"dc",
          2870 => x"c7",
          2871 => x"90",
          2872 => x"56",
          2873 => x"2e",
          2874 => x"77",
          2875 => x"81",
          2876 => x"38",
          2877 => x"98",
          2878 => x"26",
          2879 => x"56",
          2880 => x"51",
          2881 => x"80",
          2882 => x"dc",
          2883 => x"09",
          2884 => x"38",
          2885 => x"08",
          2886 => x"dc",
          2887 => x"30",
          2888 => x"80",
          2889 => x"07",
          2890 => x"08",
          2891 => x"55",
          2892 => x"ef",
          2893 => x"dc",
          2894 => x"95",
          2895 => x"08",
          2896 => x"27",
          2897 => x"98",
          2898 => x"89",
          2899 => x"85",
          2900 => x"db",
          2901 => x"81",
          2902 => x"17",
          2903 => x"89",
          2904 => x"75",
          2905 => x"ac",
          2906 => x"7a",
          2907 => x"3f",
          2908 => x"08",
          2909 => x"38",
          2910 => x"8c",
          2911 => x"2e",
          2912 => x"86",
          2913 => x"dc",
          2914 => x"8c",
          2915 => x"70",
          2916 => x"07",
          2917 => x"7c",
          2918 => x"55",
          2919 => x"f8",
          2920 => x"2e",
          2921 => x"ff",
          2922 => x"55",
          2923 => x"ff",
          2924 => x"76",
          2925 => x"3f",
          2926 => x"08",
          2927 => x"08",
          2928 => x"8c",
          2929 => x"80",
          2930 => x"55",
          2931 => x"94",
          2932 => x"2e",
          2933 => x"53",
          2934 => x"51",
          2935 => x"82",
          2936 => x"55",
          2937 => x"75",
          2938 => x"98",
          2939 => x"05",
          2940 => x"56",
          2941 => x"26",
          2942 => x"15",
          2943 => x"84",
          2944 => x"07",
          2945 => x"18",
          2946 => x"ff",
          2947 => x"2e",
          2948 => x"39",
          2949 => x"39",
          2950 => x"08",
          2951 => x"81",
          2952 => x"74",
          2953 => x"0c",
          2954 => x"04",
          2955 => x"7a",
          2956 => x"f3",
          2957 => x"8c",
          2958 => x"81",
          2959 => x"dc",
          2960 => x"38",
          2961 => x"51",
          2962 => x"82",
          2963 => x"82",
          2964 => x"b0",
          2965 => x"84",
          2966 => x"52",
          2967 => x"52",
          2968 => x"3f",
          2969 => x"39",
          2970 => x"8a",
          2971 => x"75",
          2972 => x"38",
          2973 => x"19",
          2974 => x"81",
          2975 => x"ed",
          2976 => x"8c",
          2977 => x"2e",
          2978 => x"15",
          2979 => x"70",
          2980 => x"07",
          2981 => x"53",
          2982 => x"75",
          2983 => x"0c",
          2984 => x"04",
          2985 => x"7a",
          2986 => x"58",
          2987 => x"f0",
          2988 => x"80",
          2989 => x"9f",
          2990 => x"80",
          2991 => x"90",
          2992 => x"17",
          2993 => x"aa",
          2994 => x"53",
          2995 => x"88",
          2996 => x"08",
          2997 => x"38",
          2998 => x"53",
          2999 => x"17",
          3000 => x"72",
          3001 => x"fe",
          3002 => x"08",
          3003 => x"80",
          3004 => x"16",
          3005 => x"2b",
          3006 => x"75",
          3007 => x"73",
          3008 => x"f5",
          3009 => x"8c",
          3010 => x"82",
          3011 => x"ff",
          3012 => x"81",
          3013 => x"dc",
          3014 => x"38",
          3015 => x"82",
          3016 => x"26",
          3017 => x"58",
          3018 => x"73",
          3019 => x"39",
          3020 => x"51",
          3021 => x"82",
          3022 => x"98",
          3023 => x"94",
          3024 => x"17",
          3025 => x"58",
          3026 => x"9a",
          3027 => x"81",
          3028 => x"74",
          3029 => x"98",
          3030 => x"83",
          3031 => x"b4",
          3032 => x"0c",
          3033 => x"82",
          3034 => x"8a",
          3035 => x"f8",
          3036 => x"70",
          3037 => x"08",
          3038 => x"57",
          3039 => x"0a",
          3040 => x"38",
          3041 => x"15",
          3042 => x"08",
          3043 => x"72",
          3044 => x"cb",
          3045 => x"ff",
          3046 => x"81",
          3047 => x"13",
          3048 => x"94",
          3049 => x"74",
          3050 => x"85",
          3051 => x"22",
          3052 => x"73",
          3053 => x"38",
          3054 => x"8a",
          3055 => x"05",
          3056 => x"06",
          3057 => x"8a",
          3058 => x"73",
          3059 => x"3f",
          3060 => x"08",
          3061 => x"81",
          3062 => x"dc",
          3063 => x"ff",
          3064 => x"82",
          3065 => x"ff",
          3066 => x"38",
          3067 => x"82",
          3068 => x"26",
          3069 => x"7b",
          3070 => x"98",
          3071 => x"55",
          3072 => x"94",
          3073 => x"73",
          3074 => x"3f",
          3075 => x"08",
          3076 => x"82",
          3077 => x"80",
          3078 => x"38",
          3079 => x"8c",
          3080 => x"2e",
          3081 => x"55",
          3082 => x"08",
          3083 => x"38",
          3084 => x"08",
          3085 => x"fb",
          3086 => x"8c",
          3087 => x"38",
          3088 => x"0c",
          3089 => x"51",
          3090 => x"82",
          3091 => x"98",
          3092 => x"90",
          3093 => x"16",
          3094 => x"15",
          3095 => x"74",
          3096 => x"0c",
          3097 => x"04",
          3098 => x"7b",
          3099 => x"5b",
          3100 => x"52",
          3101 => x"ac",
          3102 => x"dc",
          3103 => x"8c",
          3104 => x"ec",
          3105 => x"dc",
          3106 => x"17",
          3107 => x"51",
          3108 => x"82",
          3109 => x"54",
          3110 => x"08",
          3111 => x"82",
          3112 => x"9c",
          3113 => x"33",
          3114 => x"72",
          3115 => x"09",
          3116 => x"38",
          3117 => x"8c",
          3118 => x"72",
          3119 => x"55",
          3120 => x"53",
          3121 => x"8e",
          3122 => x"56",
          3123 => x"09",
          3124 => x"38",
          3125 => x"8c",
          3126 => x"81",
          3127 => x"fd",
          3128 => x"8c",
          3129 => x"82",
          3130 => x"80",
          3131 => x"38",
          3132 => x"09",
          3133 => x"38",
          3134 => x"82",
          3135 => x"8b",
          3136 => x"fd",
          3137 => x"9a",
          3138 => x"eb",
          3139 => x"8c",
          3140 => x"ff",
          3141 => x"70",
          3142 => x"53",
          3143 => x"09",
          3144 => x"38",
          3145 => x"eb",
          3146 => x"8c",
          3147 => x"2b",
          3148 => x"72",
          3149 => x"0c",
          3150 => x"04",
          3151 => x"77",
          3152 => x"ff",
          3153 => x"9a",
          3154 => x"55",
          3155 => x"76",
          3156 => x"53",
          3157 => x"09",
          3158 => x"38",
          3159 => x"52",
          3160 => x"eb",
          3161 => x"3d",
          3162 => x"3d",
          3163 => x"5b",
          3164 => x"08",
          3165 => x"15",
          3166 => x"81",
          3167 => x"15",
          3168 => x"51",
          3169 => x"82",
          3170 => x"58",
          3171 => x"08",
          3172 => x"9c",
          3173 => x"33",
          3174 => x"86",
          3175 => x"80",
          3176 => x"13",
          3177 => x"06",
          3178 => x"06",
          3179 => x"72",
          3180 => x"82",
          3181 => x"53",
          3182 => x"2e",
          3183 => x"53",
          3184 => x"a9",
          3185 => x"74",
          3186 => x"72",
          3187 => x"38",
          3188 => x"99",
          3189 => x"dc",
          3190 => x"06",
          3191 => x"88",
          3192 => x"06",
          3193 => x"54",
          3194 => x"a0",
          3195 => x"74",
          3196 => x"3f",
          3197 => x"08",
          3198 => x"dc",
          3199 => x"98",
          3200 => x"fa",
          3201 => x"80",
          3202 => x"0c",
          3203 => x"dc",
          3204 => x"0d",
          3205 => x"0d",
          3206 => x"57",
          3207 => x"73",
          3208 => x"3f",
          3209 => x"08",
          3210 => x"dc",
          3211 => x"98",
          3212 => x"75",
          3213 => x"3f",
          3214 => x"08",
          3215 => x"dc",
          3216 => x"a0",
          3217 => x"dc",
          3218 => x"14",
          3219 => x"db",
          3220 => x"a0",
          3221 => x"14",
          3222 => x"ac",
          3223 => x"83",
          3224 => x"82",
          3225 => x"87",
          3226 => x"fd",
          3227 => x"70",
          3228 => x"08",
          3229 => x"55",
          3230 => x"3f",
          3231 => x"08",
          3232 => x"13",
          3233 => x"73",
          3234 => x"83",
          3235 => x"3d",
          3236 => x"3d",
          3237 => x"57",
          3238 => x"89",
          3239 => x"17",
          3240 => x"81",
          3241 => x"70",
          3242 => x"55",
          3243 => x"08",
          3244 => x"81",
          3245 => x"52",
          3246 => x"a8",
          3247 => x"2e",
          3248 => x"84",
          3249 => x"52",
          3250 => x"09",
          3251 => x"38",
          3252 => x"81",
          3253 => x"81",
          3254 => x"73",
          3255 => x"55",
          3256 => x"55",
          3257 => x"c5",
          3258 => x"88",
          3259 => x"0b",
          3260 => x"9c",
          3261 => x"8b",
          3262 => x"17",
          3263 => x"08",
          3264 => x"52",
          3265 => x"82",
          3266 => x"76",
          3267 => x"51",
          3268 => x"82",
          3269 => x"86",
          3270 => x"12",
          3271 => x"3f",
          3272 => x"08",
          3273 => x"88",
          3274 => x"f3",
          3275 => x"70",
          3276 => x"80",
          3277 => x"51",
          3278 => x"af",
          3279 => x"81",
          3280 => x"dc",
          3281 => x"74",
          3282 => x"38",
          3283 => x"88",
          3284 => x"39",
          3285 => x"80",
          3286 => x"56",
          3287 => x"af",
          3288 => x"06",
          3289 => x"56",
          3290 => x"32",
          3291 => x"80",
          3292 => x"51",
          3293 => x"dc",
          3294 => x"1c",
          3295 => x"33",
          3296 => x"9f",
          3297 => x"ff",
          3298 => x"1c",
          3299 => x"7a",
          3300 => x"3f",
          3301 => x"08",
          3302 => x"39",
          3303 => x"a0",
          3304 => x"5e",
          3305 => x"52",
          3306 => x"ff",
          3307 => x"59",
          3308 => x"33",
          3309 => x"ae",
          3310 => x"06",
          3311 => x"78",
          3312 => x"81",
          3313 => x"32",
          3314 => x"9f",
          3315 => x"26",
          3316 => x"53",
          3317 => x"73",
          3318 => x"17",
          3319 => x"34",
          3320 => x"db",
          3321 => x"32",
          3322 => x"9f",
          3323 => x"54",
          3324 => x"2e",
          3325 => x"80",
          3326 => x"75",
          3327 => x"bd",
          3328 => x"7e",
          3329 => x"a0",
          3330 => x"bd",
          3331 => x"82",
          3332 => x"18",
          3333 => x"1a",
          3334 => x"a0",
          3335 => x"fc",
          3336 => x"32",
          3337 => x"80",
          3338 => x"30",
          3339 => x"71",
          3340 => x"51",
          3341 => x"55",
          3342 => x"ac",
          3343 => x"81",
          3344 => x"78",
          3345 => x"51",
          3346 => x"af",
          3347 => x"06",
          3348 => x"55",
          3349 => x"32",
          3350 => x"80",
          3351 => x"51",
          3352 => x"db",
          3353 => x"39",
          3354 => x"09",
          3355 => x"38",
          3356 => x"7c",
          3357 => x"54",
          3358 => x"a2",
          3359 => x"32",
          3360 => x"ae",
          3361 => x"72",
          3362 => x"9f",
          3363 => x"51",
          3364 => x"74",
          3365 => x"88",
          3366 => x"fe",
          3367 => x"98",
          3368 => x"80",
          3369 => x"75",
          3370 => x"81",
          3371 => x"33",
          3372 => x"51",
          3373 => x"82",
          3374 => x"80",
          3375 => x"78",
          3376 => x"81",
          3377 => x"5a",
          3378 => x"d2",
          3379 => x"dc",
          3380 => x"80",
          3381 => x"1c",
          3382 => x"27",
          3383 => x"79",
          3384 => x"74",
          3385 => x"7a",
          3386 => x"74",
          3387 => x"39",
          3388 => x"fa",
          3389 => x"fe",
          3390 => x"dc",
          3391 => x"ff",
          3392 => x"73",
          3393 => x"38",
          3394 => x"81",
          3395 => x"54",
          3396 => x"75",
          3397 => x"17",
          3398 => x"39",
          3399 => x"0c",
          3400 => x"99",
          3401 => x"54",
          3402 => x"2e",
          3403 => x"84",
          3404 => x"34",
          3405 => x"76",
          3406 => x"8b",
          3407 => x"81",
          3408 => x"56",
          3409 => x"80",
          3410 => x"1b",
          3411 => x"08",
          3412 => x"51",
          3413 => x"82",
          3414 => x"56",
          3415 => x"08",
          3416 => x"98",
          3417 => x"76",
          3418 => x"3f",
          3419 => x"08",
          3420 => x"dc",
          3421 => x"38",
          3422 => x"70",
          3423 => x"73",
          3424 => x"be",
          3425 => x"33",
          3426 => x"73",
          3427 => x"8b",
          3428 => x"83",
          3429 => x"06",
          3430 => x"73",
          3431 => x"53",
          3432 => x"51",
          3433 => x"82",
          3434 => x"80",
          3435 => x"75",
          3436 => x"f3",
          3437 => x"9f",
          3438 => x"1c",
          3439 => x"74",
          3440 => x"38",
          3441 => x"09",
          3442 => x"e7",
          3443 => x"2a",
          3444 => x"77",
          3445 => x"51",
          3446 => x"2e",
          3447 => x"81",
          3448 => x"80",
          3449 => x"38",
          3450 => x"ab",
          3451 => x"55",
          3452 => x"75",
          3453 => x"73",
          3454 => x"55",
          3455 => x"82",
          3456 => x"06",
          3457 => x"ab",
          3458 => x"33",
          3459 => x"70",
          3460 => x"55",
          3461 => x"2e",
          3462 => x"1b",
          3463 => x"06",
          3464 => x"52",
          3465 => x"db",
          3466 => x"dc",
          3467 => x"0c",
          3468 => x"74",
          3469 => x"0c",
          3470 => x"04",
          3471 => x"7c",
          3472 => x"08",
          3473 => x"55",
          3474 => x"59",
          3475 => x"81",
          3476 => x"70",
          3477 => x"33",
          3478 => x"52",
          3479 => x"2e",
          3480 => x"ee",
          3481 => x"2e",
          3482 => x"81",
          3483 => x"33",
          3484 => x"81",
          3485 => x"52",
          3486 => x"26",
          3487 => x"14",
          3488 => x"06",
          3489 => x"52",
          3490 => x"80",
          3491 => x"0b",
          3492 => x"59",
          3493 => x"7a",
          3494 => x"70",
          3495 => x"33",
          3496 => x"05",
          3497 => x"9f",
          3498 => x"53",
          3499 => x"89",
          3500 => x"70",
          3501 => x"54",
          3502 => x"12",
          3503 => x"26",
          3504 => x"12",
          3505 => x"06",
          3506 => x"30",
          3507 => x"51",
          3508 => x"2e",
          3509 => x"85",
          3510 => x"be",
          3511 => x"74",
          3512 => x"30",
          3513 => x"9f",
          3514 => x"2a",
          3515 => x"54",
          3516 => x"2e",
          3517 => x"15",
          3518 => x"55",
          3519 => x"ff",
          3520 => x"39",
          3521 => x"86",
          3522 => x"7c",
          3523 => x"51",
          3524 => x"8d",
          3525 => x"70",
          3526 => x"0c",
          3527 => x"04",
          3528 => x"78",
          3529 => x"83",
          3530 => x"0b",
          3531 => x"79",
          3532 => x"e2",
          3533 => x"55",
          3534 => x"08",
          3535 => x"84",
          3536 => x"df",
          3537 => x"8c",
          3538 => x"ff",
          3539 => x"83",
          3540 => x"d4",
          3541 => x"81",
          3542 => x"38",
          3543 => x"17",
          3544 => x"74",
          3545 => x"09",
          3546 => x"38",
          3547 => x"81",
          3548 => x"30",
          3549 => x"79",
          3550 => x"54",
          3551 => x"74",
          3552 => x"09",
          3553 => x"38",
          3554 => x"fa",
          3555 => x"ea",
          3556 => x"b1",
          3557 => x"dc",
          3558 => x"8c",
          3559 => x"2e",
          3560 => x"53",
          3561 => x"52",
          3562 => x"51",
          3563 => x"82",
          3564 => x"55",
          3565 => x"08",
          3566 => x"38",
          3567 => x"82",
          3568 => x"88",
          3569 => x"f2",
          3570 => x"02",
          3571 => x"cb",
          3572 => x"55",
          3573 => x"60",
          3574 => x"3f",
          3575 => x"08",
          3576 => x"80",
          3577 => x"dc",
          3578 => x"fc",
          3579 => x"dc",
          3580 => x"82",
          3581 => x"70",
          3582 => x"8c",
          3583 => x"2e",
          3584 => x"73",
          3585 => x"81",
          3586 => x"33",
          3587 => x"80",
          3588 => x"81",
          3589 => x"d7",
          3590 => x"8c",
          3591 => x"ff",
          3592 => x"06",
          3593 => x"98",
          3594 => x"2e",
          3595 => x"74",
          3596 => x"81",
          3597 => x"8a",
          3598 => x"ac",
          3599 => x"39",
          3600 => x"77",
          3601 => x"81",
          3602 => x"33",
          3603 => x"3f",
          3604 => x"08",
          3605 => x"70",
          3606 => x"55",
          3607 => x"86",
          3608 => x"80",
          3609 => x"74",
          3610 => x"81",
          3611 => x"8a",
          3612 => x"f4",
          3613 => x"53",
          3614 => x"fd",
          3615 => x"8c",
          3616 => x"ff",
          3617 => x"82",
          3618 => x"06",
          3619 => x"8c",
          3620 => x"58",
          3621 => x"f6",
          3622 => x"58",
          3623 => x"2e",
          3624 => x"fa",
          3625 => x"e8",
          3626 => x"dc",
          3627 => x"78",
          3628 => x"5a",
          3629 => x"90",
          3630 => x"75",
          3631 => x"38",
          3632 => x"3d",
          3633 => x"70",
          3634 => x"08",
          3635 => x"7a",
          3636 => x"38",
          3637 => x"51",
          3638 => x"82",
          3639 => x"81",
          3640 => x"81",
          3641 => x"38",
          3642 => x"83",
          3643 => x"38",
          3644 => x"84",
          3645 => x"38",
          3646 => x"81",
          3647 => x"38",
          3648 => x"db",
          3649 => x"8c",
          3650 => x"ff",
          3651 => x"72",
          3652 => x"09",
          3653 => x"d0",
          3654 => x"14",
          3655 => x"3f",
          3656 => x"08",
          3657 => x"06",
          3658 => x"38",
          3659 => x"51",
          3660 => x"82",
          3661 => x"58",
          3662 => x"0c",
          3663 => x"33",
          3664 => x"80",
          3665 => x"ff",
          3666 => x"ff",
          3667 => x"55",
          3668 => x"81",
          3669 => x"38",
          3670 => x"06",
          3671 => x"80",
          3672 => x"52",
          3673 => x"8a",
          3674 => x"80",
          3675 => x"ff",
          3676 => x"53",
          3677 => x"86",
          3678 => x"83",
          3679 => x"c5",
          3680 => x"f5",
          3681 => x"dc",
          3682 => x"8c",
          3683 => x"15",
          3684 => x"06",
          3685 => x"76",
          3686 => x"80",
          3687 => x"da",
          3688 => x"8c",
          3689 => x"ff",
          3690 => x"74",
          3691 => x"d4",
          3692 => x"dc",
          3693 => x"dc",
          3694 => x"c2",
          3695 => x"b9",
          3696 => x"dc",
          3697 => x"ff",
          3698 => x"56",
          3699 => x"83",
          3700 => x"14",
          3701 => x"71",
          3702 => x"5a",
          3703 => x"26",
          3704 => x"8a",
          3705 => x"74",
          3706 => x"ff",
          3707 => x"82",
          3708 => x"55",
          3709 => x"08",
          3710 => x"ec",
          3711 => x"dc",
          3712 => x"ff",
          3713 => x"83",
          3714 => x"74",
          3715 => x"26",
          3716 => x"57",
          3717 => x"26",
          3718 => x"57",
          3719 => x"56",
          3720 => x"82",
          3721 => x"15",
          3722 => x"0c",
          3723 => x"0c",
          3724 => x"a4",
          3725 => x"1d",
          3726 => x"54",
          3727 => x"2e",
          3728 => x"af",
          3729 => x"14",
          3730 => x"3f",
          3731 => x"08",
          3732 => x"06",
          3733 => x"72",
          3734 => x"79",
          3735 => x"80",
          3736 => x"d9",
          3737 => x"8c",
          3738 => x"15",
          3739 => x"2b",
          3740 => x"8d",
          3741 => x"2e",
          3742 => x"77",
          3743 => x"0c",
          3744 => x"76",
          3745 => x"38",
          3746 => x"70",
          3747 => x"81",
          3748 => x"53",
          3749 => x"89",
          3750 => x"56",
          3751 => x"08",
          3752 => x"38",
          3753 => x"15",
          3754 => x"8c",
          3755 => x"80",
          3756 => x"34",
          3757 => x"09",
          3758 => x"92",
          3759 => x"14",
          3760 => x"3f",
          3761 => x"08",
          3762 => x"06",
          3763 => x"2e",
          3764 => x"80",
          3765 => x"1b",
          3766 => x"db",
          3767 => x"8c",
          3768 => x"ea",
          3769 => x"dc",
          3770 => x"34",
          3771 => x"51",
          3772 => x"82",
          3773 => x"83",
          3774 => x"53",
          3775 => x"d5",
          3776 => x"06",
          3777 => x"b4",
          3778 => x"84",
          3779 => x"dc",
          3780 => x"85",
          3781 => x"09",
          3782 => x"38",
          3783 => x"51",
          3784 => x"82",
          3785 => x"86",
          3786 => x"f2",
          3787 => x"06",
          3788 => x"9c",
          3789 => x"d8",
          3790 => x"dc",
          3791 => x"0c",
          3792 => x"51",
          3793 => x"82",
          3794 => x"8c",
          3795 => x"74",
          3796 => x"9c",
          3797 => x"53",
          3798 => x"9c",
          3799 => x"15",
          3800 => x"94",
          3801 => x"56",
          3802 => x"dc",
          3803 => x"0d",
          3804 => x"0d",
          3805 => x"55",
          3806 => x"b9",
          3807 => x"53",
          3808 => x"b1",
          3809 => x"52",
          3810 => x"a9",
          3811 => x"22",
          3812 => x"57",
          3813 => x"2e",
          3814 => x"99",
          3815 => x"33",
          3816 => x"3f",
          3817 => x"08",
          3818 => x"71",
          3819 => x"74",
          3820 => x"83",
          3821 => x"78",
          3822 => x"52",
          3823 => x"dc",
          3824 => x"0d",
          3825 => x"0d",
          3826 => x"33",
          3827 => x"3d",
          3828 => x"56",
          3829 => x"8b",
          3830 => x"82",
          3831 => x"24",
          3832 => x"8c",
          3833 => x"29",
          3834 => x"05",
          3835 => x"55",
          3836 => x"84",
          3837 => x"34",
          3838 => x"80",
          3839 => x"80",
          3840 => x"75",
          3841 => x"75",
          3842 => x"38",
          3843 => x"3d",
          3844 => x"05",
          3845 => x"3f",
          3846 => x"08",
          3847 => x"8c",
          3848 => x"3d",
          3849 => x"3d",
          3850 => x"84",
          3851 => x"05",
          3852 => x"89",
          3853 => x"2e",
          3854 => x"77",
          3855 => x"54",
          3856 => x"05",
          3857 => x"84",
          3858 => x"f6",
          3859 => x"8c",
          3860 => x"82",
          3861 => x"84",
          3862 => x"5c",
          3863 => x"3d",
          3864 => x"ed",
          3865 => x"8c",
          3866 => x"82",
          3867 => x"92",
          3868 => x"d7",
          3869 => x"98",
          3870 => x"73",
          3871 => x"38",
          3872 => x"9c",
          3873 => x"80",
          3874 => x"38",
          3875 => x"95",
          3876 => x"2e",
          3877 => x"aa",
          3878 => x"ea",
          3879 => x"8c",
          3880 => x"9e",
          3881 => x"05",
          3882 => x"54",
          3883 => x"38",
          3884 => x"70",
          3885 => x"54",
          3886 => x"8e",
          3887 => x"83",
          3888 => x"88",
          3889 => x"83",
          3890 => x"83",
          3891 => x"06",
          3892 => x"80",
          3893 => x"38",
          3894 => x"51",
          3895 => x"82",
          3896 => x"56",
          3897 => x"0a",
          3898 => x"05",
          3899 => x"3f",
          3900 => x"0b",
          3901 => x"80",
          3902 => x"7a",
          3903 => x"3f",
          3904 => x"9c",
          3905 => x"d1",
          3906 => x"81",
          3907 => x"34",
          3908 => x"80",
          3909 => x"b0",
          3910 => x"54",
          3911 => x"52",
          3912 => x"05",
          3913 => x"3f",
          3914 => x"08",
          3915 => x"dc",
          3916 => x"38",
          3917 => x"82",
          3918 => x"b2",
          3919 => x"84",
          3920 => x"06",
          3921 => x"73",
          3922 => x"38",
          3923 => x"ad",
          3924 => x"2a",
          3925 => x"51",
          3926 => x"2e",
          3927 => x"81",
          3928 => x"80",
          3929 => x"87",
          3930 => x"39",
          3931 => x"51",
          3932 => x"82",
          3933 => x"7b",
          3934 => x"12",
          3935 => x"82",
          3936 => x"81",
          3937 => x"83",
          3938 => x"06",
          3939 => x"80",
          3940 => x"77",
          3941 => x"58",
          3942 => x"08",
          3943 => x"63",
          3944 => x"63",
          3945 => x"57",
          3946 => x"82",
          3947 => x"82",
          3948 => x"88",
          3949 => x"9c",
          3950 => x"d2",
          3951 => x"8c",
          3952 => x"8c",
          3953 => x"1b",
          3954 => x"0c",
          3955 => x"22",
          3956 => x"77",
          3957 => x"80",
          3958 => x"34",
          3959 => x"1a",
          3960 => x"94",
          3961 => x"85",
          3962 => x"06",
          3963 => x"80",
          3964 => x"38",
          3965 => x"08",
          3966 => x"84",
          3967 => x"dc",
          3968 => x"0c",
          3969 => x"70",
          3970 => x"52",
          3971 => x"39",
          3972 => x"51",
          3973 => x"82",
          3974 => x"57",
          3975 => x"08",
          3976 => x"38",
          3977 => x"8c",
          3978 => x"2e",
          3979 => x"83",
          3980 => x"75",
          3981 => x"74",
          3982 => x"07",
          3983 => x"54",
          3984 => x"8a",
          3985 => x"75",
          3986 => x"73",
          3987 => x"98",
          3988 => x"a9",
          3989 => x"ff",
          3990 => x"80",
          3991 => x"76",
          3992 => x"d6",
          3993 => x"8c",
          3994 => x"38",
          3995 => x"39",
          3996 => x"82",
          3997 => x"05",
          3998 => x"84",
          3999 => x"0c",
          4000 => x"82",
          4001 => x"97",
          4002 => x"f2",
          4003 => x"63",
          4004 => x"40",
          4005 => x"7e",
          4006 => x"fc",
          4007 => x"51",
          4008 => x"82",
          4009 => x"55",
          4010 => x"08",
          4011 => x"19",
          4012 => x"80",
          4013 => x"74",
          4014 => x"39",
          4015 => x"81",
          4016 => x"56",
          4017 => x"82",
          4018 => x"39",
          4019 => x"1a",
          4020 => x"82",
          4021 => x"0b",
          4022 => x"81",
          4023 => x"39",
          4024 => x"94",
          4025 => x"55",
          4026 => x"83",
          4027 => x"7b",
          4028 => x"89",
          4029 => x"08",
          4030 => x"06",
          4031 => x"81",
          4032 => x"8a",
          4033 => x"05",
          4034 => x"06",
          4035 => x"a8",
          4036 => x"38",
          4037 => x"55",
          4038 => x"19",
          4039 => x"51",
          4040 => x"82",
          4041 => x"55",
          4042 => x"ff",
          4043 => x"ff",
          4044 => x"38",
          4045 => x"0c",
          4046 => x"52",
          4047 => x"cb",
          4048 => x"dc",
          4049 => x"ff",
          4050 => x"8c",
          4051 => x"7c",
          4052 => x"57",
          4053 => x"80",
          4054 => x"1a",
          4055 => x"22",
          4056 => x"75",
          4057 => x"38",
          4058 => x"58",
          4059 => x"53",
          4060 => x"1b",
          4061 => x"88",
          4062 => x"dc",
          4063 => x"38",
          4064 => x"33",
          4065 => x"80",
          4066 => x"b0",
          4067 => x"31",
          4068 => x"27",
          4069 => x"80",
          4070 => x"52",
          4071 => x"77",
          4072 => x"7d",
          4073 => x"e0",
          4074 => x"2b",
          4075 => x"76",
          4076 => x"94",
          4077 => x"ff",
          4078 => x"71",
          4079 => x"7b",
          4080 => x"38",
          4081 => x"19",
          4082 => x"51",
          4083 => x"82",
          4084 => x"fe",
          4085 => x"53",
          4086 => x"83",
          4087 => x"b4",
          4088 => x"51",
          4089 => x"7b",
          4090 => x"08",
          4091 => x"76",
          4092 => x"08",
          4093 => x"0c",
          4094 => x"f3",
          4095 => x"75",
          4096 => x"0c",
          4097 => x"04",
          4098 => x"60",
          4099 => x"40",
          4100 => x"80",
          4101 => x"3d",
          4102 => x"77",
          4103 => x"3f",
          4104 => x"08",
          4105 => x"dc",
          4106 => x"91",
          4107 => x"74",
          4108 => x"38",
          4109 => x"b8",
          4110 => x"33",
          4111 => x"70",
          4112 => x"56",
          4113 => x"74",
          4114 => x"a4",
          4115 => x"82",
          4116 => x"34",
          4117 => x"98",
          4118 => x"91",
          4119 => x"56",
          4120 => x"94",
          4121 => x"11",
          4122 => x"76",
          4123 => x"75",
          4124 => x"80",
          4125 => x"38",
          4126 => x"70",
          4127 => x"56",
          4128 => x"fd",
          4129 => x"11",
          4130 => x"77",
          4131 => x"5c",
          4132 => x"38",
          4133 => x"88",
          4134 => x"74",
          4135 => x"52",
          4136 => x"18",
          4137 => x"51",
          4138 => x"82",
          4139 => x"55",
          4140 => x"08",
          4141 => x"ab",
          4142 => x"2e",
          4143 => x"74",
          4144 => x"95",
          4145 => x"19",
          4146 => x"08",
          4147 => x"88",
          4148 => x"55",
          4149 => x"9c",
          4150 => x"09",
          4151 => x"38",
          4152 => x"c1",
          4153 => x"dc",
          4154 => x"38",
          4155 => x"52",
          4156 => x"97",
          4157 => x"dc",
          4158 => x"fe",
          4159 => x"8c",
          4160 => x"7c",
          4161 => x"57",
          4162 => x"80",
          4163 => x"1b",
          4164 => x"22",
          4165 => x"75",
          4166 => x"38",
          4167 => x"59",
          4168 => x"53",
          4169 => x"1a",
          4170 => x"be",
          4171 => x"dc",
          4172 => x"38",
          4173 => x"08",
          4174 => x"56",
          4175 => x"9b",
          4176 => x"53",
          4177 => x"77",
          4178 => x"7d",
          4179 => x"16",
          4180 => x"3f",
          4181 => x"0b",
          4182 => x"78",
          4183 => x"80",
          4184 => x"18",
          4185 => x"08",
          4186 => x"7e",
          4187 => x"3f",
          4188 => x"08",
          4189 => x"7e",
          4190 => x"0c",
          4191 => x"19",
          4192 => x"08",
          4193 => x"84",
          4194 => x"57",
          4195 => x"27",
          4196 => x"56",
          4197 => x"52",
          4198 => x"f9",
          4199 => x"dc",
          4200 => x"38",
          4201 => x"52",
          4202 => x"83",
          4203 => x"b4",
          4204 => x"d4",
          4205 => x"81",
          4206 => x"34",
          4207 => x"7e",
          4208 => x"0c",
          4209 => x"1a",
          4210 => x"94",
          4211 => x"1b",
          4212 => x"5e",
          4213 => x"27",
          4214 => x"55",
          4215 => x"0c",
          4216 => x"90",
          4217 => x"c0",
          4218 => x"90",
          4219 => x"56",
          4220 => x"dc",
          4221 => x"0d",
          4222 => x"0d",
          4223 => x"fc",
          4224 => x"52",
          4225 => x"3f",
          4226 => x"08",
          4227 => x"dc",
          4228 => x"38",
          4229 => x"70",
          4230 => x"81",
          4231 => x"55",
          4232 => x"80",
          4233 => x"16",
          4234 => x"51",
          4235 => x"82",
          4236 => x"57",
          4237 => x"08",
          4238 => x"a4",
          4239 => x"11",
          4240 => x"55",
          4241 => x"16",
          4242 => x"08",
          4243 => x"75",
          4244 => x"e8",
          4245 => x"08",
          4246 => x"51",
          4247 => x"82",
          4248 => x"52",
          4249 => x"c9",
          4250 => x"52",
          4251 => x"c9",
          4252 => x"54",
          4253 => x"15",
          4254 => x"cc",
          4255 => x"8c",
          4256 => x"17",
          4257 => x"06",
          4258 => x"90",
          4259 => x"82",
          4260 => x"8a",
          4261 => x"fc",
          4262 => x"70",
          4263 => x"d9",
          4264 => x"dc",
          4265 => x"8c",
          4266 => x"38",
          4267 => x"05",
          4268 => x"f1",
          4269 => x"8c",
          4270 => x"82",
          4271 => x"87",
          4272 => x"dc",
          4273 => x"72",
          4274 => x"0c",
          4275 => x"04",
          4276 => x"84",
          4277 => x"e4",
          4278 => x"80",
          4279 => x"dc",
          4280 => x"38",
          4281 => x"08",
          4282 => x"34",
          4283 => x"82",
          4284 => x"83",
          4285 => x"ef",
          4286 => x"53",
          4287 => x"05",
          4288 => x"51",
          4289 => x"82",
          4290 => x"55",
          4291 => x"08",
          4292 => x"76",
          4293 => x"93",
          4294 => x"51",
          4295 => x"82",
          4296 => x"55",
          4297 => x"08",
          4298 => x"80",
          4299 => x"70",
          4300 => x"56",
          4301 => x"89",
          4302 => x"94",
          4303 => x"b2",
          4304 => x"05",
          4305 => x"2a",
          4306 => x"51",
          4307 => x"80",
          4308 => x"76",
          4309 => x"52",
          4310 => x"3f",
          4311 => x"08",
          4312 => x"8e",
          4313 => x"dc",
          4314 => x"09",
          4315 => x"38",
          4316 => x"82",
          4317 => x"93",
          4318 => x"e4",
          4319 => x"6f",
          4320 => x"7a",
          4321 => x"9e",
          4322 => x"05",
          4323 => x"51",
          4324 => x"82",
          4325 => x"57",
          4326 => x"08",
          4327 => x"7b",
          4328 => x"94",
          4329 => x"55",
          4330 => x"73",
          4331 => x"ed",
          4332 => x"93",
          4333 => x"55",
          4334 => x"82",
          4335 => x"57",
          4336 => x"08",
          4337 => x"68",
          4338 => x"c9",
          4339 => x"8c",
          4340 => x"82",
          4341 => x"82",
          4342 => x"52",
          4343 => x"a3",
          4344 => x"dc",
          4345 => x"52",
          4346 => x"b8",
          4347 => x"dc",
          4348 => x"8c",
          4349 => x"a2",
          4350 => x"74",
          4351 => x"3f",
          4352 => x"08",
          4353 => x"dc",
          4354 => x"69",
          4355 => x"d9",
          4356 => x"82",
          4357 => x"2e",
          4358 => x"52",
          4359 => x"cf",
          4360 => x"dc",
          4361 => x"8c",
          4362 => x"2e",
          4363 => x"84",
          4364 => x"06",
          4365 => x"57",
          4366 => x"76",
          4367 => x"9e",
          4368 => x"05",
          4369 => x"dc",
          4370 => x"90",
          4371 => x"81",
          4372 => x"56",
          4373 => x"80",
          4374 => x"02",
          4375 => x"81",
          4376 => x"70",
          4377 => x"56",
          4378 => x"81",
          4379 => x"78",
          4380 => x"38",
          4381 => x"99",
          4382 => x"81",
          4383 => x"18",
          4384 => x"18",
          4385 => x"58",
          4386 => x"33",
          4387 => x"ee",
          4388 => x"6f",
          4389 => x"af",
          4390 => x"8d",
          4391 => x"2e",
          4392 => x"8a",
          4393 => x"6f",
          4394 => x"af",
          4395 => x"0b",
          4396 => x"33",
          4397 => x"81",
          4398 => x"70",
          4399 => x"52",
          4400 => x"56",
          4401 => x"8d",
          4402 => x"70",
          4403 => x"51",
          4404 => x"f5",
          4405 => x"54",
          4406 => x"a7",
          4407 => x"74",
          4408 => x"38",
          4409 => x"73",
          4410 => x"81",
          4411 => x"81",
          4412 => x"39",
          4413 => x"81",
          4414 => x"74",
          4415 => x"81",
          4416 => x"91",
          4417 => x"6e",
          4418 => x"59",
          4419 => x"7a",
          4420 => x"5c",
          4421 => x"26",
          4422 => x"7a",
          4423 => x"8c",
          4424 => x"3d",
          4425 => x"3d",
          4426 => x"8d",
          4427 => x"54",
          4428 => x"55",
          4429 => x"82",
          4430 => x"53",
          4431 => x"08",
          4432 => x"91",
          4433 => x"72",
          4434 => x"8c",
          4435 => x"73",
          4436 => x"38",
          4437 => x"70",
          4438 => x"81",
          4439 => x"57",
          4440 => x"73",
          4441 => x"08",
          4442 => x"94",
          4443 => x"75",
          4444 => x"97",
          4445 => x"11",
          4446 => x"2b",
          4447 => x"73",
          4448 => x"38",
          4449 => x"16",
          4450 => x"d0",
          4451 => x"dc",
          4452 => x"78",
          4453 => x"55",
          4454 => x"c0",
          4455 => x"dc",
          4456 => x"96",
          4457 => x"70",
          4458 => x"94",
          4459 => x"71",
          4460 => x"08",
          4461 => x"53",
          4462 => x"15",
          4463 => x"a6",
          4464 => x"74",
          4465 => x"3f",
          4466 => x"08",
          4467 => x"dc",
          4468 => x"81",
          4469 => x"8c",
          4470 => x"2e",
          4471 => x"82",
          4472 => x"88",
          4473 => x"98",
          4474 => x"80",
          4475 => x"38",
          4476 => x"80",
          4477 => x"77",
          4478 => x"08",
          4479 => x"0c",
          4480 => x"70",
          4481 => x"81",
          4482 => x"5a",
          4483 => x"2e",
          4484 => x"52",
          4485 => x"f9",
          4486 => x"dc",
          4487 => x"8c",
          4488 => x"38",
          4489 => x"08",
          4490 => x"73",
          4491 => x"c7",
          4492 => x"8c",
          4493 => x"73",
          4494 => x"38",
          4495 => x"af",
          4496 => x"73",
          4497 => x"27",
          4498 => x"98",
          4499 => x"a0",
          4500 => x"08",
          4501 => x"0c",
          4502 => x"06",
          4503 => x"2e",
          4504 => x"52",
          4505 => x"a3",
          4506 => x"dc",
          4507 => x"82",
          4508 => x"34",
          4509 => x"c4",
          4510 => x"91",
          4511 => x"53",
          4512 => x"89",
          4513 => x"dc",
          4514 => x"94",
          4515 => x"8c",
          4516 => x"27",
          4517 => x"8c",
          4518 => x"15",
          4519 => x"07",
          4520 => x"16",
          4521 => x"ff",
          4522 => x"80",
          4523 => x"77",
          4524 => x"2e",
          4525 => x"9c",
          4526 => x"53",
          4527 => x"dc",
          4528 => x"0d",
          4529 => x"0d",
          4530 => x"54",
          4531 => x"81",
          4532 => x"53",
          4533 => x"05",
          4534 => x"84",
          4535 => x"e7",
          4536 => x"dc",
          4537 => x"8c",
          4538 => x"ea",
          4539 => x"0c",
          4540 => x"51",
          4541 => x"82",
          4542 => x"55",
          4543 => x"08",
          4544 => x"ab",
          4545 => x"98",
          4546 => x"80",
          4547 => x"38",
          4548 => x"70",
          4549 => x"81",
          4550 => x"57",
          4551 => x"ad",
          4552 => x"08",
          4553 => x"d3",
          4554 => x"8c",
          4555 => x"17",
          4556 => x"86",
          4557 => x"17",
          4558 => x"75",
          4559 => x"3f",
          4560 => x"08",
          4561 => x"2e",
          4562 => x"85",
          4563 => x"86",
          4564 => x"2e",
          4565 => x"76",
          4566 => x"73",
          4567 => x"0c",
          4568 => x"04",
          4569 => x"76",
          4570 => x"05",
          4571 => x"53",
          4572 => x"82",
          4573 => x"87",
          4574 => x"dc",
          4575 => x"86",
          4576 => x"fb",
          4577 => x"79",
          4578 => x"05",
          4579 => x"56",
          4580 => x"3f",
          4581 => x"08",
          4582 => x"dc",
          4583 => x"38",
          4584 => x"82",
          4585 => x"52",
          4586 => x"f8",
          4587 => x"dc",
          4588 => x"ca",
          4589 => x"dc",
          4590 => x"51",
          4591 => x"82",
          4592 => x"53",
          4593 => x"08",
          4594 => x"81",
          4595 => x"80",
          4596 => x"82",
          4597 => x"a6",
          4598 => x"73",
          4599 => x"3f",
          4600 => x"51",
          4601 => x"82",
          4602 => x"84",
          4603 => x"70",
          4604 => x"2c",
          4605 => x"dc",
          4606 => x"51",
          4607 => x"82",
          4608 => x"87",
          4609 => x"ee",
          4610 => x"57",
          4611 => x"3d",
          4612 => x"3d",
          4613 => x"af",
          4614 => x"dc",
          4615 => x"8c",
          4616 => x"38",
          4617 => x"51",
          4618 => x"82",
          4619 => x"55",
          4620 => x"08",
          4621 => x"80",
          4622 => x"70",
          4623 => x"58",
          4624 => x"85",
          4625 => x"8d",
          4626 => x"2e",
          4627 => x"52",
          4628 => x"be",
          4629 => x"8c",
          4630 => x"3d",
          4631 => x"3d",
          4632 => x"55",
          4633 => x"92",
          4634 => x"52",
          4635 => x"de",
          4636 => x"8c",
          4637 => x"82",
          4638 => x"82",
          4639 => x"74",
          4640 => x"98",
          4641 => x"11",
          4642 => x"59",
          4643 => x"75",
          4644 => x"38",
          4645 => x"81",
          4646 => x"5b",
          4647 => x"82",
          4648 => x"39",
          4649 => x"08",
          4650 => x"59",
          4651 => x"09",
          4652 => x"38",
          4653 => x"57",
          4654 => x"3d",
          4655 => x"c1",
          4656 => x"8c",
          4657 => x"2e",
          4658 => x"8c",
          4659 => x"2e",
          4660 => x"8c",
          4661 => x"70",
          4662 => x"08",
          4663 => x"7a",
          4664 => x"7f",
          4665 => x"54",
          4666 => x"77",
          4667 => x"80",
          4668 => x"15",
          4669 => x"dc",
          4670 => x"75",
          4671 => x"52",
          4672 => x"52",
          4673 => x"8d",
          4674 => x"dc",
          4675 => x"8c",
          4676 => x"d6",
          4677 => x"33",
          4678 => x"1a",
          4679 => x"54",
          4680 => x"09",
          4681 => x"38",
          4682 => x"ff",
          4683 => x"82",
          4684 => x"83",
          4685 => x"70",
          4686 => x"25",
          4687 => x"59",
          4688 => x"9b",
          4689 => x"51",
          4690 => x"3f",
          4691 => x"08",
          4692 => x"70",
          4693 => x"25",
          4694 => x"59",
          4695 => x"75",
          4696 => x"7a",
          4697 => x"ff",
          4698 => x"7c",
          4699 => x"90",
          4700 => x"11",
          4701 => x"56",
          4702 => x"15",
          4703 => x"8c",
          4704 => x"3d",
          4705 => x"3d",
          4706 => x"3d",
          4707 => x"70",
          4708 => x"dd",
          4709 => x"dc",
          4710 => x"8c",
          4711 => x"a8",
          4712 => x"33",
          4713 => x"a0",
          4714 => x"33",
          4715 => x"70",
          4716 => x"55",
          4717 => x"73",
          4718 => x"8e",
          4719 => x"08",
          4720 => x"18",
          4721 => x"80",
          4722 => x"38",
          4723 => x"08",
          4724 => x"08",
          4725 => x"c4",
          4726 => x"8c",
          4727 => x"88",
          4728 => x"80",
          4729 => x"17",
          4730 => x"51",
          4731 => x"3f",
          4732 => x"08",
          4733 => x"81",
          4734 => x"81",
          4735 => x"dc",
          4736 => x"09",
          4737 => x"38",
          4738 => x"39",
          4739 => x"77",
          4740 => x"dc",
          4741 => x"08",
          4742 => x"98",
          4743 => x"82",
          4744 => x"52",
          4745 => x"bd",
          4746 => x"dc",
          4747 => x"17",
          4748 => x"0c",
          4749 => x"80",
          4750 => x"73",
          4751 => x"75",
          4752 => x"38",
          4753 => x"34",
          4754 => x"82",
          4755 => x"89",
          4756 => x"e2",
          4757 => x"53",
          4758 => x"a4",
          4759 => x"3d",
          4760 => x"3f",
          4761 => x"08",
          4762 => x"dc",
          4763 => x"38",
          4764 => x"3d",
          4765 => x"3d",
          4766 => x"d1",
          4767 => x"8c",
          4768 => x"82",
          4769 => x"81",
          4770 => x"80",
          4771 => x"70",
          4772 => x"81",
          4773 => x"56",
          4774 => x"81",
          4775 => x"98",
          4776 => x"74",
          4777 => x"38",
          4778 => x"05",
          4779 => x"06",
          4780 => x"55",
          4781 => x"38",
          4782 => x"51",
          4783 => x"82",
          4784 => x"74",
          4785 => x"81",
          4786 => x"56",
          4787 => x"80",
          4788 => x"54",
          4789 => x"08",
          4790 => x"2e",
          4791 => x"73",
          4792 => x"dc",
          4793 => x"52",
          4794 => x"52",
          4795 => x"3f",
          4796 => x"08",
          4797 => x"dc",
          4798 => x"38",
          4799 => x"08",
          4800 => x"cc",
          4801 => x"8c",
          4802 => x"82",
          4803 => x"86",
          4804 => x"80",
          4805 => x"8c",
          4806 => x"2e",
          4807 => x"8c",
          4808 => x"c0",
          4809 => x"ce",
          4810 => x"8c",
          4811 => x"8c",
          4812 => x"70",
          4813 => x"08",
          4814 => x"51",
          4815 => x"80",
          4816 => x"73",
          4817 => x"38",
          4818 => x"52",
          4819 => x"95",
          4820 => x"dc",
          4821 => x"8c",
          4822 => x"ff",
          4823 => x"82",
          4824 => x"55",
          4825 => x"dc",
          4826 => x"0d",
          4827 => x"0d",
          4828 => x"3d",
          4829 => x"9a",
          4830 => x"cb",
          4831 => x"dc",
          4832 => x"8c",
          4833 => x"b0",
          4834 => x"69",
          4835 => x"70",
          4836 => x"97",
          4837 => x"dc",
          4838 => x"8c",
          4839 => x"38",
          4840 => x"94",
          4841 => x"dc",
          4842 => x"09",
          4843 => x"88",
          4844 => x"df",
          4845 => x"85",
          4846 => x"51",
          4847 => x"74",
          4848 => x"78",
          4849 => x"8a",
          4850 => x"57",
          4851 => x"82",
          4852 => x"75",
          4853 => x"8c",
          4854 => x"38",
          4855 => x"8c",
          4856 => x"2e",
          4857 => x"83",
          4858 => x"82",
          4859 => x"ff",
          4860 => x"06",
          4861 => x"54",
          4862 => x"73",
          4863 => x"82",
          4864 => x"52",
          4865 => x"a4",
          4866 => x"dc",
          4867 => x"8c",
          4868 => x"9a",
          4869 => x"a0",
          4870 => x"51",
          4871 => x"3f",
          4872 => x"0b",
          4873 => x"78",
          4874 => x"bf",
          4875 => x"88",
          4876 => x"80",
          4877 => x"ff",
          4878 => x"75",
          4879 => x"11",
          4880 => x"f8",
          4881 => x"78",
          4882 => x"80",
          4883 => x"ff",
          4884 => x"78",
          4885 => x"80",
          4886 => x"7f",
          4887 => x"d4",
          4888 => x"c9",
          4889 => x"54",
          4890 => x"15",
          4891 => x"cb",
          4892 => x"8c",
          4893 => x"82",
          4894 => x"b2",
          4895 => x"b2",
          4896 => x"96",
          4897 => x"b5",
          4898 => x"53",
          4899 => x"51",
          4900 => x"64",
          4901 => x"8b",
          4902 => x"54",
          4903 => x"15",
          4904 => x"ff",
          4905 => x"82",
          4906 => x"54",
          4907 => x"53",
          4908 => x"51",
          4909 => x"3f",
          4910 => x"dc",
          4911 => x"0d",
          4912 => x"0d",
          4913 => x"05",
          4914 => x"3f",
          4915 => x"3d",
          4916 => x"52",
          4917 => x"d5",
          4918 => x"8c",
          4919 => x"82",
          4920 => x"82",
          4921 => x"4d",
          4922 => x"52",
          4923 => x"52",
          4924 => x"3f",
          4925 => x"08",
          4926 => x"dc",
          4927 => x"38",
          4928 => x"05",
          4929 => x"06",
          4930 => x"73",
          4931 => x"a0",
          4932 => x"08",
          4933 => x"ff",
          4934 => x"ff",
          4935 => x"ac",
          4936 => x"92",
          4937 => x"54",
          4938 => x"3f",
          4939 => x"52",
          4940 => x"f7",
          4941 => x"dc",
          4942 => x"8c",
          4943 => x"38",
          4944 => x"09",
          4945 => x"38",
          4946 => x"08",
          4947 => x"88",
          4948 => x"39",
          4949 => x"08",
          4950 => x"81",
          4951 => x"38",
          4952 => x"b1",
          4953 => x"dc",
          4954 => x"8c",
          4955 => x"c8",
          4956 => x"93",
          4957 => x"ff",
          4958 => x"8d",
          4959 => x"b4",
          4960 => x"af",
          4961 => x"17",
          4962 => x"33",
          4963 => x"70",
          4964 => x"55",
          4965 => x"38",
          4966 => x"54",
          4967 => x"34",
          4968 => x"0b",
          4969 => x"8b",
          4970 => x"84",
          4971 => x"06",
          4972 => x"73",
          4973 => x"e5",
          4974 => x"2e",
          4975 => x"75",
          4976 => x"c6",
          4977 => x"8c",
          4978 => x"78",
          4979 => x"bb",
          4980 => x"82",
          4981 => x"80",
          4982 => x"38",
          4983 => x"08",
          4984 => x"ff",
          4985 => x"82",
          4986 => x"79",
          4987 => x"58",
          4988 => x"8c",
          4989 => x"c0",
          4990 => x"33",
          4991 => x"2e",
          4992 => x"99",
          4993 => x"75",
          4994 => x"c6",
          4995 => x"54",
          4996 => x"15",
          4997 => x"82",
          4998 => x"9c",
          4999 => x"c8",
          5000 => x"8c",
          5001 => x"82",
          5002 => x"8c",
          5003 => x"ff",
          5004 => x"82",
          5005 => x"55",
          5006 => x"dc",
          5007 => x"0d",
          5008 => x"0d",
          5009 => x"05",
          5010 => x"05",
          5011 => x"33",
          5012 => x"53",
          5013 => x"05",
          5014 => x"51",
          5015 => x"82",
          5016 => x"55",
          5017 => x"08",
          5018 => x"78",
          5019 => x"95",
          5020 => x"51",
          5021 => x"82",
          5022 => x"55",
          5023 => x"08",
          5024 => x"80",
          5025 => x"81",
          5026 => x"86",
          5027 => x"38",
          5028 => x"61",
          5029 => x"12",
          5030 => x"7a",
          5031 => x"51",
          5032 => x"74",
          5033 => x"78",
          5034 => x"83",
          5035 => x"51",
          5036 => x"3f",
          5037 => x"08",
          5038 => x"8c",
          5039 => x"3d",
          5040 => x"3d",
          5041 => x"82",
          5042 => x"d0",
          5043 => x"3d",
          5044 => x"3f",
          5045 => x"08",
          5046 => x"dc",
          5047 => x"38",
          5048 => x"52",
          5049 => x"05",
          5050 => x"3f",
          5051 => x"08",
          5052 => x"dc",
          5053 => x"02",
          5054 => x"33",
          5055 => x"54",
          5056 => x"a6",
          5057 => x"22",
          5058 => x"71",
          5059 => x"53",
          5060 => x"51",
          5061 => x"3f",
          5062 => x"0b",
          5063 => x"76",
          5064 => x"b8",
          5065 => x"dc",
          5066 => x"82",
          5067 => x"93",
          5068 => x"ea",
          5069 => x"6b",
          5070 => x"53",
          5071 => x"05",
          5072 => x"51",
          5073 => x"82",
          5074 => x"82",
          5075 => x"30",
          5076 => x"dc",
          5077 => x"25",
          5078 => x"79",
          5079 => x"85",
          5080 => x"75",
          5081 => x"73",
          5082 => x"f9",
          5083 => x"80",
          5084 => x"8d",
          5085 => x"54",
          5086 => x"3f",
          5087 => x"08",
          5088 => x"dc",
          5089 => x"38",
          5090 => x"51",
          5091 => x"82",
          5092 => x"57",
          5093 => x"08",
          5094 => x"8c",
          5095 => x"8c",
          5096 => x"5b",
          5097 => x"18",
          5098 => x"18",
          5099 => x"74",
          5100 => x"81",
          5101 => x"78",
          5102 => x"8b",
          5103 => x"54",
          5104 => x"75",
          5105 => x"38",
          5106 => x"1b",
          5107 => x"55",
          5108 => x"2e",
          5109 => x"39",
          5110 => x"09",
          5111 => x"38",
          5112 => x"80",
          5113 => x"70",
          5114 => x"25",
          5115 => x"80",
          5116 => x"38",
          5117 => x"bc",
          5118 => x"11",
          5119 => x"ff",
          5120 => x"82",
          5121 => x"57",
          5122 => x"08",
          5123 => x"70",
          5124 => x"80",
          5125 => x"83",
          5126 => x"80",
          5127 => x"84",
          5128 => x"a7",
          5129 => x"b4",
          5130 => x"ad",
          5131 => x"8c",
          5132 => x"0c",
          5133 => x"dc",
          5134 => x"0d",
          5135 => x"0d",
          5136 => x"3d",
          5137 => x"52",
          5138 => x"ce",
          5139 => x"8c",
          5140 => x"8c",
          5141 => x"54",
          5142 => x"08",
          5143 => x"8b",
          5144 => x"8b",
          5145 => x"59",
          5146 => x"3f",
          5147 => x"33",
          5148 => x"06",
          5149 => x"57",
          5150 => x"81",
          5151 => x"58",
          5152 => x"06",
          5153 => x"4e",
          5154 => x"ff",
          5155 => x"82",
          5156 => x"80",
          5157 => x"6c",
          5158 => x"53",
          5159 => x"ae",
          5160 => x"8c",
          5161 => x"2e",
          5162 => x"88",
          5163 => x"6d",
          5164 => x"55",
          5165 => x"8c",
          5166 => x"ff",
          5167 => x"83",
          5168 => x"51",
          5169 => x"26",
          5170 => x"15",
          5171 => x"ff",
          5172 => x"80",
          5173 => x"87",
          5174 => x"ec",
          5175 => x"74",
          5176 => x"38",
          5177 => x"fb",
          5178 => x"ae",
          5179 => x"8c",
          5180 => x"38",
          5181 => x"27",
          5182 => x"89",
          5183 => x"8b",
          5184 => x"27",
          5185 => x"55",
          5186 => x"81",
          5187 => x"8f",
          5188 => x"2a",
          5189 => x"70",
          5190 => x"34",
          5191 => x"74",
          5192 => x"05",
          5193 => x"17",
          5194 => x"70",
          5195 => x"52",
          5196 => x"73",
          5197 => x"c8",
          5198 => x"33",
          5199 => x"73",
          5200 => x"81",
          5201 => x"80",
          5202 => x"02",
          5203 => x"76",
          5204 => x"51",
          5205 => x"2e",
          5206 => x"87",
          5207 => x"57",
          5208 => x"79",
          5209 => x"80",
          5210 => x"70",
          5211 => x"ba",
          5212 => x"8c",
          5213 => x"82",
          5214 => x"80",
          5215 => x"52",
          5216 => x"bf",
          5217 => x"8c",
          5218 => x"82",
          5219 => x"8d",
          5220 => x"c4",
          5221 => x"e5",
          5222 => x"c6",
          5223 => x"dc",
          5224 => x"09",
          5225 => x"cc",
          5226 => x"76",
          5227 => x"c4",
          5228 => x"74",
          5229 => x"b0",
          5230 => x"dc",
          5231 => x"8c",
          5232 => x"38",
          5233 => x"8c",
          5234 => x"67",
          5235 => x"db",
          5236 => x"88",
          5237 => x"34",
          5238 => x"52",
          5239 => x"ab",
          5240 => x"54",
          5241 => x"15",
          5242 => x"ff",
          5243 => x"82",
          5244 => x"54",
          5245 => x"82",
          5246 => x"9c",
          5247 => x"f2",
          5248 => x"62",
          5249 => x"80",
          5250 => x"93",
          5251 => x"55",
          5252 => x"5e",
          5253 => x"3f",
          5254 => x"08",
          5255 => x"dc",
          5256 => x"38",
          5257 => x"58",
          5258 => x"38",
          5259 => x"97",
          5260 => x"08",
          5261 => x"38",
          5262 => x"70",
          5263 => x"81",
          5264 => x"55",
          5265 => x"87",
          5266 => x"39",
          5267 => x"90",
          5268 => x"82",
          5269 => x"8a",
          5270 => x"89",
          5271 => x"7f",
          5272 => x"56",
          5273 => x"3f",
          5274 => x"06",
          5275 => x"72",
          5276 => x"82",
          5277 => x"05",
          5278 => x"7c",
          5279 => x"55",
          5280 => x"27",
          5281 => x"16",
          5282 => x"83",
          5283 => x"76",
          5284 => x"80",
          5285 => x"79",
          5286 => x"99",
          5287 => x"7f",
          5288 => x"14",
          5289 => x"83",
          5290 => x"82",
          5291 => x"81",
          5292 => x"38",
          5293 => x"08",
          5294 => x"95",
          5295 => x"dc",
          5296 => x"81",
          5297 => x"7b",
          5298 => x"06",
          5299 => x"39",
          5300 => x"56",
          5301 => x"09",
          5302 => x"b9",
          5303 => x"80",
          5304 => x"80",
          5305 => x"78",
          5306 => x"7a",
          5307 => x"38",
          5308 => x"73",
          5309 => x"81",
          5310 => x"ff",
          5311 => x"74",
          5312 => x"ff",
          5313 => x"82",
          5314 => x"58",
          5315 => x"08",
          5316 => x"74",
          5317 => x"16",
          5318 => x"73",
          5319 => x"39",
          5320 => x"7e",
          5321 => x"0c",
          5322 => x"2e",
          5323 => x"88",
          5324 => x"8c",
          5325 => x"1a",
          5326 => x"07",
          5327 => x"1b",
          5328 => x"08",
          5329 => x"16",
          5330 => x"75",
          5331 => x"38",
          5332 => x"90",
          5333 => x"15",
          5334 => x"54",
          5335 => x"34",
          5336 => x"82",
          5337 => x"90",
          5338 => x"e9",
          5339 => x"6d",
          5340 => x"80",
          5341 => x"9d",
          5342 => x"5c",
          5343 => x"3f",
          5344 => x"0b",
          5345 => x"08",
          5346 => x"38",
          5347 => x"08",
          5348 => x"8d",
          5349 => x"08",
          5350 => x"80",
          5351 => x"80",
          5352 => x"8c",
          5353 => x"ff",
          5354 => x"52",
          5355 => x"a0",
          5356 => x"8c",
          5357 => x"ff",
          5358 => x"06",
          5359 => x"56",
          5360 => x"38",
          5361 => x"70",
          5362 => x"55",
          5363 => x"8b",
          5364 => x"3d",
          5365 => x"83",
          5366 => x"ff",
          5367 => x"82",
          5368 => x"99",
          5369 => x"74",
          5370 => x"38",
          5371 => x"80",
          5372 => x"ff",
          5373 => x"55",
          5374 => x"83",
          5375 => x"78",
          5376 => x"38",
          5377 => x"26",
          5378 => x"81",
          5379 => x"8b",
          5380 => x"79",
          5381 => x"80",
          5382 => x"93",
          5383 => x"39",
          5384 => x"6e",
          5385 => x"89",
          5386 => x"48",
          5387 => x"83",
          5388 => x"61",
          5389 => x"25",
          5390 => x"55",
          5391 => x"8a",
          5392 => x"3d",
          5393 => x"81",
          5394 => x"ff",
          5395 => x"81",
          5396 => x"dc",
          5397 => x"38",
          5398 => x"70",
          5399 => x"8c",
          5400 => x"56",
          5401 => x"38",
          5402 => x"55",
          5403 => x"75",
          5404 => x"38",
          5405 => x"70",
          5406 => x"ff",
          5407 => x"83",
          5408 => x"78",
          5409 => x"89",
          5410 => x"81",
          5411 => x"06",
          5412 => x"80",
          5413 => x"77",
          5414 => x"74",
          5415 => x"8d",
          5416 => x"06",
          5417 => x"2e",
          5418 => x"77",
          5419 => x"93",
          5420 => x"74",
          5421 => x"cb",
          5422 => x"7d",
          5423 => x"81",
          5424 => x"38",
          5425 => x"66",
          5426 => x"81",
          5427 => x"90",
          5428 => x"74",
          5429 => x"38",
          5430 => x"98",
          5431 => x"90",
          5432 => x"82",
          5433 => x"57",
          5434 => x"80",
          5435 => x"76",
          5436 => x"38",
          5437 => x"51",
          5438 => x"3f",
          5439 => x"08",
          5440 => x"87",
          5441 => x"2a",
          5442 => x"5c",
          5443 => x"8c",
          5444 => x"80",
          5445 => x"44",
          5446 => x"0a",
          5447 => x"ec",
          5448 => x"39",
          5449 => x"66",
          5450 => x"81",
          5451 => x"80",
          5452 => x"74",
          5453 => x"38",
          5454 => x"98",
          5455 => x"80",
          5456 => x"82",
          5457 => x"57",
          5458 => x"80",
          5459 => x"76",
          5460 => x"38",
          5461 => x"51",
          5462 => x"3f",
          5463 => x"08",
          5464 => x"57",
          5465 => x"08",
          5466 => x"96",
          5467 => x"82",
          5468 => x"10",
          5469 => x"08",
          5470 => x"72",
          5471 => x"59",
          5472 => x"ff",
          5473 => x"5d",
          5474 => x"44",
          5475 => x"11",
          5476 => x"70",
          5477 => x"71",
          5478 => x"06",
          5479 => x"52",
          5480 => x"40",
          5481 => x"09",
          5482 => x"38",
          5483 => x"18",
          5484 => x"39",
          5485 => x"79",
          5486 => x"70",
          5487 => x"58",
          5488 => x"76",
          5489 => x"38",
          5490 => x"7d",
          5491 => x"70",
          5492 => x"55",
          5493 => x"3f",
          5494 => x"08",
          5495 => x"2e",
          5496 => x"9b",
          5497 => x"dc",
          5498 => x"f5",
          5499 => x"38",
          5500 => x"38",
          5501 => x"59",
          5502 => x"38",
          5503 => x"7d",
          5504 => x"81",
          5505 => x"38",
          5506 => x"0b",
          5507 => x"08",
          5508 => x"78",
          5509 => x"1a",
          5510 => x"c0",
          5511 => x"74",
          5512 => x"39",
          5513 => x"55",
          5514 => x"8f",
          5515 => x"fd",
          5516 => x"8c",
          5517 => x"f5",
          5518 => x"78",
          5519 => x"79",
          5520 => x"80",
          5521 => x"f1",
          5522 => x"39",
          5523 => x"81",
          5524 => x"06",
          5525 => x"55",
          5526 => x"27",
          5527 => x"81",
          5528 => x"56",
          5529 => x"38",
          5530 => x"80",
          5531 => x"ff",
          5532 => x"8b",
          5533 => x"a8",
          5534 => x"ff",
          5535 => x"84",
          5536 => x"1b",
          5537 => x"b3",
          5538 => x"1c",
          5539 => x"ff",
          5540 => x"8e",
          5541 => x"a1",
          5542 => x"0b",
          5543 => x"7d",
          5544 => x"30",
          5545 => x"84",
          5546 => x"51",
          5547 => x"51",
          5548 => x"3f",
          5549 => x"83",
          5550 => x"90",
          5551 => x"ff",
          5552 => x"93",
          5553 => x"a0",
          5554 => x"39",
          5555 => x"1b",
          5556 => x"85",
          5557 => x"95",
          5558 => x"52",
          5559 => x"ff",
          5560 => x"81",
          5561 => x"1b",
          5562 => x"cf",
          5563 => x"9c",
          5564 => x"a0",
          5565 => x"83",
          5566 => x"06",
          5567 => x"82",
          5568 => x"52",
          5569 => x"51",
          5570 => x"3f",
          5571 => x"1b",
          5572 => x"c5",
          5573 => x"ac",
          5574 => x"a0",
          5575 => x"52",
          5576 => x"ff",
          5577 => x"86",
          5578 => x"51",
          5579 => x"3f",
          5580 => x"80",
          5581 => x"a9",
          5582 => x"1c",
          5583 => x"81",
          5584 => x"80",
          5585 => x"ae",
          5586 => x"b2",
          5587 => x"1b",
          5588 => x"85",
          5589 => x"ff",
          5590 => x"96",
          5591 => x"9f",
          5592 => x"80",
          5593 => x"34",
          5594 => x"1c",
          5595 => x"81",
          5596 => x"ab",
          5597 => x"a0",
          5598 => x"d4",
          5599 => x"fe",
          5600 => x"59",
          5601 => x"3f",
          5602 => x"53",
          5603 => x"51",
          5604 => x"3f",
          5605 => x"8c",
          5606 => x"e7",
          5607 => x"2e",
          5608 => x"80",
          5609 => x"54",
          5610 => x"53",
          5611 => x"51",
          5612 => x"3f",
          5613 => x"80",
          5614 => x"ff",
          5615 => x"84",
          5616 => x"d2",
          5617 => x"ff",
          5618 => x"86",
          5619 => x"f2",
          5620 => x"1b",
          5621 => x"81",
          5622 => x"52",
          5623 => x"51",
          5624 => x"3f",
          5625 => x"ec",
          5626 => x"9e",
          5627 => x"d4",
          5628 => x"51",
          5629 => x"3f",
          5630 => x"87",
          5631 => x"52",
          5632 => x"9a",
          5633 => x"54",
          5634 => x"7a",
          5635 => x"ff",
          5636 => x"65",
          5637 => x"7a",
          5638 => x"8f",
          5639 => x"80",
          5640 => x"2e",
          5641 => x"9a",
          5642 => x"7a",
          5643 => x"a9",
          5644 => x"84",
          5645 => x"9e",
          5646 => x"0a",
          5647 => x"51",
          5648 => x"ff",
          5649 => x"7d",
          5650 => x"38",
          5651 => x"52",
          5652 => x"9e",
          5653 => x"55",
          5654 => x"62",
          5655 => x"74",
          5656 => x"75",
          5657 => x"7e",
          5658 => x"fe",
          5659 => x"dc",
          5660 => x"38",
          5661 => x"82",
          5662 => x"52",
          5663 => x"9e",
          5664 => x"16",
          5665 => x"56",
          5666 => x"38",
          5667 => x"77",
          5668 => x"8d",
          5669 => x"7d",
          5670 => x"38",
          5671 => x"57",
          5672 => x"83",
          5673 => x"76",
          5674 => x"7a",
          5675 => x"ff",
          5676 => x"82",
          5677 => x"81",
          5678 => x"16",
          5679 => x"56",
          5680 => x"38",
          5681 => x"83",
          5682 => x"86",
          5683 => x"ff",
          5684 => x"38",
          5685 => x"82",
          5686 => x"81",
          5687 => x"06",
          5688 => x"fe",
          5689 => x"53",
          5690 => x"51",
          5691 => x"3f",
          5692 => x"52",
          5693 => x"9c",
          5694 => x"be",
          5695 => x"75",
          5696 => x"81",
          5697 => x"0b",
          5698 => x"77",
          5699 => x"75",
          5700 => x"60",
          5701 => x"80",
          5702 => x"75",
          5703 => x"bc",
          5704 => x"85",
          5705 => x"8c",
          5706 => x"2a",
          5707 => x"75",
          5708 => x"82",
          5709 => x"87",
          5710 => x"52",
          5711 => x"51",
          5712 => x"3f",
          5713 => x"ca",
          5714 => x"9c",
          5715 => x"54",
          5716 => x"52",
          5717 => x"98",
          5718 => x"56",
          5719 => x"08",
          5720 => x"53",
          5721 => x"51",
          5722 => x"3f",
          5723 => x"8c",
          5724 => x"38",
          5725 => x"56",
          5726 => x"56",
          5727 => x"8c",
          5728 => x"75",
          5729 => x"0c",
          5730 => x"04",
          5731 => x"7d",
          5732 => x"80",
          5733 => x"05",
          5734 => x"76",
          5735 => x"38",
          5736 => x"11",
          5737 => x"53",
          5738 => x"79",
          5739 => x"3f",
          5740 => x"09",
          5741 => x"38",
          5742 => x"55",
          5743 => x"db",
          5744 => x"70",
          5745 => x"34",
          5746 => x"74",
          5747 => x"81",
          5748 => x"80",
          5749 => x"55",
          5750 => x"76",
          5751 => x"8c",
          5752 => x"3d",
          5753 => x"3d",
          5754 => x"84",
          5755 => x"33",
          5756 => x"8a",
          5757 => x"06",
          5758 => x"52",
          5759 => x"3f",
          5760 => x"56",
          5761 => x"be",
          5762 => x"08",
          5763 => x"05",
          5764 => x"75",
          5765 => x"56",
          5766 => x"a1",
          5767 => x"fc",
          5768 => x"53",
          5769 => x"76",
          5770 => x"dc",
          5771 => x"32",
          5772 => x"72",
          5773 => x"70",
          5774 => x"56",
          5775 => x"18",
          5776 => x"88",
          5777 => x"3d",
          5778 => x"3d",
          5779 => x"11",
          5780 => x"80",
          5781 => x"38",
          5782 => x"05",
          5783 => x"8c",
          5784 => x"08",
          5785 => x"3f",
          5786 => x"08",
          5787 => x"16",
          5788 => x"09",
          5789 => x"38",
          5790 => x"55",
          5791 => x"55",
          5792 => x"dc",
          5793 => x"0d",
          5794 => x"0d",
          5795 => x"cc",
          5796 => x"73",
          5797 => x"93",
          5798 => x"0c",
          5799 => x"04",
          5800 => x"02",
          5801 => x"33",
          5802 => x"3d",
          5803 => x"54",
          5804 => x"52",
          5805 => x"ae",
          5806 => x"ff",
          5807 => x"3d",
          5808 => x"3d",
          5809 => x"08",
          5810 => x"59",
          5811 => x"80",
          5812 => x"39",
          5813 => x"0c",
          5814 => x"54",
          5815 => x"74",
          5816 => x"a0",
          5817 => x"06",
          5818 => x"15",
          5819 => x"80",
          5820 => x"29",
          5821 => x"05",
          5822 => x"56",
          5823 => x"3f",
          5824 => x"08",
          5825 => x"08",
          5826 => x"76",
          5827 => x"fe",
          5828 => x"82",
          5829 => x"8b",
          5830 => x"33",
          5831 => x"2e",
          5832 => x"81",
          5833 => x"ff",
          5834 => x"98",
          5835 => x"38",
          5836 => x"82",
          5837 => x"8a",
          5838 => x"ff",
          5839 => x"52",
          5840 => x"81",
          5841 => x"84",
          5842 => x"94",
          5843 => x"08",
          5844 => x"c8",
          5845 => x"39",
          5846 => x"51",
          5847 => x"81",
          5848 => x"80",
          5849 => x"fd",
          5850 => x"eb",
          5851 => x"8c",
          5852 => x"39",
          5853 => x"51",
          5854 => x"81",
          5855 => x"80",
          5856 => x"fe",
          5857 => x"cf",
          5858 => x"d8",
          5859 => x"39",
          5860 => x"51",
          5861 => x"81",
          5862 => x"bb",
          5863 => x"a4",
          5864 => x"81",
          5865 => x"af",
          5866 => x"e4",
          5867 => x"81",
          5868 => x"a3",
          5869 => x"98",
          5870 => x"82",
          5871 => x"97",
          5872 => x"c4",
          5873 => x"82",
          5874 => x"8b",
          5875 => x"f4",
          5876 => x"82",
          5877 => x"fe",
          5878 => x"83",
          5879 => x"fb",
          5880 => x"79",
          5881 => x"87",
          5882 => x"38",
          5883 => x"87",
          5884 => x"91",
          5885 => x"52",
          5886 => x"d2",
          5887 => x"8c",
          5888 => x"75",
          5889 => x"d4",
          5890 => x"dc",
          5891 => x"53",
          5892 => x"81",
          5893 => x"f7",
          5894 => x"3d",
          5895 => x"3d",
          5896 => x"84",
          5897 => x"05",
          5898 => x"80",
          5899 => x"70",
          5900 => x"25",
          5901 => x"59",
          5902 => x"87",
          5903 => x"38",
          5904 => x"76",
          5905 => x"ff",
          5906 => x"93",
          5907 => x"80",
          5908 => x"76",
          5909 => x"70",
          5910 => x"bf",
          5911 => x"8c",
          5912 => x"82",
          5913 => x"b8",
          5914 => x"dc",
          5915 => x"98",
          5916 => x"8c",
          5917 => x"96",
          5918 => x"54",
          5919 => x"77",
          5920 => x"c4",
          5921 => x"8c",
          5922 => x"82",
          5923 => x"90",
          5924 => x"74",
          5925 => x"38",
          5926 => x"19",
          5927 => x"39",
          5928 => x"05",
          5929 => x"3f",
          5930 => x"78",
          5931 => x"7b",
          5932 => x"2a",
          5933 => x"57",
          5934 => x"80",
          5935 => x"82",
          5936 => x"87",
          5937 => x"08",
          5938 => x"fe",
          5939 => x"56",
          5940 => x"dc",
          5941 => x"0d",
          5942 => x"0d",
          5943 => x"05",
          5944 => x"57",
          5945 => x"80",
          5946 => x"79",
          5947 => x"3f",
          5948 => x"08",
          5949 => x"80",
          5950 => x"75",
          5951 => x"38",
          5952 => x"55",
          5953 => x"8c",
          5954 => x"52",
          5955 => x"2d",
          5956 => x"08",
          5957 => x"77",
          5958 => x"8c",
          5959 => x"3d",
          5960 => x"3d",
          5961 => x"63",
          5962 => x"80",
          5963 => x"73",
          5964 => x"41",
          5965 => x"5e",
          5966 => x"52",
          5967 => x"51",
          5968 => x"3f",
          5969 => x"51",
          5970 => x"3f",
          5971 => x"79",
          5972 => x"38",
          5973 => x"89",
          5974 => x"2e",
          5975 => x"c6",
          5976 => x"53",
          5977 => x"8e",
          5978 => x"52",
          5979 => x"51",
          5980 => x"3f",
          5981 => x"81",
          5982 => x"ef",
          5983 => x"15",
          5984 => x"39",
          5985 => x"72",
          5986 => x"38",
          5987 => x"82",
          5988 => x"fe",
          5989 => x"89",
          5990 => x"d0",
          5991 => x"e8",
          5992 => x"55",
          5993 => x"18",
          5994 => x"27",
          5995 => x"33",
          5996 => x"dc",
          5997 => x"b4",
          5998 => x"82",
          5999 => x"fe",
          6000 => x"81",
          6001 => x"51",
          6002 => x"3f",
          6003 => x"82",
          6004 => x"fe",
          6005 => x"80",
          6006 => x"27",
          6007 => x"18",
          6008 => x"53",
          6009 => x"7a",
          6010 => x"81",
          6011 => x"9f",
          6012 => x"38",
          6013 => x"73",
          6014 => x"ff",
          6015 => x"72",
          6016 => x"38",
          6017 => x"26",
          6018 => x"51",
          6019 => x"51",
          6020 => x"3f",
          6021 => x"c1",
          6022 => x"ec",
          6023 => x"e8",
          6024 => x"79",
          6025 => x"fe",
          6026 => x"82",
          6027 => x"98",
          6028 => x"2c",
          6029 => x"a0",
          6030 => x"06",
          6031 => x"de",
          6032 => x"8c",
          6033 => x"2b",
          6034 => x"70",
          6035 => x"30",
          6036 => x"70",
          6037 => x"07",
          6038 => x"06",
          6039 => x"59",
          6040 => x"80",
          6041 => x"38",
          6042 => x"09",
          6043 => x"38",
          6044 => x"39",
          6045 => x"72",
          6046 => x"be",
          6047 => x"72",
          6048 => x"0c",
          6049 => x"04",
          6050 => x"02",
          6051 => x"82",
          6052 => x"82",
          6053 => x"55",
          6054 => x"3f",
          6055 => x"22",
          6056 => x"96",
          6057 => x"80",
          6058 => x"8c",
          6059 => x"8d",
          6060 => x"82",
          6061 => x"f2",
          6062 => x"80",
          6063 => x"fe",
          6064 => x"86",
          6065 => x"fe",
          6066 => x"c0",
          6067 => x"53",
          6068 => x"3f",
          6069 => x"d9",
          6070 => x"82",
          6071 => x"db",
          6072 => x"51",
          6073 => x"3f",
          6074 => x"70",
          6075 => x"52",
          6076 => x"95",
          6077 => x"fe",
          6078 => x"82",
          6079 => x"fe",
          6080 => x"80",
          6081 => x"8b",
          6082 => x"2a",
          6083 => x"51",
          6084 => x"2e",
          6085 => x"51",
          6086 => x"3f",
          6087 => x"51",
          6088 => x"3f",
          6089 => x"d8",
          6090 => x"83",
          6091 => x"06",
          6092 => x"80",
          6093 => x"81",
          6094 => x"d7",
          6095 => x"ec",
          6096 => x"cf",
          6097 => x"fe",
          6098 => x"72",
          6099 => x"81",
          6100 => x"71",
          6101 => x"38",
          6102 => x"d8",
          6103 => x"83",
          6104 => x"da",
          6105 => x"51",
          6106 => x"3f",
          6107 => x"70",
          6108 => x"52",
          6109 => x"95",
          6110 => x"fe",
          6111 => x"82",
          6112 => x"fe",
          6113 => x"80",
          6114 => x"87",
          6115 => x"2a",
          6116 => x"51",
          6117 => x"2e",
          6118 => x"51",
          6119 => x"3f",
          6120 => x"51",
          6121 => x"3f",
          6122 => x"d7",
          6123 => x"87",
          6124 => x"06",
          6125 => x"80",
          6126 => x"81",
          6127 => x"d3",
          6128 => x"bc",
          6129 => x"cb",
          6130 => x"fe",
          6131 => x"72",
          6132 => x"81",
          6133 => x"71",
          6134 => x"38",
          6135 => x"d7",
          6136 => x"83",
          6137 => x"d9",
          6138 => x"51",
          6139 => x"3f",
          6140 => x"3f",
          6141 => x"04",
          6142 => x"77",
          6143 => x"a3",
          6144 => x"55",
          6145 => x"52",
          6146 => x"ce",
          6147 => x"89",
          6148 => x"73",
          6149 => x"53",
          6150 => x"52",
          6151 => x"51",
          6152 => x"3f",
          6153 => x"08",
          6154 => x"8c",
          6155 => x"80",
          6156 => x"31",
          6157 => x"73",
          6158 => x"34",
          6159 => x"33",
          6160 => x"2e",
          6161 => x"ac",
          6162 => x"f4",
          6163 => x"75",
          6164 => x"3f",
          6165 => x"08",
          6166 => x"38",
          6167 => x"08",
          6168 => x"a4",
          6169 => x"82",
          6170 => x"c4",
          6171 => x"0b",
          6172 => x"34",
          6173 => x"33",
          6174 => x"2e",
          6175 => x"89",
          6176 => x"75",
          6177 => x"e4",
          6178 => x"82",
          6179 => x"87",
          6180 => x"ce",
          6181 => x"70",
          6182 => x"f0",
          6183 => x"81",
          6184 => x"ff",
          6185 => x"82",
          6186 => x"81",
          6187 => x"78",
          6188 => x"81",
          6189 => x"82",
          6190 => x"96",
          6191 => x"59",
          6192 => x"3f",
          6193 => x"52",
          6194 => x"51",
          6195 => x"3f",
          6196 => x"08",
          6197 => x"38",
          6198 => x"51",
          6199 => x"81",
          6200 => x"82",
          6201 => x"fe",
          6202 => x"96",
          6203 => x"5a",
          6204 => x"79",
          6205 => x"3f",
          6206 => x"84",
          6207 => x"c2",
          6208 => x"dc",
          6209 => x"70",
          6210 => x"59",
          6211 => x"2e",
          6212 => x"78",
          6213 => x"b2",
          6214 => x"2e",
          6215 => x"78",
          6216 => x"38",
          6217 => x"ff",
          6218 => x"bc",
          6219 => x"38",
          6220 => x"78",
          6221 => x"83",
          6222 => x"80",
          6223 => x"dd",
          6224 => x"2e",
          6225 => x"8a",
          6226 => x"80",
          6227 => x"ea",
          6228 => x"f9",
          6229 => x"78",
          6230 => x"88",
          6231 => x"80",
          6232 => x"b1",
          6233 => x"39",
          6234 => x"2e",
          6235 => x"78",
          6236 => x"8b",
          6237 => x"82",
          6238 => x"38",
          6239 => x"78",
          6240 => x"8a",
          6241 => x"93",
          6242 => x"ff",
          6243 => x"ff",
          6244 => x"fe",
          6245 => x"82",
          6246 => x"80",
          6247 => x"38",
          6248 => x"fc",
          6249 => x"84",
          6250 => x"ee",
          6251 => x"8c",
          6252 => x"2e",
          6253 => x"b4",
          6254 => x"11",
          6255 => x"05",
          6256 => x"9d",
          6257 => x"dc",
          6258 => x"82",
          6259 => x"42",
          6260 => x"51",
          6261 => x"3f",
          6262 => x"5a",
          6263 => x"81",
          6264 => x"59",
          6265 => x"84",
          6266 => x"7a",
          6267 => x"38",
          6268 => x"b4",
          6269 => x"11",
          6270 => x"05",
          6271 => x"e1",
          6272 => x"dc",
          6273 => x"fd",
          6274 => x"3d",
          6275 => x"53",
          6276 => x"51",
          6277 => x"3f",
          6278 => x"08",
          6279 => x"c3",
          6280 => x"fe",
          6281 => x"ff",
          6282 => x"fe",
          6283 => x"82",
          6284 => x"80",
          6285 => x"38",
          6286 => x"51",
          6287 => x"3f",
          6288 => x"63",
          6289 => x"38",
          6290 => x"70",
          6291 => x"33",
          6292 => x"81",
          6293 => x"39",
          6294 => x"80",
          6295 => x"84",
          6296 => x"ec",
          6297 => x"8c",
          6298 => x"2e",
          6299 => x"b4",
          6300 => x"11",
          6301 => x"05",
          6302 => x"e5",
          6303 => x"dc",
          6304 => x"fc",
          6305 => x"3d",
          6306 => x"53",
          6307 => x"51",
          6308 => x"3f",
          6309 => x"08",
          6310 => x"c7",
          6311 => x"fc",
          6312 => x"e4",
          6313 => x"79",
          6314 => x"38",
          6315 => x"7b",
          6316 => x"5b",
          6317 => x"92",
          6318 => x"7a",
          6319 => x"53",
          6320 => x"85",
          6321 => x"ea",
          6322 => x"1a",
          6323 => x"43",
          6324 => x"82",
          6325 => x"82",
          6326 => x"3d",
          6327 => x"53",
          6328 => x"51",
          6329 => x"3f",
          6330 => x"08",
          6331 => x"82",
          6332 => x"59",
          6333 => x"89",
          6334 => x"d8",
          6335 => x"cd",
          6336 => x"a1",
          6337 => x"80",
          6338 => x"82",
          6339 => x"44",
          6340 => x"88",
          6341 => x"78",
          6342 => x"38",
          6343 => x"08",
          6344 => x"82",
          6345 => x"59",
          6346 => x"88",
          6347 => x"f0",
          6348 => x"39",
          6349 => x"33",
          6350 => x"2e",
          6351 => x"87",
          6352 => x"89",
          6353 => x"88",
          6354 => x"05",
          6355 => x"fe",
          6356 => x"ff",
          6357 => x"fe",
          6358 => x"82",
          6359 => x"80",
          6360 => x"88",
          6361 => x"78",
          6362 => x"38",
          6363 => x"08",
          6364 => x"39",
          6365 => x"33",
          6366 => x"2e",
          6367 => x"87",
          6368 => x"bb",
          6369 => x"a2",
          6370 => x"80",
          6371 => x"82",
          6372 => x"43",
          6373 => x"88",
          6374 => x"78",
          6375 => x"38",
          6376 => x"08",
          6377 => x"82",
          6378 => x"59",
          6379 => x"88",
          6380 => x"fc",
          6381 => x"39",
          6382 => x"08",
          6383 => x"b4",
          6384 => x"11",
          6385 => x"05",
          6386 => x"95",
          6387 => x"dc",
          6388 => x"a7",
          6389 => x"5c",
          6390 => x"2e",
          6391 => x"5c",
          6392 => x"70",
          6393 => x"07",
          6394 => x"7f",
          6395 => x"5a",
          6396 => x"2e",
          6397 => x"a0",
          6398 => x"88",
          6399 => x"a8",
          6400 => x"84",
          6401 => x"63",
          6402 => x"62",
          6403 => x"f2",
          6404 => x"85",
          6405 => x"e1",
          6406 => x"c7",
          6407 => x"ff",
          6408 => x"ff",
          6409 => x"fe",
          6410 => x"82",
          6411 => x"80",
          6412 => x"38",
          6413 => x"fc",
          6414 => x"84",
          6415 => x"e9",
          6416 => x"8c",
          6417 => x"2e",
          6418 => x"59",
          6419 => x"05",
          6420 => x"63",
          6421 => x"b4",
          6422 => x"11",
          6423 => x"05",
          6424 => x"fd",
          6425 => x"dc",
          6426 => x"f8",
          6427 => x"70",
          6428 => x"82",
          6429 => x"fe",
          6430 => x"80",
          6431 => x"51",
          6432 => x"3f",
          6433 => x"33",
          6434 => x"2e",
          6435 => x"9f",
          6436 => x"38",
          6437 => x"fc",
          6438 => x"84",
          6439 => x"e8",
          6440 => x"8c",
          6441 => x"2e",
          6442 => x"59",
          6443 => x"05",
          6444 => x"63",
          6445 => x"ff",
          6446 => x"85",
          6447 => x"e0",
          6448 => x"aa",
          6449 => x"fe",
          6450 => x"ff",
          6451 => x"fe",
          6452 => x"82",
          6453 => x"80",
          6454 => x"38",
          6455 => x"f0",
          6456 => x"84",
          6457 => x"e9",
          6458 => x"8c",
          6459 => x"2e",
          6460 => x"59",
          6461 => x"22",
          6462 => x"05",
          6463 => x"41",
          6464 => x"f0",
          6465 => x"84",
          6466 => x"e9",
          6467 => x"8c",
          6468 => x"38",
          6469 => x"60",
          6470 => x"52",
          6471 => x"51",
          6472 => x"3f",
          6473 => x"79",
          6474 => x"9a",
          6475 => x"79",
          6476 => x"ae",
          6477 => x"38",
          6478 => x"87",
          6479 => x"05",
          6480 => x"b4",
          6481 => x"11",
          6482 => x"05",
          6483 => x"83",
          6484 => x"dc",
          6485 => x"92",
          6486 => x"02",
          6487 => x"79",
          6488 => x"5b",
          6489 => x"ff",
          6490 => x"85",
          6491 => x"df",
          6492 => x"a3",
          6493 => x"fe",
          6494 => x"ff",
          6495 => x"fe",
          6496 => x"82",
          6497 => x"80",
          6498 => x"38",
          6499 => x"f0",
          6500 => x"84",
          6501 => x"e8",
          6502 => x"8c",
          6503 => x"2e",
          6504 => x"60",
          6505 => x"60",
          6506 => x"b4",
          6507 => x"11",
          6508 => x"05",
          6509 => x"9b",
          6510 => x"dc",
          6511 => x"f6",
          6512 => x"70",
          6513 => x"82",
          6514 => x"fe",
          6515 => x"80",
          6516 => x"51",
          6517 => x"3f",
          6518 => x"33",
          6519 => x"2e",
          6520 => x"9f",
          6521 => x"38",
          6522 => x"f0",
          6523 => x"84",
          6524 => x"e7",
          6525 => x"8c",
          6526 => x"2e",
          6527 => x"60",
          6528 => x"60",
          6529 => x"ff",
          6530 => x"85",
          6531 => x"dd",
          6532 => x"ae",
          6533 => x"ff",
          6534 => x"ff",
          6535 => x"fe",
          6536 => x"82",
          6537 => x"80",
          6538 => x"38",
          6539 => x"85",
          6540 => x"e3",
          6541 => x"59",
          6542 => x"3d",
          6543 => x"53",
          6544 => x"51",
          6545 => x"3f",
          6546 => x"08",
          6547 => x"93",
          6548 => x"82",
          6549 => x"fe",
          6550 => x"63",
          6551 => x"82",
          6552 => x"80",
          6553 => x"38",
          6554 => x"08",
          6555 => x"a8",
          6556 => x"f8",
          6557 => x"39",
          6558 => x"51",
          6559 => x"3f",
          6560 => x"3f",
          6561 => x"82",
          6562 => x"fe",
          6563 => x"80",
          6564 => x"39",
          6565 => x"3f",
          6566 => x"79",
          6567 => x"59",
          6568 => x"f4",
          6569 => x"7d",
          6570 => x"80",
          6571 => x"38",
          6572 => x"84",
          6573 => x"c6",
          6574 => x"8c",
          6575 => x"81",
          6576 => x"2e",
          6577 => x"82",
          6578 => x"7a",
          6579 => x"38",
          6580 => x"7a",
          6581 => x"38",
          6582 => x"82",
          6583 => x"7b",
          6584 => x"f8",
          6585 => x"82",
          6586 => x"b4",
          6587 => x"05",
          6588 => x"8e",
          6589 => x"82",
          6590 => x"b4",
          6591 => x"05",
          6592 => x"fe",
          6593 => x"7b",
          6594 => x"f8",
          6595 => x"82",
          6596 => x"b4",
          6597 => x"05",
          6598 => x"e6",
          6599 => x"7b",
          6600 => x"82",
          6601 => x"b4",
          6602 => x"05",
          6603 => x"d2",
          6604 => x"d8",
          6605 => x"a4",
          6606 => x"64",
          6607 => x"83",
          6608 => x"83",
          6609 => x"b4",
          6610 => x"05",
          6611 => x"3f",
          6612 => x"08",
          6613 => x"08",
          6614 => x"70",
          6615 => x"25",
          6616 => x"5f",
          6617 => x"83",
          6618 => x"81",
          6619 => x"06",
          6620 => x"2e",
          6621 => x"1b",
          6622 => x"06",
          6623 => x"fe",
          6624 => x"81",
          6625 => x"32",
          6626 => x"8a",
          6627 => x"2e",
          6628 => x"f2",
          6629 => x"87",
          6630 => x"e0",
          6631 => x"c3",
          6632 => x"0d",
          6633 => x"8d",
          6634 => x"c0",
          6635 => x"08",
          6636 => x"84",
          6637 => x"51",
          6638 => x"3f",
          6639 => x"08",
          6640 => x"08",
          6641 => x"84",
          6642 => x"51",
          6643 => x"3f",
          6644 => x"dc",
          6645 => x"0c",
          6646 => x"9c",
          6647 => x"55",
          6648 => x"52",
          6649 => x"ba",
          6650 => x"8c",
          6651 => x"2b",
          6652 => x"53",
          6653 => x"52",
          6654 => x"ba",
          6655 => x"82",
          6656 => x"07",
          6657 => x"80",
          6658 => x"c0",
          6659 => x"8c",
          6660 => x"87",
          6661 => x"0c",
          6662 => x"82",
          6663 => x"ba",
          6664 => x"8c",
          6665 => x"cb",
          6666 => x"d4",
          6667 => x"87",
          6668 => x"d9",
          6669 => x"87",
          6670 => x"d9",
          6671 => x"dd",
          6672 => x"d4",
          6673 => x"51",
          6674 => x"f0",
          6675 => x"04",
          6676 => x"22",
          6677 => x"22",
          6678 => x"22",
          6679 => x"22",
          6680 => x"22",
          6681 => x"2f",
          6682 => x"30",
          6683 => x"31",
          6684 => x"31",
          6685 => x"31",
          6686 => x"32",
          6687 => x"2e",
          6688 => x"2e",
          6689 => x"32",
          6690 => x"32",
          6691 => x"33",
          6692 => x"33",
          6693 => x"6b",
          6694 => x"6b",
          6695 => x"6b",
          6696 => x"6b",
          6697 => x"6b",
          6698 => x"6b",
          6699 => x"6b",
          6700 => x"6b",
          6701 => x"6b",
          6702 => x"6b",
          6703 => x"6b",
          6704 => x"6b",
          6705 => x"6b",
          6706 => x"6b",
          6707 => x"6b",
          6708 => x"6b",
          6709 => x"6b",
          6710 => x"6b",
          6711 => x"6b",
          6712 => x"6b",
          6713 => x"2f",
          6714 => x"25",
          6715 => x"64",
          6716 => x"3a",
          6717 => x"25",
          6718 => x"0a",
          6719 => x"43",
          6720 => x"6e",
          6721 => x"75",
          6722 => x"69",
          6723 => x"00",
          6724 => x"66",
          6725 => x"20",
          6726 => x"20",
          6727 => x"66",
          6728 => x"00",
          6729 => x"44",
          6730 => x"63",
          6731 => x"69",
          6732 => x"65",
          6733 => x"74",
          6734 => x"0a",
          6735 => x"20",
          6736 => x"20",
          6737 => x"41",
          6738 => x"28",
          6739 => x"58",
          6740 => x"38",
          6741 => x"0a",
          6742 => x"20",
          6743 => x"52",
          6744 => x"20",
          6745 => x"28",
          6746 => x"58",
          6747 => x"38",
          6748 => x"0a",
          6749 => x"20",
          6750 => x"53",
          6751 => x"52",
          6752 => x"28",
          6753 => x"58",
          6754 => x"38",
          6755 => x"0a",
          6756 => x"20",
          6757 => x"41",
          6758 => x"20",
          6759 => x"28",
          6760 => x"58",
          6761 => x"38",
          6762 => x"0a",
          6763 => x"20",
          6764 => x"4d",
          6765 => x"20",
          6766 => x"28",
          6767 => x"58",
          6768 => x"38",
          6769 => x"0a",
          6770 => x"20",
          6771 => x"20",
          6772 => x"44",
          6773 => x"28",
          6774 => x"69",
          6775 => x"20",
          6776 => x"32",
          6777 => x"0a",
          6778 => x"20",
          6779 => x"4d",
          6780 => x"20",
          6781 => x"28",
          6782 => x"65",
          6783 => x"20",
          6784 => x"32",
          6785 => x"0a",
          6786 => x"20",
          6787 => x"54",
          6788 => x"54",
          6789 => x"28",
          6790 => x"6e",
          6791 => x"73",
          6792 => x"32",
          6793 => x"0a",
          6794 => x"20",
          6795 => x"53",
          6796 => x"4e",
          6797 => x"55",
          6798 => x"00",
          6799 => x"20",
          6800 => x"20",
          6801 => x"0a",
          6802 => x"20",
          6803 => x"43",
          6804 => x"00",
          6805 => x"20",
          6806 => x"32",
          6807 => x"00",
          6808 => x"20",
          6809 => x"49",
          6810 => x"00",
          6811 => x"64",
          6812 => x"73",
          6813 => x"0a",
          6814 => x"20",
          6815 => x"55",
          6816 => x"73",
          6817 => x"56",
          6818 => x"6f",
          6819 => x"64",
          6820 => x"73",
          6821 => x"20",
          6822 => x"58",
          6823 => x"00",
          6824 => x"20",
          6825 => x"55",
          6826 => x"6d",
          6827 => x"20",
          6828 => x"72",
          6829 => x"64",
          6830 => x"73",
          6831 => x"20",
          6832 => x"58",
          6833 => x"00",
          6834 => x"20",
          6835 => x"61",
          6836 => x"53",
          6837 => x"74",
          6838 => x"64",
          6839 => x"73",
          6840 => x"20",
          6841 => x"20",
          6842 => x"58",
          6843 => x"00",
          6844 => x"73",
          6845 => x"00",
          6846 => x"20",
          6847 => x"55",
          6848 => x"20",
          6849 => x"20",
          6850 => x"20",
          6851 => x"20",
          6852 => x"20",
          6853 => x"20",
          6854 => x"58",
          6855 => x"00",
          6856 => x"20",
          6857 => x"73",
          6858 => x"20",
          6859 => x"63",
          6860 => x"72",
          6861 => x"20",
          6862 => x"20",
          6863 => x"20",
          6864 => x"25",
          6865 => x"4d",
          6866 => x"00",
          6867 => x"20",
          6868 => x"52",
          6869 => x"43",
          6870 => x"6b",
          6871 => x"65",
          6872 => x"20",
          6873 => x"20",
          6874 => x"20",
          6875 => x"25",
          6876 => x"4d",
          6877 => x"00",
          6878 => x"20",
          6879 => x"73",
          6880 => x"6e",
          6881 => x"44",
          6882 => x"20",
          6883 => x"63",
          6884 => x"72",
          6885 => x"20",
          6886 => x"25",
          6887 => x"4d",
          6888 => x"00",
          6889 => x"61",
          6890 => x"00",
          6891 => x"64",
          6892 => x"00",
          6893 => x"65",
          6894 => x"00",
          6895 => x"4f",
          6896 => x"4f",
          6897 => x"00",
          6898 => x"6b",
          6899 => x"6e",
          6900 => x"73",
          6901 => x"79",
          6902 => x"74",
          6903 => x"73",
          6904 => x"79",
          6905 => x"73",
          6906 => x"00",
          6907 => x"00",
          6908 => x"34",
          6909 => x"25",
          6910 => x"00",
          6911 => x"69",
          6912 => x"20",
          6913 => x"72",
          6914 => x"74",
          6915 => x"65",
          6916 => x"73",
          6917 => x"79",
          6918 => x"6c",
          6919 => x"6f",
          6920 => x"46",
          6921 => x"00",
          6922 => x"6e",
          6923 => x"20",
          6924 => x"6e",
          6925 => x"65",
          6926 => x"20",
          6927 => x"74",
          6928 => x"20",
          6929 => x"65",
          6930 => x"69",
          6931 => x"6c",
          6932 => x"2e",
          6933 => x"00",
          6934 => x"7d",
          6935 => x"00",
          6936 => x"00",
          6937 => x"7d",
          6938 => x"00",
          6939 => x"00",
          6940 => x"7c",
          6941 => x"00",
          6942 => x"00",
          6943 => x"7c",
          6944 => x"00",
          6945 => x"00",
          6946 => x"7c",
          6947 => x"00",
          6948 => x"00",
          6949 => x"7c",
          6950 => x"00",
          6951 => x"00",
          6952 => x"7c",
          6953 => x"00",
          6954 => x"00",
          6955 => x"7c",
          6956 => x"00",
          6957 => x"00",
          6958 => x"7c",
          6959 => x"00",
          6960 => x"00",
          6961 => x"7c",
          6962 => x"00",
          6963 => x"00",
          6964 => x"7c",
          6965 => x"00",
          6966 => x"00",
          6967 => x"44",
          6968 => x"43",
          6969 => x"42",
          6970 => x"41",
          6971 => x"36",
          6972 => x"35",
          6973 => x"34",
          6974 => x"33",
          6975 => x"31",
          6976 => x"00",
          6977 => x"00",
          6978 => x"00",
          6979 => x"2b",
          6980 => x"3c",
          6981 => x"5b",
          6982 => x"00",
          6983 => x"54",
          6984 => x"54",
          6985 => x"00",
          6986 => x"90",
          6987 => x"4f",
          6988 => x"30",
          6989 => x"20",
          6990 => x"45",
          6991 => x"20",
          6992 => x"33",
          6993 => x"20",
          6994 => x"20",
          6995 => x"45",
          6996 => x"20",
          6997 => x"20",
          6998 => x"20",
          6999 => x"7d",
          7000 => x"00",
          7001 => x"00",
          7002 => x"00",
          7003 => x"45",
          7004 => x"8f",
          7005 => x"45",
          7006 => x"8e",
          7007 => x"92",
          7008 => x"55",
          7009 => x"9a",
          7010 => x"9e",
          7011 => x"4f",
          7012 => x"a6",
          7013 => x"aa",
          7014 => x"ae",
          7015 => x"b2",
          7016 => x"b6",
          7017 => x"ba",
          7018 => x"be",
          7019 => x"c2",
          7020 => x"c6",
          7021 => x"ca",
          7022 => x"ce",
          7023 => x"d2",
          7024 => x"d6",
          7025 => x"da",
          7026 => x"de",
          7027 => x"e2",
          7028 => x"e6",
          7029 => x"ea",
          7030 => x"ee",
          7031 => x"f2",
          7032 => x"f6",
          7033 => x"fa",
          7034 => x"fe",
          7035 => x"2c",
          7036 => x"5d",
          7037 => x"2a",
          7038 => x"3f",
          7039 => x"00",
          7040 => x"00",
          7041 => x"00",
          7042 => x"02",
          7043 => x"00",
          7044 => x"00",
          7045 => x"00",
          7046 => x"00",
          7047 => x"00",
          7048 => x"6e",
          7049 => x"00",
          7050 => x"6f",
          7051 => x"00",
          7052 => x"6e",
          7053 => x"00",
          7054 => x"6f",
          7055 => x"00",
          7056 => x"78",
          7057 => x"00",
          7058 => x"6c",
          7059 => x"00",
          7060 => x"6f",
          7061 => x"00",
          7062 => x"69",
          7063 => x"00",
          7064 => x"75",
          7065 => x"00",
          7066 => x"62",
          7067 => x"68",
          7068 => x"77",
          7069 => x"64",
          7070 => x"65",
          7071 => x"64",
          7072 => x"65",
          7073 => x"6c",
          7074 => x"00",
          7075 => x"70",
          7076 => x"73",
          7077 => x"74",
          7078 => x"73",
          7079 => x"00",
          7080 => x"66",
          7081 => x"00",
          7082 => x"73",
          7083 => x"00",
          7084 => x"61",
          7085 => x"00",
          7086 => x"61",
          7087 => x"00",
          7088 => x"6c",
          7089 => x"00",
          7090 => x"73",
          7091 => x"72",
          7092 => x"0a",
          7093 => x"74",
          7094 => x"61",
          7095 => x"72",
          7096 => x"2e",
          7097 => x"00",
          7098 => x"73",
          7099 => x"6f",
          7100 => x"65",
          7101 => x"2e",
          7102 => x"00",
          7103 => x"20",
          7104 => x"65",
          7105 => x"75",
          7106 => x"0a",
          7107 => x"20",
          7108 => x"68",
          7109 => x"75",
          7110 => x"0a",
          7111 => x"76",
          7112 => x"64",
          7113 => x"6c",
          7114 => x"6d",
          7115 => x"00",
          7116 => x"63",
          7117 => x"20",
          7118 => x"69",
          7119 => x"0a",
          7120 => x"6c",
          7121 => x"6c",
          7122 => x"64",
          7123 => x"78",
          7124 => x"73",
          7125 => x"00",
          7126 => x"6c",
          7127 => x"61",
          7128 => x"65",
          7129 => x"76",
          7130 => x"64",
          7131 => x"00",
          7132 => x"20",
          7133 => x"77",
          7134 => x"65",
          7135 => x"6f",
          7136 => x"74",
          7137 => x"0a",
          7138 => x"69",
          7139 => x"6e",
          7140 => x"65",
          7141 => x"73",
          7142 => x"76",
          7143 => x"64",
          7144 => x"00",
          7145 => x"73",
          7146 => x"6f",
          7147 => x"6e",
          7148 => x"65",
          7149 => x"00",
          7150 => x"20",
          7151 => x"70",
          7152 => x"62",
          7153 => x"66",
          7154 => x"73",
          7155 => x"65",
          7156 => x"6f",
          7157 => x"20",
          7158 => x"64",
          7159 => x"2e",
          7160 => x"00",
          7161 => x"72",
          7162 => x"20",
          7163 => x"72",
          7164 => x"2e",
          7165 => x"00",
          7166 => x"6d",
          7167 => x"74",
          7168 => x"70",
          7169 => x"74",
          7170 => x"20",
          7171 => x"63",
          7172 => x"65",
          7173 => x"00",
          7174 => x"6c",
          7175 => x"73",
          7176 => x"63",
          7177 => x"2e",
          7178 => x"00",
          7179 => x"73",
          7180 => x"69",
          7181 => x"6e",
          7182 => x"65",
          7183 => x"79",
          7184 => x"00",
          7185 => x"6f",
          7186 => x"6e",
          7187 => x"70",
          7188 => x"66",
          7189 => x"73",
          7190 => x"00",
          7191 => x"72",
          7192 => x"74",
          7193 => x"20",
          7194 => x"6f",
          7195 => x"63",
          7196 => x"00",
          7197 => x"63",
          7198 => x"73",
          7199 => x"00",
          7200 => x"6b",
          7201 => x"6e",
          7202 => x"72",
          7203 => x"0a",
          7204 => x"6c",
          7205 => x"79",
          7206 => x"20",
          7207 => x"61",
          7208 => x"6c",
          7209 => x"79",
          7210 => x"2f",
          7211 => x"2e",
          7212 => x"00",
          7213 => x"61",
          7214 => x"00",
          7215 => x"38",
          7216 => x"00",
          7217 => x"20",
          7218 => x"34",
          7219 => x"00",
          7220 => x"20",
          7221 => x"20",
          7222 => x"00",
          7223 => x"32",
          7224 => x"00",
          7225 => x"00",
          7226 => x"00",
          7227 => x"0a",
          7228 => x"53",
          7229 => x"2a",
          7230 => x"20",
          7231 => x"00",
          7232 => x"2f",
          7233 => x"32",
          7234 => x"00",
          7235 => x"2e",
          7236 => x"00",
          7237 => x"50",
          7238 => x"72",
          7239 => x"25",
          7240 => x"29",
          7241 => x"20",
          7242 => x"2a",
          7243 => x"00",
          7244 => x"55",
          7245 => x"74",
          7246 => x"75",
          7247 => x"48",
          7248 => x"6c",
          7249 => x"00",
          7250 => x"6d",
          7251 => x"69",
          7252 => x"72",
          7253 => x"74",
          7254 => x"00",
          7255 => x"32",
          7256 => x"74",
          7257 => x"75",
          7258 => x"00",
          7259 => x"43",
          7260 => x"52",
          7261 => x"6e",
          7262 => x"72",
          7263 => x"0a",
          7264 => x"43",
          7265 => x"57",
          7266 => x"6e",
          7267 => x"72",
          7268 => x"0a",
          7269 => x"52",
          7270 => x"52",
          7271 => x"6e",
          7272 => x"72",
          7273 => x"0a",
          7274 => x"52",
          7275 => x"54",
          7276 => x"6e",
          7277 => x"72",
          7278 => x"0a",
          7279 => x"52",
          7280 => x"52",
          7281 => x"6e",
          7282 => x"72",
          7283 => x"0a",
          7284 => x"52",
          7285 => x"54",
          7286 => x"6e",
          7287 => x"72",
          7288 => x"0a",
          7289 => x"74",
          7290 => x"67",
          7291 => x"20",
          7292 => x"65",
          7293 => x"2e",
          7294 => x"00",
          7295 => x"61",
          7296 => x"6e",
          7297 => x"69",
          7298 => x"2e",
          7299 => x"00",
          7300 => x"74",
          7301 => x"65",
          7302 => x"61",
          7303 => x"00",
          7304 => x"00",
          7305 => x"69",
          7306 => x"20",
          7307 => x"69",
          7308 => x"69",
          7309 => x"73",
          7310 => x"64",
          7311 => x"72",
          7312 => x"2c",
          7313 => x"65",
          7314 => x"20",
          7315 => x"74",
          7316 => x"6e",
          7317 => x"6c",
          7318 => x"00",
          7319 => x"00",
          7320 => x"65",
          7321 => x"6e",
          7322 => x"2e",
          7323 => x"00",
          7324 => x"70",
          7325 => x"67",
          7326 => x"00",
          7327 => x"6d",
          7328 => x"69",
          7329 => x"2e",
          7330 => x"00",
          7331 => x"38",
          7332 => x"25",
          7333 => x"29",
          7334 => x"30",
          7335 => x"28",
          7336 => x"78",
          7337 => x"00",
          7338 => x"6d",
          7339 => x"65",
          7340 => x"79",
          7341 => x"00",
          7342 => x"6f",
          7343 => x"65",
          7344 => x"0a",
          7345 => x"38",
          7346 => x"30",
          7347 => x"00",
          7348 => x"3f",
          7349 => x"00",
          7350 => x"38",
          7351 => x"30",
          7352 => x"00",
          7353 => x"38",
          7354 => x"30",
          7355 => x"00",
          7356 => x"65",
          7357 => x"69",
          7358 => x"63",
          7359 => x"20",
          7360 => x"30",
          7361 => x"2e",
          7362 => x"00",
          7363 => x"6c",
          7364 => x"67",
          7365 => x"64",
          7366 => x"20",
          7367 => x"78",
          7368 => x"2e",
          7369 => x"00",
          7370 => x"6c",
          7371 => x"65",
          7372 => x"6e",
          7373 => x"63",
          7374 => x"20",
          7375 => x"29",
          7376 => x"00",
          7377 => x"73",
          7378 => x"74",
          7379 => x"20",
          7380 => x"6c",
          7381 => x"74",
          7382 => x"2e",
          7383 => x"00",
          7384 => x"6c",
          7385 => x"65",
          7386 => x"74",
          7387 => x"2e",
          7388 => x"00",
          7389 => x"55",
          7390 => x"6e",
          7391 => x"3a",
          7392 => x"5c",
          7393 => x"25",
          7394 => x"00",
          7395 => x"3a",
          7396 => x"5c",
          7397 => x"00",
          7398 => x"3a",
          7399 => x"00",
          7400 => x"64",
          7401 => x"6d",
          7402 => x"64",
          7403 => x"00",
          7404 => x"6e",
          7405 => x"67",
          7406 => x"0a",
          7407 => x"61",
          7408 => x"6e",
          7409 => x"6e",
          7410 => x"72",
          7411 => x"73",
          7412 => x"0a",
          7413 => x"00",
          7414 => x"00",
          7415 => x"7f",
          7416 => x"00",
          7417 => x"7f",
          7418 => x"00",
          7419 => x"7f",
          7420 => x"00",
          7421 => x"00",
          7422 => x"00",
          7423 => x"ff",
          7424 => x"00",
          7425 => x"00",
          7426 => x"78",
          7427 => x"00",
          7428 => x"e1",
          7429 => x"e1",
          7430 => x"e1",
          7431 => x"00",
          7432 => x"01",
          7433 => x"01",
          7434 => x"10",
          7435 => x"00",
          7436 => x"00",
          7437 => x"00",
          7438 => x"00",
          7439 => x"84",
          7440 => x"84",
          7441 => x"84",
          7442 => x"84",
          7443 => x"7b",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"7b",
          7468 => x"00",
          7469 => x"7b",
          7470 => x"00",
          7471 => x"7b",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"7e",
          7476 => x"01",
          7477 => x"00",
          7478 => x"00",
          7479 => x"7e",
          7480 => x"01",
          7481 => x"00",
          7482 => x"00",
          7483 => x"7e",
          7484 => x"03",
          7485 => x"00",
          7486 => x"00",
          7487 => x"7e",
          7488 => x"03",
          7489 => x"00",
          7490 => x"00",
          7491 => x"7e",
          7492 => x"03",
          7493 => x"00",
          7494 => x"00",
          7495 => x"7e",
          7496 => x"04",
          7497 => x"00",
          7498 => x"00",
          7499 => x"7e",
          7500 => x"04",
          7501 => x"00",
          7502 => x"00",
          7503 => x"7e",
          7504 => x"04",
          7505 => x"00",
          7506 => x"00",
          7507 => x"7e",
          7508 => x"04",
          7509 => x"00",
          7510 => x"00",
          7511 => x"7e",
          7512 => x"04",
          7513 => x"00",
          7514 => x"00",
          7515 => x"7e",
          7516 => x"04",
          7517 => x"00",
          7518 => x"00",
          7519 => x"7e",
          7520 => x"04",
          7521 => x"00",
          7522 => x"00",
          7523 => x"7e",
          7524 => x"05",
          7525 => x"00",
          7526 => x"00",
          7527 => x"7e",
          7528 => x"05",
          7529 => x"00",
          7530 => x"00",
          7531 => x"7e",
          7532 => x"05",
          7533 => x"00",
          7534 => x"00",
          7535 => x"7e",
          7536 => x"05",
          7537 => x"00",
          7538 => x"00",
          7539 => x"7e",
          7540 => x"07",
          7541 => x"00",
          7542 => x"00",
          7543 => x"7e",
          7544 => x"07",
          7545 => x"00",
          7546 => x"00",
          7547 => x"7e",
          7548 => x"08",
          7549 => x"00",
          7550 => x"00",
          7551 => x"7e",
          7552 => x"08",
          7553 => x"00",
          7554 => x"00",
          7555 => x"7e",
          7556 => x"08",
          7557 => x"00",
          7558 => x"00",
          7559 => x"7e",
          7560 => x"08",
          7561 => x"00",
          7562 => x"00",
          7563 => x"7e",
          7564 => x"09",
          7565 => x"00",
          7566 => x"00",
          7567 => x"7e",
          7568 => x"09",
          7569 => x"00",
          7570 => x"00",
          7571 => x"7e",
          7572 => x"09",
          7573 => x"00",
          7574 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"aa",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"a4",
            11 => x"0b",
            12 => x"04",
            13 => x"a4",
            14 => x"0b",
            15 => x"04",
            16 => x"a4",
            17 => x"0b",
            18 => x"04",
            19 => x"a4",
            20 => x"0b",
            21 => x"04",
            22 => x"a5",
            23 => x"0b",
            24 => x"04",
            25 => x"a5",
            26 => x"0b",
            27 => x"04",
            28 => x"a5",
            29 => x"0b",
            30 => x"04",
            31 => x"a5",
            32 => x"0b",
            33 => x"04",
            34 => x"a6",
            35 => x"0b",
            36 => x"04",
            37 => x"a6",
            38 => x"0b",
            39 => x"04",
            40 => x"a6",
            41 => x"0b",
            42 => x"04",
            43 => x"a6",
            44 => x"0b",
            45 => x"04",
            46 => x"a6",
            47 => x"0b",
            48 => x"04",
            49 => x"a7",
            50 => x"0b",
            51 => x"04",
            52 => x"a7",
            53 => x"0b",
            54 => x"04",
            55 => x"a7",
            56 => x"0b",
            57 => x"04",
            58 => x"a7",
            59 => x"0b",
            60 => x"04",
            61 => x"a8",
            62 => x"0b",
            63 => x"04",
            64 => x"a8",
            65 => x"0b",
            66 => x"04",
            67 => x"a8",
            68 => x"0b",
            69 => x"04",
            70 => x"a8",
            71 => x"0b",
            72 => x"04",
            73 => x"a9",
            74 => x"0b",
            75 => x"04",
            76 => x"a9",
            77 => x"0b",
            78 => x"04",
            79 => x"a9",
            80 => x"0b",
            81 => x"04",
            82 => x"a9",
            83 => x"0b",
            84 => x"04",
            85 => x"aa",
            86 => x"0b",
            87 => x"04",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"a4",
           129 => x"8c",
           130 => x"a0",
           131 => x"e8",
           132 => x"90",
           133 => x"e8",
           134 => x"aa",
           135 => x"e8",
           136 => x"90",
           137 => x"e8",
           138 => x"e9",
           139 => x"e8",
           140 => x"90",
           141 => x"e8",
           142 => x"87",
           143 => x"e8",
           144 => x"90",
           145 => x"e8",
           146 => x"c5",
           147 => x"e8",
           148 => x"90",
           149 => x"e8",
           150 => x"c3",
           151 => x"e8",
           152 => x"90",
           153 => x"e8",
           154 => x"aa",
           155 => x"e8",
           156 => x"90",
           157 => x"e8",
           158 => x"e0",
           159 => x"e8",
           160 => x"90",
           161 => x"e8",
           162 => x"d2",
           163 => x"e8",
           164 => x"90",
           165 => x"e8",
           166 => x"eb",
           167 => x"e8",
           168 => x"90",
           169 => x"e8",
           170 => x"dc",
           171 => x"e8",
           172 => x"90",
           173 => x"e8",
           174 => x"81",
           175 => x"e8",
           176 => x"90",
           177 => x"e8",
           178 => x"a5",
           179 => x"e8",
           180 => x"90",
           181 => x"e8",
           182 => x"2d",
           183 => x"08",
           184 => x"04",
           185 => x"0c",
           186 => x"82",
           187 => x"83",
           188 => x"82",
           189 => x"b3",
           190 => x"8c",
           191 => x"80",
           192 => x"8c",
           193 => x"cf",
           194 => x"e8",
           195 => x"90",
           196 => x"e8",
           197 => x"2d",
           198 => x"08",
           199 => x"04",
           200 => x"0c",
           201 => x"2d",
           202 => x"08",
           203 => x"04",
           204 => x"0c",
           205 => x"2d",
           206 => x"08",
           207 => x"04",
           208 => x"0c",
           209 => x"2d",
           210 => x"08",
           211 => x"04",
           212 => x"0c",
           213 => x"2d",
           214 => x"08",
           215 => x"04",
           216 => x"0c",
           217 => x"2d",
           218 => x"08",
           219 => x"04",
           220 => x"0c",
           221 => x"2d",
           222 => x"08",
           223 => x"04",
           224 => x"0c",
           225 => x"2d",
           226 => x"08",
           227 => x"04",
           228 => x"0c",
           229 => x"2d",
           230 => x"08",
           231 => x"04",
           232 => x"0c",
           233 => x"2d",
           234 => x"08",
           235 => x"04",
           236 => x"0c",
           237 => x"2d",
           238 => x"08",
           239 => x"04",
           240 => x"0c",
           241 => x"2d",
           242 => x"08",
           243 => x"04",
           244 => x"0c",
           245 => x"2d",
           246 => x"08",
           247 => x"04",
           248 => x"0c",
           249 => x"2d",
           250 => x"08",
           251 => x"04",
           252 => x"0c",
           253 => x"2d",
           254 => x"08",
           255 => x"04",
           256 => x"0c",
           257 => x"2d",
           258 => x"08",
           259 => x"04",
           260 => x"0c",
           261 => x"2d",
           262 => x"08",
           263 => x"04",
           264 => x"0c",
           265 => x"2d",
           266 => x"08",
           267 => x"04",
           268 => x"0c",
           269 => x"2d",
           270 => x"08",
           271 => x"04",
           272 => x"0c",
           273 => x"2d",
           274 => x"08",
           275 => x"04",
           276 => x"0c",
           277 => x"2d",
           278 => x"08",
           279 => x"04",
           280 => x"0c",
           281 => x"2d",
           282 => x"08",
           283 => x"04",
           284 => x"0c",
           285 => x"2d",
           286 => x"08",
           287 => x"04",
           288 => x"0c",
           289 => x"2d",
           290 => x"08",
           291 => x"04",
           292 => x"0c",
           293 => x"2d",
           294 => x"08",
           295 => x"04",
           296 => x"0c",
           297 => x"2d",
           298 => x"08",
           299 => x"04",
           300 => x"0c",
           301 => x"2d",
           302 => x"08",
           303 => x"04",
           304 => x"0c",
           305 => x"2d",
           306 => x"08",
           307 => x"04",
           308 => x"0c",
           309 => x"2d",
           310 => x"08",
           311 => x"04",
           312 => x"0c",
           313 => x"2d",
           314 => x"08",
           315 => x"04",
           316 => x"0c",
           317 => x"2d",
           318 => x"08",
           319 => x"04",
           320 => x"0c",
           321 => x"82",
           322 => x"83",
           323 => x"82",
           324 => x"b4",
           325 => x"8c",
           326 => x"80",
           327 => x"8c",
           328 => x"92",
           329 => x"e8",
           330 => x"90",
           331 => x"e8",
           332 => x"ba",
           333 => x"e8",
           334 => x"90",
           335 => x"dc",
           336 => x"9c",
           337 => x"80",
           338 => x"05",
           339 => x"0b",
           340 => x"04",
           341 => x"81",
           342 => x"3c",
           343 => x"e8",
           344 => x"8c",
           345 => x"3d",
           346 => x"82",
           347 => x"8c",
           348 => x"82",
           349 => x"88",
           350 => x"80",
           351 => x"8c",
           352 => x"82",
           353 => x"54",
           354 => x"82",
           355 => x"04",
           356 => x"08",
           357 => x"e8",
           358 => x"0d",
           359 => x"8c",
           360 => x"05",
           361 => x"8c",
           362 => x"05",
           363 => x"3f",
           364 => x"08",
           365 => x"dc",
           366 => x"3d",
           367 => x"e8",
           368 => x"8c",
           369 => x"82",
           370 => x"fd",
           371 => x"0b",
           372 => x"08",
           373 => x"80",
           374 => x"e8",
           375 => x"0c",
           376 => x"08",
           377 => x"82",
           378 => x"88",
           379 => x"b9",
           380 => x"e8",
           381 => x"08",
           382 => x"38",
           383 => x"8c",
           384 => x"05",
           385 => x"38",
           386 => x"08",
           387 => x"10",
           388 => x"08",
           389 => x"82",
           390 => x"fc",
           391 => x"82",
           392 => x"fc",
           393 => x"b8",
           394 => x"e8",
           395 => x"08",
           396 => x"e1",
           397 => x"e8",
           398 => x"08",
           399 => x"08",
           400 => x"26",
           401 => x"8c",
           402 => x"05",
           403 => x"e8",
           404 => x"08",
           405 => x"e8",
           406 => x"0c",
           407 => x"08",
           408 => x"82",
           409 => x"fc",
           410 => x"82",
           411 => x"f8",
           412 => x"8c",
           413 => x"05",
           414 => x"82",
           415 => x"fc",
           416 => x"8c",
           417 => x"05",
           418 => x"82",
           419 => x"8c",
           420 => x"95",
           421 => x"e8",
           422 => x"08",
           423 => x"38",
           424 => x"08",
           425 => x"70",
           426 => x"08",
           427 => x"51",
           428 => x"8c",
           429 => x"05",
           430 => x"8c",
           431 => x"05",
           432 => x"8c",
           433 => x"05",
           434 => x"dc",
           435 => x"0d",
           436 => x"0c",
           437 => x"0d",
           438 => x"7b",
           439 => x"55",
           440 => x"8c",
           441 => x"07",
           442 => x"70",
           443 => x"38",
           444 => x"71",
           445 => x"38",
           446 => x"05",
           447 => x"70",
           448 => x"34",
           449 => x"71",
           450 => x"81",
           451 => x"74",
           452 => x"0c",
           453 => x"04",
           454 => x"70",
           455 => x"08",
           456 => x"05",
           457 => x"70",
           458 => x"08",
           459 => x"05",
           460 => x"70",
           461 => x"08",
           462 => x"05",
           463 => x"70",
           464 => x"08",
           465 => x"05",
           466 => x"12",
           467 => x"26",
           468 => x"72",
           469 => x"72",
           470 => x"54",
           471 => x"84",
           472 => x"fc",
           473 => x"83",
           474 => x"70",
           475 => x"39",
           476 => x"76",
           477 => x"8c",
           478 => x"33",
           479 => x"55",
           480 => x"8a",
           481 => x"06",
           482 => x"2e",
           483 => x"12",
           484 => x"2e",
           485 => x"73",
           486 => x"55",
           487 => x"52",
           488 => x"09",
           489 => x"38",
           490 => x"dc",
           491 => x"0d",
           492 => x"88",
           493 => x"70",
           494 => x"07",
           495 => x"8f",
           496 => x"38",
           497 => x"84",
           498 => x"72",
           499 => x"05",
           500 => x"71",
           501 => x"53",
           502 => x"70",
           503 => x"0c",
           504 => x"71",
           505 => x"38",
           506 => x"90",
           507 => x"70",
           508 => x"0c",
           509 => x"71",
           510 => x"38",
           511 => x"8e",
           512 => x"0d",
           513 => x"70",
           514 => x"06",
           515 => x"55",
           516 => x"38",
           517 => x"70",
           518 => x"fb",
           519 => x"06",
           520 => x"82",
           521 => x"51",
           522 => x"54",
           523 => x"84",
           524 => x"70",
           525 => x"0c",
           526 => x"09",
           527 => x"fd",
           528 => x"70",
           529 => x"81",
           530 => x"51",
           531 => x"70",
           532 => x"38",
           533 => x"70",
           534 => x"33",
           535 => x"70",
           536 => x"34",
           537 => x"74",
           538 => x"0c",
           539 => x"04",
           540 => x"75",
           541 => x"06",
           542 => x"70",
           543 => x"70",
           544 => x"f7",
           545 => x"12",
           546 => x"84",
           547 => x"06",
           548 => x"53",
           549 => x"84",
           550 => x"70",
           551 => x"fd",
           552 => x"70",
           553 => x"81",
           554 => x"51",
           555 => x"80",
           556 => x"72",
           557 => x"51",
           558 => x"8a",
           559 => x"70",
           560 => x"70",
           561 => x"74",
           562 => x"dc",
           563 => x"0d",
           564 => x"0d",
           565 => x"70",
           566 => x"52",
           567 => x"80",
           568 => x"74",
           569 => x"51",
           570 => x"80",
           571 => x"13",
           572 => x"2e",
           573 => x"33",
           574 => x"51",
           575 => x"09",
           576 => x"38",
           577 => x"81",
           578 => x"81",
           579 => x"70",
           580 => x"fe",
           581 => x"81",
           582 => x"55",
           583 => x"ff",
           584 => x"06",
           585 => x"33",
           586 => x"51",
           587 => x"06",
           588 => x"06",
           589 => x"51",
           590 => x"82",
           591 => x"88",
           592 => x"71",
           593 => x"83",
           594 => x"38",
           595 => x"08",
           596 => x"74",
           597 => x"ff",
           598 => x"13",
           599 => x"2e",
           600 => x"08",
           601 => x"fb",
           602 => x"06",
           603 => x"82",
           604 => x"51",
           605 => x"9a",
           606 => x"84",
           607 => x"83",
           608 => x"38",
           609 => x"08",
           610 => x"74",
           611 => x"fe",
           612 => x"0b",
           613 => x"0c",
           614 => x"04",
           615 => x"80",
           616 => x"71",
           617 => x"87",
           618 => x"8c",
           619 => x"ff",
           620 => x"ff",
           621 => x"72",
           622 => x"38",
           623 => x"dc",
           624 => x"0d",
           625 => x"0d",
           626 => x"70",
           627 => x"71",
           628 => x"ca",
           629 => x"51",
           630 => x"09",
           631 => x"38",
           632 => x"f1",
           633 => x"84",
           634 => x"53",
           635 => x"70",
           636 => x"53",
           637 => x"a0",
           638 => x"81",
           639 => x"2e",
           640 => x"e5",
           641 => x"ff",
           642 => x"a0",
           643 => x"06",
           644 => x"73",
           645 => x"55",
           646 => x"0c",
           647 => x"82",
           648 => x"87",
           649 => x"fc",
           650 => x"53",
           651 => x"2e",
           652 => x"3d",
           653 => x"72",
           654 => x"3f",
           655 => x"08",
           656 => x"53",
           657 => x"53",
           658 => x"dc",
           659 => x"0d",
           660 => x"0d",
           661 => x"33",
           662 => x"53",
           663 => x"8b",
           664 => x"38",
           665 => x"ff",
           666 => x"52",
           667 => x"81",
           668 => x"13",
           669 => x"52",
           670 => x"80",
           671 => x"13",
           672 => x"52",
           673 => x"80",
           674 => x"13",
           675 => x"52",
           676 => x"80",
           677 => x"13",
           678 => x"52",
           679 => x"26",
           680 => x"8a",
           681 => x"87",
           682 => x"e7",
           683 => x"38",
           684 => x"c0",
           685 => x"72",
           686 => x"98",
           687 => x"13",
           688 => x"98",
           689 => x"13",
           690 => x"98",
           691 => x"13",
           692 => x"98",
           693 => x"13",
           694 => x"98",
           695 => x"13",
           696 => x"98",
           697 => x"87",
           698 => x"0c",
           699 => x"98",
           700 => x"0b",
           701 => x"9c",
           702 => x"71",
           703 => x"0c",
           704 => x"04",
           705 => x"7f",
           706 => x"98",
           707 => x"7d",
           708 => x"98",
           709 => x"7d",
           710 => x"c0",
           711 => x"5a",
           712 => x"34",
           713 => x"b4",
           714 => x"83",
           715 => x"c0",
           716 => x"5a",
           717 => x"34",
           718 => x"ac",
           719 => x"85",
           720 => x"c0",
           721 => x"5a",
           722 => x"34",
           723 => x"a4",
           724 => x"88",
           725 => x"c0",
           726 => x"5a",
           727 => x"23",
           728 => x"79",
           729 => x"06",
           730 => x"ff",
           731 => x"86",
           732 => x"85",
           733 => x"84",
           734 => x"83",
           735 => x"82",
           736 => x"7d",
           737 => x"06",
           738 => x"e4",
           739 => x"3f",
           740 => x"04",
           741 => x"02",
           742 => x"70",
           743 => x"2a",
           744 => x"70",
           745 => x"87",
           746 => x"3d",
           747 => x"3d",
           748 => x"0b",
           749 => x"33",
           750 => x"06",
           751 => x"87",
           752 => x"51",
           753 => x"86",
           754 => x"94",
           755 => x"08",
           756 => x"70",
           757 => x"54",
           758 => x"2e",
           759 => x"91",
           760 => x"06",
           761 => x"d7",
           762 => x"32",
           763 => x"51",
           764 => x"2e",
           765 => x"93",
           766 => x"06",
           767 => x"ff",
           768 => x"81",
           769 => x"87",
           770 => x"52",
           771 => x"86",
           772 => x"94",
           773 => x"72",
           774 => x"8c",
           775 => x"3d",
           776 => x"3d",
           777 => x"05",
           778 => x"82",
           779 => x"70",
           780 => x"57",
           781 => x"c0",
           782 => x"74",
           783 => x"38",
           784 => x"94",
           785 => x"70",
           786 => x"81",
           787 => x"52",
           788 => x"8c",
           789 => x"2a",
           790 => x"51",
           791 => x"38",
           792 => x"70",
           793 => x"51",
           794 => x"8d",
           795 => x"2a",
           796 => x"51",
           797 => x"be",
           798 => x"ff",
           799 => x"c0",
           800 => x"70",
           801 => x"38",
           802 => x"90",
           803 => x"0c",
           804 => x"04",
           805 => x"79",
           806 => x"33",
           807 => x"06",
           808 => x"70",
           809 => x"fe",
           810 => x"ff",
           811 => x"0b",
           812 => x"d4",
           813 => x"ff",
           814 => x"55",
           815 => x"94",
           816 => x"80",
           817 => x"87",
           818 => x"51",
           819 => x"96",
           820 => x"06",
           821 => x"70",
           822 => x"38",
           823 => x"70",
           824 => x"51",
           825 => x"72",
           826 => x"81",
           827 => x"70",
           828 => x"38",
           829 => x"70",
           830 => x"51",
           831 => x"38",
           832 => x"06",
           833 => x"94",
           834 => x"80",
           835 => x"87",
           836 => x"52",
           837 => x"81",
           838 => x"70",
           839 => x"53",
           840 => x"ff",
           841 => x"82",
           842 => x"89",
           843 => x"fe",
           844 => x"0b",
           845 => x"33",
           846 => x"06",
           847 => x"c0",
           848 => x"72",
           849 => x"38",
           850 => x"94",
           851 => x"70",
           852 => x"81",
           853 => x"51",
           854 => x"e2",
           855 => x"ff",
           856 => x"c0",
           857 => x"70",
           858 => x"38",
           859 => x"90",
           860 => x"70",
           861 => x"82",
           862 => x"51",
           863 => x"04",
           864 => x"0b",
           865 => x"d4",
           866 => x"ff",
           867 => x"87",
           868 => x"52",
           869 => x"86",
           870 => x"94",
           871 => x"08",
           872 => x"70",
           873 => x"51",
           874 => x"70",
           875 => x"38",
           876 => x"06",
           877 => x"94",
           878 => x"80",
           879 => x"87",
           880 => x"52",
           881 => x"98",
           882 => x"2c",
           883 => x"71",
           884 => x"0c",
           885 => x"04",
           886 => x"87",
           887 => x"08",
           888 => x"8a",
           889 => x"70",
           890 => x"b4",
           891 => x"9e",
           892 => x"87",
           893 => x"c0",
           894 => x"82",
           895 => x"87",
           896 => x"08",
           897 => x"0c",
           898 => x"98",
           899 => x"e4",
           900 => x"9e",
           901 => x"87",
           902 => x"c0",
           903 => x"82",
           904 => x"87",
           905 => x"08",
           906 => x"0c",
           907 => x"b0",
           908 => x"f4",
           909 => x"9e",
           910 => x"87",
           911 => x"c0",
           912 => x"82",
           913 => x"87",
           914 => x"08",
           915 => x"0c",
           916 => x"c0",
           917 => x"84",
           918 => x"9e",
           919 => x"88",
           920 => x"c0",
           921 => x"51",
           922 => x"8c",
           923 => x"9e",
           924 => x"88",
           925 => x"c0",
           926 => x"82",
           927 => x"87",
           928 => x"08",
           929 => x"0c",
           930 => x"88",
           931 => x"0b",
           932 => x"90",
           933 => x"80",
           934 => x"52",
           935 => x"2e",
           936 => x"52",
           937 => x"9d",
           938 => x"87",
           939 => x"08",
           940 => x"0a",
           941 => x"52",
           942 => x"83",
           943 => x"71",
           944 => x"34",
           945 => x"c0",
           946 => x"70",
           947 => x"06",
           948 => x"70",
           949 => x"38",
           950 => x"82",
           951 => x"80",
           952 => x"9e",
           953 => x"88",
           954 => x"51",
           955 => x"80",
           956 => x"81",
           957 => x"88",
           958 => x"0b",
           959 => x"90",
           960 => x"80",
           961 => x"52",
           962 => x"2e",
           963 => x"52",
           964 => x"a1",
           965 => x"87",
           966 => x"08",
           967 => x"80",
           968 => x"52",
           969 => x"83",
           970 => x"71",
           971 => x"34",
           972 => x"c0",
           973 => x"70",
           974 => x"06",
           975 => x"70",
           976 => x"38",
           977 => x"82",
           978 => x"80",
           979 => x"9e",
           980 => x"82",
           981 => x"51",
           982 => x"80",
           983 => x"81",
           984 => x"88",
           985 => x"0b",
           986 => x"90",
           987 => x"80",
           988 => x"52",
           989 => x"2e",
           990 => x"52",
           991 => x"a5",
           992 => x"87",
           993 => x"08",
           994 => x"80",
           995 => x"52",
           996 => x"83",
           997 => x"71",
           998 => x"34",
           999 => x"c0",
          1000 => x"70",
          1001 => x"51",
          1002 => x"80",
          1003 => x"81",
          1004 => x"88",
          1005 => x"c0",
          1006 => x"70",
          1007 => x"70",
          1008 => x"51",
          1009 => x"88",
          1010 => x"0b",
          1011 => x"90",
          1012 => x"80",
          1013 => x"52",
          1014 => x"83",
          1015 => x"71",
          1016 => x"34",
          1017 => x"90",
          1018 => x"f0",
          1019 => x"2a",
          1020 => x"70",
          1021 => x"34",
          1022 => x"c0",
          1023 => x"70",
          1024 => x"52",
          1025 => x"2e",
          1026 => x"52",
          1027 => x"ab",
          1028 => x"9e",
          1029 => x"87",
          1030 => x"70",
          1031 => x"34",
          1032 => x"04",
          1033 => x"81",
          1034 => x"89",
          1035 => x"88",
          1036 => x"73",
          1037 => x"38",
          1038 => x"51",
          1039 => x"81",
          1040 => x"89",
          1041 => x"88",
          1042 => x"73",
          1043 => x"38",
          1044 => x"08",
          1045 => x"08",
          1046 => x"81",
          1047 => x"8f",
          1048 => x"88",
          1049 => x"73",
          1050 => x"38",
          1051 => x"08",
          1052 => x"08",
          1053 => x"81",
          1054 => x"8e",
          1055 => x"88",
          1056 => x"73",
          1057 => x"38",
          1058 => x"08",
          1059 => x"08",
          1060 => x"81",
          1061 => x"8e",
          1062 => x"88",
          1063 => x"73",
          1064 => x"38",
          1065 => x"08",
          1066 => x"08",
          1067 => x"81",
          1068 => x"8e",
          1069 => x"88",
          1070 => x"73",
          1071 => x"38",
          1072 => x"08",
          1073 => x"08",
          1074 => x"81",
          1075 => x"8e",
          1076 => x"88",
          1077 => x"73",
          1078 => x"38",
          1079 => x"33",
          1080 => x"c8",
          1081 => x"3f",
          1082 => x"33",
          1083 => x"2e",
          1084 => x"88",
          1085 => x"81",
          1086 => x"8d",
          1087 => x"88",
          1088 => x"73",
          1089 => x"38",
          1090 => x"33",
          1091 => x"88",
          1092 => x"3f",
          1093 => x"33",
          1094 => x"2e",
          1095 => x"f4",
          1096 => x"e5",
          1097 => x"9f",
          1098 => x"80",
          1099 => x"81",
          1100 => x"87",
          1101 => x"88",
          1102 => x"73",
          1103 => x"38",
          1104 => x"51",
          1105 => x"82",
          1106 => x"54",
          1107 => x"88",
          1108 => x"d4",
          1109 => x"3f",
          1110 => x"33",
          1111 => x"2e",
          1112 => x"f4",
          1113 => x"a1",
          1114 => x"ec",
          1115 => x"3f",
          1116 => x"08",
          1117 => x"f8",
          1118 => x"3f",
          1119 => x"08",
          1120 => x"a0",
          1121 => x"3f",
          1122 => x"08",
          1123 => x"c8",
          1124 => x"3f",
          1125 => x"51",
          1126 => x"82",
          1127 => x"52",
          1128 => x"51",
          1129 => x"82",
          1130 => x"56",
          1131 => x"52",
          1132 => x"a9",
          1133 => x"dc",
          1134 => x"c0",
          1135 => x"31",
          1136 => x"8c",
          1137 => x"81",
          1138 => x"8c",
          1139 => x"88",
          1140 => x"73",
          1141 => x"38",
          1142 => x"08",
          1143 => x"c0",
          1144 => x"e6",
          1145 => x"8c",
          1146 => x"84",
          1147 => x"71",
          1148 => x"82",
          1149 => x"52",
          1150 => x"51",
          1151 => x"82",
          1152 => x"54",
          1153 => x"a8",
          1154 => x"98",
          1155 => x"84",
          1156 => x"51",
          1157 => x"82",
          1158 => x"bd",
          1159 => x"76",
          1160 => x"54",
          1161 => x"08",
          1162 => x"f8",
          1163 => x"3f",
          1164 => x"51",
          1165 => x"87",
          1166 => x"fe",
          1167 => x"92",
          1168 => x"05",
          1169 => x"26",
          1170 => x"84",
          1171 => x"81",
          1172 => x"52",
          1173 => x"81",
          1174 => x"9d",
          1175 => x"ac",
          1176 => x"81",
          1177 => x"91",
          1178 => x"bc",
          1179 => x"81",
          1180 => x"85",
          1181 => x"c8",
          1182 => x"3f",
          1183 => x"04",
          1184 => x"0c",
          1185 => x"87",
          1186 => x"0c",
          1187 => x"b0",
          1188 => x"96",
          1189 => x"fe",
          1190 => x"8c",
          1191 => x"38",
          1192 => x"0b",
          1193 => x"0c",
          1194 => x"08",
          1195 => x"52",
          1196 => x"83",
          1197 => x"88",
          1198 => x"8c",
          1199 => x"53",
          1200 => x"dc",
          1201 => x"0d",
          1202 => x"0d",
          1203 => x"12",
          1204 => x"90",
          1205 => x"15",
          1206 => x"5e",
          1207 => x"59",
          1208 => x"77",
          1209 => x"75",
          1210 => x"08",
          1211 => x"71",
          1212 => x"31",
          1213 => x"80",
          1214 => x"84",
          1215 => x"8c",
          1216 => x"88",
          1217 => x"8c",
          1218 => x"88",
          1219 => x"90",
          1220 => x"94",
          1221 => x"94",
          1222 => x"90",
          1223 => x"39",
          1224 => x"73",
          1225 => x"74",
          1226 => x"77",
          1227 => x"0c",
          1228 => x"04",
          1229 => x"76",
          1230 => x"88",
          1231 => x"53",
          1232 => x"81",
          1233 => x"06",
          1234 => x"12",
          1235 => x"52",
          1236 => x"2e",
          1237 => x"94",
          1238 => x"08",
          1239 => x"0c",
          1240 => x"0c",
          1241 => x"0c",
          1242 => x"39",
          1243 => x"82",
          1244 => x"90",
          1245 => x"88",
          1246 => x"14",
          1247 => x"88",
          1248 => x"13",
          1249 => x"12",
          1250 => x"08",
          1251 => x"81",
          1252 => x"84",
          1253 => x"14",
          1254 => x"74",
          1255 => x"06",
          1256 => x"14",
          1257 => x"14",
          1258 => x"08",
          1259 => x"70",
          1260 => x"52",
          1261 => x"8c",
          1262 => x"15",
          1263 => x"13",
          1264 => x"12",
          1265 => x"8c",
          1266 => x"3d",
          1267 => x"3d",
          1268 => x"55",
          1269 => x"2e",
          1270 => x"9f",
          1271 => x"82",
          1272 => x"57",
          1273 => x"82",
          1274 => x"84",
          1275 => x"27",
          1276 => x"90",
          1277 => x"ed",
          1278 => x"ff",
          1279 => x"80",
          1280 => x"58",
          1281 => x"82",
          1282 => x"82",
          1283 => x"30",
          1284 => x"dc",
          1285 => x"25",
          1286 => x"08",
          1287 => x"70",
          1288 => x"25",
          1289 => x"58",
          1290 => x"56",
          1291 => x"74",
          1292 => x"06",
          1293 => x"88",
          1294 => x"75",
          1295 => x"39",
          1296 => x"8c",
          1297 => x"77",
          1298 => x"08",
          1299 => x"82",
          1300 => x"53",
          1301 => x"2e",
          1302 => x"73",
          1303 => x"8c",
          1304 => x"f0",
          1305 => x"08",
          1306 => x"72",
          1307 => x"75",
          1308 => x"88",
          1309 => x"8c",
          1310 => x"75",
          1311 => x"3f",
          1312 => x"8c",
          1313 => x"fc",
          1314 => x"8c",
          1315 => x"73",
          1316 => x"0c",
          1317 => x"04",
          1318 => x"73",
          1319 => x"2e",
          1320 => x"12",
          1321 => x"3f",
          1322 => x"04",
          1323 => x"02",
          1324 => x"53",
          1325 => x"09",
          1326 => x"38",
          1327 => x"3f",
          1328 => x"08",
          1329 => x"2e",
          1330 => x"72",
          1331 => x"f8",
          1332 => x"82",
          1333 => x"8f",
          1334 => x"f0",
          1335 => x"80",
          1336 => x"72",
          1337 => x"84",
          1338 => x"fe",
          1339 => x"97",
          1340 => x"8c",
          1341 => x"82",
          1342 => x"54",
          1343 => x"3f",
          1344 => x"f0",
          1345 => x"0d",
          1346 => x"0d",
          1347 => x"33",
          1348 => x"06",
          1349 => x"80",
          1350 => x"72",
          1351 => x"51",
          1352 => x"ff",
          1353 => x"39",
          1354 => x"04",
          1355 => x"77",
          1356 => x"08",
          1357 => x"f0",
          1358 => x"73",
          1359 => x"ff",
          1360 => x"71",
          1361 => x"38",
          1362 => x"06",
          1363 => x"54",
          1364 => x"e7",
          1365 => x"8c",
          1366 => x"3d",
          1367 => x"3d",
          1368 => x"59",
          1369 => x"81",
          1370 => x"56",
          1371 => x"84",
          1372 => x"a5",
          1373 => x"06",
          1374 => x"80",
          1375 => x"81",
          1376 => x"58",
          1377 => x"b0",
          1378 => x"06",
          1379 => x"5a",
          1380 => x"ad",
          1381 => x"06",
          1382 => x"5a",
          1383 => x"05",
          1384 => x"75",
          1385 => x"81",
          1386 => x"77",
          1387 => x"08",
          1388 => x"05",
          1389 => x"5d",
          1390 => x"39",
          1391 => x"72",
          1392 => x"38",
          1393 => x"7b",
          1394 => x"05",
          1395 => x"70",
          1396 => x"33",
          1397 => x"39",
          1398 => x"32",
          1399 => x"72",
          1400 => x"78",
          1401 => x"70",
          1402 => x"07",
          1403 => x"07",
          1404 => x"51",
          1405 => x"80",
          1406 => x"79",
          1407 => x"70",
          1408 => x"33",
          1409 => x"80",
          1410 => x"38",
          1411 => x"e0",
          1412 => x"38",
          1413 => x"81",
          1414 => x"53",
          1415 => x"2e",
          1416 => x"73",
          1417 => x"a2",
          1418 => x"c3",
          1419 => x"38",
          1420 => x"24",
          1421 => x"80",
          1422 => x"8c",
          1423 => x"39",
          1424 => x"2e",
          1425 => x"81",
          1426 => x"80",
          1427 => x"80",
          1428 => x"d5",
          1429 => x"73",
          1430 => x"8e",
          1431 => x"39",
          1432 => x"2e",
          1433 => x"80",
          1434 => x"84",
          1435 => x"56",
          1436 => x"74",
          1437 => x"72",
          1438 => x"38",
          1439 => x"15",
          1440 => x"54",
          1441 => x"38",
          1442 => x"56",
          1443 => x"81",
          1444 => x"72",
          1445 => x"38",
          1446 => x"90",
          1447 => x"06",
          1448 => x"2e",
          1449 => x"51",
          1450 => x"74",
          1451 => x"53",
          1452 => x"fd",
          1453 => x"51",
          1454 => x"ef",
          1455 => x"19",
          1456 => x"53",
          1457 => x"39",
          1458 => x"39",
          1459 => x"39",
          1460 => x"39",
          1461 => x"39",
          1462 => x"d0",
          1463 => x"39",
          1464 => x"70",
          1465 => x"53",
          1466 => x"88",
          1467 => x"19",
          1468 => x"39",
          1469 => x"54",
          1470 => x"74",
          1471 => x"70",
          1472 => x"07",
          1473 => x"55",
          1474 => x"80",
          1475 => x"72",
          1476 => x"38",
          1477 => x"90",
          1478 => x"80",
          1479 => x"5e",
          1480 => x"74",
          1481 => x"3f",
          1482 => x"08",
          1483 => x"7c",
          1484 => x"54",
          1485 => x"82",
          1486 => x"55",
          1487 => x"92",
          1488 => x"53",
          1489 => x"2e",
          1490 => x"14",
          1491 => x"ff",
          1492 => x"14",
          1493 => x"70",
          1494 => x"34",
          1495 => x"30",
          1496 => x"9f",
          1497 => x"57",
          1498 => x"85",
          1499 => x"b1",
          1500 => x"2a",
          1501 => x"51",
          1502 => x"2e",
          1503 => x"3d",
          1504 => x"05",
          1505 => x"34",
          1506 => x"76",
          1507 => x"54",
          1508 => x"72",
          1509 => x"54",
          1510 => x"70",
          1511 => x"56",
          1512 => x"81",
          1513 => x"7b",
          1514 => x"73",
          1515 => x"3f",
          1516 => x"53",
          1517 => x"74",
          1518 => x"53",
          1519 => x"eb",
          1520 => x"77",
          1521 => x"53",
          1522 => x"14",
          1523 => x"54",
          1524 => x"3f",
          1525 => x"74",
          1526 => x"53",
          1527 => x"fb",
          1528 => x"51",
          1529 => x"ef",
          1530 => x"0d",
          1531 => x"0d",
          1532 => x"70",
          1533 => x"08",
          1534 => x"51",
          1535 => x"85",
          1536 => x"fe",
          1537 => x"82",
          1538 => x"85",
          1539 => x"52",
          1540 => x"ca",
          1541 => x"f8",
          1542 => x"73",
          1543 => x"82",
          1544 => x"84",
          1545 => x"fd",
          1546 => x"8c",
          1547 => x"82",
          1548 => x"87",
          1549 => x"53",
          1550 => x"fa",
          1551 => x"82",
          1552 => x"85",
          1553 => x"fb",
          1554 => x"79",
          1555 => x"08",
          1556 => x"57",
          1557 => x"71",
          1558 => x"e0",
          1559 => x"f4",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"53",
          1563 => x"80",
          1564 => x"8d",
          1565 => x"72",
          1566 => x"30",
          1567 => x"51",
          1568 => x"80",
          1569 => x"71",
          1570 => x"38",
          1571 => x"97",
          1572 => x"25",
          1573 => x"16",
          1574 => x"25",
          1575 => x"14",
          1576 => x"34",
          1577 => x"72",
          1578 => x"3f",
          1579 => x"73",
          1580 => x"72",
          1581 => x"f7",
          1582 => x"53",
          1583 => x"dc",
          1584 => x"0d",
          1585 => x"0d",
          1586 => x"08",
          1587 => x"f4",
          1588 => x"76",
          1589 => x"ef",
          1590 => x"8c",
          1591 => x"3d",
          1592 => x"3d",
          1593 => x"5a",
          1594 => x"7a",
          1595 => x"08",
          1596 => x"53",
          1597 => x"09",
          1598 => x"38",
          1599 => x"0c",
          1600 => x"ad",
          1601 => x"06",
          1602 => x"76",
          1603 => x"0c",
          1604 => x"33",
          1605 => x"73",
          1606 => x"81",
          1607 => x"38",
          1608 => x"05",
          1609 => x"08",
          1610 => x"53",
          1611 => x"2e",
          1612 => x"57",
          1613 => x"2e",
          1614 => x"39",
          1615 => x"13",
          1616 => x"08",
          1617 => x"53",
          1618 => x"55",
          1619 => x"80",
          1620 => x"14",
          1621 => x"88",
          1622 => x"27",
          1623 => x"eb",
          1624 => x"53",
          1625 => x"89",
          1626 => x"38",
          1627 => x"55",
          1628 => x"8a",
          1629 => x"a0",
          1630 => x"c2",
          1631 => x"74",
          1632 => x"e0",
          1633 => x"ff",
          1634 => x"d0",
          1635 => x"ff",
          1636 => x"90",
          1637 => x"38",
          1638 => x"81",
          1639 => x"53",
          1640 => x"ca",
          1641 => x"27",
          1642 => x"77",
          1643 => x"08",
          1644 => x"0c",
          1645 => x"33",
          1646 => x"ff",
          1647 => x"80",
          1648 => x"74",
          1649 => x"79",
          1650 => x"74",
          1651 => x"0c",
          1652 => x"04",
          1653 => x"7a",
          1654 => x"80",
          1655 => x"58",
          1656 => x"33",
          1657 => x"a0",
          1658 => x"06",
          1659 => x"13",
          1660 => x"39",
          1661 => x"09",
          1662 => x"38",
          1663 => x"11",
          1664 => x"08",
          1665 => x"54",
          1666 => x"2e",
          1667 => x"80",
          1668 => x"08",
          1669 => x"0c",
          1670 => x"33",
          1671 => x"80",
          1672 => x"38",
          1673 => x"80",
          1674 => x"38",
          1675 => x"57",
          1676 => x"0c",
          1677 => x"33",
          1678 => x"39",
          1679 => x"74",
          1680 => x"38",
          1681 => x"80",
          1682 => x"89",
          1683 => x"38",
          1684 => x"d0",
          1685 => x"55",
          1686 => x"80",
          1687 => x"39",
          1688 => x"d9",
          1689 => x"80",
          1690 => x"27",
          1691 => x"80",
          1692 => x"89",
          1693 => x"70",
          1694 => x"55",
          1695 => x"70",
          1696 => x"55",
          1697 => x"27",
          1698 => x"14",
          1699 => x"06",
          1700 => x"74",
          1701 => x"73",
          1702 => x"38",
          1703 => x"14",
          1704 => x"05",
          1705 => x"08",
          1706 => x"54",
          1707 => x"39",
          1708 => x"84",
          1709 => x"55",
          1710 => x"81",
          1711 => x"8c",
          1712 => x"3d",
          1713 => x"3d",
          1714 => x"2b",
          1715 => x"79",
          1716 => x"98",
          1717 => x"13",
          1718 => x"51",
          1719 => x"51",
          1720 => x"81",
          1721 => x"33",
          1722 => x"74",
          1723 => x"81",
          1724 => x"08",
          1725 => x"05",
          1726 => x"71",
          1727 => x"52",
          1728 => x"09",
          1729 => x"38",
          1730 => x"82",
          1731 => x"85",
          1732 => x"fc",
          1733 => x"02",
          1734 => x"05",
          1735 => x"54",
          1736 => x"80",
          1737 => x"88",
          1738 => x"3f",
          1739 => x"fc",
          1740 => x"f2",
          1741 => x"33",
          1742 => x"71",
          1743 => x"81",
          1744 => x"de",
          1745 => x"f3",
          1746 => x"73",
          1747 => x"0d",
          1748 => x"0d",
          1749 => x"05",
          1750 => x"02",
          1751 => x"05",
          1752 => x"a8",
          1753 => x"29",
          1754 => x"05",
          1755 => x"59",
          1756 => x"59",
          1757 => x"86",
          1758 => x"f2",
          1759 => x"89",
          1760 => x"84",
          1761 => x"d0",
          1762 => x"70",
          1763 => x"5a",
          1764 => x"82",
          1765 => x"75",
          1766 => x"a8",
          1767 => x"29",
          1768 => x"05",
          1769 => x"56",
          1770 => x"2e",
          1771 => x"53",
          1772 => x"51",
          1773 => x"82",
          1774 => x"81",
          1775 => x"82",
          1776 => x"74",
          1777 => x"55",
          1778 => x"87",
          1779 => x"82",
          1780 => x"77",
          1781 => x"38",
          1782 => x"08",
          1783 => x"2e",
          1784 => x"89",
          1785 => x"74",
          1786 => x"3d",
          1787 => x"76",
          1788 => x"75",
          1789 => x"91",
          1790 => x"a4",
          1791 => x"51",
          1792 => x"3f",
          1793 => x"08",
          1794 => x"ee",
          1795 => x"0d",
          1796 => x"0d",
          1797 => x"52",
          1798 => x"08",
          1799 => x"87",
          1800 => x"dc",
          1801 => x"38",
          1802 => x"08",
          1803 => x"52",
          1804 => x"52",
          1805 => x"d5",
          1806 => x"dc",
          1807 => x"b8",
          1808 => x"d8",
          1809 => x"8c",
          1810 => x"80",
          1811 => x"dc",
          1812 => x"38",
          1813 => x"08",
          1814 => x"17",
          1815 => x"74",
          1816 => x"76",
          1817 => x"81",
          1818 => x"57",
          1819 => x"74",
          1820 => x"81",
          1821 => x"38",
          1822 => x"04",
          1823 => x"aa",
          1824 => x"3d",
          1825 => x"81",
          1826 => x"80",
          1827 => x"a4",
          1828 => x"d1",
          1829 => x"8c",
          1830 => x"91",
          1831 => x"82",
          1832 => x"54",
          1833 => x"52",
          1834 => x"52",
          1835 => x"dd",
          1836 => x"dc",
          1837 => x"a4",
          1838 => x"d7",
          1839 => x"8c",
          1840 => x"18",
          1841 => x"0b",
          1842 => x"08",
          1843 => x"82",
          1844 => x"ff",
          1845 => x"55",
          1846 => x"34",
          1847 => x"30",
          1848 => x"9f",
          1849 => x"55",
          1850 => x"85",
          1851 => x"ad",
          1852 => x"a4",
          1853 => x"08",
          1854 => x"d0",
          1855 => x"8c",
          1856 => x"2e",
          1857 => x"f7",
          1858 => x"fd",
          1859 => x"2e",
          1860 => x"99",
          1861 => x"79",
          1862 => x"3f",
          1863 => x"d0",
          1864 => x"08",
          1865 => x"dc",
          1866 => x"80",
          1867 => x"8c",
          1868 => x"3d",
          1869 => x"3d",
          1870 => x"71",
          1871 => x"33",
          1872 => x"58",
          1873 => x"09",
          1874 => x"38",
          1875 => x"05",
          1876 => x"27",
          1877 => x"17",
          1878 => x"71",
          1879 => x"55",
          1880 => x"09",
          1881 => x"38",
          1882 => x"ea",
          1883 => x"73",
          1884 => x"89",
          1885 => x"08",
          1886 => x"f4",
          1887 => x"dc",
          1888 => x"52",
          1889 => x"d6",
          1890 => x"8c",
          1891 => x"c4",
          1892 => x"33",
          1893 => x"2e",
          1894 => x"82",
          1895 => x"b4",
          1896 => x"3f",
          1897 => x"1a",
          1898 => x"fc",
          1899 => x"05",
          1900 => x"3f",
          1901 => x"08",
          1902 => x"38",
          1903 => x"52",
          1904 => x"b8",
          1905 => x"dc",
          1906 => x"06",
          1907 => x"38",
          1908 => x"39",
          1909 => x"81",
          1910 => x"54",
          1911 => x"ff",
          1912 => x"54",
          1913 => x"dc",
          1914 => x"0d",
          1915 => x"0d",
          1916 => x"02",
          1917 => x"c3",
          1918 => x"5a",
          1919 => x"3d",
          1920 => x"a8",
          1921 => x"89",
          1922 => x"a3",
          1923 => x"a0",
          1924 => x"81",
          1925 => x"51",
          1926 => x"82",
          1927 => x"82",
          1928 => x"82",
          1929 => x"80",
          1930 => x"38",
          1931 => x"88",
          1932 => x"82",
          1933 => x"51",
          1934 => x"82",
          1935 => x"80",
          1936 => x"81",
          1937 => x"f3",
          1938 => x"e3",
          1939 => x"a4",
          1940 => x"f8",
          1941 => x"70",
          1942 => x"f6",
          1943 => x"8c",
          1944 => x"82",
          1945 => x"74",
          1946 => x"06",
          1947 => x"82",
          1948 => x"51",
          1949 => x"82",
          1950 => x"55",
          1951 => x"8c",
          1952 => x"9a",
          1953 => x"dc",
          1954 => x"70",
          1955 => x"80",
          1956 => x"53",
          1957 => x"06",
          1958 => x"f9",
          1959 => x"ff",
          1960 => x"06",
          1961 => x"87",
          1962 => x"82",
          1963 => x"8f",
          1964 => x"cc",
          1965 => x"dc",
          1966 => x"70",
          1967 => x"59",
          1968 => x"ee",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"2b",
          1972 => x"82",
          1973 => x"70",
          1974 => x"97",
          1975 => x"2c",
          1976 => x"29",
          1977 => x"05",
          1978 => x"70",
          1979 => x"51",
          1980 => x"51",
          1981 => x"81",
          1982 => x"2e",
          1983 => x"77",
          1984 => x"38",
          1985 => x"0a",
          1986 => x"0a",
          1987 => x"2c",
          1988 => x"75",
          1989 => x"38",
          1990 => x"52",
          1991 => x"a6",
          1992 => x"dc",
          1993 => x"06",
          1994 => x"2e",
          1995 => x"82",
          1996 => x"81",
          1997 => x"74",
          1998 => x"29",
          1999 => x"05",
          2000 => x"70",
          2001 => x"56",
          2002 => x"8a",
          2003 => x"76",
          2004 => x"77",
          2005 => x"3f",
          2006 => x"08",
          2007 => x"54",
          2008 => x"d3",
          2009 => x"75",
          2010 => x"ca",
          2011 => x"55",
          2012 => x"80",
          2013 => x"2b",
          2014 => x"82",
          2015 => x"70",
          2016 => x"98",
          2017 => x"11",
          2018 => x"81",
          2019 => x"33",
          2020 => x"51",
          2021 => x"55",
          2022 => x"09",
          2023 => x"92",
          2024 => x"e0",
          2025 => x"0c",
          2026 => x"8d",
          2027 => x"0b",
          2028 => x"34",
          2029 => x"82",
          2030 => x"75",
          2031 => x"34",
          2032 => x"34",
          2033 => x"7e",
          2034 => x"26",
          2035 => x"73",
          2036 => x"f0",
          2037 => x"73",
          2038 => x"8d",
          2039 => x"73",
          2040 => x"cb",
          2041 => x"84",
          2042 => x"75",
          2043 => x"74",
          2044 => x"98",
          2045 => x"73",
          2046 => x"38",
          2047 => x"73",
          2048 => x"34",
          2049 => x"0a",
          2050 => x"0a",
          2051 => x"2c",
          2052 => x"33",
          2053 => x"df",
          2054 => x"88",
          2055 => x"56",
          2056 => x"8d",
          2057 => x"1a",
          2058 => x"33",
          2059 => x"8d",
          2060 => x"73",
          2061 => x"38",
          2062 => x"73",
          2063 => x"34",
          2064 => x"33",
          2065 => x"0a",
          2066 => x"0a",
          2067 => x"2c",
          2068 => x"33",
          2069 => x"56",
          2070 => x"a2",
          2071 => x"70",
          2072 => x"e8",
          2073 => x"81",
          2074 => x"81",
          2075 => x"70",
          2076 => x"8d",
          2077 => x"51",
          2078 => x"24",
          2079 => x"8d",
          2080 => x"98",
          2081 => x"2c",
          2082 => x"33",
          2083 => x"56",
          2084 => x"fc",
          2085 => x"51",
          2086 => x"74",
          2087 => x"29",
          2088 => x"05",
          2089 => x"82",
          2090 => x"56",
          2091 => x"75",
          2092 => x"fb",
          2093 => x"8d",
          2094 => x"81",
          2095 => x"55",
          2096 => x"fb",
          2097 => x"8d",
          2098 => x"05",
          2099 => x"8d",
          2100 => x"15",
          2101 => x"8d",
          2102 => x"51",
          2103 => x"82",
          2104 => x"70",
          2105 => x"98",
          2106 => x"84",
          2107 => x"56",
          2108 => x"25",
          2109 => x"1a",
          2110 => x"33",
          2111 => x"33",
          2112 => x"3f",
          2113 => x"0a",
          2114 => x"0a",
          2115 => x"2c",
          2116 => x"33",
          2117 => x"75",
          2118 => x"38",
          2119 => x"8c",
          2120 => x"88",
          2121 => x"2b",
          2122 => x"82",
          2123 => x"57",
          2124 => x"74",
          2125 => x"f7",
          2126 => x"e6",
          2127 => x"81",
          2128 => x"81",
          2129 => x"70",
          2130 => x"8d",
          2131 => x"51",
          2132 => x"25",
          2133 => x"d7",
          2134 => x"84",
          2135 => x"54",
          2136 => x"8a",
          2137 => x"3f",
          2138 => x"52",
          2139 => x"c6",
          2140 => x"dc",
          2141 => x"06",
          2142 => x"38",
          2143 => x"33",
          2144 => x"2e",
          2145 => x"81",
          2146 => x"79",
          2147 => x"3f",
          2148 => x"80",
          2149 => x"b7",
          2150 => x"88",
          2151 => x"80",
          2152 => x"38",
          2153 => x"84",
          2154 => x"88",
          2155 => x"54",
          2156 => x"88",
          2157 => x"ff",
          2158 => x"39",
          2159 => x"33",
          2160 => x"33",
          2161 => x"75",
          2162 => x"38",
          2163 => x"73",
          2164 => x"34",
          2165 => x"70",
          2166 => x"81",
          2167 => x"51",
          2168 => x"25",
          2169 => x"1a",
          2170 => x"33",
          2171 => x"33",
          2172 => x"3f",
          2173 => x"0a",
          2174 => x"0a",
          2175 => x"2c",
          2176 => x"33",
          2177 => x"75",
          2178 => x"38",
          2179 => x"9c",
          2180 => x"88",
          2181 => x"2b",
          2182 => x"82",
          2183 => x"57",
          2184 => x"74",
          2185 => x"87",
          2186 => x"e4",
          2187 => x"81",
          2188 => x"81",
          2189 => x"70",
          2190 => x"8d",
          2191 => x"51",
          2192 => x"25",
          2193 => x"e7",
          2194 => x"88",
          2195 => x"ff",
          2196 => x"84",
          2197 => x"54",
          2198 => x"f8",
          2199 => x"14",
          2200 => x"8d",
          2201 => x"1a",
          2202 => x"54",
          2203 => x"82",
          2204 => x"70",
          2205 => x"82",
          2206 => x"58",
          2207 => x"75",
          2208 => x"f8",
          2209 => x"ae",
          2210 => x"9c",
          2211 => x"80",
          2212 => x"74",
          2213 => x"3f",
          2214 => x"08",
          2215 => x"34",
          2216 => x"08",
          2217 => x"81",
          2218 => x"52",
          2219 => x"a5",
          2220 => x"81",
          2221 => x"84",
          2222 => x"d0",
          2223 => x"08",
          2224 => x"80",
          2225 => x"74",
          2226 => x"3f",
          2227 => x"08",
          2228 => x"34",
          2229 => x"08",
          2230 => x"81",
          2231 => x"52",
          2232 => x"f1",
          2233 => x"54",
          2234 => x"73",
          2235 => x"80",
          2236 => x"38",
          2237 => x"f8",
          2238 => x"39",
          2239 => x"09",
          2240 => x"38",
          2241 => x"08",
          2242 => x"2e",
          2243 => x"51",
          2244 => x"80",
          2245 => x"84",
          2246 => x"d0",
          2247 => x"08",
          2248 => x"80",
          2249 => x"74",
          2250 => x"3f",
          2251 => x"08",
          2252 => x"34",
          2253 => x"08",
          2254 => x"81",
          2255 => x"52",
          2256 => x"91",
          2257 => x"54",
          2258 => x"06",
          2259 => x"73",
          2260 => x"80",
          2261 => x"38",
          2262 => x"94",
          2263 => x"dc",
          2264 => x"84",
          2265 => x"dc",
          2266 => x"06",
          2267 => x"74",
          2268 => x"c6",
          2269 => x"8d",
          2270 => x"8d",
          2271 => x"79",
          2272 => x"3f",
          2273 => x"82",
          2274 => x"70",
          2275 => x"82",
          2276 => x"59",
          2277 => x"77",
          2278 => x"38",
          2279 => x"73",
          2280 => x"34",
          2281 => x"33",
          2282 => x"80",
          2283 => x"39",
          2284 => x"33",
          2285 => x"2e",
          2286 => x"88",
          2287 => x"3f",
          2288 => x"33",
          2289 => x"73",
          2290 => x"34",
          2291 => x"80",
          2292 => x"88",
          2293 => x"82",
          2294 => x"79",
          2295 => x"0c",
          2296 => x"04",
          2297 => x"02",
          2298 => x"51",
          2299 => x"72",
          2300 => x"82",
          2301 => x"33",
          2302 => x"8c",
          2303 => x"3d",
          2304 => x"3d",
          2305 => x"05",
          2306 => x"05",
          2307 => x"56",
          2308 => x"72",
          2309 => x"e0",
          2310 => x"2b",
          2311 => x"8c",
          2312 => x"88",
          2313 => x"2e",
          2314 => x"88",
          2315 => x"0c",
          2316 => x"8c",
          2317 => x"71",
          2318 => x"87",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"51",
          2322 => x"2e",
          2323 => x"c0",
          2324 => x"51",
          2325 => x"71",
          2326 => x"80",
          2327 => x"92",
          2328 => x"98",
          2329 => x"70",
          2330 => x"38",
          2331 => x"c4",
          2332 => x"89",
          2333 => x"51",
          2334 => x"dc",
          2335 => x"0d",
          2336 => x"0d",
          2337 => x"02",
          2338 => x"05",
          2339 => x"58",
          2340 => x"52",
          2341 => x"3f",
          2342 => x"08",
          2343 => x"54",
          2344 => x"be",
          2345 => x"75",
          2346 => x"c0",
          2347 => x"87",
          2348 => x"12",
          2349 => x"84",
          2350 => x"40",
          2351 => x"85",
          2352 => x"98",
          2353 => x"7d",
          2354 => x"0c",
          2355 => x"85",
          2356 => x"06",
          2357 => x"71",
          2358 => x"38",
          2359 => x"71",
          2360 => x"05",
          2361 => x"19",
          2362 => x"a2",
          2363 => x"71",
          2364 => x"38",
          2365 => x"83",
          2366 => x"38",
          2367 => x"8a",
          2368 => x"98",
          2369 => x"71",
          2370 => x"c0",
          2371 => x"52",
          2372 => x"87",
          2373 => x"80",
          2374 => x"81",
          2375 => x"c0",
          2376 => x"53",
          2377 => x"82",
          2378 => x"71",
          2379 => x"1a",
          2380 => x"84",
          2381 => x"19",
          2382 => x"06",
          2383 => x"79",
          2384 => x"38",
          2385 => x"80",
          2386 => x"87",
          2387 => x"26",
          2388 => x"73",
          2389 => x"06",
          2390 => x"2e",
          2391 => x"52",
          2392 => x"82",
          2393 => x"8f",
          2394 => x"f3",
          2395 => x"62",
          2396 => x"05",
          2397 => x"57",
          2398 => x"83",
          2399 => x"52",
          2400 => x"3f",
          2401 => x"08",
          2402 => x"54",
          2403 => x"2e",
          2404 => x"81",
          2405 => x"74",
          2406 => x"c0",
          2407 => x"87",
          2408 => x"12",
          2409 => x"84",
          2410 => x"5f",
          2411 => x"0b",
          2412 => x"8c",
          2413 => x"0c",
          2414 => x"80",
          2415 => x"70",
          2416 => x"81",
          2417 => x"54",
          2418 => x"8c",
          2419 => x"81",
          2420 => x"7c",
          2421 => x"58",
          2422 => x"70",
          2423 => x"52",
          2424 => x"8a",
          2425 => x"98",
          2426 => x"71",
          2427 => x"c0",
          2428 => x"52",
          2429 => x"87",
          2430 => x"80",
          2431 => x"81",
          2432 => x"c0",
          2433 => x"53",
          2434 => x"82",
          2435 => x"71",
          2436 => x"19",
          2437 => x"81",
          2438 => x"ff",
          2439 => x"19",
          2440 => x"78",
          2441 => x"38",
          2442 => x"80",
          2443 => x"87",
          2444 => x"26",
          2445 => x"73",
          2446 => x"06",
          2447 => x"2e",
          2448 => x"52",
          2449 => x"82",
          2450 => x"8f",
          2451 => x"fa",
          2452 => x"02",
          2453 => x"05",
          2454 => x"05",
          2455 => x"71",
          2456 => x"57",
          2457 => x"82",
          2458 => x"81",
          2459 => x"54",
          2460 => x"38",
          2461 => x"c0",
          2462 => x"81",
          2463 => x"2e",
          2464 => x"71",
          2465 => x"38",
          2466 => x"87",
          2467 => x"11",
          2468 => x"80",
          2469 => x"80",
          2470 => x"83",
          2471 => x"38",
          2472 => x"72",
          2473 => x"2a",
          2474 => x"51",
          2475 => x"80",
          2476 => x"87",
          2477 => x"08",
          2478 => x"38",
          2479 => x"8c",
          2480 => x"96",
          2481 => x"0c",
          2482 => x"8c",
          2483 => x"08",
          2484 => x"51",
          2485 => x"38",
          2486 => x"56",
          2487 => x"80",
          2488 => x"85",
          2489 => x"77",
          2490 => x"83",
          2491 => x"75",
          2492 => x"8c",
          2493 => x"3d",
          2494 => x"3d",
          2495 => x"11",
          2496 => x"71",
          2497 => x"82",
          2498 => x"53",
          2499 => x"0d",
          2500 => x"0d",
          2501 => x"33",
          2502 => x"71",
          2503 => x"88",
          2504 => x"14",
          2505 => x"07",
          2506 => x"33",
          2507 => x"8c",
          2508 => x"53",
          2509 => x"52",
          2510 => x"04",
          2511 => x"73",
          2512 => x"92",
          2513 => x"52",
          2514 => x"81",
          2515 => x"70",
          2516 => x"70",
          2517 => x"3d",
          2518 => x"3d",
          2519 => x"52",
          2520 => x"70",
          2521 => x"34",
          2522 => x"51",
          2523 => x"81",
          2524 => x"70",
          2525 => x"70",
          2526 => x"05",
          2527 => x"88",
          2528 => x"72",
          2529 => x"0d",
          2530 => x"0d",
          2531 => x"54",
          2532 => x"80",
          2533 => x"71",
          2534 => x"53",
          2535 => x"81",
          2536 => x"ff",
          2537 => x"39",
          2538 => x"04",
          2539 => x"75",
          2540 => x"52",
          2541 => x"70",
          2542 => x"34",
          2543 => x"70",
          2544 => x"3d",
          2545 => x"3d",
          2546 => x"79",
          2547 => x"74",
          2548 => x"56",
          2549 => x"81",
          2550 => x"71",
          2551 => x"16",
          2552 => x"52",
          2553 => x"86",
          2554 => x"2e",
          2555 => x"82",
          2556 => x"86",
          2557 => x"fe",
          2558 => x"76",
          2559 => x"39",
          2560 => x"8a",
          2561 => x"51",
          2562 => x"71",
          2563 => x"33",
          2564 => x"0c",
          2565 => x"04",
          2566 => x"8c",
          2567 => x"80",
          2568 => x"dc",
          2569 => x"3d",
          2570 => x"80",
          2571 => x"33",
          2572 => x"7a",
          2573 => x"38",
          2574 => x"16",
          2575 => x"16",
          2576 => x"17",
          2577 => x"fa",
          2578 => x"8c",
          2579 => x"2e",
          2580 => x"b7",
          2581 => x"dc",
          2582 => x"34",
          2583 => x"70",
          2584 => x"31",
          2585 => x"59",
          2586 => x"77",
          2587 => x"82",
          2588 => x"74",
          2589 => x"81",
          2590 => x"81",
          2591 => x"53",
          2592 => x"16",
          2593 => x"e3",
          2594 => x"81",
          2595 => x"8c",
          2596 => x"3d",
          2597 => x"3d",
          2598 => x"56",
          2599 => x"74",
          2600 => x"2e",
          2601 => x"51",
          2602 => x"82",
          2603 => x"57",
          2604 => x"08",
          2605 => x"54",
          2606 => x"16",
          2607 => x"33",
          2608 => x"3f",
          2609 => x"08",
          2610 => x"38",
          2611 => x"57",
          2612 => x"0c",
          2613 => x"dc",
          2614 => x"0d",
          2615 => x"0d",
          2616 => x"57",
          2617 => x"82",
          2618 => x"58",
          2619 => x"08",
          2620 => x"76",
          2621 => x"83",
          2622 => x"06",
          2623 => x"84",
          2624 => x"78",
          2625 => x"81",
          2626 => x"38",
          2627 => x"82",
          2628 => x"52",
          2629 => x"52",
          2630 => x"3f",
          2631 => x"52",
          2632 => x"51",
          2633 => x"84",
          2634 => x"d2",
          2635 => x"fc",
          2636 => x"8a",
          2637 => x"52",
          2638 => x"51",
          2639 => x"90",
          2640 => x"84",
          2641 => x"fc",
          2642 => x"17",
          2643 => x"a0",
          2644 => x"86",
          2645 => x"08",
          2646 => x"b0",
          2647 => x"55",
          2648 => x"81",
          2649 => x"f8",
          2650 => x"84",
          2651 => x"53",
          2652 => x"17",
          2653 => x"d7",
          2654 => x"dc",
          2655 => x"83",
          2656 => x"77",
          2657 => x"0c",
          2658 => x"04",
          2659 => x"77",
          2660 => x"12",
          2661 => x"55",
          2662 => x"56",
          2663 => x"8d",
          2664 => x"22",
          2665 => x"ac",
          2666 => x"57",
          2667 => x"8c",
          2668 => x"3d",
          2669 => x"3d",
          2670 => x"70",
          2671 => x"57",
          2672 => x"81",
          2673 => x"98",
          2674 => x"81",
          2675 => x"74",
          2676 => x"72",
          2677 => x"f5",
          2678 => x"24",
          2679 => x"81",
          2680 => x"81",
          2681 => x"83",
          2682 => x"38",
          2683 => x"76",
          2684 => x"70",
          2685 => x"16",
          2686 => x"74",
          2687 => x"96",
          2688 => x"dc",
          2689 => x"38",
          2690 => x"06",
          2691 => x"33",
          2692 => x"89",
          2693 => x"08",
          2694 => x"54",
          2695 => x"fc",
          2696 => x"8c",
          2697 => x"fe",
          2698 => x"ff",
          2699 => x"11",
          2700 => x"2b",
          2701 => x"81",
          2702 => x"2a",
          2703 => x"51",
          2704 => x"e2",
          2705 => x"ff",
          2706 => x"da",
          2707 => x"2a",
          2708 => x"05",
          2709 => x"fc",
          2710 => x"8c",
          2711 => x"c6",
          2712 => x"83",
          2713 => x"05",
          2714 => x"f9",
          2715 => x"8c",
          2716 => x"ff",
          2717 => x"ae",
          2718 => x"2a",
          2719 => x"05",
          2720 => x"fc",
          2721 => x"8c",
          2722 => x"38",
          2723 => x"83",
          2724 => x"05",
          2725 => x"f8",
          2726 => x"8c",
          2727 => x"0a",
          2728 => x"39",
          2729 => x"82",
          2730 => x"89",
          2731 => x"f8",
          2732 => x"7c",
          2733 => x"56",
          2734 => x"77",
          2735 => x"38",
          2736 => x"08",
          2737 => x"38",
          2738 => x"72",
          2739 => x"9d",
          2740 => x"24",
          2741 => x"81",
          2742 => x"82",
          2743 => x"83",
          2744 => x"38",
          2745 => x"76",
          2746 => x"70",
          2747 => x"18",
          2748 => x"76",
          2749 => x"9e",
          2750 => x"dc",
          2751 => x"8c",
          2752 => x"d9",
          2753 => x"ff",
          2754 => x"05",
          2755 => x"81",
          2756 => x"54",
          2757 => x"80",
          2758 => x"77",
          2759 => x"f0",
          2760 => x"8f",
          2761 => x"51",
          2762 => x"34",
          2763 => x"17",
          2764 => x"2a",
          2765 => x"05",
          2766 => x"fa",
          2767 => x"8c",
          2768 => x"82",
          2769 => x"81",
          2770 => x"83",
          2771 => x"b4",
          2772 => x"2a",
          2773 => x"8f",
          2774 => x"2a",
          2775 => x"f0",
          2776 => x"06",
          2777 => x"72",
          2778 => x"ec",
          2779 => x"2a",
          2780 => x"05",
          2781 => x"fa",
          2782 => x"8c",
          2783 => x"82",
          2784 => x"80",
          2785 => x"83",
          2786 => x"52",
          2787 => x"fe",
          2788 => x"b4",
          2789 => x"a4",
          2790 => x"76",
          2791 => x"17",
          2792 => x"75",
          2793 => x"3f",
          2794 => x"08",
          2795 => x"dc",
          2796 => x"77",
          2797 => x"77",
          2798 => x"fc",
          2799 => x"b4",
          2800 => x"51",
          2801 => x"c9",
          2802 => x"dc",
          2803 => x"06",
          2804 => x"72",
          2805 => x"3f",
          2806 => x"17",
          2807 => x"8c",
          2808 => x"3d",
          2809 => x"3d",
          2810 => x"7e",
          2811 => x"56",
          2812 => x"75",
          2813 => x"74",
          2814 => x"27",
          2815 => x"80",
          2816 => x"ff",
          2817 => x"75",
          2818 => x"3f",
          2819 => x"08",
          2820 => x"dc",
          2821 => x"38",
          2822 => x"54",
          2823 => x"81",
          2824 => x"39",
          2825 => x"08",
          2826 => x"39",
          2827 => x"51",
          2828 => x"82",
          2829 => x"58",
          2830 => x"08",
          2831 => x"c7",
          2832 => x"dc",
          2833 => x"d2",
          2834 => x"dc",
          2835 => x"cf",
          2836 => x"74",
          2837 => x"fc",
          2838 => x"8c",
          2839 => x"38",
          2840 => x"fe",
          2841 => x"08",
          2842 => x"74",
          2843 => x"38",
          2844 => x"17",
          2845 => x"33",
          2846 => x"73",
          2847 => x"77",
          2848 => x"26",
          2849 => x"80",
          2850 => x"8c",
          2851 => x"3d",
          2852 => x"3d",
          2853 => x"71",
          2854 => x"5b",
          2855 => x"8c",
          2856 => x"77",
          2857 => x"38",
          2858 => x"78",
          2859 => x"81",
          2860 => x"79",
          2861 => x"f9",
          2862 => x"55",
          2863 => x"dc",
          2864 => x"e0",
          2865 => x"dc",
          2866 => x"8c",
          2867 => x"2e",
          2868 => x"98",
          2869 => x"8c",
          2870 => x"82",
          2871 => x"58",
          2872 => x"70",
          2873 => x"80",
          2874 => x"38",
          2875 => x"09",
          2876 => x"e2",
          2877 => x"56",
          2878 => x"76",
          2879 => x"82",
          2880 => x"7a",
          2881 => x"3f",
          2882 => x"8c",
          2883 => x"2e",
          2884 => x"86",
          2885 => x"dc",
          2886 => x"8c",
          2887 => x"70",
          2888 => x"07",
          2889 => x"7c",
          2890 => x"dc",
          2891 => x"51",
          2892 => x"81",
          2893 => x"8c",
          2894 => x"2e",
          2895 => x"17",
          2896 => x"74",
          2897 => x"73",
          2898 => x"27",
          2899 => x"58",
          2900 => x"80",
          2901 => x"56",
          2902 => x"98",
          2903 => x"26",
          2904 => x"56",
          2905 => x"81",
          2906 => x"52",
          2907 => x"c6",
          2908 => x"dc",
          2909 => x"b8",
          2910 => x"82",
          2911 => x"81",
          2912 => x"06",
          2913 => x"8c",
          2914 => x"82",
          2915 => x"09",
          2916 => x"72",
          2917 => x"70",
          2918 => x"51",
          2919 => x"80",
          2920 => x"78",
          2921 => x"06",
          2922 => x"73",
          2923 => x"39",
          2924 => x"52",
          2925 => x"f7",
          2926 => x"dc",
          2927 => x"dc",
          2928 => x"82",
          2929 => x"07",
          2930 => x"55",
          2931 => x"2e",
          2932 => x"80",
          2933 => x"75",
          2934 => x"76",
          2935 => x"3f",
          2936 => x"08",
          2937 => x"38",
          2938 => x"0c",
          2939 => x"fe",
          2940 => x"08",
          2941 => x"74",
          2942 => x"ff",
          2943 => x"0c",
          2944 => x"81",
          2945 => x"84",
          2946 => x"39",
          2947 => x"81",
          2948 => x"8c",
          2949 => x"8c",
          2950 => x"dc",
          2951 => x"39",
          2952 => x"55",
          2953 => x"dc",
          2954 => x"0d",
          2955 => x"0d",
          2956 => x"55",
          2957 => x"82",
          2958 => x"58",
          2959 => x"8c",
          2960 => x"d8",
          2961 => x"74",
          2962 => x"3f",
          2963 => x"08",
          2964 => x"08",
          2965 => x"59",
          2966 => x"77",
          2967 => x"70",
          2968 => x"c8",
          2969 => x"84",
          2970 => x"56",
          2971 => x"58",
          2972 => x"97",
          2973 => x"75",
          2974 => x"52",
          2975 => x"51",
          2976 => x"82",
          2977 => x"80",
          2978 => x"8a",
          2979 => x"32",
          2980 => x"72",
          2981 => x"2a",
          2982 => x"56",
          2983 => x"dc",
          2984 => x"0d",
          2985 => x"0d",
          2986 => x"08",
          2987 => x"74",
          2988 => x"26",
          2989 => x"74",
          2990 => x"72",
          2991 => x"74",
          2992 => x"88",
          2993 => x"73",
          2994 => x"33",
          2995 => x"27",
          2996 => x"16",
          2997 => x"9b",
          2998 => x"2a",
          2999 => x"88",
          3000 => x"58",
          3001 => x"80",
          3002 => x"16",
          3003 => x"0c",
          3004 => x"8a",
          3005 => x"89",
          3006 => x"72",
          3007 => x"38",
          3008 => x"51",
          3009 => x"82",
          3010 => x"54",
          3011 => x"08",
          3012 => x"38",
          3013 => x"8c",
          3014 => x"8b",
          3015 => x"08",
          3016 => x"08",
          3017 => x"82",
          3018 => x"74",
          3019 => x"cb",
          3020 => x"75",
          3021 => x"3f",
          3022 => x"08",
          3023 => x"73",
          3024 => x"98",
          3025 => x"82",
          3026 => x"2e",
          3027 => x"39",
          3028 => x"39",
          3029 => x"13",
          3030 => x"74",
          3031 => x"16",
          3032 => x"18",
          3033 => x"77",
          3034 => x"0c",
          3035 => x"04",
          3036 => x"7a",
          3037 => x"12",
          3038 => x"59",
          3039 => x"80",
          3040 => x"86",
          3041 => x"98",
          3042 => x"14",
          3043 => x"55",
          3044 => x"81",
          3045 => x"83",
          3046 => x"77",
          3047 => x"81",
          3048 => x"0c",
          3049 => x"55",
          3050 => x"76",
          3051 => x"17",
          3052 => x"74",
          3053 => x"9b",
          3054 => x"39",
          3055 => x"ff",
          3056 => x"2a",
          3057 => x"81",
          3058 => x"52",
          3059 => x"e6",
          3060 => x"dc",
          3061 => x"55",
          3062 => x"8c",
          3063 => x"80",
          3064 => x"55",
          3065 => x"08",
          3066 => x"f4",
          3067 => x"08",
          3068 => x"08",
          3069 => x"38",
          3070 => x"77",
          3071 => x"84",
          3072 => x"39",
          3073 => x"52",
          3074 => x"86",
          3075 => x"dc",
          3076 => x"55",
          3077 => x"08",
          3078 => x"c4",
          3079 => x"82",
          3080 => x"81",
          3081 => x"81",
          3082 => x"dc",
          3083 => x"b0",
          3084 => x"dc",
          3085 => x"51",
          3086 => x"82",
          3087 => x"a0",
          3088 => x"15",
          3089 => x"75",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"76",
          3093 => x"77",
          3094 => x"9c",
          3095 => x"55",
          3096 => x"dc",
          3097 => x"0d",
          3098 => x"0d",
          3099 => x"08",
          3100 => x"80",
          3101 => x"fc",
          3102 => x"8c",
          3103 => x"82",
          3104 => x"80",
          3105 => x"8c",
          3106 => x"98",
          3107 => x"78",
          3108 => x"3f",
          3109 => x"08",
          3110 => x"dc",
          3111 => x"38",
          3112 => x"08",
          3113 => x"70",
          3114 => x"58",
          3115 => x"2e",
          3116 => x"83",
          3117 => x"82",
          3118 => x"55",
          3119 => x"81",
          3120 => x"07",
          3121 => x"2e",
          3122 => x"16",
          3123 => x"2e",
          3124 => x"88",
          3125 => x"82",
          3126 => x"56",
          3127 => x"51",
          3128 => x"82",
          3129 => x"54",
          3130 => x"08",
          3131 => x"9b",
          3132 => x"2e",
          3133 => x"83",
          3134 => x"73",
          3135 => x"0c",
          3136 => x"04",
          3137 => x"76",
          3138 => x"54",
          3139 => x"82",
          3140 => x"83",
          3141 => x"76",
          3142 => x"53",
          3143 => x"2e",
          3144 => x"90",
          3145 => x"51",
          3146 => x"82",
          3147 => x"90",
          3148 => x"53",
          3149 => x"dc",
          3150 => x"0d",
          3151 => x"0d",
          3152 => x"83",
          3153 => x"54",
          3154 => x"55",
          3155 => x"3f",
          3156 => x"51",
          3157 => x"2e",
          3158 => x"8b",
          3159 => x"2a",
          3160 => x"51",
          3161 => x"86",
          3162 => x"f7",
          3163 => x"7d",
          3164 => x"75",
          3165 => x"98",
          3166 => x"2e",
          3167 => x"98",
          3168 => x"78",
          3169 => x"3f",
          3170 => x"08",
          3171 => x"dc",
          3172 => x"38",
          3173 => x"70",
          3174 => x"73",
          3175 => x"58",
          3176 => x"8b",
          3177 => x"bf",
          3178 => x"ff",
          3179 => x"53",
          3180 => x"34",
          3181 => x"08",
          3182 => x"e5",
          3183 => x"81",
          3184 => x"2e",
          3185 => x"70",
          3186 => x"57",
          3187 => x"9e",
          3188 => x"2e",
          3189 => x"8c",
          3190 => x"df",
          3191 => x"72",
          3192 => x"81",
          3193 => x"76",
          3194 => x"2e",
          3195 => x"52",
          3196 => x"fc",
          3197 => x"dc",
          3198 => x"8c",
          3199 => x"38",
          3200 => x"fe",
          3201 => x"39",
          3202 => x"16",
          3203 => x"8c",
          3204 => x"3d",
          3205 => x"3d",
          3206 => x"08",
          3207 => x"52",
          3208 => x"c5",
          3209 => x"dc",
          3210 => x"8c",
          3211 => x"38",
          3212 => x"52",
          3213 => x"de",
          3214 => x"dc",
          3215 => x"8c",
          3216 => x"38",
          3217 => x"8c",
          3218 => x"9c",
          3219 => x"ea",
          3220 => x"53",
          3221 => x"9c",
          3222 => x"ea",
          3223 => x"0b",
          3224 => x"74",
          3225 => x"0c",
          3226 => x"04",
          3227 => x"75",
          3228 => x"12",
          3229 => x"53",
          3230 => x"9a",
          3231 => x"dc",
          3232 => x"9c",
          3233 => x"e5",
          3234 => x"0b",
          3235 => x"85",
          3236 => x"fa",
          3237 => x"7a",
          3238 => x"0b",
          3239 => x"98",
          3240 => x"2e",
          3241 => x"80",
          3242 => x"55",
          3243 => x"17",
          3244 => x"33",
          3245 => x"51",
          3246 => x"2e",
          3247 => x"85",
          3248 => x"06",
          3249 => x"e5",
          3250 => x"2e",
          3251 => x"8b",
          3252 => x"70",
          3253 => x"34",
          3254 => x"71",
          3255 => x"05",
          3256 => x"15",
          3257 => x"27",
          3258 => x"15",
          3259 => x"80",
          3260 => x"34",
          3261 => x"52",
          3262 => x"88",
          3263 => x"17",
          3264 => x"52",
          3265 => x"3f",
          3266 => x"08",
          3267 => x"12",
          3268 => x"3f",
          3269 => x"08",
          3270 => x"98",
          3271 => x"da",
          3272 => x"dc",
          3273 => x"23",
          3274 => x"04",
          3275 => x"7f",
          3276 => x"5b",
          3277 => x"33",
          3278 => x"73",
          3279 => x"38",
          3280 => x"80",
          3281 => x"38",
          3282 => x"8c",
          3283 => x"08",
          3284 => x"aa",
          3285 => x"41",
          3286 => x"33",
          3287 => x"73",
          3288 => x"81",
          3289 => x"81",
          3290 => x"dc",
          3291 => x"70",
          3292 => x"07",
          3293 => x"73",
          3294 => x"88",
          3295 => x"70",
          3296 => x"73",
          3297 => x"38",
          3298 => x"ab",
          3299 => x"52",
          3300 => x"91",
          3301 => x"dc",
          3302 => x"98",
          3303 => x"61",
          3304 => x"5a",
          3305 => x"a0",
          3306 => x"e7",
          3307 => x"70",
          3308 => x"79",
          3309 => x"73",
          3310 => x"81",
          3311 => x"38",
          3312 => x"33",
          3313 => x"ae",
          3314 => x"70",
          3315 => x"82",
          3316 => x"51",
          3317 => x"54",
          3318 => x"79",
          3319 => x"74",
          3320 => x"57",
          3321 => x"af",
          3322 => x"70",
          3323 => x"51",
          3324 => x"dc",
          3325 => x"73",
          3326 => x"38",
          3327 => x"82",
          3328 => x"19",
          3329 => x"54",
          3330 => x"82",
          3331 => x"54",
          3332 => x"78",
          3333 => x"81",
          3334 => x"54",
          3335 => x"81",
          3336 => x"af",
          3337 => x"77",
          3338 => x"70",
          3339 => x"25",
          3340 => x"07",
          3341 => x"51",
          3342 => x"2e",
          3343 => x"39",
          3344 => x"80",
          3345 => x"33",
          3346 => x"73",
          3347 => x"81",
          3348 => x"81",
          3349 => x"dc",
          3350 => x"70",
          3351 => x"07",
          3352 => x"73",
          3353 => x"b5",
          3354 => x"2e",
          3355 => x"83",
          3356 => x"76",
          3357 => x"07",
          3358 => x"2e",
          3359 => x"8b",
          3360 => x"77",
          3361 => x"30",
          3362 => x"71",
          3363 => x"53",
          3364 => x"55",
          3365 => x"38",
          3366 => x"5c",
          3367 => x"75",
          3368 => x"73",
          3369 => x"38",
          3370 => x"06",
          3371 => x"11",
          3372 => x"75",
          3373 => x"3f",
          3374 => x"08",
          3375 => x"38",
          3376 => x"33",
          3377 => x"54",
          3378 => x"e6",
          3379 => x"8c",
          3380 => x"2e",
          3381 => x"ff",
          3382 => x"74",
          3383 => x"38",
          3384 => x"75",
          3385 => x"17",
          3386 => x"57",
          3387 => x"a7",
          3388 => x"81",
          3389 => x"e5",
          3390 => x"8c",
          3391 => x"38",
          3392 => x"54",
          3393 => x"89",
          3394 => x"70",
          3395 => x"57",
          3396 => x"54",
          3397 => x"81",
          3398 => x"f7",
          3399 => x"7e",
          3400 => x"2e",
          3401 => x"33",
          3402 => x"e5",
          3403 => x"06",
          3404 => x"7a",
          3405 => x"a0",
          3406 => x"38",
          3407 => x"55",
          3408 => x"84",
          3409 => x"39",
          3410 => x"8b",
          3411 => x"7b",
          3412 => x"7a",
          3413 => x"3f",
          3414 => x"08",
          3415 => x"dc",
          3416 => x"38",
          3417 => x"52",
          3418 => x"aa",
          3419 => x"dc",
          3420 => x"8c",
          3421 => x"c2",
          3422 => x"08",
          3423 => x"55",
          3424 => x"ff",
          3425 => x"15",
          3426 => x"54",
          3427 => x"34",
          3428 => x"70",
          3429 => x"81",
          3430 => x"58",
          3431 => x"8b",
          3432 => x"74",
          3433 => x"3f",
          3434 => x"08",
          3435 => x"38",
          3436 => x"51",
          3437 => x"ff",
          3438 => x"ab",
          3439 => x"55",
          3440 => x"bb",
          3441 => x"2e",
          3442 => x"80",
          3443 => x"85",
          3444 => x"06",
          3445 => x"58",
          3446 => x"80",
          3447 => x"75",
          3448 => x"73",
          3449 => x"b5",
          3450 => x"0b",
          3451 => x"80",
          3452 => x"39",
          3453 => x"54",
          3454 => x"85",
          3455 => x"75",
          3456 => x"81",
          3457 => x"73",
          3458 => x"1b",
          3459 => x"2a",
          3460 => x"51",
          3461 => x"80",
          3462 => x"90",
          3463 => x"ff",
          3464 => x"05",
          3465 => x"f5",
          3466 => x"8c",
          3467 => x"1c",
          3468 => x"39",
          3469 => x"dc",
          3470 => x"0d",
          3471 => x"0d",
          3472 => x"7b",
          3473 => x"73",
          3474 => x"55",
          3475 => x"2e",
          3476 => x"75",
          3477 => x"57",
          3478 => x"26",
          3479 => x"ba",
          3480 => x"70",
          3481 => x"ba",
          3482 => x"06",
          3483 => x"73",
          3484 => x"70",
          3485 => x"51",
          3486 => x"89",
          3487 => x"82",
          3488 => x"ff",
          3489 => x"56",
          3490 => x"2e",
          3491 => x"80",
          3492 => x"dc",
          3493 => x"08",
          3494 => x"76",
          3495 => x"58",
          3496 => x"81",
          3497 => x"ff",
          3498 => x"53",
          3499 => x"26",
          3500 => x"13",
          3501 => x"06",
          3502 => x"9f",
          3503 => x"99",
          3504 => x"e0",
          3505 => x"ff",
          3506 => x"72",
          3507 => x"2a",
          3508 => x"72",
          3509 => x"06",
          3510 => x"ff",
          3511 => x"30",
          3512 => x"70",
          3513 => x"07",
          3514 => x"9f",
          3515 => x"54",
          3516 => x"80",
          3517 => x"81",
          3518 => x"59",
          3519 => x"25",
          3520 => x"8b",
          3521 => x"24",
          3522 => x"76",
          3523 => x"78",
          3524 => x"82",
          3525 => x"51",
          3526 => x"dc",
          3527 => x"0d",
          3528 => x"0d",
          3529 => x"0b",
          3530 => x"ff",
          3531 => x"0c",
          3532 => x"51",
          3533 => x"84",
          3534 => x"dc",
          3535 => x"38",
          3536 => x"51",
          3537 => x"82",
          3538 => x"83",
          3539 => x"54",
          3540 => x"82",
          3541 => x"09",
          3542 => x"e3",
          3543 => x"b4",
          3544 => x"57",
          3545 => x"2e",
          3546 => x"83",
          3547 => x"74",
          3548 => x"70",
          3549 => x"25",
          3550 => x"51",
          3551 => x"38",
          3552 => x"2e",
          3553 => x"b5",
          3554 => x"81",
          3555 => x"80",
          3556 => x"e0",
          3557 => x"8c",
          3558 => x"82",
          3559 => x"80",
          3560 => x"85",
          3561 => x"a0",
          3562 => x"16",
          3563 => x"3f",
          3564 => x"08",
          3565 => x"dc",
          3566 => x"83",
          3567 => x"74",
          3568 => x"0c",
          3569 => x"04",
          3570 => x"61",
          3571 => x"80",
          3572 => x"58",
          3573 => x"0c",
          3574 => x"e1",
          3575 => x"dc",
          3576 => x"56",
          3577 => x"8c",
          3578 => x"86",
          3579 => x"8c",
          3580 => x"29",
          3581 => x"05",
          3582 => x"53",
          3583 => x"80",
          3584 => x"38",
          3585 => x"76",
          3586 => x"74",
          3587 => x"72",
          3588 => x"38",
          3589 => x"51",
          3590 => x"82",
          3591 => x"81",
          3592 => x"81",
          3593 => x"72",
          3594 => x"80",
          3595 => x"38",
          3596 => x"70",
          3597 => x"53",
          3598 => x"86",
          3599 => x"a7",
          3600 => x"34",
          3601 => x"34",
          3602 => x"14",
          3603 => x"b2",
          3604 => x"dc",
          3605 => x"06",
          3606 => x"54",
          3607 => x"72",
          3608 => x"76",
          3609 => x"38",
          3610 => x"70",
          3611 => x"53",
          3612 => x"85",
          3613 => x"70",
          3614 => x"5b",
          3615 => x"82",
          3616 => x"81",
          3617 => x"76",
          3618 => x"81",
          3619 => x"38",
          3620 => x"56",
          3621 => x"83",
          3622 => x"70",
          3623 => x"80",
          3624 => x"83",
          3625 => x"dc",
          3626 => x"8c",
          3627 => x"76",
          3628 => x"05",
          3629 => x"16",
          3630 => x"56",
          3631 => x"d7",
          3632 => x"8d",
          3633 => x"72",
          3634 => x"54",
          3635 => x"57",
          3636 => x"95",
          3637 => x"73",
          3638 => x"3f",
          3639 => x"08",
          3640 => x"57",
          3641 => x"89",
          3642 => x"56",
          3643 => x"d7",
          3644 => x"76",
          3645 => x"f1",
          3646 => x"76",
          3647 => x"e9",
          3648 => x"51",
          3649 => x"82",
          3650 => x"83",
          3651 => x"53",
          3652 => x"2e",
          3653 => x"84",
          3654 => x"ca",
          3655 => x"da",
          3656 => x"dc",
          3657 => x"ff",
          3658 => x"8d",
          3659 => x"14",
          3660 => x"3f",
          3661 => x"08",
          3662 => x"15",
          3663 => x"14",
          3664 => x"34",
          3665 => x"33",
          3666 => x"81",
          3667 => x"54",
          3668 => x"72",
          3669 => x"91",
          3670 => x"ff",
          3671 => x"29",
          3672 => x"33",
          3673 => x"72",
          3674 => x"72",
          3675 => x"38",
          3676 => x"06",
          3677 => x"2e",
          3678 => x"56",
          3679 => x"80",
          3680 => x"da",
          3681 => x"8c",
          3682 => x"82",
          3683 => x"88",
          3684 => x"8f",
          3685 => x"56",
          3686 => x"38",
          3687 => x"51",
          3688 => x"82",
          3689 => x"83",
          3690 => x"55",
          3691 => x"80",
          3692 => x"da",
          3693 => x"8c",
          3694 => x"80",
          3695 => x"da",
          3696 => x"8c",
          3697 => x"ff",
          3698 => x"8d",
          3699 => x"2e",
          3700 => x"88",
          3701 => x"14",
          3702 => x"05",
          3703 => x"75",
          3704 => x"38",
          3705 => x"52",
          3706 => x"51",
          3707 => x"3f",
          3708 => x"08",
          3709 => x"dc",
          3710 => x"82",
          3711 => x"8c",
          3712 => x"ff",
          3713 => x"26",
          3714 => x"57",
          3715 => x"f5",
          3716 => x"82",
          3717 => x"f5",
          3718 => x"81",
          3719 => x"8d",
          3720 => x"2e",
          3721 => x"82",
          3722 => x"16",
          3723 => x"16",
          3724 => x"70",
          3725 => x"7a",
          3726 => x"0c",
          3727 => x"83",
          3728 => x"06",
          3729 => x"de",
          3730 => x"ae",
          3731 => x"dc",
          3732 => x"ff",
          3733 => x"56",
          3734 => x"38",
          3735 => x"38",
          3736 => x"51",
          3737 => x"82",
          3738 => x"a8",
          3739 => x"82",
          3740 => x"39",
          3741 => x"80",
          3742 => x"38",
          3743 => x"15",
          3744 => x"53",
          3745 => x"8d",
          3746 => x"15",
          3747 => x"76",
          3748 => x"51",
          3749 => x"13",
          3750 => x"8d",
          3751 => x"15",
          3752 => x"c5",
          3753 => x"90",
          3754 => x"0b",
          3755 => x"ff",
          3756 => x"15",
          3757 => x"2e",
          3758 => x"81",
          3759 => x"e4",
          3760 => x"b6",
          3761 => x"dc",
          3762 => x"ff",
          3763 => x"81",
          3764 => x"06",
          3765 => x"81",
          3766 => x"51",
          3767 => x"82",
          3768 => x"80",
          3769 => x"8c",
          3770 => x"15",
          3771 => x"14",
          3772 => x"3f",
          3773 => x"08",
          3774 => x"06",
          3775 => x"d4",
          3776 => x"81",
          3777 => x"38",
          3778 => x"d8",
          3779 => x"8c",
          3780 => x"8b",
          3781 => x"2e",
          3782 => x"b3",
          3783 => x"14",
          3784 => x"3f",
          3785 => x"08",
          3786 => x"e4",
          3787 => x"81",
          3788 => x"84",
          3789 => x"d7",
          3790 => x"8c",
          3791 => x"15",
          3792 => x"14",
          3793 => x"3f",
          3794 => x"08",
          3795 => x"76",
          3796 => x"8d",
          3797 => x"05",
          3798 => x"8d",
          3799 => x"86",
          3800 => x"0b",
          3801 => x"80",
          3802 => x"8c",
          3803 => x"3d",
          3804 => x"3d",
          3805 => x"89",
          3806 => x"2e",
          3807 => x"08",
          3808 => x"2e",
          3809 => x"33",
          3810 => x"2e",
          3811 => x"13",
          3812 => x"22",
          3813 => x"76",
          3814 => x"06",
          3815 => x"13",
          3816 => x"c0",
          3817 => x"dc",
          3818 => x"52",
          3819 => x"71",
          3820 => x"55",
          3821 => x"53",
          3822 => x"0c",
          3823 => x"8c",
          3824 => x"3d",
          3825 => x"3d",
          3826 => x"05",
          3827 => x"89",
          3828 => x"52",
          3829 => x"3f",
          3830 => x"0b",
          3831 => x"08",
          3832 => x"82",
          3833 => x"84",
          3834 => x"8c",
          3835 => x"55",
          3836 => x"2e",
          3837 => x"74",
          3838 => x"73",
          3839 => x"38",
          3840 => x"78",
          3841 => x"54",
          3842 => x"92",
          3843 => x"89",
          3844 => x"84",
          3845 => x"b0",
          3846 => x"dc",
          3847 => x"82",
          3848 => x"88",
          3849 => x"eb",
          3850 => x"02",
          3851 => x"e7",
          3852 => x"59",
          3853 => x"80",
          3854 => x"38",
          3855 => x"70",
          3856 => x"d0",
          3857 => x"3d",
          3858 => x"58",
          3859 => x"82",
          3860 => x"55",
          3861 => x"08",
          3862 => x"7a",
          3863 => x"8c",
          3864 => x"56",
          3865 => x"82",
          3866 => x"55",
          3867 => x"08",
          3868 => x"80",
          3869 => x"70",
          3870 => x"57",
          3871 => x"83",
          3872 => x"77",
          3873 => x"73",
          3874 => x"ab",
          3875 => x"2e",
          3876 => x"84",
          3877 => x"06",
          3878 => x"51",
          3879 => x"82",
          3880 => x"55",
          3881 => x"b2",
          3882 => x"06",
          3883 => x"b8",
          3884 => x"2a",
          3885 => x"51",
          3886 => x"2e",
          3887 => x"55",
          3888 => x"77",
          3889 => x"74",
          3890 => x"77",
          3891 => x"81",
          3892 => x"73",
          3893 => x"af",
          3894 => x"7a",
          3895 => x"3f",
          3896 => x"08",
          3897 => x"b2",
          3898 => x"8e",
          3899 => x"ea",
          3900 => x"a0",
          3901 => x"34",
          3902 => x"52",
          3903 => x"bd",
          3904 => x"62",
          3905 => x"d4",
          3906 => x"54",
          3907 => x"15",
          3908 => x"2e",
          3909 => x"7a",
          3910 => x"51",
          3911 => x"75",
          3912 => x"d4",
          3913 => x"be",
          3914 => x"dc",
          3915 => x"8c",
          3916 => x"ca",
          3917 => x"74",
          3918 => x"02",
          3919 => x"70",
          3920 => x"81",
          3921 => x"56",
          3922 => x"86",
          3923 => x"82",
          3924 => x"81",
          3925 => x"06",
          3926 => x"80",
          3927 => x"75",
          3928 => x"73",
          3929 => x"38",
          3930 => x"92",
          3931 => x"7a",
          3932 => x"3f",
          3933 => x"08",
          3934 => x"8c",
          3935 => x"55",
          3936 => x"08",
          3937 => x"77",
          3938 => x"81",
          3939 => x"73",
          3940 => x"38",
          3941 => x"07",
          3942 => x"11",
          3943 => x"0c",
          3944 => x"0c",
          3945 => x"52",
          3946 => x"3f",
          3947 => x"08",
          3948 => x"08",
          3949 => x"63",
          3950 => x"5a",
          3951 => x"82",
          3952 => x"82",
          3953 => x"8c",
          3954 => x"7a",
          3955 => x"17",
          3956 => x"23",
          3957 => x"34",
          3958 => x"1a",
          3959 => x"9c",
          3960 => x"0b",
          3961 => x"77",
          3962 => x"81",
          3963 => x"73",
          3964 => x"8d",
          3965 => x"dc",
          3966 => x"81",
          3967 => x"8c",
          3968 => x"1a",
          3969 => x"22",
          3970 => x"7b",
          3971 => x"a8",
          3972 => x"78",
          3973 => x"3f",
          3974 => x"08",
          3975 => x"dc",
          3976 => x"83",
          3977 => x"82",
          3978 => x"ff",
          3979 => x"06",
          3980 => x"55",
          3981 => x"56",
          3982 => x"76",
          3983 => x"51",
          3984 => x"27",
          3985 => x"70",
          3986 => x"5a",
          3987 => x"76",
          3988 => x"74",
          3989 => x"83",
          3990 => x"73",
          3991 => x"38",
          3992 => x"51",
          3993 => x"82",
          3994 => x"85",
          3995 => x"8e",
          3996 => x"2a",
          3997 => x"08",
          3998 => x"0c",
          3999 => x"79",
          4000 => x"73",
          4001 => x"0c",
          4002 => x"04",
          4003 => x"60",
          4004 => x"40",
          4005 => x"80",
          4006 => x"3d",
          4007 => x"78",
          4008 => x"3f",
          4009 => x"08",
          4010 => x"dc",
          4011 => x"91",
          4012 => x"74",
          4013 => x"38",
          4014 => x"c4",
          4015 => x"33",
          4016 => x"87",
          4017 => x"2e",
          4018 => x"95",
          4019 => x"91",
          4020 => x"56",
          4021 => x"81",
          4022 => x"34",
          4023 => x"a0",
          4024 => x"08",
          4025 => x"31",
          4026 => x"27",
          4027 => x"5c",
          4028 => x"82",
          4029 => x"19",
          4030 => x"ff",
          4031 => x"74",
          4032 => x"7e",
          4033 => x"ff",
          4034 => x"2a",
          4035 => x"79",
          4036 => x"87",
          4037 => x"08",
          4038 => x"98",
          4039 => x"78",
          4040 => x"3f",
          4041 => x"08",
          4042 => x"27",
          4043 => x"74",
          4044 => x"a3",
          4045 => x"1a",
          4046 => x"08",
          4047 => x"d4",
          4048 => x"8c",
          4049 => x"2e",
          4050 => x"82",
          4051 => x"1a",
          4052 => x"59",
          4053 => x"2e",
          4054 => x"77",
          4055 => x"11",
          4056 => x"55",
          4057 => x"85",
          4058 => x"31",
          4059 => x"76",
          4060 => x"81",
          4061 => x"ca",
          4062 => x"8c",
          4063 => x"d7",
          4064 => x"11",
          4065 => x"74",
          4066 => x"38",
          4067 => x"77",
          4068 => x"78",
          4069 => x"84",
          4070 => x"16",
          4071 => x"08",
          4072 => x"2b",
          4073 => x"cf",
          4074 => x"89",
          4075 => x"39",
          4076 => x"0c",
          4077 => x"83",
          4078 => x"80",
          4079 => x"55",
          4080 => x"83",
          4081 => x"9c",
          4082 => x"7e",
          4083 => x"3f",
          4084 => x"08",
          4085 => x"75",
          4086 => x"08",
          4087 => x"1f",
          4088 => x"7c",
          4089 => x"3f",
          4090 => x"7e",
          4091 => x"0c",
          4092 => x"1b",
          4093 => x"1c",
          4094 => x"fd",
          4095 => x"56",
          4096 => x"dc",
          4097 => x"0d",
          4098 => x"0d",
          4099 => x"64",
          4100 => x"58",
          4101 => x"90",
          4102 => x"52",
          4103 => x"d2",
          4104 => x"dc",
          4105 => x"8c",
          4106 => x"38",
          4107 => x"55",
          4108 => x"86",
          4109 => x"83",
          4110 => x"18",
          4111 => x"2a",
          4112 => x"51",
          4113 => x"56",
          4114 => x"83",
          4115 => x"39",
          4116 => x"19",
          4117 => x"83",
          4118 => x"0b",
          4119 => x"81",
          4120 => x"39",
          4121 => x"7c",
          4122 => x"74",
          4123 => x"38",
          4124 => x"7b",
          4125 => x"ec",
          4126 => x"08",
          4127 => x"06",
          4128 => x"81",
          4129 => x"8a",
          4130 => x"05",
          4131 => x"06",
          4132 => x"bf",
          4133 => x"38",
          4134 => x"55",
          4135 => x"7a",
          4136 => x"98",
          4137 => x"77",
          4138 => x"3f",
          4139 => x"08",
          4140 => x"dc",
          4141 => x"82",
          4142 => x"81",
          4143 => x"38",
          4144 => x"ff",
          4145 => x"98",
          4146 => x"18",
          4147 => x"74",
          4148 => x"7e",
          4149 => x"08",
          4150 => x"2e",
          4151 => x"8d",
          4152 => x"ce",
          4153 => x"8c",
          4154 => x"ee",
          4155 => x"08",
          4156 => x"d1",
          4157 => x"8c",
          4158 => x"2e",
          4159 => x"82",
          4160 => x"1b",
          4161 => x"5a",
          4162 => x"2e",
          4163 => x"78",
          4164 => x"11",
          4165 => x"55",
          4166 => x"85",
          4167 => x"31",
          4168 => x"76",
          4169 => x"81",
          4170 => x"c8",
          4171 => x"8c",
          4172 => x"a6",
          4173 => x"11",
          4174 => x"56",
          4175 => x"27",
          4176 => x"80",
          4177 => x"08",
          4178 => x"2b",
          4179 => x"b4",
          4180 => x"b5",
          4181 => x"80",
          4182 => x"34",
          4183 => x"56",
          4184 => x"8c",
          4185 => x"19",
          4186 => x"38",
          4187 => x"b6",
          4188 => x"dc",
          4189 => x"38",
          4190 => x"12",
          4191 => x"9c",
          4192 => x"18",
          4193 => x"06",
          4194 => x"31",
          4195 => x"76",
          4196 => x"7b",
          4197 => x"08",
          4198 => x"cd",
          4199 => x"8c",
          4200 => x"b6",
          4201 => x"7c",
          4202 => x"08",
          4203 => x"1f",
          4204 => x"cb",
          4205 => x"55",
          4206 => x"16",
          4207 => x"31",
          4208 => x"7f",
          4209 => x"94",
          4210 => x"70",
          4211 => x"8c",
          4212 => x"58",
          4213 => x"76",
          4214 => x"75",
          4215 => x"19",
          4216 => x"39",
          4217 => x"80",
          4218 => x"74",
          4219 => x"80",
          4220 => x"8c",
          4221 => x"3d",
          4222 => x"3d",
          4223 => x"3d",
          4224 => x"70",
          4225 => x"ea",
          4226 => x"dc",
          4227 => x"8c",
          4228 => x"fb",
          4229 => x"33",
          4230 => x"70",
          4231 => x"55",
          4232 => x"2e",
          4233 => x"a0",
          4234 => x"78",
          4235 => x"3f",
          4236 => x"08",
          4237 => x"dc",
          4238 => x"38",
          4239 => x"8b",
          4240 => x"07",
          4241 => x"8b",
          4242 => x"16",
          4243 => x"52",
          4244 => x"dd",
          4245 => x"16",
          4246 => x"15",
          4247 => x"3f",
          4248 => x"0a",
          4249 => x"51",
          4250 => x"76",
          4251 => x"51",
          4252 => x"78",
          4253 => x"83",
          4254 => x"51",
          4255 => x"82",
          4256 => x"90",
          4257 => x"bf",
          4258 => x"73",
          4259 => x"76",
          4260 => x"0c",
          4261 => x"04",
          4262 => x"76",
          4263 => x"fe",
          4264 => x"8c",
          4265 => x"82",
          4266 => x"9c",
          4267 => x"fc",
          4268 => x"51",
          4269 => x"82",
          4270 => x"53",
          4271 => x"08",
          4272 => x"8c",
          4273 => x"0c",
          4274 => x"dc",
          4275 => x"0d",
          4276 => x"0d",
          4277 => x"e6",
          4278 => x"52",
          4279 => x"8c",
          4280 => x"8b",
          4281 => x"dc",
          4282 => x"a0",
          4283 => x"71",
          4284 => x"0c",
          4285 => x"04",
          4286 => x"80",
          4287 => x"d0",
          4288 => x"3d",
          4289 => x"3f",
          4290 => x"08",
          4291 => x"dc",
          4292 => x"38",
          4293 => x"52",
          4294 => x"05",
          4295 => x"3f",
          4296 => x"08",
          4297 => x"dc",
          4298 => x"02",
          4299 => x"33",
          4300 => x"55",
          4301 => x"25",
          4302 => x"7a",
          4303 => x"54",
          4304 => x"a2",
          4305 => x"84",
          4306 => x"06",
          4307 => x"73",
          4308 => x"38",
          4309 => x"70",
          4310 => x"a8",
          4311 => x"dc",
          4312 => x"0c",
          4313 => x"8c",
          4314 => x"2e",
          4315 => x"83",
          4316 => x"74",
          4317 => x"0c",
          4318 => x"04",
          4319 => x"6f",
          4320 => x"80",
          4321 => x"53",
          4322 => x"b8",
          4323 => x"3d",
          4324 => x"3f",
          4325 => x"08",
          4326 => x"dc",
          4327 => x"38",
          4328 => x"7c",
          4329 => x"47",
          4330 => x"54",
          4331 => x"81",
          4332 => x"52",
          4333 => x"52",
          4334 => x"3f",
          4335 => x"08",
          4336 => x"dc",
          4337 => x"38",
          4338 => x"51",
          4339 => x"82",
          4340 => x"57",
          4341 => x"08",
          4342 => x"69",
          4343 => x"da",
          4344 => x"8c",
          4345 => x"76",
          4346 => x"d5",
          4347 => x"8c",
          4348 => x"82",
          4349 => x"82",
          4350 => x"52",
          4351 => x"eb",
          4352 => x"dc",
          4353 => x"8c",
          4354 => x"38",
          4355 => x"51",
          4356 => x"73",
          4357 => x"08",
          4358 => x"76",
          4359 => x"d6",
          4360 => x"8c",
          4361 => x"82",
          4362 => x"80",
          4363 => x"76",
          4364 => x"81",
          4365 => x"82",
          4366 => x"39",
          4367 => x"38",
          4368 => x"bc",
          4369 => x"51",
          4370 => x"76",
          4371 => x"11",
          4372 => x"51",
          4373 => x"73",
          4374 => x"38",
          4375 => x"55",
          4376 => x"16",
          4377 => x"56",
          4378 => x"38",
          4379 => x"73",
          4380 => x"90",
          4381 => x"2e",
          4382 => x"16",
          4383 => x"ff",
          4384 => x"ff",
          4385 => x"58",
          4386 => x"74",
          4387 => x"75",
          4388 => x"18",
          4389 => x"58",
          4390 => x"fe",
          4391 => x"7b",
          4392 => x"06",
          4393 => x"18",
          4394 => x"58",
          4395 => x"80",
          4396 => x"a0",
          4397 => x"29",
          4398 => x"05",
          4399 => x"33",
          4400 => x"56",
          4401 => x"2e",
          4402 => x"16",
          4403 => x"33",
          4404 => x"73",
          4405 => x"16",
          4406 => x"26",
          4407 => x"55",
          4408 => x"91",
          4409 => x"54",
          4410 => x"70",
          4411 => x"34",
          4412 => x"ec",
          4413 => x"70",
          4414 => x"34",
          4415 => x"09",
          4416 => x"38",
          4417 => x"39",
          4418 => x"19",
          4419 => x"33",
          4420 => x"05",
          4421 => x"78",
          4422 => x"80",
          4423 => x"82",
          4424 => x"9e",
          4425 => x"f7",
          4426 => x"7d",
          4427 => x"05",
          4428 => x"57",
          4429 => x"3f",
          4430 => x"08",
          4431 => x"dc",
          4432 => x"38",
          4433 => x"53",
          4434 => x"38",
          4435 => x"54",
          4436 => x"92",
          4437 => x"33",
          4438 => x"70",
          4439 => x"54",
          4440 => x"38",
          4441 => x"15",
          4442 => x"70",
          4443 => x"58",
          4444 => x"82",
          4445 => x"8a",
          4446 => x"89",
          4447 => x"53",
          4448 => x"b7",
          4449 => x"ff",
          4450 => x"ff",
          4451 => x"8c",
          4452 => x"15",
          4453 => x"53",
          4454 => x"ff",
          4455 => x"8c",
          4456 => x"26",
          4457 => x"30",
          4458 => x"70",
          4459 => x"77",
          4460 => x"18",
          4461 => x"51",
          4462 => x"88",
          4463 => x"73",
          4464 => x"52",
          4465 => x"ca",
          4466 => x"dc",
          4467 => x"8c",
          4468 => x"2e",
          4469 => x"82",
          4470 => x"ff",
          4471 => x"38",
          4472 => x"08",
          4473 => x"73",
          4474 => x"73",
          4475 => x"9c",
          4476 => x"27",
          4477 => x"75",
          4478 => x"16",
          4479 => x"17",
          4480 => x"33",
          4481 => x"70",
          4482 => x"55",
          4483 => x"80",
          4484 => x"73",
          4485 => x"cc",
          4486 => x"8c",
          4487 => x"82",
          4488 => x"94",
          4489 => x"dc",
          4490 => x"39",
          4491 => x"51",
          4492 => x"82",
          4493 => x"54",
          4494 => x"be",
          4495 => x"27",
          4496 => x"53",
          4497 => x"08",
          4498 => x"73",
          4499 => x"ff",
          4500 => x"15",
          4501 => x"16",
          4502 => x"ff",
          4503 => x"80",
          4504 => x"73",
          4505 => x"c6",
          4506 => x"8c",
          4507 => x"38",
          4508 => x"16",
          4509 => x"80",
          4510 => x"0b",
          4511 => x"81",
          4512 => x"75",
          4513 => x"8c",
          4514 => x"58",
          4515 => x"54",
          4516 => x"74",
          4517 => x"73",
          4518 => x"90",
          4519 => x"c0",
          4520 => x"90",
          4521 => x"83",
          4522 => x"72",
          4523 => x"38",
          4524 => x"08",
          4525 => x"77",
          4526 => x"80",
          4527 => x"8c",
          4528 => x"3d",
          4529 => x"3d",
          4530 => x"89",
          4531 => x"2e",
          4532 => x"80",
          4533 => x"fc",
          4534 => x"3d",
          4535 => x"e1",
          4536 => x"8c",
          4537 => x"82",
          4538 => x"80",
          4539 => x"76",
          4540 => x"75",
          4541 => x"3f",
          4542 => x"08",
          4543 => x"dc",
          4544 => x"38",
          4545 => x"70",
          4546 => x"57",
          4547 => x"a2",
          4548 => x"33",
          4549 => x"70",
          4550 => x"55",
          4551 => x"2e",
          4552 => x"16",
          4553 => x"51",
          4554 => x"82",
          4555 => x"88",
          4556 => x"54",
          4557 => x"84",
          4558 => x"52",
          4559 => x"e5",
          4560 => x"dc",
          4561 => x"84",
          4562 => x"06",
          4563 => x"55",
          4564 => x"80",
          4565 => x"80",
          4566 => x"54",
          4567 => x"dc",
          4568 => x"0d",
          4569 => x"0d",
          4570 => x"fc",
          4571 => x"52",
          4572 => x"3f",
          4573 => x"08",
          4574 => x"8c",
          4575 => x"0c",
          4576 => x"04",
          4577 => x"77",
          4578 => x"fc",
          4579 => x"53",
          4580 => x"de",
          4581 => x"dc",
          4582 => x"8c",
          4583 => x"df",
          4584 => x"38",
          4585 => x"08",
          4586 => x"cd",
          4587 => x"8c",
          4588 => x"80",
          4589 => x"8c",
          4590 => x"73",
          4591 => x"3f",
          4592 => x"08",
          4593 => x"dc",
          4594 => x"09",
          4595 => x"38",
          4596 => x"39",
          4597 => x"08",
          4598 => x"52",
          4599 => x"b3",
          4600 => x"73",
          4601 => x"3f",
          4602 => x"08",
          4603 => x"30",
          4604 => x"9f",
          4605 => x"8c",
          4606 => x"51",
          4607 => x"72",
          4608 => x"0c",
          4609 => x"04",
          4610 => x"65",
          4611 => x"89",
          4612 => x"96",
          4613 => x"df",
          4614 => x"8c",
          4615 => x"82",
          4616 => x"b2",
          4617 => x"75",
          4618 => x"3f",
          4619 => x"08",
          4620 => x"dc",
          4621 => x"02",
          4622 => x"33",
          4623 => x"55",
          4624 => x"25",
          4625 => x"55",
          4626 => x"80",
          4627 => x"76",
          4628 => x"d4",
          4629 => x"82",
          4630 => x"94",
          4631 => x"f0",
          4632 => x"65",
          4633 => x"53",
          4634 => x"05",
          4635 => x"51",
          4636 => x"82",
          4637 => x"5b",
          4638 => x"08",
          4639 => x"7c",
          4640 => x"08",
          4641 => x"fe",
          4642 => x"08",
          4643 => x"55",
          4644 => x"91",
          4645 => x"0c",
          4646 => x"81",
          4647 => x"39",
          4648 => x"c7",
          4649 => x"dc",
          4650 => x"55",
          4651 => x"2e",
          4652 => x"bf",
          4653 => x"5f",
          4654 => x"92",
          4655 => x"51",
          4656 => x"82",
          4657 => x"ff",
          4658 => x"82",
          4659 => x"81",
          4660 => x"82",
          4661 => x"30",
          4662 => x"dc",
          4663 => x"25",
          4664 => x"19",
          4665 => x"5a",
          4666 => x"08",
          4667 => x"38",
          4668 => x"a4",
          4669 => x"8c",
          4670 => x"58",
          4671 => x"77",
          4672 => x"7d",
          4673 => x"bf",
          4674 => x"8c",
          4675 => x"82",
          4676 => x"80",
          4677 => x"70",
          4678 => x"ff",
          4679 => x"56",
          4680 => x"2e",
          4681 => x"9e",
          4682 => x"51",
          4683 => x"3f",
          4684 => x"08",
          4685 => x"06",
          4686 => x"80",
          4687 => x"19",
          4688 => x"54",
          4689 => x"14",
          4690 => x"c5",
          4691 => x"dc",
          4692 => x"06",
          4693 => x"80",
          4694 => x"19",
          4695 => x"54",
          4696 => x"06",
          4697 => x"79",
          4698 => x"78",
          4699 => x"79",
          4700 => x"84",
          4701 => x"07",
          4702 => x"84",
          4703 => x"82",
          4704 => x"92",
          4705 => x"f9",
          4706 => x"8a",
          4707 => x"53",
          4708 => x"e3",
          4709 => x"8c",
          4710 => x"82",
          4711 => x"81",
          4712 => x"17",
          4713 => x"81",
          4714 => x"17",
          4715 => x"2a",
          4716 => x"51",
          4717 => x"55",
          4718 => x"81",
          4719 => x"17",
          4720 => x"8c",
          4721 => x"81",
          4722 => x"9b",
          4723 => x"dc",
          4724 => x"17",
          4725 => x"51",
          4726 => x"82",
          4727 => x"74",
          4728 => x"56",
          4729 => x"98",
          4730 => x"76",
          4731 => x"c6",
          4732 => x"dc",
          4733 => x"09",
          4734 => x"38",
          4735 => x"8c",
          4736 => x"2e",
          4737 => x"85",
          4738 => x"a3",
          4739 => x"38",
          4740 => x"8c",
          4741 => x"15",
          4742 => x"38",
          4743 => x"53",
          4744 => x"08",
          4745 => x"c3",
          4746 => x"8c",
          4747 => x"94",
          4748 => x"18",
          4749 => x"33",
          4750 => x"54",
          4751 => x"34",
          4752 => x"85",
          4753 => x"18",
          4754 => x"74",
          4755 => x"0c",
          4756 => x"04",
          4757 => x"82",
          4758 => x"ff",
          4759 => x"a1",
          4760 => x"e4",
          4761 => x"dc",
          4762 => x"8c",
          4763 => x"f5",
          4764 => x"a1",
          4765 => x"95",
          4766 => x"58",
          4767 => x"82",
          4768 => x"55",
          4769 => x"08",
          4770 => x"02",
          4771 => x"33",
          4772 => x"70",
          4773 => x"55",
          4774 => x"73",
          4775 => x"75",
          4776 => x"80",
          4777 => x"bd",
          4778 => x"d6",
          4779 => x"81",
          4780 => x"87",
          4781 => x"ad",
          4782 => x"78",
          4783 => x"3f",
          4784 => x"08",
          4785 => x"70",
          4786 => x"55",
          4787 => x"2e",
          4788 => x"78",
          4789 => x"dc",
          4790 => x"08",
          4791 => x"38",
          4792 => x"8c",
          4793 => x"76",
          4794 => x"70",
          4795 => x"b5",
          4796 => x"dc",
          4797 => x"8c",
          4798 => x"e9",
          4799 => x"dc",
          4800 => x"51",
          4801 => x"82",
          4802 => x"55",
          4803 => x"08",
          4804 => x"55",
          4805 => x"82",
          4806 => x"84",
          4807 => x"82",
          4808 => x"80",
          4809 => x"51",
          4810 => x"82",
          4811 => x"82",
          4812 => x"30",
          4813 => x"dc",
          4814 => x"25",
          4815 => x"75",
          4816 => x"38",
          4817 => x"8f",
          4818 => x"75",
          4819 => x"c1",
          4820 => x"8c",
          4821 => x"74",
          4822 => x"51",
          4823 => x"3f",
          4824 => x"08",
          4825 => x"8c",
          4826 => x"3d",
          4827 => x"3d",
          4828 => x"99",
          4829 => x"52",
          4830 => x"d8",
          4831 => x"8c",
          4832 => x"82",
          4833 => x"82",
          4834 => x"5e",
          4835 => x"3d",
          4836 => x"cf",
          4837 => x"8c",
          4838 => x"82",
          4839 => x"86",
          4840 => x"82",
          4841 => x"8c",
          4842 => x"2e",
          4843 => x"82",
          4844 => x"80",
          4845 => x"70",
          4846 => x"06",
          4847 => x"54",
          4848 => x"38",
          4849 => x"52",
          4850 => x"52",
          4851 => x"3f",
          4852 => x"08",
          4853 => x"82",
          4854 => x"83",
          4855 => x"82",
          4856 => x"81",
          4857 => x"06",
          4858 => x"54",
          4859 => x"08",
          4860 => x"81",
          4861 => x"81",
          4862 => x"39",
          4863 => x"38",
          4864 => x"08",
          4865 => x"c4",
          4866 => x"8c",
          4867 => x"82",
          4868 => x"81",
          4869 => x"53",
          4870 => x"19",
          4871 => x"8c",
          4872 => x"ae",
          4873 => x"34",
          4874 => x"0b",
          4875 => x"82",
          4876 => x"52",
          4877 => x"51",
          4878 => x"3f",
          4879 => x"b4",
          4880 => x"c9",
          4881 => x"53",
          4882 => x"53",
          4883 => x"51",
          4884 => x"3f",
          4885 => x"0b",
          4886 => x"34",
          4887 => x"80",
          4888 => x"51",
          4889 => x"78",
          4890 => x"83",
          4891 => x"51",
          4892 => x"82",
          4893 => x"54",
          4894 => x"08",
          4895 => x"88",
          4896 => x"64",
          4897 => x"ff",
          4898 => x"75",
          4899 => x"78",
          4900 => x"3f",
          4901 => x"0b",
          4902 => x"78",
          4903 => x"83",
          4904 => x"51",
          4905 => x"3f",
          4906 => x"08",
          4907 => x"80",
          4908 => x"76",
          4909 => x"ae",
          4910 => x"8c",
          4911 => x"3d",
          4912 => x"3d",
          4913 => x"84",
          4914 => x"f1",
          4915 => x"a8",
          4916 => x"05",
          4917 => x"51",
          4918 => x"82",
          4919 => x"55",
          4920 => x"08",
          4921 => x"78",
          4922 => x"08",
          4923 => x"70",
          4924 => x"b8",
          4925 => x"dc",
          4926 => x"8c",
          4927 => x"b9",
          4928 => x"9b",
          4929 => x"a0",
          4930 => x"55",
          4931 => x"38",
          4932 => x"3d",
          4933 => x"3d",
          4934 => x"51",
          4935 => x"3f",
          4936 => x"52",
          4937 => x"52",
          4938 => x"dd",
          4939 => x"08",
          4940 => x"cb",
          4941 => x"8c",
          4942 => x"82",
          4943 => x"95",
          4944 => x"2e",
          4945 => x"88",
          4946 => x"3d",
          4947 => x"38",
          4948 => x"e5",
          4949 => x"dc",
          4950 => x"09",
          4951 => x"b8",
          4952 => x"c9",
          4953 => x"8c",
          4954 => x"82",
          4955 => x"81",
          4956 => x"56",
          4957 => x"3d",
          4958 => x"52",
          4959 => x"ff",
          4960 => x"02",
          4961 => x"8b",
          4962 => x"16",
          4963 => x"2a",
          4964 => x"51",
          4965 => x"89",
          4966 => x"07",
          4967 => x"17",
          4968 => x"81",
          4969 => x"34",
          4970 => x"70",
          4971 => x"81",
          4972 => x"55",
          4973 => x"80",
          4974 => x"64",
          4975 => x"38",
          4976 => x"51",
          4977 => x"82",
          4978 => x"52",
          4979 => x"b7",
          4980 => x"55",
          4981 => x"08",
          4982 => x"dd",
          4983 => x"dc",
          4984 => x"51",
          4985 => x"3f",
          4986 => x"08",
          4987 => x"11",
          4988 => x"82",
          4989 => x"80",
          4990 => x"16",
          4991 => x"ae",
          4992 => x"06",
          4993 => x"53",
          4994 => x"51",
          4995 => x"78",
          4996 => x"83",
          4997 => x"39",
          4998 => x"08",
          4999 => x"51",
          5000 => x"82",
          5001 => x"55",
          5002 => x"08",
          5003 => x"51",
          5004 => x"3f",
          5005 => x"08",
          5006 => x"8c",
          5007 => x"3d",
          5008 => x"3d",
          5009 => x"db",
          5010 => x"84",
          5011 => x"05",
          5012 => x"82",
          5013 => x"d0",
          5014 => x"3d",
          5015 => x"3f",
          5016 => x"08",
          5017 => x"dc",
          5018 => x"38",
          5019 => x"52",
          5020 => x"05",
          5021 => x"3f",
          5022 => x"08",
          5023 => x"dc",
          5024 => x"02",
          5025 => x"33",
          5026 => x"54",
          5027 => x"aa",
          5028 => x"06",
          5029 => x"8b",
          5030 => x"06",
          5031 => x"07",
          5032 => x"56",
          5033 => x"34",
          5034 => x"0b",
          5035 => x"78",
          5036 => x"a9",
          5037 => x"dc",
          5038 => x"82",
          5039 => x"95",
          5040 => x"ef",
          5041 => x"56",
          5042 => x"3d",
          5043 => x"94",
          5044 => x"f4",
          5045 => x"dc",
          5046 => x"8c",
          5047 => x"cb",
          5048 => x"63",
          5049 => x"d4",
          5050 => x"c0",
          5051 => x"dc",
          5052 => x"8c",
          5053 => x"38",
          5054 => x"05",
          5055 => x"06",
          5056 => x"73",
          5057 => x"16",
          5058 => x"22",
          5059 => x"07",
          5060 => x"1f",
          5061 => x"c2",
          5062 => x"81",
          5063 => x"34",
          5064 => x"b3",
          5065 => x"8c",
          5066 => x"74",
          5067 => x"0c",
          5068 => x"04",
          5069 => x"69",
          5070 => x"80",
          5071 => x"d0",
          5072 => x"3d",
          5073 => x"3f",
          5074 => x"08",
          5075 => x"08",
          5076 => x"8c",
          5077 => x"80",
          5078 => x"57",
          5079 => x"81",
          5080 => x"70",
          5081 => x"55",
          5082 => x"80",
          5083 => x"5d",
          5084 => x"52",
          5085 => x"52",
          5086 => x"a9",
          5087 => x"dc",
          5088 => x"8c",
          5089 => x"d1",
          5090 => x"73",
          5091 => x"3f",
          5092 => x"08",
          5093 => x"dc",
          5094 => x"82",
          5095 => x"82",
          5096 => x"65",
          5097 => x"78",
          5098 => x"7b",
          5099 => x"55",
          5100 => x"34",
          5101 => x"8a",
          5102 => x"38",
          5103 => x"1a",
          5104 => x"34",
          5105 => x"9e",
          5106 => x"70",
          5107 => x"51",
          5108 => x"a0",
          5109 => x"8e",
          5110 => x"2e",
          5111 => x"86",
          5112 => x"34",
          5113 => x"30",
          5114 => x"80",
          5115 => x"7a",
          5116 => x"c1",
          5117 => x"2e",
          5118 => x"a0",
          5119 => x"51",
          5120 => x"3f",
          5121 => x"08",
          5122 => x"dc",
          5123 => x"7b",
          5124 => x"55",
          5125 => x"73",
          5126 => x"38",
          5127 => x"73",
          5128 => x"38",
          5129 => x"15",
          5130 => x"ff",
          5131 => x"82",
          5132 => x"7b",
          5133 => x"8c",
          5134 => x"3d",
          5135 => x"3d",
          5136 => x"9c",
          5137 => x"05",
          5138 => x"51",
          5139 => x"82",
          5140 => x"82",
          5141 => x"56",
          5142 => x"dc",
          5143 => x"38",
          5144 => x"52",
          5145 => x"52",
          5146 => x"c0",
          5147 => x"70",
          5148 => x"ff",
          5149 => x"55",
          5150 => x"27",
          5151 => x"78",
          5152 => x"ff",
          5153 => x"05",
          5154 => x"55",
          5155 => x"3f",
          5156 => x"08",
          5157 => x"38",
          5158 => x"70",
          5159 => x"ff",
          5160 => x"82",
          5161 => x"80",
          5162 => x"74",
          5163 => x"07",
          5164 => x"4e",
          5165 => x"82",
          5166 => x"55",
          5167 => x"70",
          5168 => x"06",
          5169 => x"99",
          5170 => x"e0",
          5171 => x"ff",
          5172 => x"54",
          5173 => x"27",
          5174 => x"f9",
          5175 => x"55",
          5176 => x"a3",
          5177 => x"81",
          5178 => x"ff",
          5179 => x"82",
          5180 => x"93",
          5181 => x"75",
          5182 => x"76",
          5183 => x"38",
          5184 => x"77",
          5185 => x"86",
          5186 => x"39",
          5187 => x"27",
          5188 => x"88",
          5189 => x"78",
          5190 => x"5a",
          5191 => x"57",
          5192 => x"81",
          5193 => x"81",
          5194 => x"33",
          5195 => x"06",
          5196 => x"57",
          5197 => x"fe",
          5198 => x"3d",
          5199 => x"55",
          5200 => x"2e",
          5201 => x"76",
          5202 => x"38",
          5203 => x"55",
          5204 => x"33",
          5205 => x"a0",
          5206 => x"06",
          5207 => x"17",
          5208 => x"38",
          5209 => x"43",
          5210 => x"3d",
          5211 => x"ff",
          5212 => x"82",
          5213 => x"54",
          5214 => x"08",
          5215 => x"81",
          5216 => x"ff",
          5217 => x"82",
          5218 => x"54",
          5219 => x"08",
          5220 => x"80",
          5221 => x"54",
          5222 => x"80",
          5223 => x"8c",
          5224 => x"2e",
          5225 => x"80",
          5226 => x"54",
          5227 => x"80",
          5228 => x"52",
          5229 => x"bd",
          5230 => x"8c",
          5231 => x"82",
          5232 => x"b1",
          5233 => x"82",
          5234 => x"52",
          5235 => x"ab",
          5236 => x"54",
          5237 => x"15",
          5238 => x"78",
          5239 => x"ff",
          5240 => x"79",
          5241 => x"83",
          5242 => x"51",
          5243 => x"3f",
          5244 => x"08",
          5245 => x"74",
          5246 => x"0c",
          5247 => x"04",
          5248 => x"60",
          5249 => x"05",
          5250 => x"33",
          5251 => x"05",
          5252 => x"40",
          5253 => x"da",
          5254 => x"dc",
          5255 => x"8c",
          5256 => x"bd",
          5257 => x"33",
          5258 => x"b5",
          5259 => x"2e",
          5260 => x"1a",
          5261 => x"90",
          5262 => x"33",
          5263 => x"70",
          5264 => x"55",
          5265 => x"38",
          5266 => x"97",
          5267 => x"82",
          5268 => x"58",
          5269 => x"7e",
          5270 => x"70",
          5271 => x"55",
          5272 => x"56",
          5273 => x"f5",
          5274 => x"7d",
          5275 => x"70",
          5276 => x"2a",
          5277 => x"08",
          5278 => x"08",
          5279 => x"5d",
          5280 => x"77",
          5281 => x"98",
          5282 => x"26",
          5283 => x"57",
          5284 => x"59",
          5285 => x"52",
          5286 => x"ae",
          5287 => x"15",
          5288 => x"98",
          5289 => x"26",
          5290 => x"55",
          5291 => x"08",
          5292 => x"99",
          5293 => x"dc",
          5294 => x"ff",
          5295 => x"8c",
          5296 => x"38",
          5297 => x"75",
          5298 => x"81",
          5299 => x"93",
          5300 => x"80",
          5301 => x"2e",
          5302 => x"ff",
          5303 => x"58",
          5304 => x"7d",
          5305 => x"38",
          5306 => x"55",
          5307 => x"b4",
          5308 => x"56",
          5309 => x"09",
          5310 => x"38",
          5311 => x"53",
          5312 => x"51",
          5313 => x"3f",
          5314 => x"08",
          5315 => x"dc",
          5316 => x"38",
          5317 => x"ff",
          5318 => x"5c",
          5319 => x"84",
          5320 => x"5c",
          5321 => x"12",
          5322 => x"80",
          5323 => x"78",
          5324 => x"7c",
          5325 => x"90",
          5326 => x"c0",
          5327 => x"90",
          5328 => x"15",
          5329 => x"90",
          5330 => x"54",
          5331 => x"91",
          5332 => x"31",
          5333 => x"84",
          5334 => x"07",
          5335 => x"16",
          5336 => x"73",
          5337 => x"0c",
          5338 => x"04",
          5339 => x"6b",
          5340 => x"05",
          5341 => x"33",
          5342 => x"5a",
          5343 => x"bd",
          5344 => x"80",
          5345 => x"dc",
          5346 => x"f8",
          5347 => x"dc",
          5348 => x"82",
          5349 => x"70",
          5350 => x"74",
          5351 => x"38",
          5352 => x"82",
          5353 => x"81",
          5354 => x"81",
          5355 => x"ff",
          5356 => x"82",
          5357 => x"81",
          5358 => x"81",
          5359 => x"83",
          5360 => x"c0",
          5361 => x"2a",
          5362 => x"51",
          5363 => x"74",
          5364 => x"99",
          5365 => x"53",
          5366 => x"51",
          5367 => x"3f",
          5368 => x"08",
          5369 => x"55",
          5370 => x"92",
          5371 => x"80",
          5372 => x"38",
          5373 => x"06",
          5374 => x"2e",
          5375 => x"48",
          5376 => x"87",
          5377 => x"79",
          5378 => x"78",
          5379 => x"26",
          5380 => x"19",
          5381 => x"74",
          5382 => x"38",
          5383 => x"e4",
          5384 => x"2a",
          5385 => x"70",
          5386 => x"59",
          5387 => x"7a",
          5388 => x"56",
          5389 => x"80",
          5390 => x"51",
          5391 => x"74",
          5392 => x"99",
          5393 => x"53",
          5394 => x"51",
          5395 => x"3f",
          5396 => x"8c",
          5397 => x"ac",
          5398 => x"2a",
          5399 => x"82",
          5400 => x"43",
          5401 => x"83",
          5402 => x"66",
          5403 => x"60",
          5404 => x"90",
          5405 => x"31",
          5406 => x"80",
          5407 => x"8a",
          5408 => x"56",
          5409 => x"26",
          5410 => x"77",
          5411 => x"81",
          5412 => x"74",
          5413 => x"38",
          5414 => x"55",
          5415 => x"83",
          5416 => x"81",
          5417 => x"80",
          5418 => x"38",
          5419 => x"55",
          5420 => x"5e",
          5421 => x"89",
          5422 => x"5a",
          5423 => x"09",
          5424 => x"e1",
          5425 => x"38",
          5426 => x"57",
          5427 => x"fc",
          5428 => x"5a",
          5429 => x"9d",
          5430 => x"26",
          5431 => x"fc",
          5432 => x"10",
          5433 => x"22",
          5434 => x"74",
          5435 => x"38",
          5436 => x"ee",
          5437 => x"66",
          5438 => x"e1",
          5439 => x"dc",
          5440 => x"84",
          5441 => x"89",
          5442 => x"a0",
          5443 => x"82",
          5444 => x"fc",
          5445 => x"56",
          5446 => x"f0",
          5447 => x"80",
          5448 => x"d3",
          5449 => x"38",
          5450 => x"57",
          5451 => x"fc",
          5452 => x"5a",
          5453 => x"9d",
          5454 => x"26",
          5455 => x"fc",
          5456 => x"10",
          5457 => x"22",
          5458 => x"74",
          5459 => x"38",
          5460 => x"ee",
          5461 => x"66",
          5462 => x"81",
          5463 => x"dc",
          5464 => x"05",
          5465 => x"dc",
          5466 => x"26",
          5467 => x"0b",
          5468 => x"08",
          5469 => x"dc",
          5470 => x"11",
          5471 => x"05",
          5472 => x"83",
          5473 => x"2a",
          5474 => x"a0",
          5475 => x"7d",
          5476 => x"69",
          5477 => x"05",
          5478 => x"72",
          5479 => x"5c",
          5480 => x"59",
          5481 => x"2e",
          5482 => x"89",
          5483 => x"60",
          5484 => x"84",
          5485 => x"5d",
          5486 => x"18",
          5487 => x"68",
          5488 => x"74",
          5489 => x"af",
          5490 => x"31",
          5491 => x"53",
          5492 => x"52",
          5493 => x"85",
          5494 => x"dc",
          5495 => x"83",
          5496 => x"06",
          5497 => x"8c",
          5498 => x"ff",
          5499 => x"dd",
          5500 => x"83",
          5501 => x"2a",
          5502 => x"be",
          5503 => x"39",
          5504 => x"09",
          5505 => x"c5",
          5506 => x"f5",
          5507 => x"dc",
          5508 => x"38",
          5509 => x"79",
          5510 => x"80",
          5511 => x"38",
          5512 => x"96",
          5513 => x"06",
          5514 => x"2e",
          5515 => x"5e",
          5516 => x"82",
          5517 => x"9f",
          5518 => x"38",
          5519 => x"38",
          5520 => x"81",
          5521 => x"fc",
          5522 => x"ab",
          5523 => x"7d",
          5524 => x"81",
          5525 => x"7d",
          5526 => x"78",
          5527 => x"74",
          5528 => x"8e",
          5529 => x"9c",
          5530 => x"53",
          5531 => x"51",
          5532 => x"3f",
          5533 => x"fa",
          5534 => x"51",
          5535 => x"3f",
          5536 => x"8b",
          5537 => x"a1",
          5538 => x"8d",
          5539 => x"83",
          5540 => x"52",
          5541 => x"ff",
          5542 => x"81",
          5543 => x"34",
          5544 => x"70",
          5545 => x"2a",
          5546 => x"54",
          5547 => x"1b",
          5548 => x"88",
          5549 => x"74",
          5550 => x"26",
          5551 => x"83",
          5552 => x"52",
          5553 => x"ff",
          5554 => x"8a",
          5555 => x"a0",
          5556 => x"a1",
          5557 => x"0b",
          5558 => x"bf",
          5559 => x"51",
          5560 => x"3f",
          5561 => x"9a",
          5562 => x"a0",
          5563 => x"52",
          5564 => x"ff",
          5565 => x"7d",
          5566 => x"81",
          5567 => x"38",
          5568 => x"0a",
          5569 => x"1b",
          5570 => x"ce",
          5571 => x"a4",
          5572 => x"a0",
          5573 => x"52",
          5574 => x"ff",
          5575 => x"81",
          5576 => x"51",
          5577 => x"3f",
          5578 => x"1b",
          5579 => x"8c",
          5580 => x"0b",
          5581 => x"34",
          5582 => x"c2",
          5583 => x"53",
          5584 => x"52",
          5585 => x"51",
          5586 => x"88",
          5587 => x"a7",
          5588 => x"a0",
          5589 => x"83",
          5590 => x"52",
          5591 => x"ff",
          5592 => x"ff",
          5593 => x"1c",
          5594 => x"a6",
          5595 => x"53",
          5596 => x"52",
          5597 => x"ff",
          5598 => x"82",
          5599 => x"83",
          5600 => x"52",
          5601 => x"b4",
          5602 => x"60",
          5603 => x"7e",
          5604 => x"d7",
          5605 => x"82",
          5606 => x"83",
          5607 => x"83",
          5608 => x"06",
          5609 => x"75",
          5610 => x"05",
          5611 => x"7e",
          5612 => x"b7",
          5613 => x"53",
          5614 => x"51",
          5615 => x"3f",
          5616 => x"a4",
          5617 => x"51",
          5618 => x"3f",
          5619 => x"e4",
          5620 => x"e4",
          5621 => x"9f",
          5622 => x"18",
          5623 => x"1b",
          5624 => x"f6",
          5625 => x"83",
          5626 => x"ff",
          5627 => x"82",
          5628 => x"78",
          5629 => x"c4",
          5630 => x"60",
          5631 => x"7a",
          5632 => x"ff",
          5633 => x"75",
          5634 => x"53",
          5635 => x"51",
          5636 => x"3f",
          5637 => x"52",
          5638 => x"9f",
          5639 => x"56",
          5640 => x"83",
          5641 => x"06",
          5642 => x"52",
          5643 => x"9e",
          5644 => x"52",
          5645 => x"ff",
          5646 => x"f0",
          5647 => x"1b",
          5648 => x"87",
          5649 => x"55",
          5650 => x"83",
          5651 => x"74",
          5652 => x"ff",
          5653 => x"7c",
          5654 => x"74",
          5655 => x"38",
          5656 => x"54",
          5657 => x"52",
          5658 => x"99",
          5659 => x"8c",
          5660 => x"87",
          5661 => x"53",
          5662 => x"08",
          5663 => x"ff",
          5664 => x"76",
          5665 => x"31",
          5666 => x"cd",
          5667 => x"58",
          5668 => x"ff",
          5669 => x"55",
          5670 => x"83",
          5671 => x"61",
          5672 => x"26",
          5673 => x"57",
          5674 => x"53",
          5675 => x"51",
          5676 => x"3f",
          5677 => x"08",
          5678 => x"76",
          5679 => x"31",
          5680 => x"db",
          5681 => x"7d",
          5682 => x"38",
          5683 => x"83",
          5684 => x"8a",
          5685 => x"7d",
          5686 => x"38",
          5687 => x"81",
          5688 => x"80",
          5689 => x"80",
          5690 => x"7a",
          5691 => x"bc",
          5692 => x"d5",
          5693 => x"ff",
          5694 => x"83",
          5695 => x"77",
          5696 => x"0b",
          5697 => x"81",
          5698 => x"34",
          5699 => x"34",
          5700 => x"34",
          5701 => x"56",
          5702 => x"52",
          5703 => x"d8",
          5704 => x"0b",
          5705 => x"82",
          5706 => x"82",
          5707 => x"56",
          5708 => x"34",
          5709 => x"08",
          5710 => x"60",
          5711 => x"1b",
          5712 => x"96",
          5713 => x"83",
          5714 => x"ff",
          5715 => x"81",
          5716 => x"7a",
          5717 => x"ff",
          5718 => x"81",
          5719 => x"dc",
          5720 => x"80",
          5721 => x"7e",
          5722 => x"e3",
          5723 => x"82",
          5724 => x"90",
          5725 => x"8e",
          5726 => x"81",
          5727 => x"82",
          5728 => x"56",
          5729 => x"dc",
          5730 => x"0d",
          5731 => x"0d",
          5732 => x"59",
          5733 => x"ff",
          5734 => x"57",
          5735 => x"b4",
          5736 => x"f8",
          5737 => x"81",
          5738 => x"52",
          5739 => x"dc",
          5740 => x"2e",
          5741 => x"9c",
          5742 => x"33",
          5743 => x"2e",
          5744 => x"76",
          5745 => x"58",
          5746 => x"57",
          5747 => x"09",
          5748 => x"38",
          5749 => x"78",
          5750 => x"38",
          5751 => x"82",
          5752 => x"8d",
          5753 => x"f7",
          5754 => x"02",
          5755 => x"05",
          5756 => x"77",
          5757 => x"81",
          5758 => x"8d",
          5759 => x"e7",
          5760 => x"08",
          5761 => x"24",
          5762 => x"17",
          5763 => x"8c",
          5764 => x"77",
          5765 => x"16",
          5766 => x"25",
          5767 => x"3d",
          5768 => x"75",
          5769 => x"52",
          5770 => x"cb",
          5771 => x"76",
          5772 => x"70",
          5773 => x"2a",
          5774 => x"51",
          5775 => x"84",
          5776 => x"19",
          5777 => x"8b",
          5778 => x"f9",
          5779 => x"84",
          5780 => x"56",
          5781 => x"a7",
          5782 => x"fc",
          5783 => x"53",
          5784 => x"75",
          5785 => x"a1",
          5786 => x"dc",
          5787 => x"84",
          5788 => x"2e",
          5789 => x"87",
          5790 => x"08",
          5791 => x"ff",
          5792 => x"8c",
          5793 => x"3d",
          5794 => x"3d",
          5795 => x"80",
          5796 => x"52",
          5797 => x"9a",
          5798 => x"74",
          5799 => x"0d",
          5800 => x"0d",
          5801 => x"05",
          5802 => x"86",
          5803 => x"54",
          5804 => x"73",
          5805 => x"fe",
          5806 => x"51",
          5807 => x"98",
          5808 => x"f8",
          5809 => x"70",
          5810 => x"56",
          5811 => x"2e",
          5812 => x"8c",
          5813 => x"79",
          5814 => x"33",
          5815 => x"39",
          5816 => x"73",
          5817 => x"81",
          5818 => x"81",
          5819 => x"39",
          5820 => x"90",
          5821 => x"cc",
          5822 => x"52",
          5823 => x"f0",
          5824 => x"dc",
          5825 => x"dc",
          5826 => x"53",
          5827 => x"58",
          5828 => x"3f",
          5829 => x"08",
          5830 => x"16",
          5831 => x"81",
          5832 => x"38",
          5833 => x"81",
          5834 => x"54",
          5835 => x"c2",
          5836 => x"73",
          5837 => x"0c",
          5838 => x"04",
          5839 => x"73",
          5840 => x"26",
          5841 => x"71",
          5842 => x"f1",
          5843 => x"71",
          5844 => x"fd",
          5845 => x"80",
          5846 => x"d4",
          5847 => x"39",
          5848 => x"51",
          5849 => x"81",
          5850 => x"80",
          5851 => x"fe",
          5852 => x"e4",
          5853 => x"9c",
          5854 => x"39",
          5855 => x"51",
          5856 => x"81",
          5857 => x"80",
          5858 => x"fe",
          5859 => x"c8",
          5860 => x"f0",
          5861 => x"39",
          5862 => x"51",
          5863 => x"ff",
          5864 => x"39",
          5865 => x"51",
          5866 => x"ff",
          5867 => x"39",
          5868 => x"51",
          5869 => x"80",
          5870 => x"39",
          5871 => x"51",
          5872 => x"80",
          5873 => x"39",
          5874 => x"51",
          5875 => x"80",
          5876 => x"39",
          5877 => x"51",
          5878 => x"3f",
          5879 => x"04",
          5880 => x"77",
          5881 => x"74",
          5882 => x"8a",
          5883 => x"75",
          5884 => x"51",
          5885 => x"e8",
          5886 => x"fe",
          5887 => x"82",
          5888 => x"52",
          5889 => x"d2",
          5890 => x"8c",
          5891 => x"79",
          5892 => x"82",
          5893 => x"fe",
          5894 => x"87",
          5895 => x"ec",
          5896 => x"02",
          5897 => x"e3",
          5898 => x"57",
          5899 => x"30",
          5900 => x"73",
          5901 => x"59",
          5902 => x"77",
          5903 => x"83",
          5904 => x"74",
          5905 => x"81",
          5906 => x"55",
          5907 => x"81",
          5908 => x"53",
          5909 => x"3d",
          5910 => x"ff",
          5911 => x"82",
          5912 => x"57",
          5913 => x"08",
          5914 => x"8c",
          5915 => x"c0",
          5916 => x"82",
          5917 => x"59",
          5918 => x"05",
          5919 => x"53",
          5920 => x"51",
          5921 => x"82",
          5922 => x"57",
          5923 => x"08",
          5924 => x"55",
          5925 => x"89",
          5926 => x"75",
          5927 => x"d8",
          5928 => x"d8",
          5929 => x"f0",
          5930 => x"70",
          5931 => x"25",
          5932 => x"9f",
          5933 => x"51",
          5934 => x"74",
          5935 => x"38",
          5936 => x"53",
          5937 => x"88",
          5938 => x"51",
          5939 => x"76",
          5940 => x"8c",
          5941 => x"3d",
          5942 => x"3d",
          5943 => x"84",
          5944 => x"33",
          5945 => x"57",
          5946 => x"52",
          5947 => x"af",
          5948 => x"dc",
          5949 => x"75",
          5950 => x"38",
          5951 => x"98",
          5952 => x"60",
          5953 => x"82",
          5954 => x"7e",
          5955 => x"77",
          5956 => x"dc",
          5957 => x"39",
          5958 => x"82",
          5959 => x"89",
          5960 => x"f3",
          5961 => x"61",
          5962 => x"05",
          5963 => x"33",
          5964 => x"68",
          5965 => x"5c",
          5966 => x"7a",
          5967 => x"bc",
          5968 => x"a9",
          5969 => x"c4",
          5970 => x"bd",
          5971 => x"74",
          5972 => x"fc",
          5973 => x"2e",
          5974 => x"a0",
          5975 => x"80",
          5976 => x"18",
          5977 => x"27",
          5978 => x"22",
          5979 => x"c8",
          5980 => x"f9",
          5981 => x"82",
          5982 => x"fe",
          5983 => x"82",
          5984 => x"c3",
          5985 => x"53",
          5986 => x"8e",
          5987 => x"52",
          5988 => x"51",
          5989 => x"3f",
          5990 => x"81",
          5991 => x"ee",
          5992 => x"15",
          5993 => x"74",
          5994 => x"7a",
          5995 => x"72",
          5996 => x"81",
          5997 => x"f4",
          5998 => x"39",
          5999 => x"51",
          6000 => x"3f",
          6001 => x"a0",
          6002 => x"e0",
          6003 => x"39",
          6004 => x"51",
          6005 => x"3f",
          6006 => x"79",
          6007 => x"74",
          6008 => x"55",
          6009 => x"72",
          6010 => x"38",
          6011 => x"53",
          6012 => x"83",
          6013 => x"75",
          6014 => x"81",
          6015 => x"53",
          6016 => x"8b",
          6017 => x"fe",
          6018 => x"73",
          6019 => x"a0",
          6020 => x"98",
          6021 => x"55",
          6022 => x"81",
          6023 => x"ed",
          6024 => x"18",
          6025 => x"58",
          6026 => x"3f",
          6027 => x"08",
          6028 => x"98",
          6029 => x"76",
          6030 => x"81",
          6031 => x"fe",
          6032 => x"82",
          6033 => x"98",
          6034 => x"2c",
          6035 => x"70",
          6036 => x"32",
          6037 => x"72",
          6038 => x"07",
          6039 => x"58",
          6040 => x"57",
          6041 => x"d7",
          6042 => x"2e",
          6043 => x"85",
          6044 => x"8c",
          6045 => x"53",
          6046 => x"fd",
          6047 => x"53",
          6048 => x"dc",
          6049 => x"0d",
          6050 => x"0d",
          6051 => x"33",
          6052 => x"53",
          6053 => x"52",
          6054 => x"d1",
          6055 => x"8c",
          6056 => x"e7",
          6057 => x"82",
          6058 => x"82",
          6059 => x"88",
          6060 => x"82",
          6061 => x"fe",
          6062 => x"74",
          6063 => x"38",
          6064 => x"3f",
          6065 => x"04",
          6066 => x"87",
          6067 => x"08",
          6068 => x"b1",
          6069 => x"fe",
          6070 => x"82",
          6071 => x"fe",
          6072 => x"80",
          6073 => x"ac",
          6074 => x"2a",
          6075 => x"51",
          6076 => x"2e",
          6077 => x"51",
          6078 => x"3f",
          6079 => x"51",
          6080 => x"3f",
          6081 => x"d9",
          6082 => x"82",
          6083 => x"06",
          6084 => x"80",
          6085 => x"81",
          6086 => x"f8",
          6087 => x"dc",
          6088 => x"f0",
          6089 => x"fe",
          6090 => x"72",
          6091 => x"81",
          6092 => x"71",
          6093 => x"38",
          6094 => x"d8",
          6095 => x"82",
          6096 => x"da",
          6097 => x"51",
          6098 => x"3f",
          6099 => x"70",
          6100 => x"52",
          6101 => x"95",
          6102 => x"fe",
          6103 => x"82",
          6104 => x"fe",
          6105 => x"80",
          6106 => x"a8",
          6107 => x"2a",
          6108 => x"51",
          6109 => x"2e",
          6110 => x"51",
          6111 => x"3f",
          6112 => x"51",
          6113 => x"3f",
          6114 => x"d8",
          6115 => x"86",
          6116 => x"06",
          6117 => x"80",
          6118 => x"81",
          6119 => x"f4",
          6120 => x"a8",
          6121 => x"ec",
          6122 => x"fe",
          6123 => x"72",
          6124 => x"81",
          6125 => x"71",
          6126 => x"38",
          6127 => x"d7",
          6128 => x"83",
          6129 => x"d9",
          6130 => x"51",
          6131 => x"3f",
          6132 => x"70",
          6133 => x"52",
          6134 => x"95",
          6135 => x"fe",
          6136 => x"82",
          6137 => x"fe",
          6138 => x"80",
          6139 => x"a4",
          6140 => x"99",
          6141 => x"0d",
          6142 => x"0d",
          6143 => x"05",
          6144 => x"70",
          6145 => x"80",
          6146 => x"fe",
          6147 => x"82",
          6148 => x"54",
          6149 => x"81",
          6150 => x"90",
          6151 => x"f4",
          6152 => x"83",
          6153 => x"dc",
          6154 => x"82",
          6155 => x"07",
          6156 => x"71",
          6157 => x"54",
          6158 => x"c8",
          6159 => x"c8",
          6160 => x"81",
          6161 => x"06",
          6162 => x"a3",
          6163 => x"52",
          6164 => x"b9",
          6165 => x"dc",
          6166 => x"8c",
          6167 => x"dc",
          6168 => x"e9",
          6169 => x"39",
          6170 => x"51",
          6171 => x"82",
          6172 => x"c8",
          6173 => x"c8",
          6174 => x"82",
          6175 => x"06",
          6176 => x"52",
          6177 => x"fa",
          6178 => x"0b",
          6179 => x"0c",
          6180 => x"04",
          6181 => x"80",
          6182 => x"a3",
          6183 => x"5d",
          6184 => x"51",
          6185 => x"3f",
          6186 => x"08",
          6187 => x"59",
          6188 => x"09",
          6189 => x"38",
          6190 => x"52",
          6191 => x"52",
          6192 => x"bf",
          6193 => x"78",
          6194 => x"a0",
          6195 => x"f6",
          6196 => x"dc",
          6197 => x"88",
          6198 => x"a4",
          6199 => x"39",
          6200 => x"5d",
          6201 => x"51",
          6202 => x"3f",
          6203 => x"46",
          6204 => x"52",
          6205 => x"81",
          6206 => x"ff",
          6207 => x"f3",
          6208 => x"8c",
          6209 => x"2b",
          6210 => x"51",
          6211 => x"c2",
          6212 => x"38",
          6213 => x"24",
          6214 => x"bd",
          6215 => x"38",
          6216 => x"90",
          6217 => x"2e",
          6218 => x"78",
          6219 => x"da",
          6220 => x"39",
          6221 => x"2e",
          6222 => x"78",
          6223 => x"85",
          6224 => x"bf",
          6225 => x"38",
          6226 => x"78",
          6227 => x"89",
          6228 => x"80",
          6229 => x"38",
          6230 => x"2e",
          6231 => x"78",
          6232 => x"89",
          6233 => x"b4",
          6234 => x"83",
          6235 => x"38",
          6236 => x"24",
          6237 => x"81",
          6238 => x"fd",
          6239 => x"39",
          6240 => x"2e",
          6241 => x"8a",
          6242 => x"3d",
          6243 => x"53",
          6244 => x"51",
          6245 => x"3f",
          6246 => x"08",
          6247 => x"c4",
          6248 => x"fe",
          6249 => x"ff",
          6250 => x"fe",
          6251 => x"82",
          6252 => x"80",
          6253 => x"38",
          6254 => x"f8",
          6255 => x"84",
          6256 => x"ee",
          6257 => x"8c",
          6258 => x"38",
          6259 => x"08",
          6260 => x"e0",
          6261 => x"b1",
          6262 => x"5c",
          6263 => x"27",
          6264 => x"61",
          6265 => x"70",
          6266 => x"0c",
          6267 => x"f5",
          6268 => x"39",
          6269 => x"80",
          6270 => x"84",
          6271 => x"ed",
          6272 => x"8c",
          6273 => x"2e",
          6274 => x"b4",
          6275 => x"11",
          6276 => x"05",
          6277 => x"ca",
          6278 => x"dc",
          6279 => x"fd",
          6280 => x"3d",
          6281 => x"53",
          6282 => x"51",
          6283 => x"3f",
          6284 => x"08",
          6285 => x"ac",
          6286 => x"f0",
          6287 => x"c9",
          6288 => x"79",
          6289 => x"8c",
          6290 => x"79",
          6291 => x"5b",
          6292 => x"61",
          6293 => x"eb",
          6294 => x"ff",
          6295 => x"ff",
          6296 => x"fe",
          6297 => x"82",
          6298 => x"80",
          6299 => x"38",
          6300 => x"fc",
          6301 => x"84",
          6302 => x"ec",
          6303 => x"8c",
          6304 => x"2e",
          6305 => x"b4",
          6306 => x"11",
          6307 => x"05",
          6308 => x"ce",
          6309 => x"dc",
          6310 => x"fc",
          6311 => x"84",
          6312 => x"e4",
          6313 => x"5a",
          6314 => x"a8",
          6315 => x"33",
          6316 => x"5a",
          6317 => x"2e",
          6318 => x"55",
          6319 => x"33",
          6320 => x"82",
          6321 => x"fe",
          6322 => x"81",
          6323 => x"05",
          6324 => x"39",
          6325 => x"51",
          6326 => x"b4",
          6327 => x"11",
          6328 => x"05",
          6329 => x"fa",
          6330 => x"dc",
          6331 => x"38",
          6332 => x"33",
          6333 => x"2e",
          6334 => x"87",
          6335 => x"80",
          6336 => x"88",
          6337 => x"78",
          6338 => x"38",
          6339 => x"08",
          6340 => x"82",
          6341 => x"59",
          6342 => x"88",
          6343 => x"e8",
          6344 => x"39",
          6345 => x"33",
          6346 => x"2e",
          6347 => x"87",
          6348 => x"9a",
          6349 => x"9e",
          6350 => x"80",
          6351 => x"82",
          6352 => x"44",
          6353 => x"88",
          6354 => x"80",
          6355 => x"3d",
          6356 => x"53",
          6357 => x"51",
          6358 => x"3f",
          6359 => x"08",
          6360 => x"82",
          6361 => x"59",
          6362 => x"89",
          6363 => x"dc",
          6364 => x"cc",
          6365 => x"a1",
          6366 => x"80",
          6367 => x"82",
          6368 => x"43",
          6369 => x"88",
          6370 => x"78",
          6371 => x"38",
          6372 => x"08",
          6373 => x"82",
          6374 => x"59",
          6375 => x"88",
          6376 => x"f4",
          6377 => x"39",
          6378 => x"33",
          6379 => x"2e",
          6380 => x"87",
          6381 => x"88",
          6382 => x"88",
          6383 => x"43",
          6384 => x"f8",
          6385 => x"84",
          6386 => x"ea",
          6387 => x"8c",
          6388 => x"2e",
          6389 => x"62",
          6390 => x"88",
          6391 => x"81",
          6392 => x"32",
          6393 => x"72",
          6394 => x"70",
          6395 => x"51",
          6396 => x"80",
          6397 => x"7a",
          6398 => x"38",
          6399 => x"85",
          6400 => x"e2",
          6401 => x"55",
          6402 => x"53",
          6403 => x"51",
          6404 => x"82",
          6405 => x"fe",
          6406 => x"f9",
          6407 => x"3d",
          6408 => x"53",
          6409 => x"51",
          6410 => x"3f",
          6411 => x"08",
          6412 => x"b0",
          6413 => x"fe",
          6414 => x"ff",
          6415 => x"fe",
          6416 => x"82",
          6417 => x"80",
          6418 => x"63",
          6419 => x"cb",
          6420 => x"34",
          6421 => x"44",
          6422 => x"fc",
          6423 => x"84",
          6424 => x"e8",
          6425 => x"8c",
          6426 => x"38",
          6427 => x"63",
          6428 => x"52",
          6429 => x"51",
          6430 => x"3f",
          6431 => x"79",
          6432 => x"c3",
          6433 => x"79",
          6434 => x"ae",
          6435 => x"38",
          6436 => x"a0",
          6437 => x"fe",
          6438 => x"ff",
          6439 => x"fe",
          6440 => x"82",
          6441 => x"80",
          6442 => x"63",
          6443 => x"cb",
          6444 => x"34",
          6445 => x"44",
          6446 => x"82",
          6447 => x"fe",
          6448 => x"ff",
          6449 => x"3d",
          6450 => x"53",
          6451 => x"51",
          6452 => x"3f",
          6453 => x"08",
          6454 => x"88",
          6455 => x"fe",
          6456 => x"ff",
          6457 => x"fe",
          6458 => x"82",
          6459 => x"80",
          6460 => x"60",
          6461 => x"05",
          6462 => x"82",
          6463 => x"78",
          6464 => x"fe",
          6465 => x"ff",
          6466 => x"fe",
          6467 => x"82",
          6468 => x"df",
          6469 => x"39",
          6470 => x"54",
          6471 => x"d8",
          6472 => x"c9",
          6473 => x"52",
          6474 => x"e6",
          6475 => x"45",
          6476 => x"78",
          6477 => x"ac",
          6478 => x"26",
          6479 => x"82",
          6480 => x"39",
          6481 => x"f0",
          6482 => x"84",
          6483 => x"e9",
          6484 => x"8c",
          6485 => x"2e",
          6486 => x"59",
          6487 => x"22",
          6488 => x"05",
          6489 => x"41",
          6490 => x"82",
          6491 => x"fe",
          6492 => x"ff",
          6493 => x"3d",
          6494 => x"53",
          6495 => x"51",
          6496 => x"3f",
          6497 => x"08",
          6498 => x"d8",
          6499 => x"fe",
          6500 => x"ff",
          6501 => x"fe",
          6502 => x"82",
          6503 => x"80",
          6504 => x"60",
          6505 => x"59",
          6506 => x"41",
          6507 => x"f0",
          6508 => x"84",
          6509 => x"e8",
          6510 => x"8c",
          6511 => x"38",
          6512 => x"60",
          6513 => x"52",
          6514 => x"51",
          6515 => x"3f",
          6516 => x"79",
          6517 => x"ef",
          6518 => x"79",
          6519 => x"ae",
          6520 => x"38",
          6521 => x"9c",
          6522 => x"fe",
          6523 => x"ff",
          6524 => x"fe",
          6525 => x"82",
          6526 => x"80",
          6527 => x"60",
          6528 => x"59",
          6529 => x"41",
          6530 => x"82",
          6531 => x"fe",
          6532 => x"ff",
          6533 => x"3d",
          6534 => x"53",
          6535 => x"51",
          6536 => x"3f",
          6537 => x"08",
          6538 => x"b8",
          6539 => x"82",
          6540 => x"fe",
          6541 => x"63",
          6542 => x"b4",
          6543 => x"11",
          6544 => x"05",
          6545 => x"9a",
          6546 => x"dc",
          6547 => x"f5",
          6548 => x"52",
          6549 => x"51",
          6550 => x"3f",
          6551 => x"2d",
          6552 => x"08",
          6553 => x"fc",
          6554 => x"dc",
          6555 => x"86",
          6556 => x"e2",
          6557 => x"ec",
          6558 => x"c4",
          6559 => x"89",
          6560 => x"b9",
          6561 => x"39",
          6562 => x"51",
          6563 => x"3f",
          6564 => x"a5",
          6565 => x"8c",
          6566 => x"39",
          6567 => x"33",
          6568 => x"2e",
          6569 => x"7d",
          6570 => x"78",
          6571 => x"d3",
          6572 => x"ff",
          6573 => x"fe",
          6574 => x"82",
          6575 => x"5c",
          6576 => x"82",
          6577 => x"7a",
          6578 => x"38",
          6579 => x"8c",
          6580 => x"39",
          6581 => x"b0",
          6582 => x"39",
          6583 => x"56",
          6584 => x"86",
          6585 => x"53",
          6586 => x"52",
          6587 => x"b0",
          6588 => x"e2",
          6589 => x"39",
          6590 => x"52",
          6591 => x"b0",
          6592 => x"e1",
          6593 => x"39",
          6594 => x"86",
          6595 => x"53",
          6596 => x"52",
          6597 => x"b0",
          6598 => x"e1",
          6599 => x"39",
          6600 => x"53",
          6601 => x"52",
          6602 => x"b0",
          6603 => x"e1",
          6604 => x"87",
          6605 => x"8d",
          6606 => x"56",
          6607 => x"54",
          6608 => x"53",
          6609 => x"52",
          6610 => x"b0",
          6611 => x"8a",
          6612 => x"dc",
          6613 => x"dc",
          6614 => x"30",
          6615 => x"80",
          6616 => x"5b",
          6617 => x"7a",
          6618 => x"38",
          6619 => x"7a",
          6620 => x"80",
          6621 => x"81",
          6622 => x"ff",
          6623 => x"7a",
          6624 => x"7d",
          6625 => x"81",
          6626 => x"78",
          6627 => x"ff",
          6628 => x"06",
          6629 => x"82",
          6630 => x"fe",
          6631 => x"f2",
          6632 => x"3d",
          6633 => x"82",
          6634 => x"87",
          6635 => x"70",
          6636 => x"87",
          6637 => x"72",
          6638 => x"a1",
          6639 => x"dc",
          6640 => x"75",
          6641 => x"87",
          6642 => x"73",
          6643 => x"8d",
          6644 => x"8c",
          6645 => x"75",
          6646 => x"94",
          6647 => x"54",
          6648 => x"80",
          6649 => x"fe",
          6650 => x"82",
          6651 => x"90",
          6652 => x"55",
          6653 => x"80",
          6654 => x"fe",
          6655 => x"72",
          6656 => x"08",
          6657 => x"8c",
          6658 => x"87",
          6659 => x"0c",
          6660 => x"0b",
          6661 => x"94",
          6662 => x"0b",
          6663 => x"0c",
          6664 => x"82",
          6665 => x"fe",
          6666 => x"fe",
          6667 => x"82",
          6668 => x"fe",
          6669 => x"82",
          6670 => x"fe",
          6671 => x"81",
          6672 => x"fe",
          6673 => x"81",
          6674 => x"3f",
          6675 => x"80",
          6676 => x"00",
          6677 => x"00",
          6678 => x"00",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"00",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"00",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"00",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"00",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"00",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"00",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"00",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"00",
          6711 => x"00",
          6712 => x"00",
          6713 => x"64",
          6714 => x"2f",
          6715 => x"25",
          6716 => x"64",
          6717 => x"2e",
          6718 => x"64",
          6719 => x"6f",
          6720 => x"6f",
          6721 => x"67",
          6722 => x"74",
          6723 => x"00",
          6724 => x"28",
          6725 => x"6d",
          6726 => x"43",
          6727 => x"6e",
          6728 => x"29",
          6729 => x"0a",
          6730 => x"69",
          6731 => x"20",
          6732 => x"6c",
          6733 => x"6e",
          6734 => x"3a",
          6735 => x"20",
          6736 => x"42",
          6737 => x"52",
          6738 => x"20",
          6739 => x"38",
          6740 => x"30",
          6741 => x"2e",
          6742 => x"20",
          6743 => x"44",
          6744 => x"20",
          6745 => x"20",
          6746 => x"38",
          6747 => x"30",
          6748 => x"2e",
          6749 => x"20",
          6750 => x"4e",
          6751 => x"42",
          6752 => x"20",
          6753 => x"38",
          6754 => x"30",
          6755 => x"2e",
          6756 => x"20",
          6757 => x"52",
          6758 => x"20",
          6759 => x"20",
          6760 => x"38",
          6761 => x"30",
          6762 => x"2e",
          6763 => x"20",
          6764 => x"41",
          6765 => x"20",
          6766 => x"20",
          6767 => x"38",
          6768 => x"30",
          6769 => x"2e",
          6770 => x"20",
          6771 => x"44",
          6772 => x"52",
          6773 => x"20",
          6774 => x"76",
          6775 => x"73",
          6776 => x"30",
          6777 => x"2e",
          6778 => x"20",
          6779 => x"49",
          6780 => x"31",
          6781 => x"20",
          6782 => x"6d",
          6783 => x"20",
          6784 => x"30",
          6785 => x"2e",
          6786 => x"20",
          6787 => x"4e",
          6788 => x"43",
          6789 => x"20",
          6790 => x"61",
          6791 => x"6c",
          6792 => x"30",
          6793 => x"2e",
          6794 => x"20",
          6795 => x"49",
          6796 => x"4f",
          6797 => x"42",
          6798 => x"00",
          6799 => x"20",
          6800 => x"42",
          6801 => x"43",
          6802 => x"20",
          6803 => x"4f",
          6804 => x"0a",
          6805 => x"20",
          6806 => x"53",
          6807 => x"00",
          6808 => x"20",
          6809 => x"50",
          6810 => x"00",
          6811 => x"64",
          6812 => x"73",
          6813 => x"3a",
          6814 => x"20",
          6815 => x"50",
          6816 => x"65",
          6817 => x"20",
          6818 => x"74",
          6819 => x"41",
          6820 => x"65",
          6821 => x"3d",
          6822 => x"38",
          6823 => x"00",
          6824 => x"20",
          6825 => x"50",
          6826 => x"65",
          6827 => x"79",
          6828 => x"61",
          6829 => x"41",
          6830 => x"65",
          6831 => x"3d",
          6832 => x"38",
          6833 => x"00",
          6834 => x"20",
          6835 => x"74",
          6836 => x"20",
          6837 => x"72",
          6838 => x"64",
          6839 => x"73",
          6840 => x"20",
          6841 => x"3d",
          6842 => x"38",
          6843 => x"00",
          6844 => x"69",
          6845 => x"0a",
          6846 => x"20",
          6847 => x"50",
          6848 => x"64",
          6849 => x"20",
          6850 => x"20",
          6851 => x"20",
          6852 => x"20",
          6853 => x"3d",
          6854 => x"34",
          6855 => x"00",
          6856 => x"20",
          6857 => x"79",
          6858 => x"6d",
          6859 => x"6f",
          6860 => x"46",
          6861 => x"20",
          6862 => x"20",
          6863 => x"3d",
          6864 => x"2e",
          6865 => x"64",
          6866 => x"0a",
          6867 => x"20",
          6868 => x"44",
          6869 => x"20",
          6870 => x"63",
          6871 => x"72",
          6872 => x"20",
          6873 => x"20",
          6874 => x"3d",
          6875 => x"2e",
          6876 => x"64",
          6877 => x"0a",
          6878 => x"20",
          6879 => x"69",
          6880 => x"6f",
          6881 => x"53",
          6882 => x"4d",
          6883 => x"6f",
          6884 => x"46",
          6885 => x"3d",
          6886 => x"2e",
          6887 => x"64",
          6888 => x"0a",
          6889 => x"6d",
          6890 => x"00",
          6891 => x"65",
          6892 => x"6d",
          6893 => x"6c",
          6894 => x"00",
          6895 => x"56",
          6896 => x"56",
          6897 => x"6e",
          6898 => x"6e",
          6899 => x"77",
          6900 => x"69",
          6901 => x"72",
          6902 => x"78",
          6903 => x"69",
          6904 => x"72",
          6905 => x"69",
          6906 => x"00",
          6907 => x"00",
          6908 => x"30",
          6909 => x"20",
          6910 => x"00",
          6911 => x"61",
          6912 => x"64",
          6913 => x"20",
          6914 => x"65",
          6915 => x"68",
          6916 => x"69",
          6917 => x"72",
          6918 => x"69",
          6919 => x"74",
          6920 => x"4f",
          6921 => x"00",
          6922 => x"61",
          6923 => x"74",
          6924 => x"65",
          6925 => x"72",
          6926 => x"65",
          6927 => x"73",
          6928 => x"79",
          6929 => x"6c",
          6930 => x"64",
          6931 => x"62",
          6932 => x"67",
          6933 => x"00",
          6934 => x"00",
          6935 => x"00",
          6936 => x"00",
          6937 => x"00",
          6938 => x"00",
          6939 => x"00",
          6940 => x"00",
          6941 => x"00",
          6942 => x"00",
          6943 => x"00",
          6944 => x"00",
          6945 => x"00",
          6946 => x"00",
          6947 => x"00",
          6948 => x"00",
          6949 => x"00",
          6950 => x"00",
          6951 => x"00",
          6952 => x"00",
          6953 => x"00",
          6954 => x"00",
          6955 => x"00",
          6956 => x"00",
          6957 => x"00",
          6958 => x"00",
          6959 => x"00",
          6960 => x"00",
          6961 => x"00",
          6962 => x"00",
          6963 => x"00",
          6964 => x"00",
          6965 => x"00",
          6966 => x"00",
          6967 => x"5b",
          6968 => x"5b",
          6969 => x"5b",
          6970 => x"5b",
          6971 => x"5b",
          6972 => x"5b",
          6973 => x"5b",
          6974 => x"5b",
          6975 => x"5b",
          6976 => x"00",
          6977 => x"00",
          6978 => x"44",
          6979 => x"2a",
          6980 => x"3b",
          6981 => x"3f",
          6982 => x"7f",
          6983 => x"41",
          6984 => x"41",
          6985 => x"00",
          6986 => x"fe",
          6987 => x"44",
          6988 => x"2e",
          6989 => x"4f",
          6990 => x"4d",
          6991 => x"20",
          6992 => x"54",
          6993 => x"20",
          6994 => x"4f",
          6995 => x"4d",
          6996 => x"20",
          6997 => x"54",
          6998 => x"20",
          6999 => x"00",
          7000 => x"00",
          7001 => x"00",
          7002 => x"00",
          7003 => x"9a",
          7004 => x"41",
          7005 => x"45",
          7006 => x"49",
          7007 => x"92",
          7008 => x"4f",
          7009 => x"99",
          7010 => x"9d",
          7011 => x"49",
          7012 => x"a5",
          7013 => x"a9",
          7014 => x"ad",
          7015 => x"b1",
          7016 => x"b5",
          7017 => x"b9",
          7018 => x"bd",
          7019 => x"c1",
          7020 => x"c5",
          7021 => x"c9",
          7022 => x"cd",
          7023 => x"d1",
          7024 => x"d5",
          7025 => x"d9",
          7026 => x"dd",
          7027 => x"e1",
          7028 => x"e5",
          7029 => x"e9",
          7030 => x"ed",
          7031 => x"f1",
          7032 => x"f5",
          7033 => x"f9",
          7034 => x"fd",
          7035 => x"2e",
          7036 => x"5b",
          7037 => x"22",
          7038 => x"3e",
          7039 => x"00",
          7040 => x"01",
          7041 => x"10",
          7042 => x"00",
          7043 => x"00",
          7044 => x"01",
          7045 => x"04",
          7046 => x"10",
          7047 => x"00",
          7048 => x"69",
          7049 => x"00",
          7050 => x"69",
          7051 => x"6c",
          7052 => x"69",
          7053 => x"00",
          7054 => x"6c",
          7055 => x"00",
          7056 => x"65",
          7057 => x"00",
          7058 => x"63",
          7059 => x"72",
          7060 => x"63",
          7061 => x"00",
          7062 => x"64",
          7063 => x"00",
          7064 => x"64",
          7065 => x"00",
          7066 => x"65",
          7067 => x"65",
          7068 => x"65",
          7069 => x"69",
          7070 => x"69",
          7071 => x"66",
          7072 => x"66",
          7073 => x"61",
          7074 => x"00",
          7075 => x"6d",
          7076 => x"65",
          7077 => x"72",
          7078 => x"65",
          7079 => x"00",
          7080 => x"6e",
          7081 => x"00",
          7082 => x"65",
          7083 => x"00",
          7084 => x"62",
          7085 => x"63",
          7086 => x"62",
          7087 => x"63",
          7088 => x"69",
          7089 => x"00",
          7090 => x"69",
          7091 => x"45",
          7092 => x"72",
          7093 => x"6e",
          7094 => x"6e",
          7095 => x"65",
          7096 => x"72",
          7097 => x"00",
          7098 => x"69",
          7099 => x"6e",
          7100 => x"72",
          7101 => x"79",
          7102 => x"00",
          7103 => x"6f",
          7104 => x"6c",
          7105 => x"6f",
          7106 => x"2e",
          7107 => x"6f",
          7108 => x"74",
          7109 => x"6f",
          7110 => x"2e",
          7111 => x"6e",
          7112 => x"69",
          7113 => x"69",
          7114 => x"61",
          7115 => x"0a",
          7116 => x"63",
          7117 => x"73",
          7118 => x"6e",
          7119 => x"2e",
          7120 => x"69",
          7121 => x"61",
          7122 => x"61",
          7123 => x"65",
          7124 => x"74",
          7125 => x"00",
          7126 => x"69",
          7127 => x"68",
          7128 => x"6c",
          7129 => x"6e",
          7130 => x"69",
          7131 => x"00",
          7132 => x"44",
          7133 => x"20",
          7134 => x"74",
          7135 => x"72",
          7136 => x"63",
          7137 => x"2e",
          7138 => x"72",
          7139 => x"20",
          7140 => x"62",
          7141 => x"69",
          7142 => x"6e",
          7143 => x"69",
          7144 => x"00",
          7145 => x"69",
          7146 => x"6e",
          7147 => x"65",
          7148 => x"6c",
          7149 => x"0a",
          7150 => x"6f",
          7151 => x"6d",
          7152 => x"69",
          7153 => x"20",
          7154 => x"65",
          7155 => x"74",
          7156 => x"66",
          7157 => x"64",
          7158 => x"20",
          7159 => x"6b",
          7160 => x"00",
          7161 => x"6f",
          7162 => x"74",
          7163 => x"6f",
          7164 => x"64",
          7165 => x"00",
          7166 => x"69",
          7167 => x"75",
          7168 => x"6f",
          7169 => x"61",
          7170 => x"6e",
          7171 => x"6e",
          7172 => x"6c",
          7173 => x"0a",
          7174 => x"69",
          7175 => x"69",
          7176 => x"6f",
          7177 => x"64",
          7178 => x"00",
          7179 => x"6e",
          7180 => x"66",
          7181 => x"65",
          7182 => x"6d",
          7183 => x"72",
          7184 => x"00",
          7185 => x"6f",
          7186 => x"61",
          7187 => x"6f",
          7188 => x"20",
          7189 => x"65",
          7190 => x"00",
          7191 => x"61",
          7192 => x"65",
          7193 => x"73",
          7194 => x"63",
          7195 => x"65",
          7196 => x"0a",
          7197 => x"75",
          7198 => x"73",
          7199 => x"00",
          7200 => x"6e",
          7201 => x"77",
          7202 => x"72",
          7203 => x"2e",
          7204 => x"25",
          7205 => x"62",
          7206 => x"73",
          7207 => x"20",
          7208 => x"25",
          7209 => x"62",
          7210 => x"73",
          7211 => x"63",
          7212 => x"00",
          7213 => x"65",
          7214 => x"00",
          7215 => x"30",
          7216 => x"00",
          7217 => x"20",
          7218 => x"30",
          7219 => x"00",
          7220 => x"20",
          7221 => x"20",
          7222 => x"00",
          7223 => x"30",
          7224 => x"00",
          7225 => x"20",
          7226 => x"7c",
          7227 => x"0d",
          7228 => x"4f",
          7229 => x"2a",
          7230 => x"73",
          7231 => x"00",
          7232 => x"37",
          7233 => x"2f",
          7234 => x"30",
          7235 => x"31",
          7236 => x"00",
          7237 => x"5a",
          7238 => x"20",
          7239 => x"20",
          7240 => x"78",
          7241 => x"73",
          7242 => x"20",
          7243 => x"0a",
          7244 => x"50",
          7245 => x"6e",
          7246 => x"72",
          7247 => x"20",
          7248 => x"64",
          7249 => x"0a",
          7250 => x"69",
          7251 => x"20",
          7252 => x"65",
          7253 => x"70",
          7254 => x"00",
          7255 => x"53",
          7256 => x"6e",
          7257 => x"72",
          7258 => x"0a",
          7259 => x"4f",
          7260 => x"20",
          7261 => x"69",
          7262 => x"72",
          7263 => x"74",
          7264 => x"4f",
          7265 => x"20",
          7266 => x"69",
          7267 => x"72",
          7268 => x"74",
          7269 => x"41",
          7270 => x"20",
          7271 => x"69",
          7272 => x"72",
          7273 => x"74",
          7274 => x"41",
          7275 => x"20",
          7276 => x"69",
          7277 => x"72",
          7278 => x"74",
          7279 => x"41",
          7280 => x"20",
          7281 => x"69",
          7282 => x"72",
          7283 => x"74",
          7284 => x"41",
          7285 => x"20",
          7286 => x"69",
          7287 => x"72",
          7288 => x"74",
          7289 => x"65",
          7290 => x"6e",
          7291 => x"70",
          7292 => x"6d",
          7293 => x"2e",
          7294 => x"00",
          7295 => x"6e",
          7296 => x"69",
          7297 => x"74",
          7298 => x"72",
          7299 => x"0a",
          7300 => x"75",
          7301 => x"78",
          7302 => x"62",
          7303 => x"00",
          7304 => x"3a",
          7305 => x"61",
          7306 => x"64",
          7307 => x"20",
          7308 => x"74",
          7309 => x"69",
          7310 => x"73",
          7311 => x"61",
          7312 => x"30",
          7313 => x"6c",
          7314 => x"65",
          7315 => x"69",
          7316 => x"61",
          7317 => x"6c",
          7318 => x"0a",
          7319 => x"20",
          7320 => x"6c",
          7321 => x"69",
          7322 => x"2e",
          7323 => x"00",
          7324 => x"6f",
          7325 => x"6e",
          7326 => x"2e",
          7327 => x"6f",
          7328 => x"72",
          7329 => x"2e",
          7330 => x"00",
          7331 => x"30",
          7332 => x"28",
          7333 => x"78",
          7334 => x"25",
          7335 => x"78",
          7336 => x"38",
          7337 => x"00",
          7338 => x"75",
          7339 => x"4d",
          7340 => x"72",
          7341 => x"00",
          7342 => x"43",
          7343 => x"6c",
          7344 => x"2e",
          7345 => x"30",
          7346 => x"25",
          7347 => x"2d",
          7348 => x"3f",
          7349 => x"00",
          7350 => x"30",
          7351 => x"25",
          7352 => x"2d",
          7353 => x"30",
          7354 => x"25",
          7355 => x"2d",
          7356 => x"78",
          7357 => x"74",
          7358 => x"20",
          7359 => x"65",
          7360 => x"25",
          7361 => x"20",
          7362 => x"0a",
          7363 => x"61",
          7364 => x"6e",
          7365 => x"6f",
          7366 => x"40",
          7367 => x"38",
          7368 => x"2e",
          7369 => x"00",
          7370 => x"61",
          7371 => x"72",
          7372 => x"72",
          7373 => x"20",
          7374 => x"65",
          7375 => x"64",
          7376 => x"00",
          7377 => x"65",
          7378 => x"72",
          7379 => x"67",
          7380 => x"70",
          7381 => x"61",
          7382 => x"6e",
          7383 => x"0a",
          7384 => x"6f",
          7385 => x"72",
          7386 => x"6f",
          7387 => x"67",
          7388 => x"0a",
          7389 => x"50",
          7390 => x"69",
          7391 => x"64",
          7392 => x"73",
          7393 => x"2e",
          7394 => x"00",
          7395 => x"64",
          7396 => x"73",
          7397 => x"00",
          7398 => x"64",
          7399 => x"73",
          7400 => x"61",
          7401 => x"6f",
          7402 => x"6e",
          7403 => x"00",
          7404 => x"75",
          7405 => x"6e",
          7406 => x"2e",
          7407 => x"6e",
          7408 => x"69",
          7409 => x"69",
          7410 => x"72",
          7411 => x"74",
          7412 => x"2e",
          7413 => x"00",
          7414 => x"00",
          7415 => x"00",
          7416 => x"00",
          7417 => x"00",
          7418 => x"01",
          7419 => x"00",
          7420 => x"01",
          7421 => x"81",
          7422 => x"00",
          7423 => x"7f",
          7424 => x"00",
          7425 => x"00",
          7426 => x"00",
          7427 => x"00",
          7428 => x"f5",
          7429 => x"f5",
          7430 => x"f5",
          7431 => x"00",
          7432 => x"01",
          7433 => x"01",
          7434 => x"01",
          7435 => x"00",
          7436 => x"00",
          7437 => x"00",
          7438 => x"00",
          7439 => x"00",
          7440 => x"00",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"00",
          7469 => x"00",
          7470 => x"00",
          7471 => x"00",
          7472 => x"00",
          7473 => x"00",
          7474 => x"00",
          7475 => x"00",
          7476 => x"02",
          7477 => x"00",
          7478 => x"00",
          7479 => x"00",
          7480 => x"04",
          7481 => x"00",
          7482 => x"00",
          7483 => x"00",
          7484 => x"14",
          7485 => x"00",
          7486 => x"00",
          7487 => x"00",
          7488 => x"2b",
          7489 => x"00",
          7490 => x"00",
          7491 => x"00",
          7492 => x"30",
          7493 => x"00",
          7494 => x"00",
          7495 => x"00",
          7496 => x"3c",
          7497 => x"00",
          7498 => x"00",
          7499 => x"00",
          7500 => x"3d",
          7501 => x"00",
          7502 => x"00",
          7503 => x"00",
          7504 => x"3f",
          7505 => x"00",
          7506 => x"00",
          7507 => x"00",
          7508 => x"40",
          7509 => x"00",
          7510 => x"00",
          7511 => x"00",
          7512 => x"41",
          7513 => x"00",
          7514 => x"00",
          7515 => x"00",
          7516 => x"42",
          7517 => x"00",
          7518 => x"00",
          7519 => x"00",
          7520 => x"43",
          7521 => x"00",
          7522 => x"00",
          7523 => x"00",
          7524 => x"50",
          7525 => x"00",
          7526 => x"00",
          7527 => x"00",
          7528 => x"51",
          7529 => x"00",
          7530 => x"00",
          7531 => x"00",
          7532 => x"54",
          7533 => x"00",
          7534 => x"00",
          7535 => x"00",
          7536 => x"55",
          7537 => x"00",
          7538 => x"00",
          7539 => x"00",
          7540 => x"79",
          7541 => x"00",
          7542 => x"00",
          7543 => x"00",
          7544 => x"78",
          7545 => x"00",
          7546 => x"00",
          7547 => x"00",
          7548 => x"82",
          7549 => x"00",
          7550 => x"00",
          7551 => x"00",
          7552 => x"83",
          7553 => x"00",
          7554 => x"00",
          7555 => x"00",
          7556 => x"85",
          7557 => x"00",
          7558 => x"00",
          7559 => x"00",
          7560 => x"87",
          7561 => x"00",
          7562 => x"00",
          7563 => x"00",
          7564 => x"8c",
          7565 => x"00",
          7566 => x"00",
          7567 => x"00",
          7568 => x"8d",
          7569 => x"00",
          7570 => x"00",
          7571 => x"00",
          7572 => x"8e",
          7573 => x"00",
          7574 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"0b",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"0b",
            11 => x"0b",
            12 => x"93",
            13 => x"0b",
            14 => x"0b",
            15 => x"b3",
            16 => x"0b",
            17 => x"0b",
            18 => x"d3",
            19 => x"0b",
            20 => x"0b",
            21 => x"f3",
            22 => x"0b",
            23 => x"0b",
            24 => x"93",
            25 => x"0b",
            26 => x"0b",
            27 => x"b3",
            28 => x"0b",
            29 => x"0b",
            30 => x"d3",
            31 => x"0b",
            32 => x"0b",
            33 => x"f1",
            34 => x"0b",
            35 => x"0b",
            36 => x"8f",
            37 => x"0b",
            38 => x"0b",
            39 => x"ae",
            40 => x"0b",
            41 => x"0b",
            42 => x"ce",
            43 => x"0b",
            44 => x"0b",
            45 => x"ee",
            46 => x"0b",
            47 => x"0b",
            48 => x"8e",
            49 => x"0b",
            50 => x"0b",
            51 => x"ae",
            52 => x"0b",
            53 => x"0b",
            54 => x"ce",
            55 => x"0b",
            56 => x"0b",
            57 => x"ee",
            58 => x"0b",
            59 => x"0b",
            60 => x"8e",
            61 => x"0b",
            62 => x"0b",
            63 => x"ae",
            64 => x"0b",
            65 => x"0b",
            66 => x"ce",
            67 => x"0b",
            68 => x"0b",
            69 => x"ee",
            70 => x"0b",
            71 => x"0b",
            72 => x"8e",
            73 => x"0b",
            74 => x"0b",
            75 => x"ae",
            76 => x"0b",
            77 => x"0b",
            78 => x"ce",
            79 => x"0b",
            80 => x"0b",
            81 => x"ee",
            82 => x"0b",
            83 => x"0b",
            84 => x"8d",
            85 => x"0b",
            86 => x"0b",
            87 => x"ab",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"82",
           130 => x"b8",
           131 => x"8c",
           132 => x"80",
           133 => x"8c",
           134 => x"c9",
           135 => x"8c",
           136 => x"80",
           137 => x"8c",
           138 => x"c9",
           139 => x"8c",
           140 => x"80",
           141 => x"8c",
           142 => x"ca",
           143 => x"8c",
           144 => x"80",
           145 => x"8c",
           146 => x"d0",
           147 => x"8c",
           148 => x"80",
           149 => x"8c",
           150 => x"d1",
           151 => x"8c",
           152 => x"80",
           153 => x"8c",
           154 => x"ca",
           155 => x"8c",
           156 => x"80",
           157 => x"8c",
           158 => x"d1",
           159 => x"8c",
           160 => x"80",
           161 => x"8c",
           162 => x"d3",
           163 => x"8c",
           164 => x"80",
           165 => x"8c",
           166 => x"cf",
           167 => x"8c",
           168 => x"80",
           169 => x"8c",
           170 => x"ca",
           171 => x"8c",
           172 => x"80",
           173 => x"8c",
           174 => x"d0",
           175 => x"8c",
           176 => x"80",
           177 => x"8c",
           178 => x"d0",
           179 => x"8c",
           180 => x"80",
           181 => x"8c",
           182 => x"ad",
           183 => x"e8",
           184 => x"90",
           185 => x"e8",
           186 => x"2d",
           187 => x"08",
           188 => x"04",
           189 => x"0c",
           190 => x"82",
           191 => x"83",
           192 => x"82",
           193 => x"b4",
           194 => x"8c",
           195 => x"80",
           196 => x"8c",
           197 => x"82",
           198 => x"e8",
           199 => x"90",
           200 => x"e8",
           201 => x"a5",
           202 => x"e8",
           203 => x"90",
           204 => x"e8",
           205 => x"96",
           206 => x"e8",
           207 => x"90",
           208 => x"e8",
           209 => x"8a",
           210 => x"e8",
           211 => x"90",
           212 => x"e8",
           213 => x"87",
           214 => x"e8",
           215 => x"90",
           216 => x"e8",
           217 => x"a5",
           218 => x"e8",
           219 => x"90",
           220 => x"e8",
           221 => x"85",
           222 => x"e8",
           223 => x"90",
           224 => x"e8",
           225 => x"f8",
           226 => x"e8",
           227 => x"90",
           228 => x"e8",
           229 => x"c4",
           230 => x"e8",
           231 => x"90",
           232 => x"e8",
           233 => x"e3",
           234 => x"e8",
           235 => x"90",
           236 => x"e8",
           237 => x"82",
           238 => x"e8",
           239 => x"90",
           240 => x"e8",
           241 => x"ec",
           242 => x"e8",
           243 => x"90",
           244 => x"e8",
           245 => x"d2",
           246 => x"e8",
           247 => x"90",
           248 => x"e8",
           249 => x"c0",
           250 => x"e8",
           251 => x"90",
           252 => x"e8",
           253 => x"86",
           254 => x"e8",
           255 => x"90",
           256 => x"e8",
           257 => x"c0",
           258 => x"e8",
           259 => x"90",
           260 => x"e8",
           261 => x"c1",
           262 => x"e8",
           263 => x"90",
           264 => x"e8",
           265 => x"f6",
           266 => x"e8",
           267 => x"90",
           268 => x"e8",
           269 => x"cf",
           270 => x"e8",
           271 => x"90",
           272 => x"e8",
           273 => x"fa",
           274 => x"e8",
           275 => x"90",
           276 => x"e8",
           277 => x"dd",
           278 => x"e8",
           279 => x"90",
           280 => x"e8",
           281 => x"b2",
           282 => x"e8",
           283 => x"90",
           284 => x"e8",
           285 => x"bc",
           286 => x"e8",
           287 => x"90",
           288 => x"e8",
           289 => x"fe",
           290 => x"e8",
           291 => x"90",
           292 => x"e8",
           293 => x"c4",
           294 => x"e8",
           295 => x"90",
           296 => x"e8",
           297 => x"ea",
           298 => x"e8",
           299 => x"90",
           300 => x"e8",
           301 => x"9f",
           302 => x"e8",
           303 => x"90",
           304 => x"e8",
           305 => x"8b",
           306 => x"e8",
           307 => x"90",
           308 => x"e8",
           309 => x"ff",
           310 => x"e8",
           311 => x"90",
           312 => x"e8",
           313 => x"e9",
           314 => x"e8",
           315 => x"90",
           316 => x"e8",
           317 => x"cd",
           318 => x"e8",
           319 => x"90",
           320 => x"e8",
           321 => x"2d",
           322 => x"08",
           323 => x"04",
           324 => x"0c",
           325 => x"82",
           326 => x"83",
           327 => x"82",
           328 => x"b7",
           329 => x"8c",
           330 => x"80",
           331 => x"8c",
           332 => x"d6",
           333 => x"8c",
           334 => x"80",
           335 => x"8c",
           336 => x"a4",
           337 => x"38",
           338 => x"84",
           339 => x"0b",
           340 => x"be",
           341 => x"51",
           342 => x"04",
           343 => x"8c",
           344 => x"82",
           345 => x"fd",
           346 => x"53",
           347 => x"08",
           348 => x"52",
           349 => x"08",
           350 => x"51",
           351 => x"82",
           352 => x"70",
           353 => x"0c",
           354 => x"0d",
           355 => x"0c",
           356 => x"e8",
           357 => x"8c",
           358 => x"3d",
           359 => x"82",
           360 => x"8c",
           361 => x"82",
           362 => x"88",
           363 => x"93",
           364 => x"dc",
           365 => x"8c",
           366 => x"85",
           367 => x"8c",
           368 => x"82",
           369 => x"02",
           370 => x"0c",
           371 => x"81",
           372 => x"e8",
           373 => x"0c",
           374 => x"8c",
           375 => x"05",
           376 => x"e8",
           377 => x"08",
           378 => x"08",
           379 => x"27",
           380 => x"8c",
           381 => x"05",
           382 => x"ae",
           383 => x"82",
           384 => x"8c",
           385 => x"a2",
           386 => x"e8",
           387 => x"08",
           388 => x"e8",
           389 => x"0c",
           390 => x"08",
           391 => x"10",
           392 => x"08",
           393 => x"ff",
           394 => x"8c",
           395 => x"05",
           396 => x"80",
           397 => x"8c",
           398 => x"05",
           399 => x"e8",
           400 => x"08",
           401 => x"82",
           402 => x"88",
           403 => x"8c",
           404 => x"05",
           405 => x"8c",
           406 => x"05",
           407 => x"e8",
           408 => x"08",
           409 => x"08",
           410 => x"07",
           411 => x"08",
           412 => x"82",
           413 => x"fc",
           414 => x"2a",
           415 => x"08",
           416 => x"82",
           417 => x"8c",
           418 => x"2a",
           419 => x"08",
           420 => x"ff",
           421 => x"8c",
           422 => x"05",
           423 => x"93",
           424 => x"e8",
           425 => x"08",
           426 => x"e8",
           427 => x"0c",
           428 => x"82",
           429 => x"f8",
           430 => x"82",
           431 => x"f4",
           432 => x"82",
           433 => x"f4",
           434 => x"8c",
           435 => x"3d",
           436 => x"e8",
           437 => x"3d",
           438 => x"79",
           439 => x"55",
           440 => x"27",
           441 => x"75",
           442 => x"51",
           443 => x"a9",
           444 => x"52",
           445 => x"98",
           446 => x"81",
           447 => x"74",
           448 => x"56",
           449 => x"52",
           450 => x"09",
           451 => x"38",
           452 => x"dc",
           453 => x"0d",
           454 => x"72",
           455 => x"54",
           456 => x"84",
           457 => x"72",
           458 => x"54",
           459 => x"84",
           460 => x"72",
           461 => x"54",
           462 => x"84",
           463 => x"72",
           464 => x"54",
           465 => x"84",
           466 => x"f0",
           467 => x"8f",
           468 => x"83",
           469 => x"38",
           470 => x"05",
           471 => x"70",
           472 => x"0c",
           473 => x"71",
           474 => x"38",
           475 => x"81",
           476 => x"0d",
           477 => x"02",
           478 => x"05",
           479 => x"53",
           480 => x"27",
           481 => x"83",
           482 => x"80",
           483 => x"ff",
           484 => x"ff",
           485 => x"73",
           486 => x"05",
           487 => x"12",
           488 => x"2e",
           489 => x"ef",
           490 => x"8c",
           491 => x"3d",
           492 => x"74",
           493 => x"07",
           494 => x"2b",
           495 => x"51",
           496 => x"a5",
           497 => x"70",
           498 => x"0c",
           499 => x"84",
           500 => x"72",
           501 => x"05",
           502 => x"71",
           503 => x"53",
           504 => x"52",
           505 => x"dd",
           506 => x"27",
           507 => x"71",
           508 => x"53",
           509 => x"52",
           510 => x"f2",
           511 => x"ff",
           512 => x"3d",
           513 => x"79",
           514 => x"83",
           515 => x"54",
           516 => x"c3",
           517 => x"08",
           518 => x"f7",
           519 => x"13",
           520 => x"84",
           521 => x"06",
           522 => x"53",
           523 => x"38",
           524 => x"74",
           525 => x"56",
           526 => x"70",
           527 => x"fb",
           528 => x"06",
           529 => x"82",
           530 => x"51",
           531 => x"54",
           532 => x"dc",
           533 => x"71",
           534 => x"53",
           535 => x"73",
           536 => x"55",
           537 => x"38",
           538 => x"dc",
           539 => x"0d",
           540 => x"0d",
           541 => x"83",
           542 => x"52",
           543 => x"71",
           544 => x"09",
           545 => x"ff",
           546 => x"f8",
           547 => x"80",
           548 => x"52",
           549 => x"38",
           550 => x"08",
           551 => x"fb",
           552 => x"06",
           553 => x"82",
           554 => x"51",
           555 => x"70",
           556 => x"38",
           557 => x"33",
           558 => x"2e",
           559 => x"12",
           560 => x"52",
           561 => x"71",
           562 => x"8c",
           563 => x"3d",
           564 => x"3d",
           565 => x"7c",
           566 => x"55",
           567 => x"2e",
           568 => x"71",
           569 => x"06",
           570 => x"2e",
           571 => x"ff",
           572 => x"ff",
           573 => x"71",
           574 => x"56",
           575 => x"2e",
           576 => x"a9",
           577 => x"2e",
           578 => x"70",
           579 => x"51",
           580 => x"80",
           581 => x"12",
           582 => x"15",
           583 => x"72",
           584 => x"81",
           585 => x"71",
           586 => x"56",
           587 => x"ff",
           588 => x"ff",
           589 => x"31",
           590 => x"70",
           591 => x"0c",
           592 => x"04",
           593 => x"55",
           594 => x"88",
           595 => x"74",
           596 => x"38",
           597 => x"52",
           598 => x"fc",
           599 => x"80",
           600 => x"74",
           601 => x"f7",
           602 => x"12",
           603 => x"84",
           604 => x"06",
           605 => x"70",
           606 => x"15",
           607 => x"55",
           608 => x"d0",
           609 => x"76",
           610 => x"38",
           611 => x"52",
           612 => x"80",
           613 => x"dc",
           614 => x"0d",
           615 => x"0d",
           616 => x"53",
           617 => x"52",
           618 => x"82",
           619 => x"81",
           620 => x"07",
           621 => x"52",
           622 => x"e8",
           623 => x"8c",
           624 => x"3d",
           625 => x"3d",
           626 => x"08",
           627 => x"56",
           628 => x"80",
           629 => x"33",
           630 => x"2e",
           631 => x"86",
           632 => x"52",
           633 => x"53",
           634 => x"13",
           635 => x"33",
           636 => x"06",
           637 => x"70",
           638 => x"38",
           639 => x"80",
           640 => x"74",
           641 => x"81",
           642 => x"70",
           643 => x"81",
           644 => x"80",
           645 => x"05",
           646 => x"76",
           647 => x"70",
           648 => x"0c",
           649 => x"04",
           650 => x"76",
           651 => x"80",
           652 => x"86",
           653 => x"52",
           654 => x"99",
           655 => x"dc",
           656 => x"80",
           657 => x"74",
           658 => x"8c",
           659 => x"3d",
           660 => x"3d",
           661 => x"11",
           662 => x"52",
           663 => x"70",
           664 => x"98",
           665 => x"33",
           666 => x"82",
           667 => x"26",
           668 => x"84",
           669 => x"83",
           670 => x"26",
           671 => x"85",
           672 => x"84",
           673 => x"26",
           674 => x"86",
           675 => x"85",
           676 => x"26",
           677 => x"88",
           678 => x"86",
           679 => x"e7",
           680 => x"38",
           681 => x"54",
           682 => x"87",
           683 => x"cc",
           684 => x"87",
           685 => x"0c",
           686 => x"c0",
           687 => x"82",
           688 => x"c0",
           689 => x"83",
           690 => x"c0",
           691 => x"84",
           692 => x"c0",
           693 => x"85",
           694 => x"c0",
           695 => x"86",
           696 => x"c0",
           697 => x"74",
           698 => x"a4",
           699 => x"c0",
           700 => x"80",
           701 => x"98",
           702 => x"52",
           703 => x"dc",
           704 => x"0d",
           705 => x"0d",
           706 => x"c0",
           707 => x"81",
           708 => x"c0",
           709 => x"5e",
           710 => x"87",
           711 => x"08",
           712 => x"1c",
           713 => x"98",
           714 => x"79",
           715 => x"87",
           716 => x"08",
           717 => x"1c",
           718 => x"98",
           719 => x"79",
           720 => x"87",
           721 => x"08",
           722 => x"1c",
           723 => x"98",
           724 => x"7b",
           725 => x"87",
           726 => x"08",
           727 => x"1c",
           728 => x"0c",
           729 => x"ff",
           730 => x"83",
           731 => x"58",
           732 => x"57",
           733 => x"56",
           734 => x"55",
           735 => x"54",
           736 => x"53",
           737 => x"ff",
           738 => x"f1",
           739 => x"de",
           740 => x"0d",
           741 => x"0d",
           742 => x"33",
           743 => x"9f",
           744 => x"52",
           745 => x"82",
           746 => x"83",
           747 => x"fb",
           748 => x"0b",
           749 => x"d4",
           750 => x"ff",
           751 => x"56",
           752 => x"84",
           753 => x"2e",
           754 => x"c0",
           755 => x"70",
           756 => x"2a",
           757 => x"53",
           758 => x"80",
           759 => x"71",
           760 => x"81",
           761 => x"70",
           762 => x"81",
           763 => x"06",
           764 => x"80",
           765 => x"71",
           766 => x"81",
           767 => x"70",
           768 => x"73",
           769 => x"51",
           770 => x"80",
           771 => x"2e",
           772 => x"c0",
           773 => x"75",
           774 => x"82",
           775 => x"87",
           776 => x"fb",
           777 => x"9f",
           778 => x"0b",
           779 => x"33",
           780 => x"06",
           781 => x"87",
           782 => x"51",
           783 => x"86",
           784 => x"94",
           785 => x"08",
           786 => x"70",
           787 => x"54",
           788 => x"2e",
           789 => x"91",
           790 => x"06",
           791 => x"d7",
           792 => x"32",
           793 => x"51",
           794 => x"2e",
           795 => x"93",
           796 => x"06",
           797 => x"ff",
           798 => x"81",
           799 => x"87",
           800 => x"52",
           801 => x"86",
           802 => x"94",
           803 => x"72",
           804 => x"0d",
           805 => x"0d",
           806 => x"74",
           807 => x"ff",
           808 => x"57",
           809 => x"80",
           810 => x"81",
           811 => x"15",
           812 => x"87",
           813 => x"81",
           814 => x"57",
           815 => x"c0",
           816 => x"75",
           817 => x"38",
           818 => x"94",
           819 => x"70",
           820 => x"81",
           821 => x"52",
           822 => x"8c",
           823 => x"2a",
           824 => x"51",
           825 => x"38",
           826 => x"70",
           827 => x"51",
           828 => x"8d",
           829 => x"2a",
           830 => x"51",
           831 => x"be",
           832 => x"ff",
           833 => x"c0",
           834 => x"70",
           835 => x"38",
           836 => x"90",
           837 => x"0c",
           838 => x"33",
           839 => x"06",
           840 => x"70",
           841 => x"76",
           842 => x"0c",
           843 => x"04",
           844 => x"0b",
           845 => x"d4",
           846 => x"ff",
           847 => x"87",
           848 => x"51",
           849 => x"86",
           850 => x"94",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"2e",
           855 => x"81",
           856 => x"87",
           857 => x"52",
           858 => x"86",
           859 => x"94",
           860 => x"08",
           861 => x"06",
           862 => x"0c",
           863 => x"0d",
           864 => x"0d",
           865 => x"87",
           866 => x"81",
           867 => x"53",
           868 => x"84",
           869 => x"2e",
           870 => x"c0",
           871 => x"71",
           872 => x"2a",
           873 => x"51",
           874 => x"52",
           875 => x"a0",
           876 => x"ff",
           877 => x"c0",
           878 => x"70",
           879 => x"38",
           880 => x"90",
           881 => x"70",
           882 => x"98",
           883 => x"51",
           884 => x"dc",
           885 => x"0d",
           886 => x"0d",
           887 => x"80",
           888 => x"2a",
           889 => x"51",
           890 => x"84",
           891 => x"c0",
           892 => x"82",
           893 => x"87",
           894 => x"08",
           895 => x"0c",
           896 => x"94",
           897 => x"e0",
           898 => x"9e",
           899 => x"87",
           900 => x"c0",
           901 => x"82",
           902 => x"87",
           903 => x"08",
           904 => x"0c",
           905 => x"ac",
           906 => x"f0",
           907 => x"9e",
           908 => x"87",
           909 => x"c0",
           910 => x"82",
           911 => x"87",
           912 => x"08",
           913 => x"0c",
           914 => x"bc",
           915 => x"80",
           916 => x"9e",
           917 => x"88",
           918 => x"c0",
           919 => x"82",
           920 => x"87",
           921 => x"08",
           922 => x"88",
           923 => x"c0",
           924 => x"82",
           925 => x"87",
           926 => x"08",
           927 => x"0c",
           928 => x"8c",
           929 => x"98",
           930 => x"82",
           931 => x"80",
           932 => x"9e",
           933 => x"84",
           934 => x"51",
           935 => x"80",
           936 => x"81",
           937 => x"88",
           938 => x"0b",
           939 => x"90",
           940 => x"80",
           941 => x"52",
           942 => x"2e",
           943 => x"52",
           944 => x"9e",
           945 => x"87",
           946 => x"08",
           947 => x"0a",
           948 => x"52",
           949 => x"83",
           950 => x"71",
           951 => x"34",
           952 => x"c0",
           953 => x"70",
           954 => x"06",
           955 => x"70",
           956 => x"38",
           957 => x"82",
           958 => x"80",
           959 => x"9e",
           960 => x"a0",
           961 => x"51",
           962 => x"80",
           963 => x"81",
           964 => x"88",
           965 => x"0b",
           966 => x"90",
           967 => x"80",
           968 => x"52",
           969 => x"2e",
           970 => x"52",
           971 => x"a2",
           972 => x"87",
           973 => x"08",
           974 => x"80",
           975 => x"52",
           976 => x"83",
           977 => x"71",
           978 => x"34",
           979 => x"c0",
           980 => x"70",
           981 => x"06",
           982 => x"70",
           983 => x"38",
           984 => x"82",
           985 => x"80",
           986 => x"9e",
           987 => x"81",
           988 => x"51",
           989 => x"80",
           990 => x"81",
           991 => x"88",
           992 => x"0b",
           993 => x"90",
           994 => x"c0",
           995 => x"52",
           996 => x"2e",
           997 => x"52",
           998 => x"a6",
           999 => x"87",
          1000 => x"08",
          1001 => x"06",
          1002 => x"70",
          1003 => x"38",
          1004 => x"82",
          1005 => x"87",
          1006 => x"08",
          1007 => x"06",
          1008 => x"51",
          1009 => x"82",
          1010 => x"80",
          1011 => x"9e",
          1012 => x"84",
          1013 => x"52",
          1014 => x"2e",
          1015 => x"52",
          1016 => x"a9",
          1017 => x"9e",
          1018 => x"83",
          1019 => x"84",
          1020 => x"51",
          1021 => x"aa",
          1022 => x"87",
          1023 => x"08",
          1024 => x"51",
          1025 => x"80",
          1026 => x"81",
          1027 => x"88",
          1028 => x"c0",
          1029 => x"70",
          1030 => x"51",
          1031 => x"ac",
          1032 => x"0d",
          1033 => x"0d",
          1034 => x"51",
          1035 => x"82",
          1036 => x"54",
          1037 => x"88",
          1038 => x"90",
          1039 => x"3f",
          1040 => x"51",
          1041 => x"82",
          1042 => x"54",
          1043 => x"93",
          1044 => x"f8",
          1045 => x"fc",
          1046 => x"52",
          1047 => x"51",
          1048 => x"82",
          1049 => x"54",
          1050 => x"93",
          1051 => x"f0",
          1052 => x"f4",
          1053 => x"52",
          1054 => x"51",
          1055 => x"82",
          1056 => x"54",
          1057 => x"93",
          1058 => x"d8",
          1059 => x"dc",
          1060 => x"52",
          1061 => x"51",
          1062 => x"82",
          1063 => x"54",
          1064 => x"93",
          1065 => x"e0",
          1066 => x"e4",
          1067 => x"52",
          1068 => x"51",
          1069 => x"82",
          1070 => x"54",
          1071 => x"93",
          1072 => x"e8",
          1073 => x"ec",
          1074 => x"52",
          1075 => x"51",
          1076 => x"82",
          1077 => x"54",
          1078 => x"8d",
          1079 => x"a8",
          1080 => x"f3",
          1081 => x"86",
          1082 => x"ab",
          1083 => x"80",
          1084 => x"82",
          1085 => x"52",
          1086 => x"51",
          1087 => x"82",
          1088 => x"54",
          1089 => x"8d",
          1090 => x"aa",
          1091 => x"f4",
          1092 => x"da",
          1093 => x"9d",
          1094 => x"80",
          1095 => x"81",
          1096 => x"87",
          1097 => x"88",
          1098 => x"73",
          1099 => x"38",
          1100 => x"51",
          1101 => x"82",
          1102 => x"54",
          1103 => x"88",
          1104 => x"c8",
          1105 => x"3f",
          1106 => x"33",
          1107 => x"2e",
          1108 => x"f4",
          1109 => x"b2",
          1110 => x"a6",
          1111 => x"80",
          1112 => x"81",
          1113 => x"87",
          1114 => x"f4",
          1115 => x"9a",
          1116 => x"80",
          1117 => x"f4",
          1118 => x"f2",
          1119 => x"84",
          1120 => x"f5",
          1121 => x"e6",
          1122 => x"88",
          1123 => x"f5",
          1124 => x"da",
          1125 => x"f0",
          1126 => x"3f",
          1127 => x"22",
          1128 => x"f8",
          1129 => x"3f",
          1130 => x"08",
          1131 => x"c0",
          1132 => x"e7",
          1133 => x"8c",
          1134 => x"84",
          1135 => x"71",
          1136 => x"82",
          1137 => x"52",
          1138 => x"51",
          1139 => x"82",
          1140 => x"54",
          1141 => x"a8",
          1142 => x"94",
          1143 => x"84",
          1144 => x"51",
          1145 => x"82",
          1146 => x"bd",
          1147 => x"76",
          1148 => x"54",
          1149 => x"08",
          1150 => x"cc",
          1151 => x"3f",
          1152 => x"33",
          1153 => x"2e",
          1154 => x"88",
          1155 => x"bd",
          1156 => x"75",
          1157 => x"3f",
          1158 => x"08",
          1159 => x"29",
          1160 => x"54",
          1161 => x"dc",
          1162 => x"f6",
          1163 => x"be",
          1164 => x"a4",
          1165 => x"3f",
          1166 => x"04",
          1167 => x"02",
          1168 => x"ff",
          1169 => x"84",
          1170 => x"71",
          1171 => x"0b",
          1172 => x"05",
          1173 => x"04",
          1174 => x"51",
          1175 => x"f7",
          1176 => x"39",
          1177 => x"51",
          1178 => x"f7",
          1179 => x"39",
          1180 => x"51",
          1181 => x"f7",
          1182 => x"8e",
          1183 => x"0d",
          1184 => x"80",
          1185 => x"0b",
          1186 => x"84",
          1187 => x"88",
          1188 => x"c0",
          1189 => x"04",
          1190 => x"82",
          1191 => x"89",
          1192 => x"9c",
          1193 => x"ec",
          1194 => x"ec",
          1195 => x"52",
          1196 => x"70",
          1197 => x"26",
          1198 => x"82",
          1199 => x"71",
          1200 => x"8c",
          1201 => x"3d",
          1202 => x"3d",
          1203 => x"84",
          1204 => x"12",
          1205 => x"94",
          1206 => x"16",
          1207 => x"54",
          1208 => x"70",
          1209 => x"38",
          1210 => x"14",
          1211 => x"81",
          1212 => x"76",
          1213 => x"0c",
          1214 => x"75",
          1215 => x"72",
          1216 => x"71",
          1217 => x"70",
          1218 => x"70",
          1219 => x"73",
          1220 => x"74",
          1221 => x"70",
          1222 => x"70",
          1223 => x"8c",
          1224 => x"0c",
          1225 => x"0c",
          1226 => x"0c",
          1227 => x"dc",
          1228 => x"0d",
          1229 => x"0d",
          1230 => x"08",
          1231 => x"56",
          1232 => x"08",
          1233 => x"81",
          1234 => x"84",
          1235 => x"13",
          1236 => x"73",
          1237 => x"06",
          1238 => x"13",
          1239 => x"13",
          1240 => x"13",
          1241 => x"15",
          1242 => x"9f",
          1243 => x"0c",
          1244 => x"08",
          1245 => x"82",
          1246 => x"94",
          1247 => x"82",
          1248 => x"90",
          1249 => x"94",
          1250 => x"73",
          1251 => x"09",
          1252 => x"38",
          1253 => x"70",
          1254 => x"70",
          1255 => x"81",
          1256 => x"84",
          1257 => x"84",
          1258 => x"14",
          1259 => x"08",
          1260 => x"0c",
          1261 => x"0c",
          1262 => x"88",
          1263 => x"88",
          1264 => x"8c",
          1265 => x"82",
          1266 => x"86",
          1267 => x"f9",
          1268 => x"70",
          1269 => x"80",
          1270 => x"38",
          1271 => x"06",
          1272 => x"08",
          1273 => x"08",
          1274 => x"38",
          1275 => x"77",
          1276 => x"38",
          1277 => x"56",
          1278 => x"ff",
          1279 => x"80",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"08",
          1283 => x"08",
          1284 => x"8c",
          1285 => x"80",
          1286 => x"dc",
          1287 => x"30",
          1288 => x"80",
          1289 => x"53",
          1290 => x"54",
          1291 => x"72",
          1292 => x"81",
          1293 => x"38",
          1294 => x"52",
          1295 => x"c8",
          1296 => x"82",
          1297 => x"0c",
          1298 => x"dc",
          1299 => x"0c",
          1300 => x"08",
          1301 => x"82",
          1302 => x"75",
          1303 => x"38",
          1304 => x"53",
          1305 => x"13",
          1306 => x"0c",
          1307 => x"0c",
          1308 => x"0c",
          1309 => x"76",
          1310 => x"53",
          1311 => x"b5",
          1312 => x"82",
          1313 => x"51",
          1314 => x"82",
          1315 => x"54",
          1316 => x"dc",
          1317 => x"0d",
          1318 => x"0d",
          1319 => x"80",
          1320 => x"f0",
          1321 => x"8d",
          1322 => x"0d",
          1323 => x"0d",
          1324 => x"33",
          1325 => x"2e",
          1326 => x"85",
          1327 => x"ed",
          1328 => x"f8",
          1329 => x"80",
          1330 => x"72",
          1331 => x"8c",
          1332 => x"05",
          1333 => x"0c",
          1334 => x"8c",
          1335 => x"71",
          1336 => x"38",
          1337 => x"2d",
          1338 => x"04",
          1339 => x"02",
          1340 => x"82",
          1341 => x"76",
          1342 => x"0c",
          1343 => x"ad",
          1344 => x"8c",
          1345 => x"3d",
          1346 => x"3d",
          1347 => x"73",
          1348 => x"ff",
          1349 => x"71",
          1350 => x"38",
          1351 => x"06",
          1352 => x"54",
          1353 => x"e7",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"f0",
          1357 => x"8c",
          1358 => x"54",
          1359 => x"81",
          1360 => x"53",
          1361 => x"8e",
          1362 => x"ff",
          1363 => x"14",
          1364 => x"3f",
          1365 => x"82",
          1366 => x"86",
          1367 => x"ec",
          1368 => x"68",
          1369 => x"70",
          1370 => x"33",
          1371 => x"2e",
          1372 => x"75",
          1373 => x"81",
          1374 => x"38",
          1375 => x"70",
          1376 => x"33",
          1377 => x"75",
          1378 => x"81",
          1379 => x"81",
          1380 => x"75",
          1381 => x"81",
          1382 => x"82",
          1383 => x"81",
          1384 => x"56",
          1385 => x"09",
          1386 => x"38",
          1387 => x"71",
          1388 => x"81",
          1389 => x"59",
          1390 => x"9d",
          1391 => x"53",
          1392 => x"95",
          1393 => x"29",
          1394 => x"76",
          1395 => x"79",
          1396 => x"5b",
          1397 => x"e5",
          1398 => x"ec",
          1399 => x"70",
          1400 => x"25",
          1401 => x"32",
          1402 => x"72",
          1403 => x"73",
          1404 => x"58",
          1405 => x"73",
          1406 => x"38",
          1407 => x"79",
          1408 => x"5b",
          1409 => x"75",
          1410 => x"de",
          1411 => x"80",
          1412 => x"89",
          1413 => x"70",
          1414 => x"55",
          1415 => x"cf",
          1416 => x"38",
          1417 => x"24",
          1418 => x"80",
          1419 => x"8e",
          1420 => x"c3",
          1421 => x"73",
          1422 => x"81",
          1423 => x"99",
          1424 => x"c4",
          1425 => x"38",
          1426 => x"73",
          1427 => x"81",
          1428 => x"80",
          1429 => x"38",
          1430 => x"2e",
          1431 => x"f9",
          1432 => x"d8",
          1433 => x"38",
          1434 => x"77",
          1435 => x"08",
          1436 => x"80",
          1437 => x"55",
          1438 => x"8d",
          1439 => x"70",
          1440 => x"51",
          1441 => x"f5",
          1442 => x"2a",
          1443 => x"74",
          1444 => x"53",
          1445 => x"8f",
          1446 => x"fc",
          1447 => x"81",
          1448 => x"80",
          1449 => x"73",
          1450 => x"3f",
          1451 => x"56",
          1452 => x"27",
          1453 => x"a0",
          1454 => x"3f",
          1455 => x"84",
          1456 => x"33",
          1457 => x"93",
          1458 => x"95",
          1459 => x"91",
          1460 => x"8d",
          1461 => x"89",
          1462 => x"fb",
          1463 => x"86",
          1464 => x"2a",
          1465 => x"51",
          1466 => x"2e",
          1467 => x"84",
          1468 => x"86",
          1469 => x"78",
          1470 => x"08",
          1471 => x"32",
          1472 => x"72",
          1473 => x"51",
          1474 => x"74",
          1475 => x"38",
          1476 => x"88",
          1477 => x"7a",
          1478 => x"55",
          1479 => x"3d",
          1480 => x"52",
          1481 => x"e9",
          1482 => x"dc",
          1483 => x"06",
          1484 => x"52",
          1485 => x"3f",
          1486 => x"08",
          1487 => x"27",
          1488 => x"14",
          1489 => x"f8",
          1490 => x"87",
          1491 => x"81",
          1492 => x"b0",
          1493 => x"7d",
          1494 => x"5f",
          1495 => x"75",
          1496 => x"07",
          1497 => x"54",
          1498 => x"26",
          1499 => x"ff",
          1500 => x"84",
          1501 => x"06",
          1502 => x"80",
          1503 => x"96",
          1504 => x"e0",
          1505 => x"73",
          1506 => x"57",
          1507 => x"06",
          1508 => x"54",
          1509 => x"a0",
          1510 => x"2a",
          1511 => x"54",
          1512 => x"38",
          1513 => x"76",
          1514 => x"38",
          1515 => x"fd",
          1516 => x"06",
          1517 => x"38",
          1518 => x"56",
          1519 => x"26",
          1520 => x"3d",
          1521 => x"05",
          1522 => x"ff",
          1523 => x"53",
          1524 => x"d9",
          1525 => x"38",
          1526 => x"56",
          1527 => x"27",
          1528 => x"a0",
          1529 => x"3f",
          1530 => x"3d",
          1531 => x"3d",
          1532 => x"70",
          1533 => x"52",
          1534 => x"73",
          1535 => x"3f",
          1536 => x"04",
          1537 => x"74",
          1538 => x"0c",
          1539 => x"05",
          1540 => x"fa",
          1541 => x"8c",
          1542 => x"80",
          1543 => x"0b",
          1544 => x"0c",
          1545 => x"04",
          1546 => x"82",
          1547 => x"76",
          1548 => x"0c",
          1549 => x"05",
          1550 => x"53",
          1551 => x"72",
          1552 => x"0c",
          1553 => x"04",
          1554 => x"77",
          1555 => x"f4",
          1556 => x"54",
          1557 => x"54",
          1558 => x"80",
          1559 => x"8c",
          1560 => x"71",
          1561 => x"dc",
          1562 => x"06",
          1563 => x"2e",
          1564 => x"72",
          1565 => x"38",
          1566 => x"70",
          1567 => x"25",
          1568 => x"73",
          1569 => x"38",
          1570 => x"86",
          1571 => x"54",
          1572 => x"73",
          1573 => x"ff",
          1574 => x"72",
          1575 => x"74",
          1576 => x"72",
          1577 => x"54",
          1578 => x"81",
          1579 => x"39",
          1580 => x"80",
          1581 => x"51",
          1582 => x"81",
          1583 => x"8c",
          1584 => x"3d",
          1585 => x"3d",
          1586 => x"f4",
          1587 => x"8c",
          1588 => x"53",
          1589 => x"fe",
          1590 => x"82",
          1591 => x"84",
          1592 => x"f8",
          1593 => x"7c",
          1594 => x"70",
          1595 => x"75",
          1596 => x"55",
          1597 => x"2e",
          1598 => x"87",
          1599 => x"76",
          1600 => x"73",
          1601 => x"81",
          1602 => x"81",
          1603 => x"77",
          1604 => x"70",
          1605 => x"58",
          1606 => x"09",
          1607 => x"c2",
          1608 => x"81",
          1609 => x"75",
          1610 => x"55",
          1611 => x"e2",
          1612 => x"90",
          1613 => x"f8",
          1614 => x"8f",
          1615 => x"81",
          1616 => x"75",
          1617 => x"55",
          1618 => x"81",
          1619 => x"27",
          1620 => x"d0",
          1621 => x"55",
          1622 => x"73",
          1623 => x"80",
          1624 => x"14",
          1625 => x"72",
          1626 => x"e0",
          1627 => x"80",
          1628 => x"39",
          1629 => x"55",
          1630 => x"80",
          1631 => x"e0",
          1632 => x"38",
          1633 => x"81",
          1634 => x"53",
          1635 => x"81",
          1636 => x"53",
          1637 => x"8e",
          1638 => x"70",
          1639 => x"55",
          1640 => x"27",
          1641 => x"77",
          1642 => x"74",
          1643 => x"76",
          1644 => x"77",
          1645 => x"70",
          1646 => x"55",
          1647 => x"77",
          1648 => x"38",
          1649 => x"74",
          1650 => x"55",
          1651 => x"dc",
          1652 => x"0d",
          1653 => x"0d",
          1654 => x"56",
          1655 => x"0c",
          1656 => x"70",
          1657 => x"73",
          1658 => x"81",
          1659 => x"81",
          1660 => x"ed",
          1661 => x"2e",
          1662 => x"8e",
          1663 => x"08",
          1664 => x"76",
          1665 => x"56",
          1666 => x"b0",
          1667 => x"06",
          1668 => x"75",
          1669 => x"76",
          1670 => x"70",
          1671 => x"73",
          1672 => x"8b",
          1673 => x"73",
          1674 => x"85",
          1675 => x"82",
          1676 => x"76",
          1677 => x"70",
          1678 => x"ac",
          1679 => x"a0",
          1680 => x"fa",
          1681 => x"53",
          1682 => x"57",
          1683 => x"98",
          1684 => x"39",
          1685 => x"80",
          1686 => x"26",
          1687 => x"86",
          1688 => x"80",
          1689 => x"57",
          1690 => x"74",
          1691 => x"38",
          1692 => x"27",
          1693 => x"14",
          1694 => x"06",
          1695 => x"14",
          1696 => x"06",
          1697 => x"74",
          1698 => x"f9",
          1699 => x"ff",
          1700 => x"89",
          1701 => x"38",
          1702 => x"c5",
          1703 => x"29",
          1704 => x"81",
          1705 => x"76",
          1706 => x"56",
          1707 => x"ba",
          1708 => x"2e",
          1709 => x"30",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"8a",
          1713 => x"fd",
          1714 => x"98",
          1715 => x"2c",
          1716 => x"70",
          1717 => x"10",
          1718 => x"2b",
          1719 => x"54",
          1720 => x"0b",
          1721 => x"12",
          1722 => x"71",
          1723 => x"38",
          1724 => x"11",
          1725 => x"84",
          1726 => x"33",
          1727 => x"52",
          1728 => x"2e",
          1729 => x"83",
          1730 => x"72",
          1731 => x"0c",
          1732 => x"04",
          1733 => x"78",
          1734 => x"9f",
          1735 => x"33",
          1736 => x"71",
          1737 => x"38",
          1738 => x"81",
          1739 => x"f2",
          1740 => x"51",
          1741 => x"72",
          1742 => x"52",
          1743 => x"71",
          1744 => x"52",
          1745 => x"51",
          1746 => x"73",
          1747 => x"3d",
          1748 => x"3d",
          1749 => x"84",
          1750 => x"33",
          1751 => x"bb",
          1752 => x"89",
          1753 => x"84",
          1754 => x"d0",
          1755 => x"51",
          1756 => x"58",
          1757 => x"2e",
          1758 => x"51",
          1759 => x"82",
          1760 => x"70",
          1761 => x"88",
          1762 => x"19",
          1763 => x"56",
          1764 => x"3f",
          1765 => x"08",
          1766 => x"89",
          1767 => x"84",
          1768 => x"d0",
          1769 => x"51",
          1770 => x"80",
          1771 => x"75",
          1772 => x"74",
          1773 => x"3f",
          1774 => x"33",
          1775 => x"74",
          1776 => x"34",
          1777 => x"06",
          1778 => x"27",
          1779 => x"0b",
          1780 => x"34",
          1781 => x"b6",
          1782 => x"a4",
          1783 => x"80",
          1784 => x"82",
          1785 => x"55",
          1786 => x"8c",
          1787 => x"54",
          1788 => x"52",
          1789 => x"c8",
          1790 => x"89",
          1791 => x"8a",
          1792 => x"9e",
          1793 => x"a4",
          1794 => x"cb",
          1795 => x"3d",
          1796 => x"3d",
          1797 => x"80",
          1798 => x"a4",
          1799 => x"d2",
          1800 => x"8c",
          1801 => x"d1",
          1802 => x"a4",
          1803 => x"f8",
          1804 => x"70",
          1805 => x"fa",
          1806 => x"8c",
          1807 => x"2e",
          1808 => x"51",
          1809 => x"82",
          1810 => x"55",
          1811 => x"8c",
          1812 => x"9c",
          1813 => x"dc",
          1814 => x"70",
          1815 => x"80",
          1816 => x"53",
          1817 => x"17",
          1818 => x"52",
          1819 => x"3f",
          1820 => x"09",
          1821 => x"b1",
          1822 => x"0d",
          1823 => x"0d",
          1824 => x"ad",
          1825 => x"5a",
          1826 => x"58",
          1827 => x"89",
          1828 => x"80",
          1829 => x"82",
          1830 => x"81",
          1831 => x"0b",
          1832 => x"08",
          1833 => x"f8",
          1834 => x"70",
          1835 => x"f9",
          1836 => x"8c",
          1837 => x"2e",
          1838 => x"51",
          1839 => x"82",
          1840 => x"81",
          1841 => x"80",
          1842 => x"dc",
          1843 => x"38",
          1844 => x"08",
          1845 => x"17",
          1846 => x"74",
          1847 => x"70",
          1848 => x"07",
          1849 => x"55",
          1850 => x"2e",
          1851 => x"ff",
          1852 => x"89",
          1853 => x"11",
          1854 => x"80",
          1855 => x"82",
          1856 => x"80",
          1857 => x"81",
          1858 => x"ef",
          1859 => x"77",
          1860 => x"06",
          1861 => x"52",
          1862 => x"e6",
          1863 => x"d6",
          1864 => x"3d",
          1865 => x"8c",
          1866 => x"34",
          1867 => x"82",
          1868 => x"a9",
          1869 => x"f6",
          1870 => x"7e",
          1871 => x"72",
          1872 => x"5a",
          1873 => x"2e",
          1874 => x"a2",
          1875 => x"78",
          1876 => x"76",
          1877 => x"81",
          1878 => x"70",
          1879 => x"58",
          1880 => x"2e",
          1881 => x"86",
          1882 => x"26",
          1883 => x"54",
          1884 => x"82",
          1885 => x"70",
          1886 => x"d5",
          1887 => x"8c",
          1888 => x"79",
          1889 => x"51",
          1890 => x"82",
          1891 => x"80",
          1892 => x"15",
          1893 => x"81",
          1894 => x"74",
          1895 => x"38",
          1896 => x"ee",
          1897 => x"81",
          1898 => x"3d",
          1899 => x"f8",
          1900 => x"af",
          1901 => x"dc",
          1902 => x"99",
          1903 => x"78",
          1904 => x"fd",
          1905 => x"8c",
          1906 => x"ff",
          1907 => x"85",
          1908 => x"91",
          1909 => x"70",
          1910 => x"51",
          1911 => x"27",
          1912 => x"80",
          1913 => x"8c",
          1914 => x"3d",
          1915 => x"3d",
          1916 => x"08",
          1917 => x"81",
          1918 => x"5f",
          1919 => x"af",
          1920 => x"89",
          1921 => x"82",
          1922 => x"81",
          1923 => x"89",
          1924 => x"73",
          1925 => x"a8",
          1926 => x"3f",
          1927 => x"08",
          1928 => x"0c",
          1929 => x"08",
          1930 => x"fe",
          1931 => x"82",
          1932 => x"52",
          1933 => x"08",
          1934 => x"3f",
          1935 => x"08",
          1936 => x"38",
          1937 => x"51",
          1938 => x"80",
          1939 => x"89",
          1940 => x"80",
          1941 => x"3d",
          1942 => x"80",
          1943 => x"82",
          1944 => x"56",
          1945 => x"08",
          1946 => x"81",
          1947 => x"38",
          1948 => x"08",
          1949 => x"3f",
          1950 => x"08",
          1951 => x"82",
          1952 => x"25",
          1953 => x"8c",
          1954 => x"05",
          1955 => x"55",
          1956 => x"80",
          1957 => x"ff",
          1958 => x"51",
          1959 => x"74",
          1960 => x"81",
          1961 => x"38",
          1962 => x"0b",
          1963 => x"34",
          1964 => x"dd",
          1965 => x"8c",
          1966 => x"2b",
          1967 => x"51",
          1968 => x"2e",
          1969 => x"81",
          1970 => x"8d",
          1971 => x"98",
          1972 => x"2c",
          1973 => x"33",
          1974 => x"70",
          1975 => x"98",
          1976 => x"84",
          1977 => x"d8",
          1978 => x"15",
          1979 => x"51",
          1980 => x"59",
          1981 => x"58",
          1982 => x"78",
          1983 => x"38",
          1984 => x"b4",
          1985 => x"80",
          1986 => x"ff",
          1987 => x"98",
          1988 => x"80",
          1989 => x"ce",
          1990 => x"74",
          1991 => x"f7",
          1992 => x"8c",
          1993 => x"ff",
          1994 => x"80",
          1995 => x"74",
          1996 => x"34",
          1997 => x"39",
          1998 => x"0a",
          1999 => x"0a",
          2000 => x"2c",
          2001 => x"06",
          2002 => x"73",
          2003 => x"38",
          2004 => x"52",
          2005 => x"ef",
          2006 => x"dc",
          2007 => x"06",
          2008 => x"38",
          2009 => x"56",
          2010 => x"80",
          2011 => x"1c",
          2012 => x"8d",
          2013 => x"98",
          2014 => x"2c",
          2015 => x"33",
          2016 => x"70",
          2017 => x"10",
          2018 => x"2b",
          2019 => x"11",
          2020 => x"51",
          2021 => x"51",
          2022 => x"2e",
          2023 => x"fe",
          2024 => x"f8",
          2025 => x"7d",
          2026 => x"82",
          2027 => x"80",
          2028 => x"fc",
          2029 => x"75",
          2030 => x"34",
          2031 => x"fc",
          2032 => x"3d",
          2033 => x"0c",
          2034 => x"8b",
          2035 => x"38",
          2036 => x"81",
          2037 => x"54",
          2038 => x"82",
          2039 => x"54",
          2040 => x"fd",
          2041 => x"8d",
          2042 => x"73",
          2043 => x"38",
          2044 => x"70",
          2045 => x"55",
          2046 => x"9e",
          2047 => x"54",
          2048 => x"15",
          2049 => x"80",
          2050 => x"ff",
          2051 => x"98",
          2052 => x"88",
          2053 => x"55",
          2054 => x"8d",
          2055 => x"11",
          2056 => x"82",
          2057 => x"73",
          2058 => x"3d",
          2059 => x"82",
          2060 => x"54",
          2061 => x"89",
          2062 => x"54",
          2063 => x"84",
          2064 => x"88",
          2065 => x"80",
          2066 => x"ff",
          2067 => x"98",
          2068 => x"84",
          2069 => x"56",
          2070 => x"25",
          2071 => x"1a",
          2072 => x"54",
          2073 => x"74",
          2074 => x"29",
          2075 => x"05",
          2076 => x"82",
          2077 => x"56",
          2078 => x"75",
          2079 => x"82",
          2080 => x"70",
          2081 => x"98",
          2082 => x"84",
          2083 => x"56",
          2084 => x"25",
          2085 => x"88",
          2086 => x"3f",
          2087 => x"0a",
          2088 => x"0a",
          2089 => x"2c",
          2090 => x"33",
          2091 => x"73",
          2092 => x"38",
          2093 => x"82",
          2094 => x"70",
          2095 => x"55",
          2096 => x"2e",
          2097 => x"82",
          2098 => x"ff",
          2099 => x"82",
          2100 => x"ff",
          2101 => x"82",
          2102 => x"88",
          2103 => x"3f",
          2104 => x"33",
          2105 => x"70",
          2106 => x"8d",
          2107 => x"51",
          2108 => x"74",
          2109 => x"74",
          2110 => x"14",
          2111 => x"73",
          2112 => x"a9",
          2113 => x"80",
          2114 => x"80",
          2115 => x"98",
          2116 => x"84",
          2117 => x"55",
          2118 => x"db",
          2119 => x"e7",
          2120 => x"8d",
          2121 => x"98",
          2122 => x"2c",
          2123 => x"33",
          2124 => x"57",
          2125 => x"fa",
          2126 => x"51",
          2127 => x"74",
          2128 => x"29",
          2129 => x"05",
          2130 => x"82",
          2131 => x"58",
          2132 => x"75",
          2133 => x"fa",
          2134 => x"8d",
          2135 => x"05",
          2136 => x"34",
          2137 => x"c5",
          2138 => x"84",
          2139 => x"f7",
          2140 => x"8c",
          2141 => x"ff",
          2142 => x"98",
          2143 => x"84",
          2144 => x"80",
          2145 => x"38",
          2146 => x"52",
          2147 => x"c2",
          2148 => x"39",
          2149 => x"84",
          2150 => x"8d",
          2151 => x"73",
          2152 => x"8c",
          2153 => x"e6",
          2154 => x"8d",
          2155 => x"05",
          2156 => x"8d",
          2157 => x"81",
          2158 => x"e3",
          2159 => x"88",
          2160 => x"84",
          2161 => x"73",
          2162 => x"e4",
          2163 => x"54",
          2164 => x"84",
          2165 => x"2b",
          2166 => x"75",
          2167 => x"56",
          2168 => x"74",
          2169 => x"74",
          2170 => x"14",
          2171 => x"73",
          2172 => x"b9",
          2173 => x"80",
          2174 => x"80",
          2175 => x"98",
          2176 => x"84",
          2177 => x"55",
          2178 => x"db",
          2179 => x"e5",
          2180 => x"8d",
          2181 => x"98",
          2182 => x"2c",
          2183 => x"33",
          2184 => x"57",
          2185 => x"f9",
          2186 => x"51",
          2187 => x"74",
          2188 => x"29",
          2189 => x"05",
          2190 => x"82",
          2191 => x"58",
          2192 => x"75",
          2193 => x"f8",
          2194 => x"8d",
          2195 => x"81",
          2196 => x"8d",
          2197 => x"56",
          2198 => x"27",
          2199 => x"81",
          2200 => x"82",
          2201 => x"74",
          2202 => x"52",
          2203 => x"3f",
          2204 => x"33",
          2205 => x"06",
          2206 => x"33",
          2207 => x"75",
          2208 => x"38",
          2209 => x"7a",
          2210 => x"89",
          2211 => x"74",
          2212 => x"38",
          2213 => x"d9",
          2214 => x"dc",
          2215 => x"84",
          2216 => x"dc",
          2217 => x"06",
          2218 => x"74",
          2219 => x"c8",
          2220 => x"5b",
          2221 => x"7a",
          2222 => x"88",
          2223 => x"11",
          2224 => x"74",
          2225 => x"38",
          2226 => x"a5",
          2227 => x"dc",
          2228 => x"84",
          2229 => x"dc",
          2230 => x"06",
          2231 => x"74",
          2232 => x"c7",
          2233 => x"1b",
          2234 => x"39",
          2235 => x"74",
          2236 => x"bc",
          2237 => x"ca",
          2238 => x"e2",
          2239 => x"2e",
          2240 => x"93",
          2241 => x"d0",
          2242 => x"80",
          2243 => x"74",
          2244 => x"3f",
          2245 => x"7a",
          2246 => x"88",
          2247 => x"11",
          2248 => x"74",
          2249 => x"38",
          2250 => x"c5",
          2251 => x"dc",
          2252 => x"84",
          2253 => x"dc",
          2254 => x"06",
          2255 => x"74",
          2256 => x"c7",
          2257 => x"1b",
          2258 => x"ff",
          2259 => x"39",
          2260 => x"74",
          2261 => x"d8",
          2262 => x"ca",
          2263 => x"8c",
          2264 => x"8d",
          2265 => x"8c",
          2266 => x"ff",
          2267 => x"53",
          2268 => x"51",
          2269 => x"82",
          2270 => x"82",
          2271 => x"52",
          2272 => x"90",
          2273 => x"39",
          2274 => x"33",
          2275 => x"06",
          2276 => x"33",
          2277 => x"74",
          2278 => x"94",
          2279 => x"54",
          2280 => x"88",
          2281 => x"70",
          2282 => x"e2",
          2283 => x"80",
          2284 => x"88",
          2285 => x"80",
          2286 => x"38",
          2287 => x"ed",
          2288 => x"88",
          2289 => x"54",
          2290 => x"88",
          2291 => x"39",
          2292 => x"8d",
          2293 => x"0b",
          2294 => x"34",
          2295 => x"dc",
          2296 => x"0d",
          2297 => x"0d",
          2298 => x"33",
          2299 => x"70",
          2300 => x"38",
          2301 => x"11",
          2302 => x"82",
          2303 => x"83",
          2304 => x"fc",
          2305 => x"9b",
          2306 => x"84",
          2307 => x"33",
          2308 => x"51",
          2309 => x"80",
          2310 => x"84",
          2311 => x"92",
          2312 => x"51",
          2313 => x"80",
          2314 => x"81",
          2315 => x"72",
          2316 => x"92",
          2317 => x"81",
          2318 => x"0b",
          2319 => x"8c",
          2320 => x"71",
          2321 => x"06",
          2322 => x"80",
          2323 => x"87",
          2324 => x"08",
          2325 => x"38",
          2326 => x"80",
          2327 => x"71",
          2328 => x"c0",
          2329 => x"51",
          2330 => x"87",
          2331 => x"89",
          2332 => x"82",
          2333 => x"33",
          2334 => x"8c",
          2335 => x"3d",
          2336 => x"3d",
          2337 => x"64",
          2338 => x"bf",
          2339 => x"40",
          2340 => x"74",
          2341 => x"cd",
          2342 => x"dc",
          2343 => x"7a",
          2344 => x"81",
          2345 => x"72",
          2346 => x"87",
          2347 => x"11",
          2348 => x"8c",
          2349 => x"92",
          2350 => x"5a",
          2351 => x"58",
          2352 => x"c0",
          2353 => x"76",
          2354 => x"76",
          2355 => x"70",
          2356 => x"81",
          2357 => x"54",
          2358 => x"8e",
          2359 => x"52",
          2360 => x"81",
          2361 => x"81",
          2362 => x"74",
          2363 => x"53",
          2364 => x"83",
          2365 => x"78",
          2366 => x"8f",
          2367 => x"2e",
          2368 => x"c0",
          2369 => x"52",
          2370 => x"87",
          2371 => x"08",
          2372 => x"2e",
          2373 => x"84",
          2374 => x"38",
          2375 => x"87",
          2376 => x"15",
          2377 => x"70",
          2378 => x"52",
          2379 => x"ff",
          2380 => x"39",
          2381 => x"81",
          2382 => x"ff",
          2383 => x"57",
          2384 => x"90",
          2385 => x"80",
          2386 => x"71",
          2387 => x"78",
          2388 => x"38",
          2389 => x"80",
          2390 => x"80",
          2391 => x"81",
          2392 => x"72",
          2393 => x"0c",
          2394 => x"04",
          2395 => x"60",
          2396 => x"8c",
          2397 => x"33",
          2398 => x"5b",
          2399 => x"74",
          2400 => x"e1",
          2401 => x"dc",
          2402 => x"79",
          2403 => x"78",
          2404 => x"06",
          2405 => x"77",
          2406 => x"87",
          2407 => x"11",
          2408 => x"8c",
          2409 => x"92",
          2410 => x"59",
          2411 => x"85",
          2412 => x"98",
          2413 => x"7d",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"70",
          2417 => x"53",
          2418 => x"2e",
          2419 => x"70",
          2420 => x"33",
          2421 => x"18",
          2422 => x"2a",
          2423 => x"51",
          2424 => x"2e",
          2425 => x"c0",
          2426 => x"52",
          2427 => x"87",
          2428 => x"08",
          2429 => x"2e",
          2430 => x"84",
          2431 => x"38",
          2432 => x"87",
          2433 => x"15",
          2434 => x"70",
          2435 => x"52",
          2436 => x"ff",
          2437 => x"39",
          2438 => x"81",
          2439 => x"80",
          2440 => x"52",
          2441 => x"90",
          2442 => x"80",
          2443 => x"71",
          2444 => x"7a",
          2445 => x"38",
          2446 => x"80",
          2447 => x"80",
          2448 => x"81",
          2449 => x"72",
          2450 => x"0c",
          2451 => x"04",
          2452 => x"7a",
          2453 => x"a3",
          2454 => x"88",
          2455 => x"33",
          2456 => x"56",
          2457 => x"3f",
          2458 => x"08",
          2459 => x"83",
          2460 => x"fe",
          2461 => x"87",
          2462 => x"0c",
          2463 => x"76",
          2464 => x"38",
          2465 => x"93",
          2466 => x"2b",
          2467 => x"8c",
          2468 => x"71",
          2469 => x"38",
          2470 => x"71",
          2471 => x"c6",
          2472 => x"39",
          2473 => x"81",
          2474 => x"06",
          2475 => x"71",
          2476 => x"38",
          2477 => x"8c",
          2478 => x"e8",
          2479 => x"98",
          2480 => x"71",
          2481 => x"73",
          2482 => x"92",
          2483 => x"72",
          2484 => x"06",
          2485 => x"f7",
          2486 => x"80",
          2487 => x"88",
          2488 => x"0c",
          2489 => x"80",
          2490 => x"56",
          2491 => x"56",
          2492 => x"82",
          2493 => x"88",
          2494 => x"fe",
          2495 => x"81",
          2496 => x"33",
          2497 => x"07",
          2498 => x"0c",
          2499 => x"3d",
          2500 => x"3d",
          2501 => x"11",
          2502 => x"33",
          2503 => x"71",
          2504 => x"81",
          2505 => x"72",
          2506 => x"75",
          2507 => x"82",
          2508 => x"52",
          2509 => x"54",
          2510 => x"0d",
          2511 => x"0d",
          2512 => x"05",
          2513 => x"52",
          2514 => x"70",
          2515 => x"34",
          2516 => x"51",
          2517 => x"83",
          2518 => x"ff",
          2519 => x"75",
          2520 => x"72",
          2521 => x"54",
          2522 => x"2a",
          2523 => x"70",
          2524 => x"34",
          2525 => x"51",
          2526 => x"81",
          2527 => x"70",
          2528 => x"70",
          2529 => x"3d",
          2530 => x"3d",
          2531 => x"77",
          2532 => x"70",
          2533 => x"38",
          2534 => x"05",
          2535 => x"70",
          2536 => x"34",
          2537 => x"eb",
          2538 => x"0d",
          2539 => x"0d",
          2540 => x"54",
          2541 => x"72",
          2542 => x"54",
          2543 => x"51",
          2544 => x"84",
          2545 => x"fc",
          2546 => x"77",
          2547 => x"53",
          2548 => x"05",
          2549 => x"70",
          2550 => x"33",
          2551 => x"ff",
          2552 => x"52",
          2553 => x"2e",
          2554 => x"80",
          2555 => x"71",
          2556 => x"0c",
          2557 => x"04",
          2558 => x"74",
          2559 => x"89",
          2560 => x"2e",
          2561 => x"11",
          2562 => x"52",
          2563 => x"70",
          2564 => x"dc",
          2565 => x"0d",
          2566 => x"82",
          2567 => x"04",
          2568 => x"8c",
          2569 => x"f7",
          2570 => x"56",
          2571 => x"17",
          2572 => x"74",
          2573 => x"d6",
          2574 => x"b0",
          2575 => x"b4",
          2576 => x"81",
          2577 => x"59",
          2578 => x"82",
          2579 => x"7a",
          2580 => x"06",
          2581 => x"8c",
          2582 => x"17",
          2583 => x"08",
          2584 => x"08",
          2585 => x"08",
          2586 => x"74",
          2587 => x"38",
          2588 => x"55",
          2589 => x"09",
          2590 => x"38",
          2591 => x"18",
          2592 => x"81",
          2593 => x"f9",
          2594 => x"39",
          2595 => x"82",
          2596 => x"8b",
          2597 => x"fa",
          2598 => x"7a",
          2599 => x"57",
          2600 => x"08",
          2601 => x"75",
          2602 => x"3f",
          2603 => x"08",
          2604 => x"dc",
          2605 => x"81",
          2606 => x"b4",
          2607 => x"16",
          2608 => x"be",
          2609 => x"dc",
          2610 => x"85",
          2611 => x"81",
          2612 => x"17",
          2613 => x"8c",
          2614 => x"3d",
          2615 => x"3d",
          2616 => x"52",
          2617 => x"3f",
          2618 => x"08",
          2619 => x"dc",
          2620 => x"38",
          2621 => x"74",
          2622 => x"81",
          2623 => x"38",
          2624 => x"59",
          2625 => x"09",
          2626 => x"e3",
          2627 => x"53",
          2628 => x"08",
          2629 => x"70",
          2630 => x"91",
          2631 => x"d5",
          2632 => x"17",
          2633 => x"3f",
          2634 => x"a4",
          2635 => x"51",
          2636 => x"86",
          2637 => x"f2",
          2638 => x"17",
          2639 => x"3f",
          2640 => x"52",
          2641 => x"51",
          2642 => x"8c",
          2643 => x"84",
          2644 => x"fc",
          2645 => x"17",
          2646 => x"70",
          2647 => x"79",
          2648 => x"52",
          2649 => x"51",
          2650 => x"77",
          2651 => x"80",
          2652 => x"81",
          2653 => x"f9",
          2654 => x"8c",
          2655 => x"2e",
          2656 => x"58",
          2657 => x"dc",
          2658 => x"0d",
          2659 => x"0d",
          2660 => x"98",
          2661 => x"05",
          2662 => x"80",
          2663 => x"27",
          2664 => x"14",
          2665 => x"29",
          2666 => x"05",
          2667 => x"82",
          2668 => x"87",
          2669 => x"f9",
          2670 => x"7a",
          2671 => x"54",
          2672 => x"27",
          2673 => x"76",
          2674 => x"27",
          2675 => x"ff",
          2676 => x"58",
          2677 => x"80",
          2678 => x"82",
          2679 => x"72",
          2680 => x"38",
          2681 => x"72",
          2682 => x"8e",
          2683 => x"39",
          2684 => x"17",
          2685 => x"a4",
          2686 => x"53",
          2687 => x"fd",
          2688 => x"8c",
          2689 => x"9f",
          2690 => x"ff",
          2691 => x"11",
          2692 => x"70",
          2693 => x"18",
          2694 => x"76",
          2695 => x"53",
          2696 => x"82",
          2697 => x"80",
          2698 => x"83",
          2699 => x"b4",
          2700 => x"88",
          2701 => x"79",
          2702 => x"84",
          2703 => x"58",
          2704 => x"80",
          2705 => x"9f",
          2706 => x"80",
          2707 => x"88",
          2708 => x"08",
          2709 => x"51",
          2710 => x"82",
          2711 => x"80",
          2712 => x"10",
          2713 => x"74",
          2714 => x"51",
          2715 => x"82",
          2716 => x"83",
          2717 => x"58",
          2718 => x"87",
          2719 => x"08",
          2720 => x"51",
          2721 => x"82",
          2722 => x"9b",
          2723 => x"2b",
          2724 => x"74",
          2725 => x"51",
          2726 => x"82",
          2727 => x"f0",
          2728 => x"83",
          2729 => x"77",
          2730 => x"0c",
          2731 => x"04",
          2732 => x"7a",
          2733 => x"58",
          2734 => x"81",
          2735 => x"9e",
          2736 => x"17",
          2737 => x"96",
          2738 => x"53",
          2739 => x"81",
          2740 => x"79",
          2741 => x"72",
          2742 => x"38",
          2743 => x"72",
          2744 => x"b8",
          2745 => x"39",
          2746 => x"17",
          2747 => x"a4",
          2748 => x"53",
          2749 => x"fb",
          2750 => x"8c",
          2751 => x"82",
          2752 => x"81",
          2753 => x"83",
          2754 => x"b4",
          2755 => x"78",
          2756 => x"56",
          2757 => x"76",
          2758 => x"38",
          2759 => x"9f",
          2760 => x"33",
          2761 => x"07",
          2762 => x"74",
          2763 => x"83",
          2764 => x"89",
          2765 => x"08",
          2766 => x"51",
          2767 => x"82",
          2768 => x"59",
          2769 => x"08",
          2770 => x"74",
          2771 => x"16",
          2772 => x"84",
          2773 => x"76",
          2774 => x"88",
          2775 => x"81",
          2776 => x"8f",
          2777 => x"53",
          2778 => x"80",
          2779 => x"88",
          2780 => x"08",
          2781 => x"51",
          2782 => x"82",
          2783 => x"59",
          2784 => x"08",
          2785 => x"77",
          2786 => x"06",
          2787 => x"83",
          2788 => x"05",
          2789 => x"f7",
          2790 => x"39",
          2791 => x"a4",
          2792 => x"52",
          2793 => x"ef",
          2794 => x"dc",
          2795 => x"8c",
          2796 => x"38",
          2797 => x"06",
          2798 => x"83",
          2799 => x"18",
          2800 => x"54",
          2801 => x"f6",
          2802 => x"8c",
          2803 => x"0a",
          2804 => x"52",
          2805 => x"83",
          2806 => x"83",
          2807 => x"82",
          2808 => x"8a",
          2809 => x"f8",
          2810 => x"7c",
          2811 => x"59",
          2812 => x"81",
          2813 => x"38",
          2814 => x"08",
          2815 => x"73",
          2816 => x"38",
          2817 => x"52",
          2818 => x"a4",
          2819 => x"dc",
          2820 => x"8c",
          2821 => x"f2",
          2822 => x"82",
          2823 => x"39",
          2824 => x"e6",
          2825 => x"dc",
          2826 => x"de",
          2827 => x"78",
          2828 => x"3f",
          2829 => x"08",
          2830 => x"dc",
          2831 => x"80",
          2832 => x"8c",
          2833 => x"2e",
          2834 => x"8c",
          2835 => x"2e",
          2836 => x"53",
          2837 => x"51",
          2838 => x"82",
          2839 => x"c5",
          2840 => x"08",
          2841 => x"18",
          2842 => x"57",
          2843 => x"90",
          2844 => x"90",
          2845 => x"16",
          2846 => x"54",
          2847 => x"34",
          2848 => x"78",
          2849 => x"38",
          2850 => x"82",
          2851 => x"8a",
          2852 => x"f6",
          2853 => x"7e",
          2854 => x"5b",
          2855 => x"38",
          2856 => x"58",
          2857 => x"88",
          2858 => x"08",
          2859 => x"38",
          2860 => x"39",
          2861 => x"51",
          2862 => x"81",
          2863 => x"8c",
          2864 => x"82",
          2865 => x"8c",
          2866 => x"82",
          2867 => x"ff",
          2868 => x"38",
          2869 => x"82",
          2870 => x"26",
          2871 => x"79",
          2872 => x"08",
          2873 => x"73",
          2874 => x"b9",
          2875 => x"2e",
          2876 => x"80",
          2877 => x"1a",
          2878 => x"08",
          2879 => x"38",
          2880 => x"52",
          2881 => x"af",
          2882 => x"82",
          2883 => x"81",
          2884 => x"06",
          2885 => x"8c",
          2886 => x"82",
          2887 => x"09",
          2888 => x"72",
          2889 => x"70",
          2890 => x"8c",
          2891 => x"51",
          2892 => x"73",
          2893 => x"82",
          2894 => x"80",
          2895 => x"8c",
          2896 => x"81",
          2897 => x"38",
          2898 => x"08",
          2899 => x"73",
          2900 => x"75",
          2901 => x"77",
          2902 => x"56",
          2903 => x"76",
          2904 => x"82",
          2905 => x"26",
          2906 => x"75",
          2907 => x"f8",
          2908 => x"8c",
          2909 => x"2e",
          2910 => x"59",
          2911 => x"08",
          2912 => x"81",
          2913 => x"82",
          2914 => x"59",
          2915 => x"08",
          2916 => x"70",
          2917 => x"25",
          2918 => x"51",
          2919 => x"73",
          2920 => x"75",
          2921 => x"81",
          2922 => x"38",
          2923 => x"f5",
          2924 => x"75",
          2925 => x"f9",
          2926 => x"8c",
          2927 => x"8c",
          2928 => x"70",
          2929 => x"08",
          2930 => x"51",
          2931 => x"80",
          2932 => x"73",
          2933 => x"38",
          2934 => x"52",
          2935 => x"d0",
          2936 => x"dc",
          2937 => x"a5",
          2938 => x"18",
          2939 => x"08",
          2940 => x"18",
          2941 => x"74",
          2942 => x"38",
          2943 => x"18",
          2944 => x"33",
          2945 => x"73",
          2946 => x"97",
          2947 => x"74",
          2948 => x"38",
          2949 => x"55",
          2950 => x"8c",
          2951 => x"85",
          2952 => x"75",
          2953 => x"8c",
          2954 => x"3d",
          2955 => x"3d",
          2956 => x"52",
          2957 => x"3f",
          2958 => x"08",
          2959 => x"82",
          2960 => x"80",
          2961 => x"52",
          2962 => x"c1",
          2963 => x"dc",
          2964 => x"dc",
          2965 => x"0c",
          2966 => x"53",
          2967 => x"15",
          2968 => x"f2",
          2969 => x"56",
          2970 => x"16",
          2971 => x"22",
          2972 => x"27",
          2973 => x"54",
          2974 => x"76",
          2975 => x"33",
          2976 => x"3f",
          2977 => x"08",
          2978 => x"38",
          2979 => x"76",
          2980 => x"70",
          2981 => x"9f",
          2982 => x"56",
          2983 => x"8c",
          2984 => x"3d",
          2985 => x"3d",
          2986 => x"71",
          2987 => x"57",
          2988 => x"0a",
          2989 => x"38",
          2990 => x"53",
          2991 => x"38",
          2992 => x"0c",
          2993 => x"54",
          2994 => x"75",
          2995 => x"73",
          2996 => x"a8",
          2997 => x"73",
          2998 => x"85",
          2999 => x"0b",
          3000 => x"5a",
          3001 => x"27",
          3002 => x"a8",
          3003 => x"18",
          3004 => x"39",
          3005 => x"70",
          3006 => x"58",
          3007 => x"b2",
          3008 => x"76",
          3009 => x"3f",
          3010 => x"08",
          3011 => x"dc",
          3012 => x"bd",
          3013 => x"82",
          3014 => x"27",
          3015 => x"16",
          3016 => x"dc",
          3017 => x"38",
          3018 => x"39",
          3019 => x"55",
          3020 => x"52",
          3021 => x"d5",
          3022 => x"dc",
          3023 => x"0c",
          3024 => x"0c",
          3025 => x"53",
          3026 => x"80",
          3027 => x"85",
          3028 => x"94",
          3029 => x"2a",
          3030 => x"0c",
          3031 => x"06",
          3032 => x"9c",
          3033 => x"58",
          3034 => x"dc",
          3035 => x"0d",
          3036 => x"0d",
          3037 => x"90",
          3038 => x"05",
          3039 => x"f0",
          3040 => x"27",
          3041 => x"0b",
          3042 => x"98",
          3043 => x"84",
          3044 => x"2e",
          3045 => x"76",
          3046 => x"58",
          3047 => x"38",
          3048 => x"15",
          3049 => x"08",
          3050 => x"38",
          3051 => x"88",
          3052 => x"53",
          3053 => x"81",
          3054 => x"c0",
          3055 => x"22",
          3056 => x"89",
          3057 => x"72",
          3058 => x"74",
          3059 => x"f3",
          3060 => x"8c",
          3061 => x"82",
          3062 => x"82",
          3063 => x"27",
          3064 => x"81",
          3065 => x"dc",
          3066 => x"80",
          3067 => x"16",
          3068 => x"dc",
          3069 => x"ca",
          3070 => x"38",
          3071 => x"0c",
          3072 => x"dd",
          3073 => x"08",
          3074 => x"f9",
          3075 => x"8c",
          3076 => x"87",
          3077 => x"dc",
          3078 => x"80",
          3079 => x"55",
          3080 => x"08",
          3081 => x"38",
          3082 => x"8c",
          3083 => x"2e",
          3084 => x"8c",
          3085 => x"75",
          3086 => x"3f",
          3087 => x"08",
          3088 => x"94",
          3089 => x"52",
          3090 => x"c1",
          3091 => x"dc",
          3092 => x"0c",
          3093 => x"0c",
          3094 => x"05",
          3095 => x"80",
          3096 => x"8c",
          3097 => x"3d",
          3098 => x"3d",
          3099 => x"71",
          3100 => x"57",
          3101 => x"51",
          3102 => x"82",
          3103 => x"54",
          3104 => x"08",
          3105 => x"82",
          3106 => x"56",
          3107 => x"52",
          3108 => x"83",
          3109 => x"dc",
          3110 => x"8c",
          3111 => x"d2",
          3112 => x"dc",
          3113 => x"08",
          3114 => x"54",
          3115 => x"e5",
          3116 => x"06",
          3117 => x"58",
          3118 => x"08",
          3119 => x"38",
          3120 => x"75",
          3121 => x"80",
          3122 => x"81",
          3123 => x"7a",
          3124 => x"06",
          3125 => x"39",
          3126 => x"08",
          3127 => x"76",
          3128 => x"3f",
          3129 => x"08",
          3130 => x"dc",
          3131 => x"ff",
          3132 => x"84",
          3133 => x"06",
          3134 => x"54",
          3135 => x"dc",
          3136 => x"0d",
          3137 => x"0d",
          3138 => x"52",
          3139 => x"3f",
          3140 => x"08",
          3141 => x"06",
          3142 => x"51",
          3143 => x"83",
          3144 => x"06",
          3145 => x"14",
          3146 => x"3f",
          3147 => x"08",
          3148 => x"07",
          3149 => x"8c",
          3150 => x"3d",
          3151 => x"3d",
          3152 => x"70",
          3153 => x"06",
          3154 => x"53",
          3155 => x"ed",
          3156 => x"33",
          3157 => x"83",
          3158 => x"06",
          3159 => x"90",
          3160 => x"15",
          3161 => x"3f",
          3162 => x"04",
          3163 => x"7b",
          3164 => x"84",
          3165 => x"58",
          3166 => x"80",
          3167 => x"38",
          3168 => x"52",
          3169 => x"8f",
          3170 => x"dc",
          3171 => x"8c",
          3172 => x"f5",
          3173 => x"08",
          3174 => x"53",
          3175 => x"84",
          3176 => x"39",
          3177 => x"70",
          3178 => x"81",
          3179 => x"51",
          3180 => x"16",
          3181 => x"dc",
          3182 => x"81",
          3183 => x"38",
          3184 => x"ae",
          3185 => x"81",
          3186 => x"54",
          3187 => x"2e",
          3188 => x"8f",
          3189 => x"82",
          3190 => x"76",
          3191 => x"54",
          3192 => x"09",
          3193 => x"38",
          3194 => x"7a",
          3195 => x"80",
          3196 => x"fa",
          3197 => x"8c",
          3198 => x"82",
          3199 => x"89",
          3200 => x"08",
          3201 => x"86",
          3202 => x"98",
          3203 => x"82",
          3204 => x"8b",
          3205 => x"fb",
          3206 => x"70",
          3207 => x"81",
          3208 => x"fc",
          3209 => x"8c",
          3210 => x"82",
          3211 => x"b4",
          3212 => x"08",
          3213 => x"ec",
          3214 => x"8c",
          3215 => x"82",
          3216 => x"a0",
          3217 => x"82",
          3218 => x"52",
          3219 => x"51",
          3220 => x"8b",
          3221 => x"52",
          3222 => x"51",
          3223 => x"81",
          3224 => x"34",
          3225 => x"dc",
          3226 => x"0d",
          3227 => x"0d",
          3228 => x"98",
          3229 => x"70",
          3230 => x"ec",
          3231 => x"8c",
          3232 => x"38",
          3233 => x"53",
          3234 => x"81",
          3235 => x"34",
          3236 => x"04",
          3237 => x"78",
          3238 => x"80",
          3239 => x"34",
          3240 => x"80",
          3241 => x"38",
          3242 => x"18",
          3243 => x"9c",
          3244 => x"70",
          3245 => x"56",
          3246 => x"a0",
          3247 => x"71",
          3248 => x"81",
          3249 => x"81",
          3250 => x"89",
          3251 => x"06",
          3252 => x"73",
          3253 => x"55",
          3254 => x"55",
          3255 => x"81",
          3256 => x"81",
          3257 => x"74",
          3258 => x"75",
          3259 => x"52",
          3260 => x"13",
          3261 => x"08",
          3262 => x"33",
          3263 => x"9c",
          3264 => x"11",
          3265 => x"8a",
          3266 => x"dc",
          3267 => x"96",
          3268 => x"e7",
          3269 => x"dc",
          3270 => x"23",
          3271 => x"e7",
          3272 => x"8c",
          3273 => x"17",
          3274 => x"0d",
          3275 => x"0d",
          3276 => x"5e",
          3277 => x"70",
          3278 => x"55",
          3279 => x"83",
          3280 => x"73",
          3281 => x"91",
          3282 => x"2e",
          3283 => x"1d",
          3284 => x"0c",
          3285 => x"15",
          3286 => x"70",
          3287 => x"56",
          3288 => x"09",
          3289 => x"38",
          3290 => x"80",
          3291 => x"30",
          3292 => x"78",
          3293 => x"54",
          3294 => x"73",
          3295 => x"60",
          3296 => x"54",
          3297 => x"96",
          3298 => x"0b",
          3299 => x"80",
          3300 => x"f6",
          3301 => x"8c",
          3302 => x"85",
          3303 => x"3d",
          3304 => x"5c",
          3305 => x"53",
          3306 => x"51",
          3307 => x"80",
          3308 => x"88",
          3309 => x"5c",
          3310 => x"09",
          3311 => x"d4",
          3312 => x"70",
          3313 => x"71",
          3314 => x"30",
          3315 => x"73",
          3316 => x"51",
          3317 => x"57",
          3318 => x"38",
          3319 => x"75",
          3320 => x"17",
          3321 => x"75",
          3322 => x"30",
          3323 => x"51",
          3324 => x"80",
          3325 => x"38",
          3326 => x"87",
          3327 => x"26",
          3328 => x"77",
          3329 => x"a4",
          3330 => x"27",
          3331 => x"a0",
          3332 => x"39",
          3333 => x"33",
          3334 => x"57",
          3335 => x"27",
          3336 => x"75",
          3337 => x"30",
          3338 => x"32",
          3339 => x"80",
          3340 => x"25",
          3341 => x"56",
          3342 => x"80",
          3343 => x"84",
          3344 => x"58",
          3345 => x"70",
          3346 => x"55",
          3347 => x"09",
          3348 => x"38",
          3349 => x"80",
          3350 => x"30",
          3351 => x"77",
          3352 => x"54",
          3353 => x"81",
          3354 => x"ae",
          3355 => x"06",
          3356 => x"54",
          3357 => x"74",
          3358 => x"80",
          3359 => x"7b",
          3360 => x"30",
          3361 => x"70",
          3362 => x"25",
          3363 => x"07",
          3364 => x"51",
          3365 => x"a7",
          3366 => x"8b",
          3367 => x"39",
          3368 => x"54",
          3369 => x"8c",
          3370 => x"ff",
          3371 => x"ec",
          3372 => x"54",
          3373 => x"e1",
          3374 => x"dc",
          3375 => x"b2",
          3376 => x"70",
          3377 => x"71",
          3378 => x"54",
          3379 => x"82",
          3380 => x"80",
          3381 => x"38",
          3382 => x"76",
          3383 => x"df",
          3384 => x"54",
          3385 => x"81",
          3386 => x"55",
          3387 => x"34",
          3388 => x"52",
          3389 => x"51",
          3390 => x"82",
          3391 => x"bf",
          3392 => x"16",
          3393 => x"26",
          3394 => x"16",
          3395 => x"06",
          3396 => x"17",
          3397 => x"34",
          3398 => x"fd",
          3399 => x"19",
          3400 => x"80",
          3401 => x"79",
          3402 => x"81",
          3403 => x"81",
          3404 => x"85",
          3405 => x"54",
          3406 => x"8f",
          3407 => x"86",
          3408 => x"39",
          3409 => x"f3",
          3410 => x"73",
          3411 => x"80",
          3412 => x"52",
          3413 => x"ce",
          3414 => x"dc",
          3415 => x"8c",
          3416 => x"d7",
          3417 => x"08",
          3418 => x"e6",
          3419 => x"8c",
          3420 => x"82",
          3421 => x"80",
          3422 => x"1b",
          3423 => x"55",
          3424 => x"2e",
          3425 => x"8b",
          3426 => x"06",
          3427 => x"1c",
          3428 => x"33",
          3429 => x"70",
          3430 => x"55",
          3431 => x"38",
          3432 => x"52",
          3433 => x"9f",
          3434 => x"dc",
          3435 => x"8b",
          3436 => x"7a",
          3437 => x"3f",
          3438 => x"75",
          3439 => x"57",
          3440 => x"2e",
          3441 => x"84",
          3442 => x"06",
          3443 => x"75",
          3444 => x"81",
          3445 => x"2a",
          3446 => x"73",
          3447 => x"38",
          3448 => x"54",
          3449 => x"fb",
          3450 => x"80",
          3451 => x"34",
          3452 => x"c1",
          3453 => x"06",
          3454 => x"38",
          3455 => x"39",
          3456 => x"70",
          3457 => x"54",
          3458 => x"86",
          3459 => x"84",
          3460 => x"06",
          3461 => x"73",
          3462 => x"38",
          3463 => x"83",
          3464 => x"b4",
          3465 => x"51",
          3466 => x"82",
          3467 => x"88",
          3468 => x"ea",
          3469 => x"8c",
          3470 => x"3d",
          3471 => x"3d",
          3472 => x"ff",
          3473 => x"71",
          3474 => x"5c",
          3475 => x"80",
          3476 => x"38",
          3477 => x"05",
          3478 => x"a0",
          3479 => x"71",
          3480 => x"38",
          3481 => x"71",
          3482 => x"81",
          3483 => x"38",
          3484 => x"11",
          3485 => x"06",
          3486 => x"70",
          3487 => x"38",
          3488 => x"81",
          3489 => x"05",
          3490 => x"76",
          3491 => x"38",
          3492 => x"fa",
          3493 => x"77",
          3494 => x"57",
          3495 => x"05",
          3496 => x"70",
          3497 => x"33",
          3498 => x"53",
          3499 => x"99",
          3500 => x"e0",
          3501 => x"ff",
          3502 => x"ff",
          3503 => x"70",
          3504 => x"38",
          3505 => x"81",
          3506 => x"51",
          3507 => x"9f",
          3508 => x"72",
          3509 => x"81",
          3510 => x"70",
          3511 => x"72",
          3512 => x"32",
          3513 => x"72",
          3514 => x"73",
          3515 => x"53",
          3516 => x"70",
          3517 => x"38",
          3518 => x"19",
          3519 => x"75",
          3520 => x"38",
          3521 => x"83",
          3522 => x"74",
          3523 => x"59",
          3524 => x"39",
          3525 => x"33",
          3526 => x"8c",
          3527 => x"3d",
          3528 => x"3d",
          3529 => x"80",
          3530 => x"34",
          3531 => x"17",
          3532 => x"75",
          3533 => x"3f",
          3534 => x"8c",
          3535 => x"80",
          3536 => x"16",
          3537 => x"3f",
          3538 => x"08",
          3539 => x"06",
          3540 => x"73",
          3541 => x"2e",
          3542 => x"80",
          3543 => x"0b",
          3544 => x"56",
          3545 => x"e9",
          3546 => x"06",
          3547 => x"57",
          3548 => x"32",
          3549 => x"80",
          3550 => x"51",
          3551 => x"8a",
          3552 => x"e8",
          3553 => x"06",
          3554 => x"53",
          3555 => x"52",
          3556 => x"51",
          3557 => x"82",
          3558 => x"55",
          3559 => x"08",
          3560 => x"38",
          3561 => x"fa",
          3562 => x"86",
          3563 => x"97",
          3564 => x"dc",
          3565 => x"8c",
          3566 => x"2e",
          3567 => x"55",
          3568 => x"dc",
          3569 => x"0d",
          3570 => x"0d",
          3571 => x"05",
          3572 => x"33",
          3573 => x"75",
          3574 => x"fc",
          3575 => x"8c",
          3576 => x"8b",
          3577 => x"82",
          3578 => x"24",
          3579 => x"82",
          3580 => x"84",
          3581 => x"8c",
          3582 => x"55",
          3583 => x"73",
          3584 => x"e6",
          3585 => x"0c",
          3586 => x"06",
          3587 => x"57",
          3588 => x"ae",
          3589 => x"33",
          3590 => x"3f",
          3591 => x"08",
          3592 => x"70",
          3593 => x"55",
          3594 => x"76",
          3595 => x"b8",
          3596 => x"2a",
          3597 => x"51",
          3598 => x"72",
          3599 => x"86",
          3600 => x"74",
          3601 => x"15",
          3602 => x"81",
          3603 => x"d7",
          3604 => x"8c",
          3605 => x"ff",
          3606 => x"06",
          3607 => x"56",
          3608 => x"38",
          3609 => x"8f",
          3610 => x"2a",
          3611 => x"51",
          3612 => x"72",
          3613 => x"80",
          3614 => x"52",
          3615 => x"3f",
          3616 => x"08",
          3617 => x"57",
          3618 => x"09",
          3619 => x"e2",
          3620 => x"74",
          3621 => x"56",
          3622 => x"33",
          3623 => x"72",
          3624 => x"38",
          3625 => x"51",
          3626 => x"82",
          3627 => x"57",
          3628 => x"84",
          3629 => x"ff",
          3630 => x"56",
          3631 => x"25",
          3632 => x"0b",
          3633 => x"56",
          3634 => x"05",
          3635 => x"83",
          3636 => x"2e",
          3637 => x"52",
          3638 => x"c6",
          3639 => x"dc",
          3640 => x"06",
          3641 => x"27",
          3642 => x"16",
          3643 => x"27",
          3644 => x"56",
          3645 => x"84",
          3646 => x"56",
          3647 => x"84",
          3648 => x"14",
          3649 => x"3f",
          3650 => x"08",
          3651 => x"06",
          3652 => x"80",
          3653 => x"06",
          3654 => x"80",
          3655 => x"db",
          3656 => x"8c",
          3657 => x"ff",
          3658 => x"77",
          3659 => x"d8",
          3660 => x"de",
          3661 => x"dc",
          3662 => x"9c",
          3663 => x"c4",
          3664 => x"15",
          3665 => x"14",
          3666 => x"70",
          3667 => x"51",
          3668 => x"56",
          3669 => x"84",
          3670 => x"81",
          3671 => x"71",
          3672 => x"16",
          3673 => x"53",
          3674 => x"23",
          3675 => x"8b",
          3676 => x"73",
          3677 => x"80",
          3678 => x"8d",
          3679 => x"39",
          3680 => x"51",
          3681 => x"82",
          3682 => x"53",
          3683 => x"08",
          3684 => x"72",
          3685 => x"8d",
          3686 => x"ce",
          3687 => x"14",
          3688 => x"3f",
          3689 => x"08",
          3690 => x"06",
          3691 => x"38",
          3692 => x"51",
          3693 => x"82",
          3694 => x"55",
          3695 => x"51",
          3696 => x"82",
          3697 => x"83",
          3698 => x"53",
          3699 => x"80",
          3700 => x"38",
          3701 => x"78",
          3702 => x"2a",
          3703 => x"78",
          3704 => x"86",
          3705 => x"22",
          3706 => x"31",
          3707 => x"ee",
          3708 => x"dc",
          3709 => x"8c",
          3710 => x"2e",
          3711 => x"82",
          3712 => x"80",
          3713 => x"f5",
          3714 => x"83",
          3715 => x"ff",
          3716 => x"38",
          3717 => x"9f",
          3718 => x"38",
          3719 => x"39",
          3720 => x"80",
          3721 => x"38",
          3722 => x"98",
          3723 => x"a0",
          3724 => x"1c",
          3725 => x"0c",
          3726 => x"17",
          3727 => x"76",
          3728 => x"81",
          3729 => x"80",
          3730 => x"d9",
          3731 => x"8c",
          3732 => x"ff",
          3733 => x"8d",
          3734 => x"8e",
          3735 => x"8a",
          3736 => x"14",
          3737 => x"3f",
          3738 => x"08",
          3739 => x"74",
          3740 => x"a2",
          3741 => x"79",
          3742 => x"ee",
          3743 => x"a8",
          3744 => x"15",
          3745 => x"2e",
          3746 => x"10",
          3747 => x"2a",
          3748 => x"05",
          3749 => x"ff",
          3750 => x"53",
          3751 => x"9c",
          3752 => x"81",
          3753 => x"0b",
          3754 => x"ff",
          3755 => x"0c",
          3756 => x"84",
          3757 => x"83",
          3758 => x"06",
          3759 => x"80",
          3760 => x"d8",
          3761 => x"8c",
          3762 => x"ff",
          3763 => x"72",
          3764 => x"81",
          3765 => x"38",
          3766 => x"73",
          3767 => x"3f",
          3768 => x"08",
          3769 => x"82",
          3770 => x"84",
          3771 => x"b2",
          3772 => x"87",
          3773 => x"dc",
          3774 => x"ff",
          3775 => x"82",
          3776 => x"09",
          3777 => x"c8",
          3778 => x"51",
          3779 => x"82",
          3780 => x"84",
          3781 => x"d2",
          3782 => x"06",
          3783 => x"98",
          3784 => x"ee",
          3785 => x"dc",
          3786 => x"85",
          3787 => x"09",
          3788 => x"38",
          3789 => x"51",
          3790 => x"82",
          3791 => x"90",
          3792 => x"a0",
          3793 => x"ca",
          3794 => x"dc",
          3795 => x"0c",
          3796 => x"82",
          3797 => x"81",
          3798 => x"82",
          3799 => x"72",
          3800 => x"80",
          3801 => x"0c",
          3802 => x"82",
          3803 => x"90",
          3804 => x"fb",
          3805 => x"54",
          3806 => x"80",
          3807 => x"73",
          3808 => x"80",
          3809 => x"72",
          3810 => x"80",
          3811 => x"86",
          3812 => x"15",
          3813 => x"71",
          3814 => x"81",
          3815 => x"81",
          3816 => x"d0",
          3817 => x"8c",
          3818 => x"06",
          3819 => x"38",
          3820 => x"54",
          3821 => x"80",
          3822 => x"71",
          3823 => x"82",
          3824 => x"87",
          3825 => x"fa",
          3826 => x"ab",
          3827 => x"58",
          3828 => x"05",
          3829 => x"e6",
          3830 => x"80",
          3831 => x"dc",
          3832 => x"38",
          3833 => x"08",
          3834 => x"8d",
          3835 => x"08",
          3836 => x"80",
          3837 => x"80",
          3838 => x"54",
          3839 => x"84",
          3840 => x"34",
          3841 => x"75",
          3842 => x"2e",
          3843 => x"53",
          3844 => x"53",
          3845 => x"f7",
          3846 => x"8c",
          3847 => x"73",
          3848 => x"0c",
          3849 => x"04",
          3850 => x"67",
          3851 => x"80",
          3852 => x"59",
          3853 => x"78",
          3854 => x"c8",
          3855 => x"06",
          3856 => x"3d",
          3857 => x"99",
          3858 => x"52",
          3859 => x"3f",
          3860 => x"08",
          3861 => x"dc",
          3862 => x"38",
          3863 => x"52",
          3864 => x"52",
          3865 => x"3f",
          3866 => x"08",
          3867 => x"dc",
          3868 => x"02",
          3869 => x"33",
          3870 => x"55",
          3871 => x"25",
          3872 => x"55",
          3873 => x"54",
          3874 => x"81",
          3875 => x"80",
          3876 => x"74",
          3877 => x"81",
          3878 => x"75",
          3879 => x"3f",
          3880 => x"08",
          3881 => x"02",
          3882 => x"91",
          3883 => x"81",
          3884 => x"82",
          3885 => x"06",
          3886 => x"80",
          3887 => x"88",
          3888 => x"39",
          3889 => x"58",
          3890 => x"38",
          3891 => x"70",
          3892 => x"54",
          3893 => x"81",
          3894 => x"52",
          3895 => x"a5",
          3896 => x"dc",
          3897 => x"88",
          3898 => x"62",
          3899 => x"d4",
          3900 => x"54",
          3901 => x"15",
          3902 => x"62",
          3903 => x"e8",
          3904 => x"52",
          3905 => x"51",
          3906 => x"7a",
          3907 => x"83",
          3908 => x"80",
          3909 => x"38",
          3910 => x"08",
          3911 => x"53",
          3912 => x"3d",
          3913 => x"dd",
          3914 => x"8c",
          3915 => x"82",
          3916 => x"82",
          3917 => x"39",
          3918 => x"38",
          3919 => x"33",
          3920 => x"70",
          3921 => x"55",
          3922 => x"2e",
          3923 => x"55",
          3924 => x"77",
          3925 => x"81",
          3926 => x"73",
          3927 => x"38",
          3928 => x"54",
          3929 => x"a0",
          3930 => x"82",
          3931 => x"52",
          3932 => x"a3",
          3933 => x"dc",
          3934 => x"18",
          3935 => x"55",
          3936 => x"dc",
          3937 => x"38",
          3938 => x"70",
          3939 => x"54",
          3940 => x"86",
          3941 => x"c0",
          3942 => x"b0",
          3943 => x"1b",
          3944 => x"1b",
          3945 => x"70",
          3946 => x"d9",
          3947 => x"dc",
          3948 => x"dc",
          3949 => x"0c",
          3950 => x"52",
          3951 => x"3f",
          3952 => x"08",
          3953 => x"08",
          3954 => x"77",
          3955 => x"86",
          3956 => x"1a",
          3957 => x"1a",
          3958 => x"91",
          3959 => x"0b",
          3960 => x"80",
          3961 => x"0c",
          3962 => x"70",
          3963 => x"54",
          3964 => x"81",
          3965 => x"8c",
          3966 => x"2e",
          3967 => x"82",
          3968 => x"94",
          3969 => x"17",
          3970 => x"2b",
          3971 => x"57",
          3972 => x"52",
          3973 => x"9f",
          3974 => x"dc",
          3975 => x"8c",
          3976 => x"26",
          3977 => x"55",
          3978 => x"08",
          3979 => x"81",
          3980 => x"79",
          3981 => x"31",
          3982 => x"70",
          3983 => x"25",
          3984 => x"76",
          3985 => x"81",
          3986 => x"55",
          3987 => x"38",
          3988 => x"0c",
          3989 => x"75",
          3990 => x"54",
          3991 => x"a2",
          3992 => x"7a",
          3993 => x"3f",
          3994 => x"08",
          3995 => x"55",
          3996 => x"89",
          3997 => x"dc",
          3998 => x"1a",
          3999 => x"80",
          4000 => x"54",
          4001 => x"dc",
          4002 => x"0d",
          4003 => x"0d",
          4004 => x"64",
          4005 => x"59",
          4006 => x"90",
          4007 => x"52",
          4008 => x"cf",
          4009 => x"dc",
          4010 => x"8c",
          4011 => x"38",
          4012 => x"55",
          4013 => x"86",
          4014 => x"82",
          4015 => x"19",
          4016 => x"55",
          4017 => x"80",
          4018 => x"38",
          4019 => x"0b",
          4020 => x"82",
          4021 => x"39",
          4022 => x"1a",
          4023 => x"82",
          4024 => x"19",
          4025 => x"08",
          4026 => x"7c",
          4027 => x"74",
          4028 => x"2e",
          4029 => x"94",
          4030 => x"83",
          4031 => x"56",
          4032 => x"38",
          4033 => x"22",
          4034 => x"89",
          4035 => x"55",
          4036 => x"75",
          4037 => x"19",
          4038 => x"39",
          4039 => x"52",
          4040 => x"93",
          4041 => x"dc",
          4042 => x"75",
          4043 => x"38",
          4044 => x"ff",
          4045 => x"98",
          4046 => x"19",
          4047 => x"51",
          4048 => x"82",
          4049 => x"80",
          4050 => x"38",
          4051 => x"08",
          4052 => x"2a",
          4053 => x"80",
          4054 => x"38",
          4055 => x"8a",
          4056 => x"5c",
          4057 => x"27",
          4058 => x"7a",
          4059 => x"54",
          4060 => x"52",
          4061 => x"51",
          4062 => x"82",
          4063 => x"fe",
          4064 => x"83",
          4065 => x"56",
          4066 => x"9f",
          4067 => x"08",
          4068 => x"74",
          4069 => x"38",
          4070 => x"b4",
          4071 => x"16",
          4072 => x"89",
          4073 => x"51",
          4074 => x"77",
          4075 => x"b9",
          4076 => x"1a",
          4077 => x"08",
          4078 => x"84",
          4079 => x"57",
          4080 => x"27",
          4081 => x"56",
          4082 => x"52",
          4083 => x"c7",
          4084 => x"dc",
          4085 => x"38",
          4086 => x"19",
          4087 => x"06",
          4088 => x"52",
          4089 => x"a2",
          4090 => x"31",
          4091 => x"7f",
          4092 => x"94",
          4093 => x"94",
          4094 => x"5c",
          4095 => x"80",
          4096 => x"8c",
          4097 => x"3d",
          4098 => x"3d",
          4099 => x"65",
          4100 => x"5d",
          4101 => x"0c",
          4102 => x"05",
          4103 => x"f6",
          4104 => x"8c",
          4105 => x"82",
          4106 => x"8a",
          4107 => x"33",
          4108 => x"2e",
          4109 => x"56",
          4110 => x"90",
          4111 => x"81",
          4112 => x"06",
          4113 => x"87",
          4114 => x"2e",
          4115 => x"95",
          4116 => x"91",
          4117 => x"56",
          4118 => x"81",
          4119 => x"34",
          4120 => x"8e",
          4121 => x"08",
          4122 => x"56",
          4123 => x"84",
          4124 => x"5c",
          4125 => x"82",
          4126 => x"18",
          4127 => x"ff",
          4128 => x"74",
          4129 => x"7e",
          4130 => x"ff",
          4131 => x"2a",
          4132 => x"7a",
          4133 => x"8c",
          4134 => x"08",
          4135 => x"38",
          4136 => x"39",
          4137 => x"52",
          4138 => x"e7",
          4139 => x"dc",
          4140 => x"8c",
          4141 => x"2e",
          4142 => x"74",
          4143 => x"91",
          4144 => x"2e",
          4145 => x"74",
          4146 => x"88",
          4147 => x"38",
          4148 => x"0c",
          4149 => x"15",
          4150 => x"08",
          4151 => x"06",
          4152 => x"51",
          4153 => x"82",
          4154 => x"fe",
          4155 => x"18",
          4156 => x"51",
          4157 => x"82",
          4158 => x"80",
          4159 => x"38",
          4160 => x"08",
          4161 => x"2a",
          4162 => x"80",
          4163 => x"38",
          4164 => x"8a",
          4165 => x"5b",
          4166 => x"27",
          4167 => x"7b",
          4168 => x"54",
          4169 => x"52",
          4170 => x"51",
          4171 => x"82",
          4172 => x"fe",
          4173 => x"b0",
          4174 => x"31",
          4175 => x"79",
          4176 => x"84",
          4177 => x"16",
          4178 => x"89",
          4179 => x"52",
          4180 => x"cc",
          4181 => x"55",
          4182 => x"16",
          4183 => x"2b",
          4184 => x"39",
          4185 => x"94",
          4186 => x"93",
          4187 => x"cd",
          4188 => x"8c",
          4189 => x"e3",
          4190 => x"b0",
          4191 => x"76",
          4192 => x"94",
          4193 => x"ff",
          4194 => x"71",
          4195 => x"7b",
          4196 => x"38",
          4197 => x"18",
          4198 => x"51",
          4199 => x"82",
          4200 => x"fd",
          4201 => x"53",
          4202 => x"18",
          4203 => x"06",
          4204 => x"51",
          4205 => x"7e",
          4206 => x"83",
          4207 => x"76",
          4208 => x"17",
          4209 => x"1e",
          4210 => x"18",
          4211 => x"0c",
          4212 => x"58",
          4213 => x"74",
          4214 => x"38",
          4215 => x"8c",
          4216 => x"90",
          4217 => x"33",
          4218 => x"55",
          4219 => x"34",
          4220 => x"82",
          4221 => x"90",
          4222 => x"f8",
          4223 => x"8b",
          4224 => x"53",
          4225 => x"f2",
          4226 => x"8c",
          4227 => x"82",
          4228 => x"80",
          4229 => x"16",
          4230 => x"2a",
          4231 => x"51",
          4232 => x"80",
          4233 => x"38",
          4234 => x"52",
          4235 => x"e7",
          4236 => x"dc",
          4237 => x"8c",
          4238 => x"d4",
          4239 => x"08",
          4240 => x"a0",
          4241 => x"73",
          4242 => x"88",
          4243 => x"74",
          4244 => x"51",
          4245 => x"8c",
          4246 => x"9c",
          4247 => x"fb",
          4248 => x"b2",
          4249 => x"15",
          4250 => x"3f",
          4251 => x"15",
          4252 => x"3f",
          4253 => x"0b",
          4254 => x"78",
          4255 => x"3f",
          4256 => x"08",
          4257 => x"81",
          4258 => x"57",
          4259 => x"34",
          4260 => x"dc",
          4261 => x"0d",
          4262 => x"0d",
          4263 => x"54",
          4264 => x"82",
          4265 => x"53",
          4266 => x"08",
          4267 => x"3d",
          4268 => x"73",
          4269 => x"3f",
          4270 => x"08",
          4271 => x"dc",
          4272 => x"82",
          4273 => x"74",
          4274 => x"8c",
          4275 => x"3d",
          4276 => x"3d",
          4277 => x"51",
          4278 => x"8b",
          4279 => x"82",
          4280 => x"24",
          4281 => x"8c",
          4282 => x"8d",
          4283 => x"52",
          4284 => x"dc",
          4285 => x"0d",
          4286 => x"0d",
          4287 => x"3d",
          4288 => x"94",
          4289 => x"c1",
          4290 => x"dc",
          4291 => x"8c",
          4292 => x"e0",
          4293 => x"63",
          4294 => x"d4",
          4295 => x"8d",
          4296 => x"dc",
          4297 => x"8c",
          4298 => x"38",
          4299 => x"05",
          4300 => x"2b",
          4301 => x"80",
          4302 => x"76",
          4303 => x"0c",
          4304 => x"02",
          4305 => x"70",
          4306 => x"81",
          4307 => x"56",
          4308 => x"9e",
          4309 => x"53",
          4310 => x"db",
          4311 => x"8c",
          4312 => x"15",
          4313 => x"82",
          4314 => x"84",
          4315 => x"06",
          4316 => x"55",
          4317 => x"dc",
          4318 => x"0d",
          4319 => x"0d",
          4320 => x"5b",
          4321 => x"80",
          4322 => x"ff",
          4323 => x"9f",
          4324 => x"b5",
          4325 => x"dc",
          4326 => x"8c",
          4327 => x"fc",
          4328 => x"7a",
          4329 => x"08",
          4330 => x"64",
          4331 => x"2e",
          4332 => x"a0",
          4333 => x"70",
          4334 => x"ea",
          4335 => x"dc",
          4336 => x"8c",
          4337 => x"d4",
          4338 => x"7b",
          4339 => x"3f",
          4340 => x"08",
          4341 => x"dc",
          4342 => x"38",
          4343 => x"51",
          4344 => x"82",
          4345 => x"45",
          4346 => x"51",
          4347 => x"82",
          4348 => x"57",
          4349 => x"08",
          4350 => x"80",
          4351 => x"da",
          4352 => x"8c",
          4353 => x"82",
          4354 => x"a4",
          4355 => x"7b",
          4356 => x"3f",
          4357 => x"dc",
          4358 => x"38",
          4359 => x"51",
          4360 => x"82",
          4361 => x"57",
          4362 => x"08",
          4363 => x"38",
          4364 => x"09",
          4365 => x"38",
          4366 => x"e0",
          4367 => x"dc",
          4368 => x"ff",
          4369 => x"74",
          4370 => x"3f",
          4371 => x"78",
          4372 => x"33",
          4373 => x"56",
          4374 => x"91",
          4375 => x"05",
          4376 => x"81",
          4377 => x"56",
          4378 => x"f5",
          4379 => x"54",
          4380 => x"81",
          4381 => x"80",
          4382 => x"78",
          4383 => x"55",
          4384 => x"11",
          4385 => x"18",
          4386 => x"58",
          4387 => x"34",
          4388 => x"ff",
          4389 => x"55",
          4390 => x"34",
          4391 => x"77",
          4392 => x"81",
          4393 => x"ff",
          4394 => x"55",
          4395 => x"34",
          4396 => x"8d",
          4397 => x"84",
          4398 => x"dc",
          4399 => x"70",
          4400 => x"56",
          4401 => x"76",
          4402 => x"81",
          4403 => x"70",
          4404 => x"56",
          4405 => x"82",
          4406 => x"78",
          4407 => x"80",
          4408 => x"27",
          4409 => x"19",
          4410 => x"7a",
          4411 => x"5c",
          4412 => x"55",
          4413 => x"7a",
          4414 => x"5c",
          4415 => x"2e",
          4416 => x"85",
          4417 => x"94",
          4418 => x"81",
          4419 => x"73",
          4420 => x"81",
          4421 => x"7a",
          4422 => x"38",
          4423 => x"76",
          4424 => x"0c",
          4425 => x"04",
          4426 => x"7b",
          4427 => x"fc",
          4428 => x"53",
          4429 => x"bb",
          4430 => x"dc",
          4431 => x"8c",
          4432 => x"fa",
          4433 => x"33",
          4434 => x"f2",
          4435 => x"08",
          4436 => x"27",
          4437 => x"15",
          4438 => x"2a",
          4439 => x"51",
          4440 => x"83",
          4441 => x"94",
          4442 => x"80",
          4443 => x"0c",
          4444 => x"2e",
          4445 => x"79",
          4446 => x"70",
          4447 => x"51",
          4448 => x"2e",
          4449 => x"52",
          4450 => x"fe",
          4451 => x"82",
          4452 => x"ff",
          4453 => x"70",
          4454 => x"fe",
          4455 => x"82",
          4456 => x"73",
          4457 => x"76",
          4458 => x"06",
          4459 => x"0c",
          4460 => x"98",
          4461 => x"58",
          4462 => x"39",
          4463 => x"54",
          4464 => x"73",
          4465 => x"cd",
          4466 => x"8c",
          4467 => x"82",
          4468 => x"81",
          4469 => x"38",
          4470 => x"08",
          4471 => x"9b",
          4472 => x"dc",
          4473 => x"0c",
          4474 => x"0c",
          4475 => x"81",
          4476 => x"76",
          4477 => x"38",
          4478 => x"94",
          4479 => x"94",
          4480 => x"16",
          4481 => x"2a",
          4482 => x"51",
          4483 => x"72",
          4484 => x"38",
          4485 => x"51",
          4486 => x"82",
          4487 => x"54",
          4488 => x"08",
          4489 => x"8c",
          4490 => x"a7",
          4491 => x"74",
          4492 => x"3f",
          4493 => x"08",
          4494 => x"2e",
          4495 => x"74",
          4496 => x"79",
          4497 => x"14",
          4498 => x"38",
          4499 => x"0c",
          4500 => x"94",
          4501 => x"94",
          4502 => x"83",
          4503 => x"72",
          4504 => x"38",
          4505 => x"51",
          4506 => x"82",
          4507 => x"94",
          4508 => x"91",
          4509 => x"53",
          4510 => x"81",
          4511 => x"34",
          4512 => x"39",
          4513 => x"82",
          4514 => x"05",
          4515 => x"08",
          4516 => x"08",
          4517 => x"38",
          4518 => x"0c",
          4519 => x"80",
          4520 => x"72",
          4521 => x"73",
          4522 => x"53",
          4523 => x"8c",
          4524 => x"16",
          4525 => x"38",
          4526 => x"0c",
          4527 => x"82",
          4528 => x"8b",
          4529 => x"f9",
          4530 => x"56",
          4531 => x"80",
          4532 => x"38",
          4533 => x"3d",
          4534 => x"8a",
          4535 => x"51",
          4536 => x"82",
          4537 => x"55",
          4538 => x"08",
          4539 => x"77",
          4540 => x"52",
          4541 => x"b5",
          4542 => x"dc",
          4543 => x"8c",
          4544 => x"c3",
          4545 => x"33",
          4546 => x"55",
          4547 => x"24",
          4548 => x"16",
          4549 => x"2a",
          4550 => x"51",
          4551 => x"80",
          4552 => x"9c",
          4553 => x"77",
          4554 => x"3f",
          4555 => x"08",
          4556 => x"77",
          4557 => x"22",
          4558 => x"74",
          4559 => x"ce",
          4560 => x"8c",
          4561 => x"74",
          4562 => x"81",
          4563 => x"85",
          4564 => x"74",
          4565 => x"38",
          4566 => x"74",
          4567 => x"8c",
          4568 => x"3d",
          4569 => x"3d",
          4570 => x"3d",
          4571 => x"70",
          4572 => x"ff",
          4573 => x"dc",
          4574 => x"82",
          4575 => x"73",
          4576 => x"0d",
          4577 => x"0d",
          4578 => x"3d",
          4579 => x"71",
          4580 => x"e7",
          4581 => x"8c",
          4582 => x"82",
          4583 => x"80",
          4584 => x"93",
          4585 => x"dc",
          4586 => x"51",
          4587 => x"82",
          4588 => x"53",
          4589 => x"82",
          4590 => x"52",
          4591 => x"ac",
          4592 => x"dc",
          4593 => x"8c",
          4594 => x"2e",
          4595 => x"85",
          4596 => x"87",
          4597 => x"dc",
          4598 => x"74",
          4599 => x"d5",
          4600 => x"52",
          4601 => x"89",
          4602 => x"dc",
          4603 => x"70",
          4604 => x"07",
          4605 => x"82",
          4606 => x"06",
          4607 => x"54",
          4608 => x"dc",
          4609 => x"0d",
          4610 => x"0d",
          4611 => x"53",
          4612 => x"53",
          4613 => x"56",
          4614 => x"82",
          4615 => x"55",
          4616 => x"08",
          4617 => x"52",
          4618 => x"81",
          4619 => x"dc",
          4620 => x"8c",
          4621 => x"38",
          4622 => x"05",
          4623 => x"2b",
          4624 => x"80",
          4625 => x"86",
          4626 => x"76",
          4627 => x"38",
          4628 => x"51",
          4629 => x"74",
          4630 => x"0c",
          4631 => x"04",
          4632 => x"63",
          4633 => x"80",
          4634 => x"ec",
          4635 => x"3d",
          4636 => x"3f",
          4637 => x"08",
          4638 => x"dc",
          4639 => x"38",
          4640 => x"73",
          4641 => x"08",
          4642 => x"13",
          4643 => x"58",
          4644 => x"26",
          4645 => x"7c",
          4646 => x"39",
          4647 => x"cc",
          4648 => x"81",
          4649 => x"8c",
          4650 => x"33",
          4651 => x"81",
          4652 => x"06",
          4653 => x"75",
          4654 => x"52",
          4655 => x"05",
          4656 => x"3f",
          4657 => x"08",
          4658 => x"38",
          4659 => x"08",
          4660 => x"38",
          4661 => x"08",
          4662 => x"8c",
          4663 => x"80",
          4664 => x"81",
          4665 => x"59",
          4666 => x"14",
          4667 => x"ca",
          4668 => x"39",
          4669 => x"82",
          4670 => x"57",
          4671 => x"38",
          4672 => x"18",
          4673 => x"ff",
          4674 => x"82",
          4675 => x"5b",
          4676 => x"08",
          4677 => x"7c",
          4678 => x"12",
          4679 => x"52",
          4680 => x"82",
          4681 => x"06",
          4682 => x"14",
          4683 => x"cb",
          4684 => x"dc",
          4685 => x"ff",
          4686 => x"70",
          4687 => x"82",
          4688 => x"51",
          4689 => x"b4",
          4690 => x"bb",
          4691 => x"8c",
          4692 => x"0a",
          4693 => x"70",
          4694 => x"84",
          4695 => x"51",
          4696 => x"ff",
          4697 => x"56",
          4698 => x"38",
          4699 => x"7c",
          4700 => x"0c",
          4701 => x"81",
          4702 => x"74",
          4703 => x"7a",
          4704 => x"0c",
          4705 => x"04",
          4706 => x"79",
          4707 => x"05",
          4708 => x"57",
          4709 => x"82",
          4710 => x"56",
          4711 => x"08",
          4712 => x"91",
          4713 => x"75",
          4714 => x"90",
          4715 => x"81",
          4716 => x"06",
          4717 => x"87",
          4718 => x"2e",
          4719 => x"94",
          4720 => x"73",
          4721 => x"27",
          4722 => x"73",
          4723 => x"8c",
          4724 => x"88",
          4725 => x"76",
          4726 => x"3f",
          4727 => x"08",
          4728 => x"0c",
          4729 => x"39",
          4730 => x"52",
          4731 => x"bf",
          4732 => x"8c",
          4733 => x"2e",
          4734 => x"83",
          4735 => x"82",
          4736 => x"81",
          4737 => x"06",
          4738 => x"56",
          4739 => x"a0",
          4740 => x"82",
          4741 => x"98",
          4742 => x"94",
          4743 => x"08",
          4744 => x"dc",
          4745 => x"51",
          4746 => x"82",
          4747 => x"56",
          4748 => x"8c",
          4749 => x"17",
          4750 => x"07",
          4751 => x"18",
          4752 => x"2e",
          4753 => x"91",
          4754 => x"55",
          4755 => x"dc",
          4756 => x"0d",
          4757 => x"0d",
          4758 => x"3d",
          4759 => x"52",
          4760 => x"da",
          4761 => x"8c",
          4762 => x"82",
          4763 => x"81",
          4764 => x"45",
          4765 => x"52",
          4766 => x"52",
          4767 => x"3f",
          4768 => x"08",
          4769 => x"dc",
          4770 => x"38",
          4771 => x"05",
          4772 => x"2a",
          4773 => x"51",
          4774 => x"55",
          4775 => x"38",
          4776 => x"54",
          4777 => x"81",
          4778 => x"80",
          4779 => x"70",
          4780 => x"54",
          4781 => x"81",
          4782 => x"52",
          4783 => x"c5",
          4784 => x"dc",
          4785 => x"2a",
          4786 => x"51",
          4787 => x"80",
          4788 => x"38",
          4789 => x"8c",
          4790 => x"15",
          4791 => x"86",
          4792 => x"82",
          4793 => x"5c",
          4794 => x"3d",
          4795 => x"c7",
          4796 => x"8c",
          4797 => x"82",
          4798 => x"80",
          4799 => x"8c",
          4800 => x"73",
          4801 => x"3f",
          4802 => x"08",
          4803 => x"dc",
          4804 => x"87",
          4805 => x"39",
          4806 => x"08",
          4807 => x"38",
          4808 => x"08",
          4809 => x"77",
          4810 => x"3f",
          4811 => x"08",
          4812 => x"08",
          4813 => x"8c",
          4814 => x"80",
          4815 => x"55",
          4816 => x"94",
          4817 => x"2e",
          4818 => x"53",
          4819 => x"51",
          4820 => x"82",
          4821 => x"55",
          4822 => x"78",
          4823 => x"fe",
          4824 => x"dc",
          4825 => x"82",
          4826 => x"a0",
          4827 => x"e9",
          4828 => x"53",
          4829 => x"05",
          4830 => x"51",
          4831 => x"82",
          4832 => x"54",
          4833 => x"08",
          4834 => x"78",
          4835 => x"8e",
          4836 => x"58",
          4837 => x"82",
          4838 => x"54",
          4839 => x"08",
          4840 => x"54",
          4841 => x"82",
          4842 => x"84",
          4843 => x"06",
          4844 => x"02",
          4845 => x"33",
          4846 => x"81",
          4847 => x"86",
          4848 => x"f6",
          4849 => x"74",
          4850 => x"70",
          4851 => x"c3",
          4852 => x"dc",
          4853 => x"56",
          4854 => x"08",
          4855 => x"54",
          4856 => x"08",
          4857 => x"81",
          4858 => x"82",
          4859 => x"dc",
          4860 => x"09",
          4861 => x"38",
          4862 => x"b4",
          4863 => x"b0",
          4864 => x"dc",
          4865 => x"51",
          4866 => x"82",
          4867 => x"54",
          4868 => x"08",
          4869 => x"8b",
          4870 => x"b4",
          4871 => x"b7",
          4872 => x"54",
          4873 => x"15",
          4874 => x"90",
          4875 => x"34",
          4876 => x"0a",
          4877 => x"19",
          4878 => x"9f",
          4879 => x"78",
          4880 => x"51",
          4881 => x"a0",
          4882 => x"11",
          4883 => x"05",
          4884 => x"b6",
          4885 => x"ae",
          4886 => x"15",
          4887 => x"78",
          4888 => x"53",
          4889 => x"3f",
          4890 => x"0b",
          4891 => x"77",
          4892 => x"3f",
          4893 => x"08",
          4894 => x"dc",
          4895 => x"82",
          4896 => x"52",
          4897 => x"51",
          4898 => x"3f",
          4899 => x"52",
          4900 => x"aa",
          4901 => x"90",
          4902 => x"34",
          4903 => x"0b",
          4904 => x"78",
          4905 => x"b6",
          4906 => x"dc",
          4907 => x"39",
          4908 => x"52",
          4909 => x"be",
          4910 => x"82",
          4911 => x"99",
          4912 => x"da",
          4913 => x"3d",
          4914 => x"d2",
          4915 => x"53",
          4916 => x"84",
          4917 => x"3d",
          4918 => x"3f",
          4919 => x"08",
          4920 => x"dc",
          4921 => x"38",
          4922 => x"3d",
          4923 => x"3d",
          4924 => x"cc",
          4925 => x"8c",
          4926 => x"82",
          4927 => x"82",
          4928 => x"81",
          4929 => x"81",
          4930 => x"86",
          4931 => x"aa",
          4932 => x"a4",
          4933 => x"a8",
          4934 => x"05",
          4935 => x"ea",
          4936 => x"77",
          4937 => x"70",
          4938 => x"b4",
          4939 => x"3d",
          4940 => x"51",
          4941 => x"82",
          4942 => x"55",
          4943 => x"08",
          4944 => x"6f",
          4945 => x"06",
          4946 => x"a2",
          4947 => x"92",
          4948 => x"81",
          4949 => x"8c",
          4950 => x"2e",
          4951 => x"81",
          4952 => x"51",
          4953 => x"82",
          4954 => x"55",
          4955 => x"08",
          4956 => x"68",
          4957 => x"a8",
          4958 => x"05",
          4959 => x"51",
          4960 => x"3f",
          4961 => x"33",
          4962 => x"8b",
          4963 => x"84",
          4964 => x"06",
          4965 => x"73",
          4966 => x"a0",
          4967 => x"8b",
          4968 => x"54",
          4969 => x"15",
          4970 => x"33",
          4971 => x"70",
          4972 => x"55",
          4973 => x"2e",
          4974 => x"6e",
          4975 => x"df",
          4976 => x"78",
          4977 => x"3f",
          4978 => x"08",
          4979 => x"ff",
          4980 => x"82",
          4981 => x"dc",
          4982 => x"80",
          4983 => x"8c",
          4984 => x"78",
          4985 => x"af",
          4986 => x"dc",
          4987 => x"d4",
          4988 => x"55",
          4989 => x"08",
          4990 => x"81",
          4991 => x"73",
          4992 => x"81",
          4993 => x"63",
          4994 => x"76",
          4995 => x"3f",
          4996 => x"0b",
          4997 => x"87",
          4998 => x"dc",
          4999 => x"77",
          5000 => x"3f",
          5001 => x"08",
          5002 => x"dc",
          5003 => x"78",
          5004 => x"aa",
          5005 => x"dc",
          5006 => x"82",
          5007 => x"a8",
          5008 => x"ed",
          5009 => x"80",
          5010 => x"02",
          5011 => x"df",
          5012 => x"57",
          5013 => x"3d",
          5014 => x"96",
          5015 => x"e9",
          5016 => x"dc",
          5017 => x"8c",
          5018 => x"cf",
          5019 => x"65",
          5020 => x"d4",
          5021 => x"b5",
          5022 => x"dc",
          5023 => x"8c",
          5024 => x"38",
          5025 => x"05",
          5026 => x"06",
          5027 => x"73",
          5028 => x"a7",
          5029 => x"09",
          5030 => x"71",
          5031 => x"06",
          5032 => x"55",
          5033 => x"15",
          5034 => x"81",
          5035 => x"34",
          5036 => x"b4",
          5037 => x"8c",
          5038 => x"74",
          5039 => x"0c",
          5040 => x"04",
          5041 => x"64",
          5042 => x"93",
          5043 => x"52",
          5044 => x"d1",
          5045 => x"8c",
          5046 => x"82",
          5047 => x"80",
          5048 => x"58",
          5049 => x"3d",
          5050 => x"c8",
          5051 => x"8c",
          5052 => x"82",
          5053 => x"b4",
          5054 => x"c7",
          5055 => x"a0",
          5056 => x"55",
          5057 => x"84",
          5058 => x"17",
          5059 => x"2b",
          5060 => x"96",
          5061 => x"b0",
          5062 => x"54",
          5063 => x"15",
          5064 => x"ff",
          5065 => x"82",
          5066 => x"55",
          5067 => x"dc",
          5068 => x"0d",
          5069 => x"0d",
          5070 => x"5a",
          5071 => x"3d",
          5072 => x"99",
          5073 => x"81",
          5074 => x"dc",
          5075 => x"dc",
          5076 => x"82",
          5077 => x"07",
          5078 => x"55",
          5079 => x"2e",
          5080 => x"81",
          5081 => x"55",
          5082 => x"2e",
          5083 => x"7b",
          5084 => x"80",
          5085 => x"70",
          5086 => x"be",
          5087 => x"8c",
          5088 => x"82",
          5089 => x"80",
          5090 => x"52",
          5091 => x"dc",
          5092 => x"dc",
          5093 => x"8c",
          5094 => x"38",
          5095 => x"08",
          5096 => x"08",
          5097 => x"56",
          5098 => x"19",
          5099 => x"59",
          5100 => x"74",
          5101 => x"56",
          5102 => x"ec",
          5103 => x"75",
          5104 => x"74",
          5105 => x"2e",
          5106 => x"16",
          5107 => x"33",
          5108 => x"73",
          5109 => x"38",
          5110 => x"84",
          5111 => x"06",
          5112 => x"7a",
          5113 => x"76",
          5114 => x"07",
          5115 => x"54",
          5116 => x"80",
          5117 => x"80",
          5118 => x"7b",
          5119 => x"53",
          5120 => x"93",
          5121 => x"dc",
          5122 => x"8c",
          5123 => x"38",
          5124 => x"55",
          5125 => x"56",
          5126 => x"8b",
          5127 => x"56",
          5128 => x"83",
          5129 => x"75",
          5130 => x"51",
          5131 => x"3f",
          5132 => x"08",
          5133 => x"82",
          5134 => x"98",
          5135 => x"e6",
          5136 => x"53",
          5137 => x"b8",
          5138 => x"3d",
          5139 => x"3f",
          5140 => x"08",
          5141 => x"08",
          5142 => x"8c",
          5143 => x"98",
          5144 => x"a0",
          5145 => x"70",
          5146 => x"ae",
          5147 => x"6d",
          5148 => x"81",
          5149 => x"57",
          5150 => x"74",
          5151 => x"38",
          5152 => x"81",
          5153 => x"81",
          5154 => x"52",
          5155 => x"89",
          5156 => x"dc",
          5157 => x"a5",
          5158 => x"33",
          5159 => x"54",
          5160 => x"3f",
          5161 => x"08",
          5162 => x"38",
          5163 => x"76",
          5164 => x"05",
          5165 => x"39",
          5166 => x"08",
          5167 => x"15",
          5168 => x"ff",
          5169 => x"73",
          5170 => x"38",
          5171 => x"83",
          5172 => x"56",
          5173 => x"75",
          5174 => x"81",
          5175 => x"33",
          5176 => x"2e",
          5177 => x"52",
          5178 => x"51",
          5179 => x"3f",
          5180 => x"08",
          5181 => x"ff",
          5182 => x"38",
          5183 => x"88",
          5184 => x"8a",
          5185 => x"38",
          5186 => x"ec",
          5187 => x"75",
          5188 => x"74",
          5189 => x"73",
          5190 => x"05",
          5191 => x"17",
          5192 => x"70",
          5193 => x"34",
          5194 => x"70",
          5195 => x"ff",
          5196 => x"55",
          5197 => x"26",
          5198 => x"8b",
          5199 => x"86",
          5200 => x"e5",
          5201 => x"38",
          5202 => x"99",
          5203 => x"05",
          5204 => x"70",
          5205 => x"73",
          5206 => x"81",
          5207 => x"ff",
          5208 => x"ed",
          5209 => x"80",
          5210 => x"91",
          5211 => x"55",
          5212 => x"3f",
          5213 => x"08",
          5214 => x"dc",
          5215 => x"38",
          5216 => x"51",
          5217 => x"3f",
          5218 => x"08",
          5219 => x"dc",
          5220 => x"76",
          5221 => x"67",
          5222 => x"34",
          5223 => x"82",
          5224 => x"84",
          5225 => x"06",
          5226 => x"80",
          5227 => x"2e",
          5228 => x"81",
          5229 => x"ff",
          5230 => x"82",
          5231 => x"54",
          5232 => x"08",
          5233 => x"53",
          5234 => x"08",
          5235 => x"ff",
          5236 => x"67",
          5237 => x"8b",
          5238 => x"53",
          5239 => x"51",
          5240 => x"3f",
          5241 => x"0b",
          5242 => x"79",
          5243 => x"ee",
          5244 => x"dc",
          5245 => x"55",
          5246 => x"dc",
          5247 => x"0d",
          5248 => x"0d",
          5249 => x"88",
          5250 => x"05",
          5251 => x"fc",
          5252 => x"54",
          5253 => x"d2",
          5254 => x"8c",
          5255 => x"82",
          5256 => x"82",
          5257 => x"1a",
          5258 => x"82",
          5259 => x"80",
          5260 => x"8c",
          5261 => x"78",
          5262 => x"1a",
          5263 => x"2a",
          5264 => x"51",
          5265 => x"90",
          5266 => x"82",
          5267 => x"58",
          5268 => x"81",
          5269 => x"39",
          5270 => x"22",
          5271 => x"70",
          5272 => x"56",
          5273 => x"e5",
          5274 => x"14",
          5275 => x"30",
          5276 => x"9f",
          5277 => x"dc",
          5278 => x"19",
          5279 => x"5a",
          5280 => x"81",
          5281 => x"38",
          5282 => x"77",
          5283 => x"82",
          5284 => x"56",
          5285 => x"74",
          5286 => x"ff",
          5287 => x"81",
          5288 => x"55",
          5289 => x"75",
          5290 => x"82",
          5291 => x"dc",
          5292 => x"ff",
          5293 => x"8c",
          5294 => x"2e",
          5295 => x"82",
          5296 => x"8e",
          5297 => x"56",
          5298 => x"09",
          5299 => x"38",
          5300 => x"59",
          5301 => x"77",
          5302 => x"06",
          5303 => x"87",
          5304 => x"39",
          5305 => x"ba",
          5306 => x"55",
          5307 => x"2e",
          5308 => x"15",
          5309 => x"2e",
          5310 => x"83",
          5311 => x"75",
          5312 => x"7e",
          5313 => x"a8",
          5314 => x"dc",
          5315 => x"8c",
          5316 => x"ce",
          5317 => x"16",
          5318 => x"56",
          5319 => x"38",
          5320 => x"19",
          5321 => x"8c",
          5322 => x"7d",
          5323 => x"38",
          5324 => x"0c",
          5325 => x"0c",
          5326 => x"80",
          5327 => x"73",
          5328 => x"98",
          5329 => x"05",
          5330 => x"57",
          5331 => x"26",
          5332 => x"7b",
          5333 => x"0c",
          5334 => x"81",
          5335 => x"84",
          5336 => x"54",
          5337 => x"dc",
          5338 => x"0d",
          5339 => x"0d",
          5340 => x"88",
          5341 => x"05",
          5342 => x"54",
          5343 => x"c5",
          5344 => x"56",
          5345 => x"8c",
          5346 => x"8b",
          5347 => x"8c",
          5348 => x"29",
          5349 => x"05",
          5350 => x"55",
          5351 => x"84",
          5352 => x"34",
          5353 => x"08",
          5354 => x"5f",
          5355 => x"51",
          5356 => x"3f",
          5357 => x"08",
          5358 => x"70",
          5359 => x"57",
          5360 => x"8b",
          5361 => x"82",
          5362 => x"06",
          5363 => x"56",
          5364 => x"38",
          5365 => x"05",
          5366 => x"7e",
          5367 => x"f0",
          5368 => x"dc",
          5369 => x"67",
          5370 => x"2e",
          5371 => x"82",
          5372 => x"8b",
          5373 => x"75",
          5374 => x"80",
          5375 => x"81",
          5376 => x"2e",
          5377 => x"80",
          5378 => x"38",
          5379 => x"0a",
          5380 => x"ff",
          5381 => x"55",
          5382 => x"86",
          5383 => x"8a",
          5384 => x"89",
          5385 => x"2a",
          5386 => x"77",
          5387 => x"59",
          5388 => x"81",
          5389 => x"70",
          5390 => x"07",
          5391 => x"56",
          5392 => x"38",
          5393 => x"05",
          5394 => x"7e",
          5395 => x"80",
          5396 => x"82",
          5397 => x"8a",
          5398 => x"83",
          5399 => x"06",
          5400 => x"08",
          5401 => x"74",
          5402 => x"41",
          5403 => x"56",
          5404 => x"8a",
          5405 => x"61",
          5406 => x"55",
          5407 => x"27",
          5408 => x"93",
          5409 => x"80",
          5410 => x"38",
          5411 => x"70",
          5412 => x"43",
          5413 => x"95",
          5414 => x"06",
          5415 => x"2e",
          5416 => x"77",
          5417 => x"74",
          5418 => x"83",
          5419 => x"06",
          5420 => x"82",
          5421 => x"2e",
          5422 => x"78",
          5423 => x"2e",
          5424 => x"80",
          5425 => x"ae",
          5426 => x"2a",
          5427 => x"81",
          5428 => x"56",
          5429 => x"2e",
          5430 => x"77",
          5431 => x"81",
          5432 => x"79",
          5433 => x"70",
          5434 => x"5a",
          5435 => x"86",
          5436 => x"27",
          5437 => x"52",
          5438 => x"e0",
          5439 => x"8c",
          5440 => x"29",
          5441 => x"70",
          5442 => x"55",
          5443 => x"0b",
          5444 => x"08",
          5445 => x"05",
          5446 => x"ff",
          5447 => x"27",
          5448 => x"88",
          5449 => x"ae",
          5450 => x"2a",
          5451 => x"81",
          5452 => x"56",
          5453 => x"2e",
          5454 => x"77",
          5455 => x"81",
          5456 => x"79",
          5457 => x"70",
          5458 => x"5a",
          5459 => x"86",
          5460 => x"27",
          5461 => x"52",
          5462 => x"e0",
          5463 => x"8c",
          5464 => x"84",
          5465 => x"8c",
          5466 => x"f5",
          5467 => x"81",
          5468 => x"dc",
          5469 => x"8c",
          5470 => x"71",
          5471 => x"83",
          5472 => x"5e",
          5473 => x"89",
          5474 => x"5c",
          5475 => x"1c",
          5476 => x"05",
          5477 => x"ff",
          5478 => x"70",
          5479 => x"31",
          5480 => x"57",
          5481 => x"83",
          5482 => x"06",
          5483 => x"1c",
          5484 => x"5c",
          5485 => x"1d",
          5486 => x"29",
          5487 => x"31",
          5488 => x"55",
          5489 => x"87",
          5490 => x"7c",
          5491 => x"7a",
          5492 => x"31",
          5493 => x"df",
          5494 => x"8c",
          5495 => x"7d",
          5496 => x"81",
          5497 => x"82",
          5498 => x"83",
          5499 => x"80",
          5500 => x"87",
          5501 => x"81",
          5502 => x"fd",
          5503 => x"f8",
          5504 => x"2e",
          5505 => x"80",
          5506 => x"ff",
          5507 => x"8c",
          5508 => x"a0",
          5509 => x"38",
          5510 => x"74",
          5511 => x"86",
          5512 => x"fd",
          5513 => x"81",
          5514 => x"80",
          5515 => x"83",
          5516 => x"39",
          5517 => x"08",
          5518 => x"92",
          5519 => x"b8",
          5520 => x"59",
          5521 => x"27",
          5522 => x"86",
          5523 => x"55",
          5524 => x"09",
          5525 => x"38",
          5526 => x"f5",
          5527 => x"38",
          5528 => x"55",
          5529 => x"86",
          5530 => x"80",
          5531 => x"7a",
          5532 => x"b9",
          5533 => x"81",
          5534 => x"7a",
          5535 => x"8a",
          5536 => x"52",
          5537 => x"ff",
          5538 => x"79",
          5539 => x"7b",
          5540 => x"06",
          5541 => x"51",
          5542 => x"3f",
          5543 => x"1c",
          5544 => x"32",
          5545 => x"96",
          5546 => x"06",
          5547 => x"91",
          5548 => x"a1",
          5549 => x"55",
          5550 => x"ff",
          5551 => x"74",
          5552 => x"06",
          5553 => x"51",
          5554 => x"3f",
          5555 => x"52",
          5556 => x"ff",
          5557 => x"f8",
          5558 => x"34",
          5559 => x"1b",
          5560 => x"d9",
          5561 => x"52",
          5562 => x"ff",
          5563 => x"60",
          5564 => x"51",
          5565 => x"3f",
          5566 => x"09",
          5567 => x"cb",
          5568 => x"b2",
          5569 => x"c3",
          5570 => x"a0",
          5571 => x"52",
          5572 => x"ff",
          5573 => x"82",
          5574 => x"51",
          5575 => x"3f",
          5576 => x"1b",
          5577 => x"95",
          5578 => x"b2",
          5579 => x"a0",
          5580 => x"80",
          5581 => x"1c",
          5582 => x"80",
          5583 => x"93",
          5584 => x"b4",
          5585 => x"1b",
          5586 => x"82",
          5587 => x"52",
          5588 => x"ff",
          5589 => x"7c",
          5590 => x"06",
          5591 => x"51",
          5592 => x"3f",
          5593 => x"a4",
          5594 => x"0b",
          5595 => x"93",
          5596 => x"c8",
          5597 => x"51",
          5598 => x"3f",
          5599 => x"52",
          5600 => x"70",
          5601 => x"9f",
          5602 => x"54",
          5603 => x"52",
          5604 => x"9b",
          5605 => x"56",
          5606 => x"08",
          5607 => x"7d",
          5608 => x"81",
          5609 => x"38",
          5610 => x"86",
          5611 => x"52",
          5612 => x"9b",
          5613 => x"80",
          5614 => x"7a",
          5615 => x"ed",
          5616 => x"85",
          5617 => x"7a",
          5618 => x"8f",
          5619 => x"85",
          5620 => x"83",
          5621 => x"ff",
          5622 => x"ff",
          5623 => x"e8",
          5624 => x"9e",
          5625 => x"52",
          5626 => x"51",
          5627 => x"3f",
          5628 => x"52",
          5629 => x"9e",
          5630 => x"54",
          5631 => x"53",
          5632 => x"51",
          5633 => x"3f",
          5634 => x"16",
          5635 => x"7e",
          5636 => x"d8",
          5637 => x"80",
          5638 => x"ff",
          5639 => x"7f",
          5640 => x"7d",
          5641 => x"81",
          5642 => x"f8",
          5643 => x"ff",
          5644 => x"ff",
          5645 => x"51",
          5646 => x"3f",
          5647 => x"88",
          5648 => x"39",
          5649 => x"f8",
          5650 => x"2e",
          5651 => x"55",
          5652 => x"51",
          5653 => x"3f",
          5654 => x"57",
          5655 => x"83",
          5656 => x"76",
          5657 => x"7a",
          5658 => x"ff",
          5659 => x"82",
          5660 => x"82",
          5661 => x"80",
          5662 => x"dc",
          5663 => x"51",
          5664 => x"3f",
          5665 => x"78",
          5666 => x"74",
          5667 => x"18",
          5668 => x"2e",
          5669 => x"79",
          5670 => x"2e",
          5671 => x"55",
          5672 => x"62",
          5673 => x"74",
          5674 => x"75",
          5675 => x"7e",
          5676 => x"b8",
          5677 => x"dc",
          5678 => x"38",
          5679 => x"78",
          5680 => x"74",
          5681 => x"56",
          5682 => x"93",
          5683 => x"66",
          5684 => x"26",
          5685 => x"56",
          5686 => x"83",
          5687 => x"64",
          5688 => x"77",
          5689 => x"84",
          5690 => x"52",
          5691 => x"9d",
          5692 => x"d4",
          5693 => x"51",
          5694 => x"3f",
          5695 => x"55",
          5696 => x"81",
          5697 => x"34",
          5698 => x"16",
          5699 => x"16",
          5700 => x"16",
          5701 => x"05",
          5702 => x"c1",
          5703 => x"fe",
          5704 => x"fe",
          5705 => x"34",
          5706 => x"08",
          5707 => x"07",
          5708 => x"16",
          5709 => x"dc",
          5710 => x"34",
          5711 => x"c6",
          5712 => x"9c",
          5713 => x"52",
          5714 => x"51",
          5715 => x"3f",
          5716 => x"53",
          5717 => x"51",
          5718 => x"3f",
          5719 => x"8c",
          5720 => x"38",
          5721 => x"52",
          5722 => x"99",
          5723 => x"56",
          5724 => x"08",
          5725 => x"39",
          5726 => x"39",
          5727 => x"39",
          5728 => x"08",
          5729 => x"8c",
          5730 => x"3d",
          5731 => x"3d",
          5732 => x"5b",
          5733 => x"60",
          5734 => x"57",
          5735 => x"25",
          5736 => x"3d",
          5737 => x"55",
          5738 => x"15",
          5739 => x"c9",
          5740 => x"81",
          5741 => x"06",
          5742 => x"3d",
          5743 => x"8d",
          5744 => x"74",
          5745 => x"05",
          5746 => x"17",
          5747 => x"2e",
          5748 => x"c9",
          5749 => x"34",
          5750 => x"83",
          5751 => x"74",
          5752 => x"0c",
          5753 => x"04",
          5754 => x"7b",
          5755 => x"b3",
          5756 => x"57",
          5757 => x"09",
          5758 => x"38",
          5759 => x"51",
          5760 => x"17",
          5761 => x"76",
          5762 => x"88",
          5763 => x"17",
          5764 => x"59",
          5765 => x"81",
          5766 => x"76",
          5767 => x"8b",
          5768 => x"54",
          5769 => x"17",
          5770 => x"51",
          5771 => x"79",
          5772 => x"30",
          5773 => x"9f",
          5774 => x"53",
          5775 => x"75",
          5776 => x"81",
          5777 => x"0c",
          5778 => x"04",
          5779 => x"79",
          5780 => x"56",
          5781 => x"24",
          5782 => x"3d",
          5783 => x"74",
          5784 => x"52",
          5785 => x"cb",
          5786 => x"8c",
          5787 => x"38",
          5788 => x"78",
          5789 => x"06",
          5790 => x"16",
          5791 => x"39",
          5792 => x"82",
          5793 => x"89",
          5794 => x"fd",
          5795 => x"54",
          5796 => x"80",
          5797 => x"ff",
          5798 => x"76",
          5799 => x"3d",
          5800 => x"3d",
          5801 => x"e3",
          5802 => x"53",
          5803 => x"53",
          5804 => x"3f",
          5805 => x"51",
          5806 => x"72",
          5807 => x"3f",
          5808 => x"04",
          5809 => x"7a",
          5810 => x"56",
          5811 => x"80",
          5812 => x"38",
          5813 => x"15",
          5814 => x"16",
          5815 => x"d4",
          5816 => x"54",
          5817 => x"09",
          5818 => x"38",
          5819 => x"f1",
          5820 => x"76",
          5821 => x"89",
          5822 => x"08",
          5823 => x"da",
          5824 => x"8c",
          5825 => x"8c",
          5826 => x"75",
          5827 => x"52",
          5828 => x"be",
          5829 => x"dc",
          5830 => x"84",
          5831 => x"73",
          5832 => x"b2",
          5833 => x"70",
          5834 => x"58",
          5835 => x"27",
          5836 => x"54",
          5837 => x"dc",
          5838 => x"0d",
          5839 => x"0d",
          5840 => x"93",
          5841 => x"38",
          5842 => x"81",
          5843 => x"52",
          5844 => x"81",
          5845 => x"81",
          5846 => x"fd",
          5847 => x"f9",
          5848 => x"e8",
          5849 => x"39",
          5850 => x"51",
          5851 => x"81",
          5852 => x"80",
          5853 => x"fe",
          5854 => x"dd",
          5855 => x"b0",
          5856 => x"39",
          5857 => x"51",
          5858 => x"81",
          5859 => x"80",
          5860 => x"fe",
          5861 => x"c1",
          5862 => x"88",
          5863 => x"81",
          5864 => x"b5",
          5865 => x"b8",
          5866 => x"81",
          5867 => x"a9",
          5868 => x"f8",
          5869 => x"82",
          5870 => x"9d",
          5871 => x"ac",
          5872 => x"82",
          5873 => x"91",
          5874 => x"dc",
          5875 => x"82",
          5876 => x"85",
          5877 => x"80",
          5878 => x"ae",
          5879 => x"0d",
          5880 => x"0d",
          5881 => x"56",
          5882 => x"26",
          5883 => x"52",
          5884 => x"29",
          5885 => x"87",
          5886 => x"51",
          5887 => x"3f",
          5888 => x"08",
          5889 => x"fe",
          5890 => x"82",
          5891 => x"54",
          5892 => x"52",
          5893 => x"51",
          5894 => x"3f",
          5895 => x"04",
          5896 => x"66",
          5897 => x"80",
          5898 => x"5b",
          5899 => x"78",
          5900 => x"07",
          5901 => x"57",
          5902 => x"56",
          5903 => x"26",
          5904 => x"56",
          5905 => x"70",
          5906 => x"51",
          5907 => x"74",
          5908 => x"81",
          5909 => x"8c",
          5910 => x"56",
          5911 => x"3f",
          5912 => x"08",
          5913 => x"dc",
          5914 => x"82",
          5915 => x"87",
          5916 => x"0c",
          5917 => x"08",
          5918 => x"d4",
          5919 => x"80",
          5920 => x"75",
          5921 => x"3f",
          5922 => x"08",
          5923 => x"dc",
          5924 => x"7a",
          5925 => x"2e",
          5926 => x"19",
          5927 => x"59",
          5928 => x"3d",
          5929 => x"cb",
          5930 => x"30",
          5931 => x"80",
          5932 => x"70",
          5933 => x"06",
          5934 => x"56",
          5935 => x"90",
          5936 => x"b4",
          5937 => x"98",
          5938 => x"78",
          5939 => x"3f",
          5940 => x"82",
          5941 => x"96",
          5942 => x"f9",
          5943 => x"02",
          5944 => x"05",
          5945 => x"ff",
          5946 => x"7a",
          5947 => x"fe",
          5948 => x"8c",
          5949 => x"38",
          5950 => x"88",
          5951 => x"2e",
          5952 => x"39",
          5953 => x"54",
          5954 => x"53",
          5955 => x"51",
          5956 => x"8c",
          5957 => x"83",
          5958 => x"76",
          5959 => x"0c",
          5960 => x"04",
          5961 => x"7f",
          5962 => x"8c",
          5963 => x"05",
          5964 => x"15",
          5965 => x"5c",
          5966 => x"5e",
          5967 => x"81",
          5968 => x"f5",
          5969 => x"81",
          5970 => x"ef",
          5971 => x"55",
          5972 => x"80",
          5973 => x"90",
          5974 => x"7b",
          5975 => x"38",
          5976 => x"74",
          5977 => x"7a",
          5978 => x"72",
          5979 => x"81",
          5980 => x"f4",
          5981 => x"39",
          5982 => x"51",
          5983 => x"3f",
          5984 => x"80",
          5985 => x"18",
          5986 => x"27",
          5987 => x"08",
          5988 => x"bc",
          5989 => x"d6",
          5990 => x"82",
          5991 => x"fe",
          5992 => x"84",
          5993 => x"39",
          5994 => x"72",
          5995 => x"38",
          5996 => x"82",
          5997 => x"fe",
          5998 => x"89",
          5999 => x"e4",
          6000 => x"c6",
          6001 => x"55",
          6002 => x"ed",
          6003 => x"80",
          6004 => x"e8",
          6005 => x"b2",
          6006 => x"74",
          6007 => x"38",
          6008 => x"33",
          6009 => x"56",
          6010 => x"83",
          6011 => x"80",
          6012 => x"27",
          6013 => x"53",
          6014 => x"70",
          6015 => x"51",
          6016 => x"2e",
          6017 => x"80",
          6018 => x"38",
          6019 => x"39",
          6020 => x"ed",
          6021 => x"15",
          6022 => x"82",
          6023 => x"fe",
          6024 => x"78",
          6025 => x"5c",
          6026 => x"d5",
          6027 => x"dc",
          6028 => x"70",
          6029 => x"57",
          6030 => x"09",
          6031 => x"38",
          6032 => x"3f",
          6033 => x"08",
          6034 => x"98",
          6035 => x"32",
          6036 => x"9b",
          6037 => x"70",
          6038 => x"75",
          6039 => x"58",
          6040 => x"51",
          6041 => x"24",
          6042 => x"9b",
          6043 => x"06",
          6044 => x"53",
          6045 => x"1e",
          6046 => x"26",
          6047 => x"ff",
          6048 => x"8c",
          6049 => x"3d",
          6050 => x"3d",
          6051 => x"05",
          6052 => x"f0",
          6053 => x"f4",
          6054 => x"f2",
          6055 => x"88",
          6056 => x"fe",
          6057 => x"82",
          6058 => x"82",
          6059 => x"82",
          6060 => x"52",
          6061 => x"51",
          6062 => x"3f",
          6063 => x"85",
          6064 => x"e1",
          6065 => x"0d",
          6066 => x"0d",
          6067 => x"80",
          6068 => x"e7",
          6069 => x"51",
          6070 => x"3f",
          6071 => x"51",
          6072 => x"3f",
          6073 => x"d9",
          6074 => x"81",
          6075 => x"06",
          6076 => x"80",
          6077 => x"81",
          6078 => x"99",
          6079 => x"c8",
          6080 => x"91",
          6081 => x"fe",
          6082 => x"72",
          6083 => x"81",
          6084 => x"71",
          6085 => x"38",
          6086 => x"d8",
          6087 => x"82",
          6088 => x"da",
          6089 => x"51",
          6090 => x"3f",
          6091 => x"70",
          6092 => x"52",
          6093 => x"95",
          6094 => x"fe",
          6095 => x"82",
          6096 => x"fe",
          6097 => x"80",
          6098 => x"c9",
          6099 => x"2a",
          6100 => x"51",
          6101 => x"2e",
          6102 => x"51",
          6103 => x"3f",
          6104 => x"51",
          6105 => x"3f",
          6106 => x"d8",
          6107 => x"85",
          6108 => x"06",
          6109 => x"80",
          6110 => x"81",
          6111 => x"95",
          6112 => x"94",
          6113 => x"8d",
          6114 => x"fe",
          6115 => x"72",
          6116 => x"81",
          6117 => x"71",
          6118 => x"38",
          6119 => x"d7",
          6120 => x"83",
          6121 => x"d9",
          6122 => x"51",
          6123 => x"3f",
          6124 => x"70",
          6125 => x"52",
          6126 => x"95",
          6127 => x"fe",
          6128 => x"82",
          6129 => x"fe",
          6130 => x"80",
          6131 => x"c5",
          6132 => x"2a",
          6133 => x"51",
          6134 => x"2e",
          6135 => x"51",
          6136 => x"3f",
          6137 => x"51",
          6138 => x"3f",
          6139 => x"d7",
          6140 => x"e5",
          6141 => x"3d",
          6142 => x"3d",
          6143 => x"84",
          6144 => x"33",
          6145 => x"56",
          6146 => x"51",
          6147 => x"3f",
          6148 => x"33",
          6149 => x"38",
          6150 => x"84",
          6151 => x"a3",
          6152 => x"b8",
          6153 => x"8c",
          6154 => x"70",
          6155 => x"08",
          6156 => x"82",
          6157 => x"51",
          6158 => x"89",
          6159 => x"89",
          6160 => x"73",
          6161 => x"81",
          6162 => x"82",
          6163 => x"74",
          6164 => x"f2",
          6165 => x"8c",
          6166 => x"2e",
          6167 => x"8c",
          6168 => x"fe",
          6169 => x"8e",
          6170 => x"f4",
          6171 => x"3f",
          6172 => x"89",
          6173 => x"89",
          6174 => x"73",
          6175 => x"81",
          6176 => x"74",
          6177 => x"fe",
          6178 => x"80",
          6179 => x"dc",
          6180 => x"0d",
          6181 => x"0d",
          6182 => x"82",
          6183 => x"5f",
          6184 => x"7c",
          6185 => x"db",
          6186 => x"dc",
          6187 => x"06",
          6188 => x"2e",
          6189 => x"a2",
          6190 => x"a0",
          6191 => x"70",
          6192 => x"ee",
          6193 => x"53",
          6194 => x"8e",
          6195 => x"b5",
          6196 => x"8c",
          6197 => x"2e",
          6198 => x"84",
          6199 => x"bc",
          6200 => x"5f",
          6201 => x"dc",
          6202 => x"9e",
          6203 => x"70",
          6204 => x"f8",
          6205 => x"fe",
          6206 => x"3d",
          6207 => x"51",
          6208 => x"82",
          6209 => x"90",
          6210 => x"2c",
          6211 => x"80",
          6212 => x"b3",
          6213 => x"c2",
          6214 => x"78",
          6215 => x"d5",
          6216 => x"24",
          6217 => x"80",
          6218 => x"38",
          6219 => x"80",
          6220 => x"e9",
          6221 => x"c0",
          6222 => x"38",
          6223 => x"24",
          6224 => x"78",
          6225 => x"92",
          6226 => x"39",
          6227 => x"2e",
          6228 => x"78",
          6229 => x"92",
          6230 => x"c3",
          6231 => x"38",
          6232 => x"2e",
          6233 => x"8a",
          6234 => x"81",
          6235 => x"99",
          6236 => x"83",
          6237 => x"78",
          6238 => x"89",
          6239 => x"9d",
          6240 => x"85",
          6241 => x"38",
          6242 => x"b4",
          6243 => x"11",
          6244 => x"05",
          6245 => x"cb",
          6246 => x"dc",
          6247 => x"fe",
          6248 => x"3d",
          6249 => x"53",
          6250 => x"51",
          6251 => x"3f",
          6252 => x"08",
          6253 => x"ad",
          6254 => x"fe",
          6255 => x"ff",
          6256 => x"fe",
          6257 => x"82",
          6258 => x"86",
          6259 => x"dc",
          6260 => x"84",
          6261 => x"e6",
          6262 => x"63",
          6263 => x"7b",
          6264 => x"38",
          6265 => x"7a",
          6266 => x"5c",
          6267 => x"26",
          6268 => x"e1",
          6269 => x"ff",
          6270 => x"ff",
          6271 => x"fe",
          6272 => x"82",
          6273 => x"80",
          6274 => x"38",
          6275 => x"fc",
          6276 => x"84",
          6277 => x"ed",
          6278 => x"8c",
          6279 => x"2e",
          6280 => x"b4",
          6281 => x"11",
          6282 => x"05",
          6283 => x"b3",
          6284 => x"dc",
          6285 => x"fd",
          6286 => x"84",
          6287 => x"e5",
          6288 => x"5a",
          6289 => x"81",
          6290 => x"59",
          6291 => x"05",
          6292 => x"34",
          6293 => x"42",
          6294 => x"3d",
          6295 => x"53",
          6296 => x"51",
          6297 => x"3f",
          6298 => x"08",
          6299 => x"f5",
          6300 => x"fe",
          6301 => x"ff",
          6302 => x"fe",
          6303 => x"82",
          6304 => x"80",
          6305 => x"38",
          6306 => x"f8",
          6307 => x"84",
          6308 => x"ec",
          6309 => x"8c",
          6310 => x"2e",
          6311 => x"82",
          6312 => x"fe",
          6313 => x"63",
          6314 => x"27",
          6315 => x"70",
          6316 => x"5e",
          6317 => x"7c",
          6318 => x"78",
          6319 => x"79",
          6320 => x"52",
          6321 => x"51",
          6322 => x"3f",
          6323 => x"81",
          6324 => x"d5",
          6325 => x"a4",
          6326 => x"39",
          6327 => x"80",
          6328 => x"84",
          6329 => x"eb",
          6330 => x"8c",
          6331 => x"df",
          6332 => x"a0",
          6333 => x"80",
          6334 => x"82",
          6335 => x"44",
          6336 => x"82",
          6337 => x"59",
          6338 => x"88",
          6339 => x"e0",
          6340 => x"39",
          6341 => x"33",
          6342 => x"2e",
          6343 => x"87",
          6344 => x"ab",
          6345 => x"a3",
          6346 => x"80",
          6347 => x"82",
          6348 => x"44",
          6349 => x"88",
          6350 => x"78",
          6351 => x"38",
          6352 => x"08",
          6353 => x"82",
          6354 => x"fc",
          6355 => x"b4",
          6356 => x"11",
          6357 => x"05",
          6358 => x"87",
          6359 => x"dc",
          6360 => x"38",
          6361 => x"33",
          6362 => x"2e",
          6363 => x"87",
          6364 => x"80",
          6365 => x"88",
          6366 => x"78",
          6367 => x"38",
          6368 => x"08",
          6369 => x"82",
          6370 => x"59",
          6371 => x"88",
          6372 => x"ec",
          6373 => x"39",
          6374 => x"33",
          6375 => x"2e",
          6376 => x"87",
          6377 => x"99",
          6378 => x"9e",
          6379 => x"80",
          6380 => x"82",
          6381 => x"43",
          6382 => x"88",
          6383 => x"05",
          6384 => x"fe",
          6385 => x"ff",
          6386 => x"fe",
          6387 => x"82",
          6388 => x"80",
          6389 => x"80",
          6390 => x"7a",
          6391 => x"38",
          6392 => x"90",
          6393 => x"70",
          6394 => x"2a",
          6395 => x"51",
          6396 => x"78",
          6397 => x"38",
          6398 => x"83",
          6399 => x"82",
          6400 => x"fe",
          6401 => x"a0",
          6402 => x"61",
          6403 => x"63",
          6404 => x"3f",
          6405 => x"51",
          6406 => x"3f",
          6407 => x"b4",
          6408 => x"11",
          6409 => x"05",
          6410 => x"b7",
          6411 => x"dc",
          6412 => x"f9",
          6413 => x"3d",
          6414 => x"53",
          6415 => x"51",
          6416 => x"3f",
          6417 => x"08",
          6418 => x"38",
          6419 => x"80",
          6420 => x"79",
          6421 => x"05",
          6422 => x"fe",
          6423 => x"ff",
          6424 => x"fe",
          6425 => x"82",
          6426 => x"e0",
          6427 => x"39",
          6428 => x"54",
          6429 => x"c4",
          6430 => x"f2",
          6431 => x"52",
          6432 => x"e7",
          6433 => x"45",
          6434 => x"78",
          6435 => x"d5",
          6436 => x"27",
          6437 => x"3d",
          6438 => x"53",
          6439 => x"51",
          6440 => x"3f",
          6441 => x"08",
          6442 => x"38",
          6443 => x"80",
          6444 => x"79",
          6445 => x"05",
          6446 => x"39",
          6447 => x"51",
          6448 => x"3f",
          6449 => x"b4",
          6450 => x"11",
          6451 => x"05",
          6452 => x"81",
          6453 => x"dc",
          6454 => x"f8",
          6455 => x"3d",
          6456 => x"53",
          6457 => x"51",
          6458 => x"3f",
          6459 => x"08",
          6460 => x"38",
          6461 => x"be",
          6462 => x"70",
          6463 => x"23",
          6464 => x"3d",
          6465 => x"53",
          6466 => x"51",
          6467 => x"3f",
          6468 => x"08",
          6469 => x"cd",
          6470 => x"22",
          6471 => x"85",
          6472 => x"e5",
          6473 => x"f8",
          6474 => x"fe",
          6475 => x"79",
          6476 => x"59",
          6477 => x"f7",
          6478 => x"9f",
          6479 => x"60",
          6480 => x"d5",
          6481 => x"fe",
          6482 => x"ff",
          6483 => x"fe",
          6484 => x"82",
          6485 => x"80",
          6486 => x"60",
          6487 => x"05",
          6488 => x"82",
          6489 => x"78",
          6490 => x"39",
          6491 => x"51",
          6492 => x"3f",
          6493 => x"b4",
          6494 => x"11",
          6495 => x"05",
          6496 => x"d1",
          6497 => x"dc",
          6498 => x"f6",
          6499 => x"3d",
          6500 => x"53",
          6501 => x"51",
          6502 => x"3f",
          6503 => x"08",
          6504 => x"38",
          6505 => x"0c",
          6506 => x"05",
          6507 => x"fe",
          6508 => x"ff",
          6509 => x"fe",
          6510 => x"82",
          6511 => x"e4",
          6512 => x"39",
          6513 => x"54",
          6514 => x"e4",
          6515 => x"9e",
          6516 => x"52",
          6517 => x"e4",
          6518 => x"45",
          6519 => x"78",
          6520 => x"81",
          6521 => x"27",
          6522 => x"3d",
          6523 => x"53",
          6524 => x"51",
          6525 => x"3f",
          6526 => x"08",
          6527 => x"38",
          6528 => x"0c",
          6529 => x"05",
          6530 => x"39",
          6531 => x"51",
          6532 => x"3f",
          6533 => x"b4",
          6534 => x"11",
          6535 => x"05",
          6536 => x"bf",
          6537 => x"dc",
          6538 => x"f5",
          6539 => x"52",
          6540 => x"51",
          6541 => x"3f",
          6542 => x"04",
          6543 => x"80",
          6544 => x"84",
          6545 => x"e5",
          6546 => x"8c",
          6547 => x"2e",
          6548 => x"63",
          6549 => x"8c",
          6550 => x"92",
          6551 => x"78",
          6552 => x"dc",
          6553 => x"f4",
          6554 => x"8c",
          6555 => x"82",
          6556 => x"fe",
          6557 => x"f4",
          6558 => x"86",
          6559 => x"dd",
          6560 => x"bd",
          6561 => x"dd",
          6562 => x"e0",
          6563 => x"fa",
          6564 => x"ff",
          6565 => x"d3",
          6566 => x"c9",
          6567 => x"79",
          6568 => x"80",
          6569 => x"38",
          6570 => x"59",
          6571 => x"81",
          6572 => x"3d",
          6573 => x"51",
          6574 => x"3f",
          6575 => x"08",
          6576 => x"7a",
          6577 => x"38",
          6578 => x"89",
          6579 => x"2e",
          6580 => x"cd",
          6581 => x"2e",
          6582 => x"c5",
          6583 => x"f4",
          6584 => x"82",
          6585 => x"80",
          6586 => x"fc",
          6587 => x"ff",
          6588 => x"fe",
          6589 => x"bb",
          6590 => x"9c",
          6591 => x"ff",
          6592 => x"fe",
          6593 => x"ab",
          6594 => x"82",
          6595 => x"80",
          6596 => x"8c",
          6597 => x"ff",
          6598 => x"fe",
          6599 => x"93",
          6600 => x"80",
          6601 => x"98",
          6602 => x"ff",
          6603 => x"fe",
          6604 => x"82",
          6605 => x"82",
          6606 => x"80",
          6607 => x"80",
          6608 => x"80",
          6609 => x"80",
          6610 => x"ff",
          6611 => x"eb",
          6612 => x"8c",
          6613 => x"8c",
          6614 => x"70",
          6615 => x"07",
          6616 => x"5b",
          6617 => x"5a",
          6618 => x"83",
          6619 => x"78",
          6620 => x"78",
          6621 => x"38",
          6622 => x"81",
          6623 => x"59",
          6624 => x"38",
          6625 => x"7d",
          6626 => x"59",
          6627 => x"7e",
          6628 => x"81",
          6629 => x"38",
          6630 => x"51",
          6631 => x"3f",
          6632 => x"fc",
          6633 => x"0b",
          6634 => x"34",
          6635 => x"8c",
          6636 => x"55",
          6637 => x"52",
          6638 => x"bb",
          6639 => x"8c",
          6640 => x"2b",
          6641 => x"53",
          6642 => x"52",
          6643 => x"bb",
          6644 => x"82",
          6645 => x"07",
          6646 => x"c0",
          6647 => x"08",
          6648 => x"84",
          6649 => x"51",
          6650 => x"3f",
          6651 => x"08",
          6652 => x"08",
          6653 => x"84",
          6654 => x"51",
          6655 => x"3f",
          6656 => x"dc",
          6657 => x"0c",
          6658 => x"0b",
          6659 => x"84",
          6660 => x"83",
          6661 => x"94",
          6662 => x"ac",
          6663 => x"f0",
          6664 => x"0b",
          6665 => x"0c",
          6666 => x"3f",
          6667 => x"3f",
          6668 => x"51",
          6669 => x"3f",
          6670 => x"51",
          6671 => x"3f",
          6672 => x"51",
          6673 => x"3f",
          6674 => x"be",
          6675 => x"3f",
          6676 => x"00",
          6677 => x"00",
          6678 => x"00",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"00",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"00",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"00",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"00",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"00",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"00",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"00",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"00",
          6711 => x"00",
          6712 => x"00",
          6713 => x"25",
          6714 => x"64",
          6715 => x"20",
          6716 => x"25",
          6717 => x"64",
          6718 => x"25",
          6719 => x"53",
          6720 => x"43",
          6721 => x"69",
          6722 => x"61",
          6723 => x"6e",
          6724 => x"20",
          6725 => x"6f",
          6726 => x"6f",
          6727 => x"6f",
          6728 => x"67",
          6729 => x"3a",
          6730 => x"76",
          6731 => x"73",
          6732 => x"70",
          6733 => x"65",
          6734 => x"64",
          6735 => x"20",
          6736 => x"57",
          6737 => x"44",
          6738 => x"20",
          6739 => x"30",
          6740 => x"25",
          6741 => x"29",
          6742 => x"20",
          6743 => x"53",
          6744 => x"4d",
          6745 => x"20",
          6746 => x"30",
          6747 => x"25",
          6748 => x"29",
          6749 => x"20",
          6750 => x"49",
          6751 => x"20",
          6752 => x"4d",
          6753 => x"30",
          6754 => x"25",
          6755 => x"29",
          6756 => x"20",
          6757 => x"42",
          6758 => x"20",
          6759 => x"20",
          6760 => x"30",
          6761 => x"25",
          6762 => x"29",
          6763 => x"20",
          6764 => x"52",
          6765 => x"20",
          6766 => x"20",
          6767 => x"30",
          6768 => x"25",
          6769 => x"29",
          6770 => x"20",
          6771 => x"53",
          6772 => x"41",
          6773 => x"20",
          6774 => x"65",
          6775 => x"65",
          6776 => x"25",
          6777 => x"29",
          6778 => x"20",
          6779 => x"54",
          6780 => x"52",
          6781 => x"20",
          6782 => x"69",
          6783 => x"73",
          6784 => x"25",
          6785 => x"29",
          6786 => x"20",
          6787 => x"49",
          6788 => x"20",
          6789 => x"4c",
          6790 => x"68",
          6791 => x"65",
          6792 => x"25",
          6793 => x"29",
          6794 => x"20",
          6795 => x"57",
          6796 => x"42",
          6797 => x"20",
          6798 => x"0a",
          6799 => x"20",
          6800 => x"57",
          6801 => x"32",
          6802 => x"20",
          6803 => x"49",
          6804 => x"4c",
          6805 => x"20",
          6806 => x"50",
          6807 => x"00",
          6808 => x"20",
          6809 => x"53",
          6810 => x"00",
          6811 => x"41",
          6812 => x"65",
          6813 => x"73",
          6814 => x"20",
          6815 => x"43",
          6816 => x"52",
          6817 => x"74",
          6818 => x"63",
          6819 => x"20",
          6820 => x"72",
          6821 => x"20",
          6822 => x"30",
          6823 => x"00",
          6824 => x"20",
          6825 => x"43",
          6826 => x"4d",
          6827 => x"72",
          6828 => x"74",
          6829 => x"20",
          6830 => x"72",
          6831 => x"20",
          6832 => x"30",
          6833 => x"00",
          6834 => x"20",
          6835 => x"53",
          6836 => x"6b",
          6837 => x"61",
          6838 => x"41",
          6839 => x"65",
          6840 => x"20",
          6841 => x"20",
          6842 => x"30",
          6843 => x"00",
          6844 => x"4d",
          6845 => x"3a",
          6846 => x"20",
          6847 => x"5a",
          6848 => x"49",
          6849 => x"20",
          6850 => x"20",
          6851 => x"20",
          6852 => x"20",
          6853 => x"20",
          6854 => x"30",
          6855 => x"00",
          6856 => x"20",
          6857 => x"53",
          6858 => x"65",
          6859 => x"6c",
          6860 => x"20",
          6861 => x"71",
          6862 => x"20",
          6863 => x"20",
          6864 => x"64",
          6865 => x"34",
          6866 => x"7a",
          6867 => x"20",
          6868 => x"53",
          6869 => x"4d",
          6870 => x"6f",
          6871 => x"46",
          6872 => x"20",
          6873 => x"20",
          6874 => x"20",
          6875 => x"64",
          6876 => x"34",
          6877 => x"7a",
          6878 => x"20",
          6879 => x"57",
          6880 => x"62",
          6881 => x"20",
          6882 => x"41",
          6883 => x"6c",
          6884 => x"20",
          6885 => x"71",
          6886 => x"64",
          6887 => x"34",
          6888 => x"7a",
          6889 => x"53",
          6890 => x"6c",
          6891 => x"4d",
          6892 => x"75",
          6893 => x"46",
          6894 => x"00",
          6895 => x"45",
          6896 => x"45",
          6897 => x"69",
          6898 => x"55",
          6899 => x"6f",
          6900 => x"68",
          6901 => x"6f",
          6902 => x"74",
          6903 => x"68",
          6904 => x"6f",
          6905 => x"68",
          6906 => x"00",
          6907 => x"21",
          6908 => x"25",
          6909 => x"20",
          6910 => x"0a",
          6911 => x"46",
          6912 => x"65",
          6913 => x"6f",
          6914 => x"73",
          6915 => x"74",
          6916 => x"68",
          6917 => x"6f",
          6918 => x"66",
          6919 => x"20",
          6920 => x"45",
          6921 => x"0a",
          6922 => x"43",
          6923 => x"6f",
          6924 => x"70",
          6925 => x"63",
          6926 => x"74",
          6927 => x"69",
          6928 => x"72",
          6929 => x"69",
          6930 => x"20",
          6931 => x"61",
          6932 => x"6e",
          6933 => x"00",
          6934 => x"00",
          6935 => x"01",
          6936 => x"00",
          6937 => x"00",
          6938 => x"01",
          6939 => x"00",
          6940 => x"00",
          6941 => x"04",
          6942 => x"00",
          6943 => x"00",
          6944 => x"04",
          6945 => x"00",
          6946 => x"00",
          6947 => x"04",
          6948 => x"00",
          6949 => x"00",
          6950 => x"04",
          6951 => x"00",
          6952 => x"00",
          6953 => x"04",
          6954 => x"00",
          6955 => x"00",
          6956 => x"03",
          6957 => x"00",
          6958 => x"00",
          6959 => x"03",
          6960 => x"00",
          6961 => x"00",
          6962 => x"03",
          6963 => x"00",
          6964 => x"00",
          6965 => x"03",
          6966 => x"00",
          6967 => x"1b",
          6968 => x"1b",
          6969 => x"1b",
          6970 => x"1b",
          6971 => x"1b",
          6972 => x"1b",
          6973 => x"1b",
          6974 => x"1b",
          6975 => x"1b",
          6976 => x"0d",
          6977 => x"08",
          6978 => x"53",
          6979 => x"22",
          6980 => x"3a",
          6981 => x"3e",
          6982 => x"7c",
          6983 => x"46",
          6984 => x"46",
          6985 => x"32",
          6986 => x"eb",
          6987 => x"53",
          6988 => x"35",
          6989 => x"4e",
          6990 => x"41",
          6991 => x"20",
          6992 => x"41",
          6993 => x"20",
          6994 => x"4e",
          6995 => x"41",
          6996 => x"20",
          6997 => x"41",
          6998 => x"20",
          6999 => x"00",
          7000 => x"00",
          7001 => x"00",
          7002 => x"00",
          7003 => x"80",
          7004 => x"8e",
          7005 => x"45",
          7006 => x"49",
          7007 => x"90",
          7008 => x"99",
          7009 => x"59",
          7010 => x"9c",
          7011 => x"41",
          7012 => x"a5",
          7013 => x"a8",
          7014 => x"ac",
          7015 => x"b0",
          7016 => x"b4",
          7017 => x"b8",
          7018 => x"bc",
          7019 => x"c0",
          7020 => x"c4",
          7021 => x"c8",
          7022 => x"cc",
          7023 => x"d0",
          7024 => x"d4",
          7025 => x"d8",
          7026 => x"dc",
          7027 => x"e0",
          7028 => x"e4",
          7029 => x"e8",
          7030 => x"ec",
          7031 => x"f0",
          7032 => x"f4",
          7033 => x"f8",
          7034 => x"fc",
          7035 => x"2b",
          7036 => x"3d",
          7037 => x"5c",
          7038 => x"3c",
          7039 => x"7f",
          7040 => x"00",
          7041 => x"00",
          7042 => x"01",
          7043 => x"00",
          7044 => x"00",
          7045 => x"00",
          7046 => x"00",
          7047 => x"00",
          7048 => x"64",
          7049 => x"74",
          7050 => x"64",
          7051 => x"74",
          7052 => x"66",
          7053 => x"74",
          7054 => x"66",
          7055 => x"64",
          7056 => x"66",
          7057 => x"63",
          7058 => x"6d",
          7059 => x"61",
          7060 => x"6d",
          7061 => x"79",
          7062 => x"6d",
          7063 => x"66",
          7064 => x"6d",
          7065 => x"70",
          7066 => x"6d",
          7067 => x"6d",
          7068 => x"6d",
          7069 => x"68",
          7070 => x"68",
          7071 => x"68",
          7072 => x"68",
          7073 => x"63",
          7074 => x"00",
          7075 => x"6a",
          7076 => x"72",
          7077 => x"61",
          7078 => x"72",
          7079 => x"74",
          7080 => x"69",
          7081 => x"00",
          7082 => x"74",
          7083 => x"00",
          7084 => x"74",
          7085 => x"69",
          7086 => x"6d",
          7087 => x"69",
          7088 => x"6b",
          7089 => x"00",
          7090 => x"44",
          7091 => x"20",
          7092 => x"6f",
          7093 => x"49",
          7094 => x"72",
          7095 => x"20",
          7096 => x"6f",
          7097 => x"00",
          7098 => x"44",
          7099 => x"20",
          7100 => x"20",
          7101 => x"64",
          7102 => x"00",
          7103 => x"4e",
          7104 => x"69",
          7105 => x"66",
          7106 => x"64",
          7107 => x"4e",
          7108 => x"61",
          7109 => x"66",
          7110 => x"64",
          7111 => x"49",
          7112 => x"6c",
          7113 => x"66",
          7114 => x"6e",
          7115 => x"2e",
          7116 => x"41",
          7117 => x"73",
          7118 => x"65",
          7119 => x"64",
          7120 => x"46",
          7121 => x"20",
          7122 => x"65",
          7123 => x"20",
          7124 => x"73",
          7125 => x"0a",
          7126 => x"46",
          7127 => x"20",
          7128 => x"64",
          7129 => x"69",
          7130 => x"6c",
          7131 => x"0a",
          7132 => x"53",
          7133 => x"73",
          7134 => x"69",
          7135 => x"70",
          7136 => x"65",
          7137 => x"64",
          7138 => x"44",
          7139 => x"65",
          7140 => x"6d",
          7141 => x"20",
          7142 => x"69",
          7143 => x"6c",
          7144 => x"0a",
          7145 => x"44",
          7146 => x"20",
          7147 => x"20",
          7148 => x"62",
          7149 => x"2e",
          7150 => x"4e",
          7151 => x"6f",
          7152 => x"74",
          7153 => x"65",
          7154 => x"6c",
          7155 => x"73",
          7156 => x"20",
          7157 => x"6e",
          7158 => x"6e",
          7159 => x"73",
          7160 => x"00",
          7161 => x"46",
          7162 => x"61",
          7163 => x"62",
          7164 => x"65",
          7165 => x"00",
          7166 => x"54",
          7167 => x"6f",
          7168 => x"20",
          7169 => x"72",
          7170 => x"6f",
          7171 => x"61",
          7172 => x"6c",
          7173 => x"2e",
          7174 => x"46",
          7175 => x"20",
          7176 => x"6c",
          7177 => x"65",
          7178 => x"00",
          7179 => x"49",
          7180 => x"66",
          7181 => x"69",
          7182 => x"20",
          7183 => x"6f",
          7184 => x"0a",
          7185 => x"54",
          7186 => x"6d",
          7187 => x"20",
          7188 => x"6e",
          7189 => x"6c",
          7190 => x"0a",
          7191 => x"50",
          7192 => x"6d",
          7193 => x"72",
          7194 => x"6e",
          7195 => x"72",
          7196 => x"2e",
          7197 => x"53",
          7198 => x"65",
          7199 => x"0a",
          7200 => x"55",
          7201 => x"6f",
          7202 => x"65",
          7203 => x"72",
          7204 => x"0a",
          7205 => x"20",
          7206 => x"65",
          7207 => x"73",
          7208 => x"20",
          7209 => x"20",
          7210 => x"65",
          7211 => x"65",
          7212 => x"00",
          7213 => x"72",
          7214 => x"00",
          7215 => x"25",
          7216 => x"00",
          7217 => x"3a",
          7218 => x"25",
          7219 => x"00",
          7220 => x"20",
          7221 => x"20",
          7222 => x"00",
          7223 => x"25",
          7224 => x"00",
          7225 => x"20",
          7226 => x"20",
          7227 => x"7c",
          7228 => x"7a",
          7229 => x"0a",
          7230 => x"25",
          7231 => x"00",
          7232 => x"31",
          7233 => x"34",
          7234 => x"32",
          7235 => x"76",
          7236 => x"31",
          7237 => x"20",
          7238 => x"2c",
          7239 => x"76",
          7240 => x"32",
          7241 => x"25",
          7242 => x"73",
          7243 => x"0a",
          7244 => x"5a",
          7245 => x"49",
          7246 => x"72",
          7247 => x"74",
          7248 => x"6e",
          7249 => x"72",
          7250 => x"54",
          7251 => x"72",
          7252 => x"74",
          7253 => x"75",
          7254 => x"00",
          7255 => x"50",
          7256 => x"69",
          7257 => x"72",
          7258 => x"74",
          7259 => x"49",
          7260 => x"4c",
          7261 => x"20",
          7262 => x"65",
          7263 => x"70",
          7264 => x"49",
          7265 => x"4c",
          7266 => x"20",
          7267 => x"65",
          7268 => x"70",
          7269 => x"55",
          7270 => x"30",
          7271 => x"20",
          7272 => x"65",
          7273 => x"70",
          7274 => x"55",
          7275 => x"30",
          7276 => x"20",
          7277 => x"65",
          7278 => x"70",
          7279 => x"55",
          7280 => x"31",
          7281 => x"20",
          7282 => x"65",
          7283 => x"70",
          7284 => x"55",
          7285 => x"31",
          7286 => x"20",
          7287 => x"65",
          7288 => x"70",
          7289 => x"53",
          7290 => x"69",
          7291 => x"75",
          7292 => x"69",
          7293 => x"2e",
          7294 => x"00",
          7295 => x"45",
          7296 => x"6c",
          7297 => x"20",
          7298 => x"65",
          7299 => x"2e",
          7300 => x"61",
          7301 => x"65",
          7302 => x"2e",
          7303 => x"00",
          7304 => x"30",
          7305 => x"46",
          7306 => x"65",
          7307 => x"6f",
          7308 => x"69",
          7309 => x"6c",
          7310 => x"20",
          7311 => x"63",
          7312 => x"20",
          7313 => x"70",
          7314 => x"73",
          7315 => x"6e",
          7316 => x"6d",
          7317 => x"61",
          7318 => x"2e",
          7319 => x"2a",
          7320 => x"43",
          7321 => x"72",
          7322 => x"2e",
          7323 => x"00",
          7324 => x"43",
          7325 => x"69",
          7326 => x"2e",
          7327 => x"43",
          7328 => x"61",
          7329 => x"67",
          7330 => x"00",
          7331 => x"25",
          7332 => x"78",
          7333 => x"38",
          7334 => x"3e",
          7335 => x"6c",
          7336 => x"30",
          7337 => x"0a",
          7338 => x"44",
          7339 => x"20",
          7340 => x"6f",
          7341 => x"00",
          7342 => x"0a",
          7343 => x"70",
          7344 => x"65",
          7345 => x"25",
          7346 => x"20",
          7347 => x"58",
          7348 => x"3f",
          7349 => x"00",
          7350 => x"25",
          7351 => x"20",
          7352 => x"58",
          7353 => x"25",
          7354 => x"20",
          7355 => x"58",
          7356 => x"45",
          7357 => x"75",
          7358 => x"67",
          7359 => x"64",
          7360 => x"20",
          7361 => x"78",
          7362 => x"2e",
          7363 => x"43",
          7364 => x"69",
          7365 => x"63",
          7366 => x"20",
          7367 => x"30",
          7368 => x"2e",
          7369 => x"00",
          7370 => x"43",
          7371 => x"20",
          7372 => x"75",
          7373 => x"64",
          7374 => x"64",
          7375 => x"25",
          7376 => x"0a",
          7377 => x"52",
          7378 => x"61",
          7379 => x"6e",
          7380 => x"70",
          7381 => x"63",
          7382 => x"6f",
          7383 => x"2e",
          7384 => x"43",
          7385 => x"20",
          7386 => x"6f",
          7387 => x"6e",
          7388 => x"2e",
          7389 => x"5a",
          7390 => x"62",
          7391 => x"25",
          7392 => x"25",
          7393 => x"73",
          7394 => x"00",
          7395 => x"25",
          7396 => x"25",
          7397 => x"73",
          7398 => x"25",
          7399 => x"25",
          7400 => x"42",
          7401 => x"63",
          7402 => x"61",
          7403 => x"0a",
          7404 => x"52",
          7405 => x"69",
          7406 => x"2e",
          7407 => x"45",
          7408 => x"6c",
          7409 => x"20",
          7410 => x"65",
          7411 => x"70",
          7412 => x"2e",
          7413 => x"00",
          7414 => x"00",
          7415 => x"00",
          7416 => x"00",
          7417 => x"00",
          7418 => x"00",
          7419 => x"00",
          7420 => x"00",
          7421 => x"00",
          7422 => x"01",
          7423 => x"01",
          7424 => x"00",
          7425 => x"00",
          7426 => x"00",
          7427 => x"00",
          7428 => x"05",
          7429 => x"05",
          7430 => x"05",
          7431 => x"00",
          7432 => x"01",
          7433 => x"01",
          7434 => x"01",
          7435 => x"01",
          7436 => x"00",
          7437 => x"00",
          7438 => x"00",
          7439 => x"00",
          7440 => x"00",
          7441 => x"00",
          7442 => x"00",
          7443 => x"00",
          7444 => x"00",
          7445 => x"00",
          7446 => x"00",
          7447 => x"00",
          7448 => x"00",
          7449 => x"00",
          7450 => x"00",
          7451 => x"00",
          7452 => x"00",
          7453 => x"00",
          7454 => x"00",
          7455 => x"00",
          7456 => x"00",
          7457 => x"00",
          7458 => x"00",
          7459 => x"00",
          7460 => x"00",
          7461 => x"00",
          7462 => x"00",
          7463 => x"00",
          7464 => x"00",
          7465 => x"00",
          7466 => x"00",
          7467 => x"00",
          7468 => x"01",
          7469 => x"00",
          7470 => x"01",
          7471 => x"00",
          7472 => x"02",
          7473 => x"01",
          7474 => x"00",
          7475 => x"00",
          7476 => x"01",
          7477 => x"00",
          7478 => x"00",
          7479 => x"00",
          7480 => x"01",
          7481 => x"00",
          7482 => x"00",
          7483 => x"00",
          7484 => x"01",
          7485 => x"00",
          7486 => x"00",
          7487 => x"00",
          7488 => x"01",
          7489 => x"00",
          7490 => x"00",
          7491 => x"00",
          7492 => x"01",
          7493 => x"00",
          7494 => x"00",
          7495 => x"00",
          7496 => x"01",
          7497 => x"00",
          7498 => x"00",
          7499 => x"00",
          7500 => x"01",
          7501 => x"00",
          7502 => x"00",
          7503 => x"00",
          7504 => x"01",
          7505 => x"00",
          7506 => x"00",
          7507 => x"00",
          7508 => x"01",
          7509 => x"00",
          7510 => x"00",
          7511 => x"00",
          7512 => x"01",
          7513 => x"00",
          7514 => x"00",
          7515 => x"00",
          7516 => x"01",
          7517 => x"00",
          7518 => x"00",
          7519 => x"00",
          7520 => x"01",
          7521 => x"00",
          7522 => x"00",
          7523 => x"00",
          7524 => x"01",
          7525 => x"00",
          7526 => x"00",
          7527 => x"00",
          7528 => x"01",
          7529 => x"00",
          7530 => x"00",
          7531 => x"00",
          7532 => x"01",
          7533 => x"00",
          7534 => x"00",
          7535 => x"00",
          7536 => x"01",
          7537 => x"00",
          7538 => x"00",
          7539 => x"00",
          7540 => x"01",
          7541 => x"00",
          7542 => x"00",
          7543 => x"00",
          7544 => x"01",
          7545 => x"00",
          7546 => x"00",
          7547 => x"00",
          7548 => x"01",
          7549 => x"00",
          7550 => x"00",
          7551 => x"00",
          7552 => x"01",
          7553 => x"00",
          7554 => x"00",
          7555 => x"00",
          7556 => x"01",
          7557 => x"00",
          7558 => x"00",
          7559 => x"00",
          7560 => x"01",
          7561 => x"00",
          7562 => x"00",
          7563 => x"00",
          7564 => x"01",
          7565 => x"00",
          7566 => x"00",
          7567 => x"00",
          7568 => x"01",
          7569 => x"00",
          7570 => x"00",
          7571 => x"00",
          7572 => x"01",
          7573 => x"00",
          7574 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
