-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use pkgs.config_pkg.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b80c4",
             1 => x"800b0b0b",
             2 => x"80ca9504",
             3 => x"ffffffff",
             4 => x"ffffffff",
             5 => x"ffffffff",
             6 => x"ffffffff",
             7 => x"ffffffff",
             8 => x"0b0b80c4",
             9 => x"80040b0b",
            10 => x"80c48504",
            11 => x"0b0b80c4",
            12 => x"95040b0b",
            13 => x"80c4a504",
            14 => x"0b0b80c4",
            15 => x"b5040b0b",
            16 => x"80c4c504",
            17 => x"0b0b80c4",
            18 => x"d5040b0b",
            19 => x"80c4e504",
            20 => x"0b0b80c4",
            21 => x"f5040b0b",
            22 => x"80c58504",
            23 => x"0b0b80c5",
            24 => x"95040b0b",
            25 => x"80c5a504",
            26 => x"0b0b80c5",
            27 => x"b5040b0b",
            28 => x"80c5c504",
            29 => x"0b0b80c5",
            30 => x"d5040b0b",
            31 => x"80c5e504",
            32 => x"0b0b80c5",
            33 => x"f5040b0b",
            34 => x"80c68504",
            35 => x"0b0b80c6",
            36 => x"95040b0b",
            37 => x"80c6a504",
            38 => x"0b0b80c6",
            39 => x"b5040b0b",
            40 => x"80c6c504",
            41 => x"0b0b80c6",
            42 => x"d5040b0b",
            43 => x"80c6e504",
            44 => x"0b0b80c6",
            45 => x"f5040b0b",
            46 => x"80c78504",
            47 => x"0b0b80c7",
            48 => x"95040b0b",
            49 => x"80c7a504",
            50 => x"0b0b80c7",
            51 => x"b5040b0b",
            52 => x"80c7c504",
            53 => x"0b0b80c7",
            54 => x"d5040b0b",
            55 => x"80c7e504",
            56 => x"0b0b80c7",
            57 => x"f5040b0b",
            58 => x"80c88504",
            59 => x"0b0b80c8",
            60 => x"95040b0b",
            61 => x"80c8a504",
            62 => x"0b0b80c8",
            63 => x"b5040b0b",
            64 => x"80c8c504",
            65 => x"0b0b80c8",
            66 => x"d5040b0b",
            67 => x"80c8e504",
            68 => x"0b0b80c8",
            69 => x"f5040b0b",
            70 => x"80c98504",
            71 => x"0b0b80c9",
            72 => x"95040b0b",
            73 => x"80c9a504",
            74 => x"0b0b80c9",
            75 => x"b5040b0b",
            76 => x"80c9c504",
            77 => x"0b0b80c9",
            78 => x"d5040b0b",
            79 => x"80c9e504",
            80 => x"0b0b80c9",
            81 => x"f5040b0b",
            82 => x"80ca8504",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"00000000",
            89 => x"00000000",
            90 => x"00000000",
            91 => x"00000000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"00000000",
            97 => x"00000000",
            98 => x"00000000",
            99 => x"00000000",
           100 => x"00000000",
           101 => x"00000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"00000000",
           105 => x"00000000",
           106 => x"00000000",
           107 => x"00000000",
           108 => x"00000000",
           109 => x"00000000",
           110 => x"00000000",
           111 => x"00000000",
           112 => x"00000000",
           113 => x"00000000",
           114 => x"00000000",
           115 => x"00000000",
           116 => x"00000000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"00000000",
           121 => x"00000000",
           122 => x"00000000",
           123 => x"00000000",
           124 => x"00000000",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"0080c480",
           129 => x"048293d4",
           130 => x"0c80d580",
           131 => x"2d8293d4",
           132 => x"08838090",
           133 => x"048293d4",
           134 => x"0c80dfc0",
           135 => x"2d8293d4",
           136 => x"08838090",
           137 => x"048293d4",
           138 => x"0c80e085",
           139 => x"2d8293d4",
           140 => x"08838090",
           141 => x"048293d4",
           142 => x"0c80e0a3",
           143 => x"2d8293d4",
           144 => x"08838090",
           145 => x"048293d4",
           146 => x"0c80e6f7",
           147 => x"2d8293d4",
           148 => x"08838090",
           149 => x"048293d4",
           150 => x"0c80e88b",
           151 => x"2d8293d4",
           152 => x"08838090",
           153 => x"048293d4",
           154 => x"0c80e0c4",
           155 => x"2d8293d4",
           156 => x"08838090",
           157 => x"048293d4",
           158 => x"0c80e8a8",
           159 => x"2d8293d4",
           160 => x"08838090",
           161 => x"048293d4",
           162 => x"0c80eabe",
           163 => x"2d8293d4",
           164 => x"08838090",
           165 => x"048293d4",
           166 => x"0c80e69d",
           167 => x"2d8293d4",
           168 => x"08838090",
           169 => x"048293d4",
           170 => x"0c80e6b3",
           171 => x"2d8293d4",
           172 => x"08838090",
           173 => x"048293d4",
           174 => x"0c80e6d7",
           175 => x"2d8293d4",
           176 => x"08838090",
           177 => x"048293d4",
           178 => x"0c80d780",
           179 => x"2d8293d4",
           180 => x"08838090",
           181 => x"048293d4",
           182 => x"0c80d7ce",
           183 => x"2d8293d4",
           184 => x"08838090",
           185 => x"048293d4",
           186 => x"0c80cfd8",
           187 => x"2d8293d4",
           188 => x"08838090",
           189 => x"048293d4",
           190 => x"0c80d190",
           191 => x"2d8293d4",
           192 => x"08838090",
           193 => x"048293d4",
           194 => x"0c80d2ea",
           195 => x"2d8293d4",
           196 => x"08838090",
           197 => x"048293d4",
           198 => x"0c819ef2",
           199 => x"2d8293d4",
           200 => x"08838090",
           201 => x"048293d4",
           202 => x"0c81ade9",
           203 => x"2d8293d4",
           204 => x"08838090",
           205 => x"048293d4",
           206 => x"0c81a3f8",
           207 => x"2d8293d4",
           208 => x"08838090",
           209 => x"048293d4",
           210 => x"0c81a7df",
           211 => x"2d8293d4",
           212 => x"08838090",
           213 => x"048293d4",
           214 => x"0c81b392",
           215 => x"2d8293d4",
           216 => x"08838090",
           217 => x"048293d4",
           218 => x"0c81bd86",
           219 => x"2d8293d4",
           220 => x"08838090",
           221 => x"048293d4",
           222 => x"0c81ac9a",
           223 => x"2d8293d4",
           224 => x"08838090",
           225 => x"048293d4",
           226 => x"0c81b7bd",
           227 => x"2d8293d4",
           228 => x"08838090",
           229 => x"048293d4",
           230 => x"0c81b8e1",
           231 => x"2d8293d4",
           232 => x"08838090",
           233 => x"048293d4",
           234 => x"0c81b98a",
           235 => x"2d8293d4",
           236 => x"08838090",
           237 => x"048293d4",
           238 => x"0c81c29a",
           239 => x"2d8293d4",
           240 => x"08838090",
           241 => x"048293d4",
           242 => x"0c81bf92",
           243 => x"2d8293d4",
           244 => x"08838090",
           245 => x"048293d4",
           246 => x"0c81c4f3",
           247 => x"2d8293d4",
           248 => x"08838090",
           249 => x"048293d4",
           250 => x"0c81ba80",
           251 => x"2d8293d4",
           252 => x"08838090",
           253 => x"048293d4",
           254 => x"0c81c7f7",
           255 => x"2d8293d4",
           256 => x"08838090",
           257 => x"048293d4",
           258 => x"0c81c8fd",
           259 => x"2d8293d4",
           260 => x"08838090",
           261 => x"048293d4",
           262 => x"0c81aec9",
           263 => x"2d8293d4",
           264 => x"08838090",
           265 => x"048293d4",
           266 => x"0c81aea2",
           267 => x"2d8293d4",
           268 => x"08838090",
           269 => x"048293d4",
           270 => x"0c81afcc",
           271 => x"2d8293d4",
           272 => x"08838090",
           273 => x"048293d4",
           274 => x"0c81bada",
           275 => x"2d8293d4",
           276 => x"08838090",
           277 => x"048293d4",
           278 => x"0c81c9f6",
           279 => x"2d8293d4",
           280 => x"08838090",
           281 => x"048293d4",
           282 => x"0c81cc81",
           283 => x"2d8293d4",
           284 => x"08838090",
           285 => x"048293d4",
           286 => x"0c81cfee",
           287 => x"2d8293d4",
           288 => x"08838090",
           289 => x"048293d4",
           290 => x"0c819e83",
           291 => x"2d8293d4",
           292 => x"08838090",
           293 => x"048293d4",
           294 => x"0c81d2df",
           295 => x"2d8293d4",
           296 => x"08838090",
           297 => x"048293d4",
           298 => x"0c80edfe",
           299 => x"2d8293d4",
           300 => x"08838090",
           301 => x"048293d4",
           302 => x"0c80efd7",
           303 => x"2d8293d4",
           304 => x"08838090",
           305 => x"048293d4",
           306 => x"0c80f1b1",
           307 => x"2d8293d4",
           308 => x"08838090",
           309 => x"048293d4",
           310 => x"0c80d081",
           311 => x"2d8293d4",
           312 => x"08838090",
           313 => x"048293d4",
           314 => x"0c80d0e6",
           315 => x"2d8293d4",
           316 => x"08838090",
           317 => x"048293d4",
           318 => x"0c80d3f3",
           319 => x"2d8293d4",
           320 => x"08838090",
           321 => x"048293d4",
           322 => x"0c81dfdd",
           323 => x"2d8293d4",
           324 => x"08838090",
           325 => x"048293c8",
           326 => x"7082b6cc",
           327 => x"278e3880",
           328 => x"71708405",
           329 => x"530c0b0b",
           330 => x"80ca9804",
           331 => x"80c48051",
           332 => x"81efda04",
           333 => x"3c048293",
           334 => x"d4080282",
           335 => x"93d40cfd",
           336 => x"3d0d8053",
           337 => x"8293d408",
           338 => x"8c050852",
           339 => x"8293d408",
           340 => x"88050851",
           341 => x"80c53f82",
           342 => x"93c80870",
           343 => x"8293c80c",
           344 => x"54853d0d",
           345 => x"8293d40c",
           346 => x"048293d4",
           347 => x"08028293",
           348 => x"d40cfd3d",
           349 => x"0d815382",
           350 => x"93d4088c",
           351 => x"05085282",
           352 => x"93d40888",
           353 => x"05085193",
           354 => x"3f8293c8",
           355 => x"08708293",
           356 => x"c80c5485",
           357 => x"3d0d8293",
           358 => x"d40c0482",
           359 => x"93d40802",
           360 => x"8293d40c",
           361 => x"fd3d0d81",
           362 => x"0b8293d4",
           363 => x"08fc050c",
           364 => x"800b8293",
           365 => x"d408f805",
           366 => x"0c8293d4",
           367 => x"088c0508",
           368 => x"8293d408",
           369 => x"88050827",
           370 => x"b9388293",
           371 => x"d408fc05",
           372 => x"08802eae",
           373 => x"38800b82",
           374 => x"93d4088c",
           375 => x"050824a2",
           376 => x"388293d4",
           377 => x"088c0508",
           378 => x"108293d4",
           379 => x"088c050c",
           380 => x"8293d408",
           381 => x"fc050810",
           382 => x"8293d408",
           383 => x"fc050cff",
           384 => x"b8398293",
           385 => x"d408fc05",
           386 => x"08802e80",
           387 => x"e1388293",
           388 => x"d4088c05",
           389 => x"088293d4",
           390 => x"08880508",
           391 => x"26ad3882",
           392 => x"93d40888",
           393 => x"05088293",
           394 => x"d4088c05",
           395 => x"08318293",
           396 => x"d4088805",
           397 => x"0c8293d4",
           398 => x"08f80508",
           399 => x"8293d408",
           400 => x"fc050807",
           401 => x"8293d408",
           402 => x"f8050c82",
           403 => x"93d408fc",
           404 => x"0508812a",
           405 => x"8293d408",
           406 => x"fc050c82",
           407 => x"93d4088c",
           408 => x"0508812a",
           409 => x"8293d408",
           410 => x"8c050cff",
           411 => x"95398293",
           412 => x"d4089005",
           413 => x"08802e93",
           414 => x"388293d4",
           415 => x"08880508",
           416 => x"708293d4",
           417 => x"08f4050c",
           418 => x"51913982",
           419 => x"93d408f8",
           420 => x"05087082",
           421 => x"93d408f4",
           422 => x"050c5182",
           423 => x"93d408f4",
           424 => x"05088293",
           425 => x"c80c853d",
           426 => x"0d8293d4",
           427 => x"0c04fc3d",
           428 => x"0d767971",
           429 => x"028c059f",
           430 => x"05335755",
           431 => x"53558372",
           432 => x"278a3874",
           433 => x"83065170",
           434 => x"802ea438",
           435 => x"ff125271",
           436 => x"ff2e9338",
           437 => x"73737081",
           438 => x"055534ff",
           439 => x"125271ff",
           440 => x"2e098106",
           441 => x"ef387482",
           442 => x"93c80c86",
           443 => x"3d0d0474",
           444 => x"74882b75",
           445 => x"07707190",
           446 => x"2b075154",
           447 => x"518f7227",
           448 => x"a5387271",
           449 => x"70840553",
           450 => x"0c727170",
           451 => x"8405530c",
           452 => x"72717084",
           453 => x"05530c72",
           454 => x"71708405",
           455 => x"530cf012",
           456 => x"52718f26",
           457 => x"dd388372",
           458 => x"27903872",
           459 => x"71708405",
           460 => x"530cfc12",
           461 => x"52718326",
           462 => x"f2387053",
           463 => x"ff8e39fb",
           464 => x"3d0d7779",
           465 => x"70720783",
           466 => x"06535452",
           467 => x"70933871",
           468 => x"73730854",
           469 => x"56547173",
           470 => x"082e80c6",
           471 => x"38737554",
           472 => x"52713370",
           473 => x"81ff0652",
           474 => x"5470802e",
           475 => x"9d387233",
           476 => x"5570752e",
           477 => x"09810695",
           478 => x"38811281",
           479 => x"14713370",
           480 => x"81ff0654",
           481 => x"56545270",
           482 => x"e5387233",
           483 => x"557381ff",
           484 => x"067581ff",
           485 => x"06717131",
           486 => x"8293c80c",
           487 => x"5252873d",
           488 => x"0d047109",
           489 => x"70f7fbfd",
           490 => x"ff140670",
           491 => x"f8848281",
           492 => x"80065151",
           493 => x"51709738",
           494 => x"84148416",
           495 => x"71085456",
           496 => x"54717508",
           497 => x"2edc3873",
           498 => x"755452ff",
           499 => x"9439800b",
           500 => x"8293c80c",
           501 => x"873d0d04",
           502 => x"fe3d0d80",
           503 => x"70545271",
           504 => x"882b5287",
           505 => x"9b3f8293",
           506 => x"c80881ff",
           507 => x"06720781",
           508 => x"14545283",
           509 => x"7325e838",
           510 => x"718293c8",
           511 => x"0c843d0d",
           512 => x"04fc3d0d",
           513 => x"76700870",
           514 => x"53555573",
           515 => x"802e80cd",
           516 => x"38733351",
           517 => x"70a02e09",
           518 => x"81068c38",
           519 => x"81147033",
           520 => x"525470a0",
           521 => x"2ef63873",
           522 => x"52843981",
           523 => x"12528072",
           524 => x"33525370",
           525 => x"a02e8338",
           526 => x"81537030",
           527 => x"709f2a74",
           528 => x"06515170",
           529 => x"e6387133",
           530 => x"5170a02e",
           531 => x"09810688",
           532 => x"38807270",
           533 => x"81055434",
           534 => x"71750c73",
           535 => x"51708293",
           536 => x"c80c863d",
           537 => x"0d04fc3d",
           538 => x"0d765372",
           539 => x"08802e91",
           540 => x"38863dfc",
           541 => x"05527251",
           542 => x"99c43f82",
           543 => x"93c80885",
           544 => x"38805383",
           545 => x"39745372",
           546 => x"8293c80c",
           547 => x"863d0d04",
           548 => x"f53d0d7d",
           549 => x"821133ff",
           550 => x"055b5c81",
           551 => x"5b798b26",
           552 => x"81bf3883",
           553 => x"1c33ff05",
           554 => x"5a825b79",
           555 => x"9e2681b1",
           556 => x"38841c33",
           557 => x"5a835b79",
           558 => x"972681a5",
           559 => x"38851c33",
           560 => x"5a845b79",
           561 => x"bb268199",
           562 => x"38861c33",
           563 => x"5a855b79",
           564 => x"bb26818d",
           565 => x"38881c22",
           566 => x"5a865b79",
           567 => x"87e72681",
           568 => x"80388a1c",
           569 => x"225a875b",
           570 => x"7987e726",
           571 => x"80f3388a",
           572 => x"1c225988",
           573 => x"1c225886",
           574 => x"1c335785",
           575 => x"1c335684",
           576 => x"1c335583",
           577 => x"1c335482",
           578 => x"1c33537b",
           579 => x"225281f6",
           580 => x"a8519489",
           581 => x"3f87c098",
           582 => x"9c5b817b",
           583 => x"0c7b2287",
           584 => x"c098bc0c",
           585 => x"821c3387",
           586 => x"c098b80c",
           587 => x"831c3387",
           588 => x"c098b40c",
           589 => x"841c3387",
           590 => x"c098b00c",
           591 => x"851c3387",
           592 => x"c098ac0c",
           593 => x"861c3387",
           594 => x"c098a80c",
           595 => x"881c2287",
           596 => x"c098a40c",
           597 => x"8a1c2287",
           598 => x"c098a00c",
           599 => x"807b0c80",
           600 => x"5b7a8293",
           601 => x"c80c8d3d",
           602 => x"0d04f53d",
           603 => x"0d7d5a87",
           604 => x"c0989c5c",
           605 => x"817c0c87",
           606 => x"c098bc08",
           607 => x"5b7a7a23",
           608 => x"87c098b8",
           609 => x"085b7a82",
           610 => x"1b3487c0",
           611 => x"98b4085b",
           612 => x"7a831b34",
           613 => x"87c098b0",
           614 => x"085b7a84",
           615 => x"1b3487c0",
           616 => x"98ac085b",
           617 => x"7a851b34",
           618 => x"87c098a8",
           619 => x"085b7a86",
           620 => x"1b3487c0",
           621 => x"98a4085b",
           622 => x"7a881b23",
           623 => x"87c098a0",
           624 => x"085b7a8a",
           625 => x"1b23807c",
           626 => x"0c8a1a22",
           627 => x"59881a22",
           628 => x"58861a33",
           629 => x"57851a33",
           630 => x"56841a33",
           631 => x"55831a33",
           632 => x"54821a33",
           633 => x"53792252",
           634 => x"81f6a851",
           635 => x"92af3f8d",
           636 => x"3d0d0480",
           637 => x"3d0d028b",
           638 => x"05337030",
           639 => x"709f2a51",
           640 => x"5151700b",
           641 => x"0b828bc0",
           642 => x"34823d0d",
           643 => x"04fd3d0d",
           644 => x"750b0b82",
           645 => x"8bc03354",
           646 => x"5487c094",
           647 => x"84517280",
           648 => x"2e863887",
           649 => x"c0949451",
           650 => x"70087096",
           651 => x"2a708106",
           652 => x"51525270",
           653 => x"802e8c38",
           654 => x"71912a70",
           655 => x"81065151",
           656 => x"70d73871",
           657 => x"962a8132",
           658 => x"70810651",
           659 => x"5170802e",
           660 => x"8d387193",
           661 => x"2a708106",
           662 => x"515170ff",
           663 => x"bc380b0b",
           664 => x"828bc033",
           665 => x"5187c094",
           666 => x"80527080",
           667 => x"2e863887",
           668 => x"c0949052",
           669 => x"73720c73",
           670 => x"8293c80c",
           671 => x"853d0d04",
           672 => x"fd3d0d02",
           673 => x"9705330b",
           674 => x"0b828bc0",
           675 => x"33545487",
           676 => x"c0948451",
           677 => x"72802e86",
           678 => x"3887c094",
           679 => x"94517008",
           680 => x"70962a70",
           681 => x"81065152",
           682 => x"5270802e",
           683 => x"8c387191",
           684 => x"2a708106",
           685 => x"515170d7",
           686 => x"3871962a",
           687 => x"81327081",
           688 => x"06515170",
           689 => x"802e8d38",
           690 => x"71932a70",
           691 => x"81065151",
           692 => x"70ffbc38",
           693 => x"0b0b828b",
           694 => x"c0335187",
           695 => x"c0948052",
           696 => x"70802e86",
           697 => x"3887c094",
           698 => x"90527372",
           699 => x"0c853d0d",
           700 => x"04fb3d0d",
           701 => x"77548074",
           702 => x"33525670",
           703 => x"762e80f7",
           704 => x"38737081",
           705 => x"0555330b",
           706 => x"0b828bc0",
           707 => x"33545587",
           708 => x"c0948451",
           709 => x"72802e86",
           710 => x"3887c094",
           711 => x"94517008",
           712 => x"70962a70",
           713 => x"81065152",
           714 => x"5270802e",
           715 => x"8c387191",
           716 => x"2a708106",
           717 => x"515170d7",
           718 => x"3871962a",
           719 => x"81327081",
           720 => x"06515170",
           721 => x"802e8d38",
           722 => x"71932a70",
           723 => x"81065151",
           724 => x"70ffbc38",
           725 => x"0b0b828b",
           726 => x"c0335187",
           727 => x"c0948052",
           728 => x"70802e86",
           729 => x"3887c094",
           730 => x"90527472",
           731 => x"0c811674",
           732 => x"33525670",
           733 => x"ff8b3875",
           734 => x"8293c80c",
           735 => x"873d0d04",
           736 => x"ff3d0d0b",
           737 => x"0b828bc0",
           738 => x"335287c0",
           739 => x"94845171",
           740 => x"802e8638",
           741 => x"87c09494",
           742 => x"51700870",
           743 => x"822a7081",
           744 => x"06515151",
           745 => x"70802ee2",
           746 => x"380b0b82",
           747 => x"8bc03351",
           748 => x"87c09480",
           749 => x"5270802e",
           750 => x"863887c0",
           751 => x"94905271",
           752 => x"087081ff",
           753 => x"068293c8",
           754 => x"0c51833d",
           755 => x"0d04ff3d",
           756 => x"0d0b0b82",
           757 => x"8bc03351",
           758 => x"87c09484",
           759 => x"5270802e",
           760 => x"863887c0",
           761 => x"94945271",
           762 => x"0870822a",
           763 => x"70810651",
           764 => x"5151ff52",
           765 => x"70802ea2",
           766 => x"380b0b82",
           767 => x"8bc03351",
           768 => x"87c09480",
           769 => x"5270802e",
           770 => x"863887c0",
           771 => x"94905271",
           772 => x"0870982b",
           773 => x"70982c51",
           774 => x"53517182",
           775 => x"93c80c83",
           776 => x"3d0d04fd",
           777 => x"3d0d87c0",
           778 => x"9e807008",
           779 => x"709c2a8a",
           780 => x"06515253",
           781 => x"70802e83",
           782 => x"9f38828b",
           783 => x"c40b87c0",
           784 => x"9e9c0871",
           785 => x"0c841187",
           786 => x"c09ea008",
           787 => x"710c5288",
           788 => x"1187c09e",
           789 => x"8c08710c",
           790 => x"528c1187",
           791 => x"c09e9008",
           792 => x"710c5290",
           793 => x"1187c09e",
           794 => x"9408710c",
           795 => x"52941187",
           796 => x"c09e9808",
           797 => x"710c5298",
           798 => x"1187c09e",
           799 => x"a408710c",
           800 => x"529c1187",
           801 => x"c09ea808",
           802 => x"710c52a0",
           803 => x"1187c09e",
           804 => x"ac08710c",
           805 => x"52730852",
           806 => x"5270a413",
           807 => x"23a81287",
           808 => x"c09e8408",
           809 => x"710c5181",
           810 => x"0bac1334",
           811 => x"ad125280",
           812 => x"0b87c09e",
           813 => x"880870a0",
           814 => x"80065152",
           815 => x"5370802e",
           816 => x"83388153",
           817 => x"72723480",
           818 => x"0b87c09e",
           819 => x"88087081",
           820 => x"80800651",
           821 => x"52527080",
           822 => x"2e833881",
           823 => x"5271828b",
           824 => x"f234800b",
           825 => x"87c09e88",
           826 => x"087080c0",
           827 => x"80065152",
           828 => x"5270802e",
           829 => x"83388152",
           830 => x"71828bf3",
           831 => x"34800b87",
           832 => x"c09e8808",
           833 => x"70908006",
           834 => x"51525270",
           835 => x"802e8338",
           836 => x"81527182",
           837 => x"8bf43480",
           838 => x"0b87c09e",
           839 => x"88087088",
           840 => x"80065152",
           841 => x"5270802e",
           842 => x"83388152",
           843 => x"71828bf5",
           844 => x"34800b87",
           845 => x"c09e8808",
           846 => x"70848006",
           847 => x"51525270",
           848 => x"802e8338",
           849 => x"81527182",
           850 => x"8bf63480",
           851 => x"0b87c09e",
           852 => x"88087082",
           853 => x"80065152",
           854 => x"5270802e",
           855 => x"83388152",
           856 => x"71828bf7",
           857 => x"34800b87",
           858 => x"c09e8808",
           859 => x"70818006",
           860 => x"51525270",
           861 => x"802e8338",
           862 => x"81527182",
           863 => x"8bf83482",
           864 => x"8bf95287",
           865 => x"c09e8870",
           866 => x"087080e0",
           867 => x"0670862c",
           868 => x"51515253",
           869 => x"70727081",
           870 => x"05543471",
           871 => x"54807308",
           872 => x"70900651",
           873 => x"52527080",
           874 => x"2e833881",
           875 => x"52717434",
           876 => x"800b87c0",
           877 => x"9e880870",
           878 => x"88065152",
           879 => x"5270802e",
           880 => x"83388152",
           881 => x"71828bfb",
           882 => x"3487c09e",
           883 => x"88087087",
           884 => x"06515170",
           885 => x"828bfc34",
           886 => x"853d0d04",
           887 => x"fc3d0d81",
           888 => x"f6c05184",
           889 => x"be3f828b",
           890 => x"f0335473",
           891 => x"802e8838",
           892 => x"81f6d451",
           893 => x"84ad3f81",
           894 => x"f6e85184",
           895 => x"a63f828b",
           896 => x"f1703355",
           897 => x"5573802e",
           898 => x"9138d715",
           899 => x"0853828b",
           900 => x"c4085281",
           901 => x"f780518a",
           902 => x"843f828b",
           903 => x"f2703355",
           904 => x"5573802e",
           905 => x"9038de15",
           906 => x"0853da15",
           907 => x"085281f7",
           908 => x"a85189e9",
           909 => x"3f828bf3",
           910 => x"70335555",
           911 => x"738a3881",
           912 => x"15335473",
           913 => x"802e9338",
           914 => x"828bd870",
           915 => x"0854fc11",
           916 => x"08535481",
           917 => x"f7cc5189",
           918 => x"c43f828b",
           919 => x"f5335473",
           920 => x"802e8838",
           921 => x"81f7f051",
           922 => x"83b93f82",
           923 => x"8bf63354",
           924 => x"73802e88",
           925 => x"3881f7fc",
           926 => x"5183a83f",
           927 => x"828bf733",
           928 => x"5473802e",
           929 => x"883881f8",
           930 => x"88518397",
           931 => x"3f828bf8",
           932 => x"70335555",
           933 => x"73802e8c",
           934 => x"38811533",
           935 => x"5281f894",
           936 => x"5188fa3f",
           937 => x"828bfa33",
           938 => x"5473802e",
           939 => x"883881f8",
           940 => x"b45182ef",
           941 => x"3f828bfb",
           942 => x"70335555",
           943 => x"73802e8c",
           944 => x"38811533",
           945 => x"5281f8d0",
           946 => x"5188d23f",
           947 => x"81f8ec51",
           948 => x"82d13f82",
           949 => x"8bdc7070",
           950 => x"70840552",
           951 => x"085481f8",
           952 => x"f8535555",
           953 => x"88b73f73",
           954 => x"085281f9",
           955 => x"a05188ad",
           956 => x"3f881508",
           957 => x"5281f9c8",
           958 => x"5188a23f",
           959 => x"8c152252",
           960 => x"81f9f051",
           961 => x"88973f90",
           962 => x"15085281",
           963 => x"fa985188",
           964 => x"8c3f863d",
           965 => x"0d04ff3d",
           966 => x"0d028e05",
           967 => x"33527185",
           968 => x"26bb3871",
           969 => x"10100b0b",
           970 => x"81f0c405",
           971 => x"52710804",
           972 => x"81fac051",
           973 => x"f7bb3fac",
           974 => x"3981fac8",
           975 => x"51f7b23f",
           976 => x"a33981fa",
           977 => x"d051f7a9",
           978 => x"3f9a3981",
           979 => x"fad851f7",
           980 => x"a03f9139",
           981 => x"81fadc51",
           982 => x"f7973f88",
           983 => x"3981fae4",
           984 => x"51f78e3f",
           985 => x"833d0d04",
           986 => x"7188800c",
           987 => x"04800b87",
           988 => x"c096840c",
           989 => x"04ff3d0d",
           990 => x"87c09684",
           991 => x"70085252",
           992 => x"80720c70",
           993 => x"74077082",
           994 => x"8c800c72",
           995 => x"0c833d0d",
           996 => x"04ff3d0d",
           997 => x"87c09684",
           998 => x"7008828c",
           999 => x"800c5280",
          1000 => x"720c7309",
          1001 => x"70828c80",
          1002 => x"08067082",
          1003 => x"8c800c73",
          1004 => x"0c51833d",
          1005 => x"0d04828c",
          1006 => x"800887c0",
          1007 => x"96840c04",
          1008 => x"fe3d0d02",
          1009 => x"93053353",
          1010 => x"728a2e09",
          1011 => x"81068538",
          1012 => x"8d51ed3f",
          1013 => x"8293e008",
          1014 => x"802e9538",
          1015 => x"8293e008",
          1016 => x"52727234",
          1017 => x"8293e008",
          1018 => x"81058293",
          1019 => x"e00c9239",
          1020 => x"8293d808",
          1021 => x"802e8a38",
          1022 => x"72518293",
          1023 => x"d8085271",
          1024 => x"2d843d0d",
          1025 => x"04fe3d0d",
          1026 => x"02970533",
          1027 => x"8293d808",
          1028 => x"768293d8",
          1029 => x"0c5451ff",
          1030 => x"a73f7282",
          1031 => x"93d80c84",
          1032 => x"3d0d04fe",
          1033 => x"3d0d7470",
          1034 => x"33535371",
          1035 => x"802e9138",
          1036 => x"72708105",
          1037 => x"543351ff",
          1038 => x"873f7233",
          1039 => x"5271f138",
          1040 => x"843d0d04",
          1041 => x"fd3d0d76",
          1042 => x"8293d808",
          1043 => x"778293d8",
          1044 => x"0c713354",
          1045 => x"55537180",
          1046 => x"2e913872",
          1047 => x"70810554",
          1048 => x"3351fedc",
          1049 => x"3f723352",
          1050 => x"71f13873",
          1051 => x"8293d80c",
          1052 => x"853d0d04",
          1053 => x"ec3d0d66",
          1054 => x"685d5978",
          1055 => x"7081055a",
          1056 => x"33567580",
          1057 => x"2e859238",
          1058 => x"75a52e88",
          1059 => x"387551fe",
          1060 => x"af3fe839",
          1061 => x"80707a70",
          1062 => x"81055c33",
          1063 => x"585e5a75",
          1064 => x"b02e0981",
          1065 => x"068c3881",
          1066 => x"79708105",
          1067 => x"5b33575d",
          1068 => x"923975ad",
          1069 => x"2e098106",
          1070 => x"8a388279",
          1071 => x"7081055b",
          1072 => x"33575d75",
          1073 => x"aa2e0981",
          1074 => x"0692387b",
          1075 => x"841d7108",
          1076 => x"7b708105",
          1077 => x"5d33595c",
          1078 => x"5d539f39",
          1079 => x"d0165372",
          1080 => x"89269738",
          1081 => x"798a2916",
          1082 => x"d0057970",
          1083 => x"81055b33",
          1084 => x"d0115557",
          1085 => x"5a897327",
          1086 => x"eb387580",
          1087 => x"ec327030",
          1088 => x"70720780",
          1089 => x"257880cc",
          1090 => x"32703070",
          1091 => x"72078025",
          1092 => x"73075359",
          1093 => x"52525454",
          1094 => x"73802e8c",
          1095 => x"387c8407",
          1096 => x"79708105",
          1097 => x"5b33575d",
          1098 => x"75802e83",
          1099 => x"ec387555",
          1100 => x"80e07627",
          1101 => x"8938e016",
          1102 => x"7081ff06",
          1103 => x"5653ffbe",
          1104 => x"15537296",
          1105 => x"26819838",
          1106 => x"72101081",
          1107 => x"f0dc0553",
          1108 => x"7208047b",
          1109 => x"841d7108",
          1110 => x"575d5380",
          1111 => x"75335454",
          1112 => x"72742e8d",
          1113 => x"38811470",
          1114 => x"16703351",
          1115 => x"545472f5",
          1116 => x"387c812a",
          1117 => x"70810651",
          1118 => x"5372a338",
          1119 => x"73811555",
          1120 => x"53727a27",
          1121 => x"99387c81",
          1122 => x"2a810656",
          1123 => x"a051fcb0",
          1124 => x"3f758b38",
          1125 => x"73811555",
          1126 => x"53797326",
          1127 => x"ef387451",
          1128 => x"fd813f73",
          1129 => x"81155553",
          1130 => x"727a27fd",
          1131 => x"ce38a051",
          1132 => x"fc8e3f73",
          1133 => x"81155553",
          1134 => x"797326f2",
          1135 => x"38fdbc39",
          1136 => x"7b841d83",
          1137 => x"1233535d",
          1138 => x"53fbf53f",
          1139 => x"fdad3982",
          1140 => x"5b953988",
          1141 => x"5b91398a",
          1142 => x"5b8d3990",
          1143 => x"5b893975",
          1144 => x"51fbdd3f",
          1145 => x"fd95397c",
          1146 => x"822a7081",
          1147 => x"06515372",
          1148 => x"802e8b38",
          1149 => x"7b841d71",
          1150 => x"08595d53",
          1151 => x"9c397480",
          1152 => x"c42e0981",
          1153 => x"068b387b",
          1154 => x"841d7108",
          1155 => x"595d5389",
          1156 => x"397b841d",
          1157 => x"7108595d",
          1158 => x"537480c4",
          1159 => x"32703070",
          1160 => x"72078025",
          1161 => x"70807b24",
          1162 => x"06515255",
          1163 => x"5372802e",
          1164 => x"88387630",
          1165 => x"7d90075e",
          1166 => x"5780587a",
          1167 => x"527651e6",
          1168 => x"a83f8293",
          1169 => x"c80881ff",
          1170 => x"067b5377",
          1171 => x"5255e5e6",
          1172 => x"3f8293c8",
          1173 => x"08578975",
          1174 => x"27993874",
          1175 => x"a7167081",
          1176 => x"ff065754",
          1177 => x"547580f8",
          1178 => x"2e893887",
          1179 => x"147081ff",
          1180 => x"06565396",
          1181 => x"3d7805e0",
          1182 => x"05b01654",
          1183 => x"54727434",
          1184 => x"81187730",
          1185 => x"7079079f",
          1186 => x"2a709f74",
          1187 => x"27065151",
          1188 => x"545872ff",
          1189 => x"a6387c84",
          1190 => x"2a708106",
          1191 => x"51537280",
          1192 => x"2e8e3896",
          1193 => x"3d7805e0",
          1194 => x"0553ad73",
          1195 => x"34811858",
          1196 => x"777d8106",
          1197 => x"5454b055",
          1198 => x"728338a0",
          1199 => x"557c812a",
          1200 => x"70810651",
          1201 => x"5372a338",
          1202 => x"73811555",
          1203 => x"53727a27",
          1204 => x"99387c81",
          1205 => x"2a810656",
          1206 => x"7451f9e4",
          1207 => x"3f758b38",
          1208 => x"73811555",
          1209 => x"53797326",
          1210 => x"ef38ff18",
          1211 => x"973de005",
          1212 => x"11703353",
          1213 => x"5458f9c8",
          1214 => x"3f77ef38",
          1215 => x"73811555",
          1216 => x"53727a27",
          1217 => x"faf538a0",
          1218 => x"51f9b53f",
          1219 => x"73811555",
          1220 => x"53797326",
          1221 => x"f238fae3",
          1222 => x"39963d0d",
          1223 => x"04fd3d0d",
          1224 => x"863d7070",
          1225 => x"84055208",
          1226 => x"55527351",
          1227 => x"fac63f85",
          1228 => x"3d0d04fe",
          1229 => x"3d0d7482",
          1230 => x"93e00c85",
          1231 => x"3d880552",
          1232 => x"7551fab0",
          1233 => x"3f8293e0",
          1234 => x"08538073",
          1235 => x"34800b82",
          1236 => x"93e00c84",
          1237 => x"3d0d04fd",
          1238 => x"3d0d8293",
          1239 => x"d8087682",
          1240 => x"93d80c87",
          1241 => x"3d880553",
          1242 => x"775253fa",
          1243 => x"873f7282",
          1244 => x"93d80c85",
          1245 => x"3d0d04fa",
          1246 => x"3d0d787a",
          1247 => x"57578053",
          1248 => x"8293dc08",
          1249 => x"732e80fa",
          1250 => x"38863973",
          1251 => x"5380f339",
          1252 => x"80558293",
          1253 => x"dc085271",
          1254 => x"2d8293c8",
          1255 => x"0881ff06",
          1256 => x"5473802e",
          1257 => x"e638738d",
          1258 => x"2e80ca38",
          1259 => x"73883270",
          1260 => x"30763070",
          1261 => x"78079f2a",
          1262 => x"72802506",
          1263 => x"52545153",
          1264 => x"72802e8e",
          1265 => x"38ff1574",
          1266 => x"81ff0652",
          1267 => x"55f7f13f",
          1268 => x"c1399f74",
          1269 => x"25ffbb38",
          1270 => x"ff165274",
          1271 => x"7225ffb2",
          1272 => x"38761552",
          1273 => x"73723481",
          1274 => x"157481ff",
          1275 => x"065255f7",
          1276 => x"cf3fff9e",
          1277 => x"39741752",
          1278 => x"8072348a",
          1279 => x"51f7c13f",
          1280 => x"81537282",
          1281 => x"93c80c88",
          1282 => x"3d0d04fe",
          1283 => x"3d0d8293",
          1284 => x"dc087582",
          1285 => x"93dc0c77",
          1286 => x"53765253",
          1287 => x"fed93f72",
          1288 => x"8293dc0c",
          1289 => x"843d0d04",
          1290 => x"f83d0d7a",
          1291 => x"7c5a5580",
          1292 => x"707a0c75",
          1293 => x"08703356",
          1294 => x"545873a0",
          1295 => x"2e098106",
          1296 => x"92387408",
          1297 => x"8105750c",
          1298 => x"74087033",
          1299 => x"555373a0",
          1300 => x"2ef03873",
          1301 => x"ad2e0981",
          1302 => x"068e3881",
          1303 => x"75081176",
          1304 => x"0c750870",
          1305 => x"33565458",
          1306 => x"73b02e09",
          1307 => x"810680d3",
          1308 => x"38740881",
          1309 => x"05750c74",
          1310 => x"08703355",
          1311 => x"537380e2",
          1312 => x"2e9a3873",
          1313 => x"80f82e09",
          1314 => x"8106a138",
          1315 => x"900b8114",
          1316 => x"760c7508",
          1317 => x"70335654",
          1318 => x"5780c139",
          1319 => x"82750881",
          1320 => x"05760c75",
          1321 => x"08703356",
          1322 => x"5457b139",
          1323 => x"8156a074",
          1324 => x"27818238",
          1325 => x"d0145380",
          1326 => x"56885789",
          1327 => x"73279d38",
          1328 => x"80f339d0",
          1329 => x"14538056",
          1330 => x"72892680",
          1331 => x"e8388b39",
          1332 => x"805680e1",
          1333 => x"39805680",
          1334 => x"dc398a57",
          1335 => x"8056a074",
          1336 => x"2780c538",
          1337 => x"80e07427",
          1338 => x"8938e014",
          1339 => x"7081ff06",
          1340 => x"5553d014",
          1341 => x"7081ff06",
          1342 => x"55539074",
          1343 => x"278e38f9",
          1344 => x"147081ff",
          1345 => x"06555389",
          1346 => x"7427c538",
          1347 => x"737727c5",
          1348 => x"38767629",
          1349 => x"14750881",
          1350 => x"05760c75",
          1351 => x"08703356",
          1352 => x"545673a0",
          1353 => x"26ffbd38",
          1354 => x"77802e84",
          1355 => x"38753056",
          1356 => x"75790c81",
          1357 => x"56758293",
          1358 => x"c80c8a3d",
          1359 => x"0d04f83d",
          1360 => x"0d7a7c5a",
          1361 => x"5580707a",
          1362 => x"0c750870",
          1363 => x"33565458",
          1364 => x"73a02e09",
          1365 => x"81069238",
          1366 => x"74088105",
          1367 => x"750c7408",
          1368 => x"70335553",
          1369 => x"73a02ef0",
          1370 => x"3873ad2e",
          1371 => x"0981068e",
          1372 => x"38817508",
          1373 => x"11760c75",
          1374 => x"08703356",
          1375 => x"545873b0",
          1376 => x"2e098106",
          1377 => x"80d33874",
          1378 => x"08810575",
          1379 => x"0c740870",
          1380 => x"33555373",
          1381 => x"80e22e9a",
          1382 => x"387380f8",
          1383 => x"2e098106",
          1384 => x"a138900b",
          1385 => x"8114760c",
          1386 => x"75087033",
          1387 => x"56545780",
          1388 => x"c1398275",
          1389 => x"08810576",
          1390 => x"0c750870",
          1391 => x"33565457",
          1392 => x"b1398156",
          1393 => x"a0742781",
          1394 => x"8238d014",
          1395 => x"53805688",
          1396 => x"57897327",
          1397 => x"9d3880f3",
          1398 => x"39d01453",
          1399 => x"80567289",
          1400 => x"2680e838",
          1401 => x"8b398056",
          1402 => x"80e13980",
          1403 => x"5680dc39",
          1404 => x"8a578056",
          1405 => x"a0742780",
          1406 => x"c53880e0",
          1407 => x"74278938",
          1408 => x"e0147081",
          1409 => x"ff065553",
          1410 => x"d0147081",
          1411 => x"ff065553",
          1412 => x"9074278e",
          1413 => x"38f91470",
          1414 => x"81ff0655",
          1415 => x"53897427",
          1416 => x"c5387377",
          1417 => x"27c53876",
          1418 => x"76291475",
          1419 => x"08810576",
          1420 => x"0c750870",
          1421 => x"33565456",
          1422 => x"73a026ff",
          1423 => x"bd387780",
          1424 => x"2e843875",
          1425 => x"30567579",
          1426 => x"0c815675",
          1427 => x"8293c80c",
          1428 => x"8a3d0d04",
          1429 => x"ff3d0d02",
          1430 => x"8f053351",
          1431 => x"81527072",
          1432 => x"26873882",
          1433 => x"8c841133",
          1434 => x"52718293",
          1435 => x"c80c833d",
          1436 => x"0d04fd3d",
          1437 => x"0d029705",
          1438 => x"33028405",
          1439 => x"9b053355",
          1440 => x"53835172",
          1441 => x"812680ed",
          1442 => x"38729029",
          1443 => x"87c0928c",
          1444 => x"05518852",
          1445 => x"73802e84",
          1446 => x"38818852",
          1447 => x"71710c72",
          1448 => x"902987c0",
          1449 => x"928c0551",
          1450 => x"81710c85",
          1451 => x"0b87c098",
          1452 => x"8c0c7052",
          1453 => x"87c0988c",
          1454 => x"54710870",
          1455 => x"82065151",
          1456 => x"70802e87",
          1457 => x"38730851",
          1458 => x"70ef3872",
          1459 => x"902987c0",
          1460 => x"928c0570",
          1461 => x"08fc8080",
          1462 => x"06535171",
          1463 => x"923887c0",
          1464 => x"988c0851",
          1465 => x"70802e87",
          1466 => x"3871828c",
          1467 => x"84143482",
          1468 => x"8c841333",
          1469 => x"51708293",
          1470 => x"c80c853d",
          1471 => x"0d04f23d",
          1472 => x"0d616365",
          1473 => x"028c0580",
          1474 => x"c3053356",
          1475 => x"415d5883",
          1476 => x"73525bfe",
          1477 => x"bf3f8293",
          1478 => x"c8088106",
          1479 => x"7b555271",
          1480 => x"81ac3880",
          1481 => x"70585d87",
          1482 => x"c0988c73",
          1483 => x"842b87c0",
          1484 => x"928c1187",
          1485 => x"c0928412",
          1486 => x"72425c57",
          1487 => x"5b568576",
          1488 => x"0c87c092",
          1489 => x"801a7c71",
          1490 => x"0c528475",
          1491 => x"0c740870",
          1492 => x"852a7081",
          1493 => x"06515354",
          1494 => x"71802e8e",
          1495 => x"38780852",
          1496 => x"71787081",
          1497 => x"055a3481",
          1498 => x"175773a2",
          1499 => x"06527180",
          1500 => x"2e873875",
          1501 => x"085271d5",
          1502 => x"38750852",
          1503 => x"71802e87",
          1504 => x"38768480",
          1505 => x"2e993881",
          1506 => x"750c87c0",
          1507 => x"928c1e53",
          1508 => x"72087082",
          1509 => x"06515271",
          1510 => x"f738ff1b",
          1511 => x"5b8d3984",
          1512 => x"801c811e",
          1513 => x"7081ff06",
          1514 => x"5f535c7a",
          1515 => x"802e9038",
          1516 => x"73fc8080",
          1517 => x"06527187",
          1518 => x"387e7d26",
          1519 => x"ff803873",
          1520 => x"fc808006",
          1521 => x"5271802e",
          1522 => x"83388152",
          1523 => x"71547382",
          1524 => x"93c80c90",
          1525 => x"3d0d04f3",
          1526 => x"3d0d6062",
          1527 => x"64028c05",
          1528 => x"bf053356",
          1529 => x"405c5783",
          1530 => x"73525afc",
          1531 => x"e73f8293",
          1532 => x"c8088106",
          1533 => x"7a555271",
          1534 => x"81ae3880",
          1535 => x"5c87c098",
          1536 => x"8c73842b",
          1537 => x"87c0928c",
          1538 => x"1187c092",
          1539 => x"84127241",
          1540 => x"5b575a56",
          1541 => x"85760c87",
          1542 => x"c0928019",
          1543 => x"7b710c52",
          1544 => x"82750c80",
          1545 => x"53740870",
          1546 => x"842a7081",
          1547 => x"06515354",
          1548 => x"71802e8c",
          1549 => x"38767081",
          1550 => x"05583378",
          1551 => x"0c811353",
          1552 => x"73812a70",
          1553 => x"81065152",
          1554 => x"71802e87",
          1555 => x"38750852",
          1556 => x"71d33875",
          1557 => x"08527180",
          1558 => x"2e873872",
          1559 => x"84802e99",
          1560 => x"3881750c",
          1561 => x"87c0928c",
          1562 => x"1d537208",
          1563 => x"70820651",
          1564 => x"5271f738",
          1565 => x"ff1a5a8d",
          1566 => x"39811c70",
          1567 => x"81ff0684",
          1568 => x"801d5d5d",
          1569 => x"5279802e",
          1570 => x"903873fc",
          1571 => x"80800652",
          1572 => x"7187387d",
          1573 => x"7c26fefc",
          1574 => x"3873fc80",
          1575 => x"80065271",
          1576 => x"802e8338",
          1577 => x"81527154",
          1578 => x"738293c8",
          1579 => x"0c8f3d0d",
          1580 => x"04f73d0d",
          1581 => x"7d028405",
          1582 => x"af053302",
          1583 => x"8805b305",
          1584 => x"33715455",
          1585 => x"5656fb8c",
          1586 => x"3f8293c8",
          1587 => x"08810652",
          1588 => x"835471bc",
          1589 => x"38815472",
          1590 => x"742ea238",
          1591 => x"72742488",
          1592 => x"3872802e",
          1593 => x"8a38a739",
          1594 => x"72832e9a",
          1595 => x"38a03974",
          1596 => x"902987c0",
          1597 => x"928c0570",
          1598 => x"08515294",
          1599 => x"3988800a",
          1600 => x"760c8054",
          1601 => x"8b398180",
          1602 => x"760c8054",
          1603 => x"83398454",
          1604 => x"738293c8",
          1605 => x"0c8b3d0d",
          1606 => x"04ff3d0d",
          1607 => x"73703381",
          1608 => x"12337088",
          1609 => x"2b720782",
          1610 => x"93c80c52",
          1611 => x"5252833d",
          1612 => x"0d04fd3d",
          1613 => x"0d758311",
          1614 => x"33821233",
          1615 => x"71902b71",
          1616 => x"882b0781",
          1617 => x"14337107",
          1618 => x"74337188",
          1619 => x"2b078293",
          1620 => x"c80c5154",
          1621 => x"56545285",
          1622 => x"3d0d04ff",
          1623 => x"3d0d7302",
          1624 => x"84059205",
          1625 => x"22525270",
          1626 => x"72708105",
          1627 => x"54347088",
          1628 => x"2a517072",
          1629 => x"34833d0d",
          1630 => x"04ff3d0d",
          1631 => x"73755252",
          1632 => x"70727081",
          1633 => x"05543470",
          1634 => x"882a5170",
          1635 => x"72708105",
          1636 => x"54347088",
          1637 => x"2a517072",
          1638 => x"70810554",
          1639 => x"3470882a",
          1640 => x"51707234",
          1641 => x"833d0d04",
          1642 => x"fe3d0d76",
          1643 => x"75775454",
          1644 => x"5170802e",
          1645 => x"93387170",
          1646 => x"81055333",
          1647 => x"73708105",
          1648 => x"5534ff11",
          1649 => x"5170ef38",
          1650 => x"843d0d04",
          1651 => x"fe3d0d75",
          1652 => x"77765452",
          1653 => x"53727270",
          1654 => x"81055434",
          1655 => x"ff115170",
          1656 => x"f438843d",
          1657 => x"0d04fc3d",
          1658 => x"0d787779",
          1659 => x"56565374",
          1660 => x"70810556",
          1661 => x"33747081",
          1662 => x"05563371",
          1663 => x"7131ff16",
          1664 => x"56525252",
          1665 => x"72802e86",
          1666 => x"3871802e",
          1667 => x"e2387182",
          1668 => x"93c80c86",
          1669 => x"3d0d04fe",
          1670 => x"3d0d7476",
          1671 => x"71335354",
          1672 => x"5270802e",
          1673 => x"99387073",
          1674 => x"2e943881",
          1675 => x"12703352",
          1676 => x"5270802e",
          1677 => x"89387073",
          1678 => x"2e098106",
          1679 => x"ee387133",
          1680 => x"8293c80c",
          1681 => x"843d0d04",
          1682 => x"800b8293",
          1683 => x"c80c0480",
          1684 => x"0b8293c8",
          1685 => x"0c04f93d",
          1686 => x"0d795680",
          1687 => x"0b831733",
          1688 => x"56587478",
          1689 => x"2e80d738",
          1690 => x"8154b016",
          1691 => x"0853b416",
          1692 => x"70538117",
          1693 => x"335257fa",
          1694 => x"de3f8293",
          1695 => x"c808782e",
          1696 => x"098106b8",
          1697 => x"388293c8",
          1698 => x"08831734",
          1699 => x"b01608a4",
          1700 => x"17083155",
          1701 => x"749c1708",
          1702 => x"27a43882",
          1703 => x"16335574",
          1704 => x"822e0981",
          1705 => x"06983881",
          1706 => x"54b01608",
          1707 => x"9c170805",
          1708 => x"53765281",
          1709 => x"163351fa",
          1710 => x"9e3f8339",
          1711 => x"81587782",
          1712 => x"93c80c89",
          1713 => x"3d0d04fa",
          1714 => x"3d0d787a",
          1715 => x"56578056",
          1716 => x"b0170875",
          1717 => x"2eaf3876",
          1718 => x"51fefb3f",
          1719 => x"8293c808",
          1720 => x"568293c8",
          1721 => x"089f3881",
          1722 => x"547453b4",
          1723 => x"17528117",
          1724 => x"3351f88a",
          1725 => x"3f8293c8",
          1726 => x"08802e85",
          1727 => x"38ff5581",
          1728 => x"5674b018",
          1729 => x"0c758293",
          1730 => x"c80c883d",
          1731 => x"0d04f83d",
          1732 => x"0d7a7052",
          1733 => x"57febf3f",
          1734 => x"8293c808",
          1735 => x"588293c8",
          1736 => x"08819138",
          1737 => x"76335574",
          1738 => x"832e0981",
          1739 => x"0680f038",
          1740 => x"84173359",
          1741 => x"78812e09",
          1742 => x"810680e3",
          1743 => x"38848053",
          1744 => x"8293c808",
          1745 => x"52b41770",
          1746 => x"5256fd80",
          1747 => x"3f82d4d5",
          1748 => x"5284b217",
          1749 => x"51fc843f",
          1750 => x"848b85a4",
          1751 => x"d2527551",
          1752 => x"fc973f86",
          1753 => x"8a85e4f2",
          1754 => x"52849817",
          1755 => x"51fc8a3f",
          1756 => x"90170852",
          1757 => x"849c1751",
          1758 => x"fbff3f8c",
          1759 => x"17085284",
          1760 => x"a01751fb",
          1761 => x"f43fa017",
          1762 => x"08810570",
          1763 => x"b0190c79",
          1764 => x"55537552",
          1765 => x"81173351",
          1766 => x"f8bd3f77",
          1767 => x"84183480",
          1768 => x"53805281",
          1769 => x"173351fa",
          1770 => x"883f8293",
          1771 => x"c808802e",
          1772 => x"83388158",
          1773 => x"778293c8",
          1774 => x"0c8a3d0d",
          1775 => x"04fb3d0d",
          1776 => x"77fe1a98",
          1777 => x"1208fe05",
          1778 => x"55565480",
          1779 => x"56747327",
          1780 => x"8d388a14",
          1781 => x"22707629",
          1782 => x"ac160805",
          1783 => x"57537582",
          1784 => x"93c80c87",
          1785 => x"3d0d04f9",
          1786 => x"3d0d7a7a",
          1787 => x"70085654",
          1788 => x"55817527",
          1789 => x"88389814",
          1790 => x"08752686",
          1791 => x"38815681",
          1792 => x"d939ff74",
          1793 => x"33545672",
          1794 => x"822e80f5",
          1795 => x"38728224",
          1796 => x"89387281",
          1797 => x"2e8d3881",
          1798 => x"bf397283",
          1799 => x"2e818e38",
          1800 => x"81b63974",
          1801 => x"812a1570",
          1802 => x"892aa416",
          1803 => x"08055374",
          1804 => x"5257fd93",
          1805 => x"3f8293c8",
          1806 => x"08819f38",
          1807 => x"7683ff06",
          1808 => x"14b41133",
          1809 => x"81197089",
          1810 => x"2aa41808",
          1811 => x"05557654",
          1812 => x"595953fc",
          1813 => x"f23f8293",
          1814 => x"c80880fe",
          1815 => x"387683ff",
          1816 => x"0614b411",
          1817 => x"3370882b",
          1818 => x"7a077781",
          1819 => x"0671842a",
          1820 => x"5a525a51",
          1821 => x"537280e2",
          1822 => x"38779fff",
          1823 => x"065680da",
          1824 => x"3974882a",
          1825 => x"a4150805",
          1826 => x"527351fc",
          1827 => x"ba3f8293",
          1828 => x"c80880c6",
          1829 => x"38741583",
          1830 => x"ff067405",
          1831 => x"b40551f8",
          1832 => x"f83f8293",
          1833 => x"c80883ff",
          1834 => x"ff0656ae",
          1835 => x"3974872a",
          1836 => x"a4150805",
          1837 => x"527351fc",
          1838 => x"8e3f8293",
          1839 => x"c8089b38",
          1840 => x"74822b83",
          1841 => x"fc067405",
          1842 => x"b40551f8",
          1843 => x"e53f8293",
          1844 => x"c808f00a",
          1845 => x"06568339",
          1846 => x"81567582",
          1847 => x"93c80c89",
          1848 => x"3d0d04f7",
          1849 => x"3d0d7b7d",
          1850 => x"7f585555",
          1851 => x"82578174",
          1852 => x"2782af38",
          1853 => x"73981608",
          1854 => x"2782a738",
          1855 => x"74335372",
          1856 => x"772e81a8",
          1857 => x"38727724",
          1858 => x"89387281",
          1859 => x"2e8d3882",
          1860 => x"91397283",
          1861 => x"2e81c938",
          1862 => x"82883973",
          1863 => x"812a1470",
          1864 => x"892aa417",
          1865 => x"08055375",
          1866 => x"5259fb9b",
          1867 => x"3f8293c8",
          1868 => x"08578293",
          1869 => x"c80881ea",
          1870 => x"387883ff",
          1871 => x"0615b411",
          1872 => x"811b7681",
          1873 => x"06565b51",
          1874 => x"58755772",
          1875 => x"802e8f38",
          1876 => x"75842b9f",
          1877 => x"f0067833",
          1878 => x"8f067107",
          1879 => x"58537678",
          1880 => x"34810b83",
          1881 => x"16347889",
          1882 => x"2aa41608",
          1883 => x"05527451",
          1884 => x"fad53f82",
          1885 => x"93c80857",
          1886 => x"8293c808",
          1887 => x"81a43878",
          1888 => x"83ff0615",
          1889 => x"b4117581",
          1890 => x"0678842a",
          1891 => x"57555158",
          1892 => x"728f3875",
          1893 => x"882a7833",
          1894 => x"578f0676",
          1895 => x"81f00607",
          1896 => x"54737834",
          1897 => x"810b8316",
          1898 => x"3480f739",
          1899 => x"73882aa4",
          1900 => x"16080552",
          1901 => x"7451fa8f",
          1902 => x"3f8293c8",
          1903 => x"08578293",
          1904 => x"c80880de",
          1905 => x"387583ff",
          1906 => x"ff065273",
          1907 => x"1483ff06",
          1908 => x"7505b405",
          1909 => x"51f7843f",
          1910 => x"810b8316",
          1911 => x"3480c339",
          1912 => x"73872aa4",
          1913 => x"16080552",
          1914 => x"7451f9db",
          1915 => x"3f8293c8",
          1916 => x"08578293",
          1917 => x"c808ab38",
          1918 => x"75f00a06",
          1919 => x"74822b83",
          1920 => x"fc067611",
          1921 => x"b4057054",
          1922 => x"515456f6",
          1923 => x"a53f8293",
          1924 => x"c8088f0a",
          1925 => x"06760752",
          1926 => x"7251f6dd",
          1927 => x"3f810b83",
          1928 => x"16347682",
          1929 => x"93c80c8b",
          1930 => x"3d0d04f9",
          1931 => x"3d0d797b",
          1932 => x"7d720858",
          1933 => x"58555781",
          1934 => x"74278838",
          1935 => x"98150874",
          1936 => x"26863882",
          1937 => x"56818e39",
          1938 => x"75802eaa",
          1939 => x"38ff5375",
          1940 => x"527451fd",
          1941 => x"8e3f8293",
          1942 => x"c8085682",
          1943 => x"93c80880",
          1944 => x"f4389339",
          1945 => x"825680ed",
          1946 => x"39815680",
          1947 => x"e8398293",
          1948 => x"c8085680",
          1949 => x"e0397352",
          1950 => x"7651faeb",
          1951 => x"3f8293c8",
          1952 => x"08568293",
          1953 => x"c808802e",
          1954 => x"80c93882",
          1955 => x"93c80881",
          1956 => x"2ed23882",
          1957 => x"93c808ff",
          1958 => x"2ecf3880",
          1959 => x"53735274",
          1960 => x"51fcc03f",
          1961 => x"8293c808",
          1962 => x"c5389815",
          1963 => x"08fe0554",
          1964 => x"90150874",
          1965 => x"27933890",
          1966 => x"15088105",
          1967 => x"90160c84",
          1968 => x"15338107",
          1969 => x"54738416",
          1970 => x"34755498",
          1971 => x"15087626",
          1972 => x"ffa43880",
          1973 => x"56758293",
          1974 => x"c80c893d",
          1975 => x"0d04f53d",
          1976 => x"0d7d7f71",
          1977 => x"085b5c5c",
          1978 => x"7a95388c",
          1979 => x"19085877",
          1980 => x"802e8838",
          1981 => x"98190878",
          1982 => x"26b73881",
          1983 => x"58b3397a",
          1984 => x"527b51f9",
          1985 => x"e23f8155",
          1986 => x"748293c8",
          1987 => x"082782e9",
          1988 => x"388293c8",
          1989 => x"08558293",
          1990 => x"c808ff2e",
          1991 => x"82db3882",
          1992 => x"93c80855",
          1993 => x"98190882",
          1994 => x"93c80826",
          1995 => x"82cb387a",
          1996 => x"58805590",
          1997 => x"1908752e",
          1998 => x"82bf3880",
          1999 => x"57777b2e",
          2000 => x"09810680",
          2001 => x"db38811b",
          2002 => x"57981908",
          2003 => x"77268338",
          2004 => x"82577652",
          2005 => x"7b51f98f",
          2006 => x"3f8293c8",
          2007 => x"0856805a",
          2008 => x"8293c808",
          2009 => x"812e0981",
          2010 => x"06863882",
          2011 => x"93c8085a",
          2012 => x"75ff3270",
          2013 => x"30707207",
          2014 => x"8025707d",
          2015 => x"07795351",
          2016 => x"52565473",
          2017 => x"81f33875",
          2018 => x"802e9538",
          2019 => x"8c190856",
          2020 => x"8176278a",
          2021 => x"3875981a",
          2022 => x"08278338",
          2023 => x"75588057",
          2024 => x"7680de38",
          2025 => x"77578117",
          2026 => x"57981908",
          2027 => x"77268938",
          2028 => x"82577678",
          2029 => x"2681b638",
          2030 => x"76527b51",
          2031 => x"f8a93f82",
          2032 => x"93c80856",
          2033 => x"8293c808",
          2034 => x"802eb638",
          2035 => x"805a8293",
          2036 => x"c808812e",
          2037 => x"09810686",
          2038 => x"388293c8",
          2039 => x"085a75ff",
          2040 => x"32703070",
          2041 => x"72078025",
          2042 => x"707d0751",
          2043 => x"52565473",
          2044 => x"80ff3876",
          2045 => x"782e0981",
          2046 => x"06ffab38",
          2047 => x"805580f9",
          2048 => x"39ff5376",
          2049 => x"527851f9",
          2050 => x"da3f8293",
          2051 => x"c8088293",
          2052 => x"c8083070",
          2053 => x"8293c808",
          2054 => x"0780257d",
          2055 => x"30707f07",
          2056 => x"9f2a7206",
          2057 => x"52575156",
          2058 => x"5674802e",
          2059 => x"8f387653",
          2060 => x"7a527851",
          2061 => x"f9ad3f82",
          2062 => x"93c80856",
          2063 => x"75a63876",
          2064 => x"8c1a0c98",
          2065 => x"1908fe05",
          2066 => x"54901908",
          2067 => x"74268938",
          2068 => x"901908ff",
          2069 => x"05901a0c",
          2070 => x"84193381",
          2071 => x"07547384",
          2072 => x"1a349439",
          2073 => x"ff577581",
          2074 => x"2e8d3889",
          2075 => x"39805589",
          2076 => x"39755585",
          2077 => x"39815776",
          2078 => x"55748293",
          2079 => x"c80c8d3d",
          2080 => x"0d04f73d",
          2081 => x"0d7b7052",
          2082 => x"57f3cb3f",
          2083 => x"81558293",
          2084 => x"c80880db",
          2085 => x"387c5276",
          2086 => x"51f6a23f",
          2087 => x"8293c808",
          2088 => x"8293c808",
          2089 => x"b0190c5a",
          2090 => x"84805380",
          2091 => x"52b41770",
          2092 => x"5255f298",
          2093 => x"3f745981",
          2094 => x"58805684",
          2095 => x"39771656",
          2096 => x"8a172255",
          2097 => x"75752797",
          2098 => x"38775475",
          2099 => x"1a537852",
          2100 => x"81173351",
          2101 => x"ee813f82",
          2102 => x"93c80880",
          2103 => x"2edf3880",
          2104 => x"0b8a1822",
          2105 => x"56587476",
          2106 => x"2e833881",
          2107 => x"58775574",
          2108 => x"8293c80c",
          2109 => x"8b3d0d04",
          2110 => x"f83d0d7a",
          2111 => x"7c710858",
          2112 => x"565774f0",
          2113 => x"800a268a",
          2114 => x"38749f06",
          2115 => x"5372802e",
          2116 => x"86388258",
          2117 => x"81ae3974",
          2118 => x"90180c88",
          2119 => x"17085473",
          2120 => x"aa387533",
          2121 => x"53827327",
          2122 => x"8538a816",
          2123 => x"0854739b",
          2124 => x"3874852a",
          2125 => x"53820b88",
          2126 => x"17225a58",
          2127 => x"72792781",
          2128 => x"8338a816",
          2129 => x"0898180c",
          2130 => x"80d1398a",
          2131 => x"16227089",
          2132 => x"2b545872",
          2133 => x"7526b638",
          2134 => x"73527651",
          2135 => x"f5893f82",
          2136 => x"93c80854",
          2137 => x"8293c808",
          2138 => x"ff2ebf38",
          2139 => x"810b8293",
          2140 => x"c808278b",
          2141 => x"38981608",
          2142 => x"8293c808",
          2143 => x"26863882",
          2144 => x"5880c139",
          2145 => x"74733155",
          2146 => x"747327cc",
          2147 => x"38735275",
          2148 => x"51f4aa3f",
          2149 => x"8293c808",
          2150 => x"98180c73",
          2151 => x"94180c82",
          2152 => x"58981708",
          2153 => x"802e9d38",
          2154 => x"85398158",
          2155 => x"97397489",
          2156 => x"2a981808",
          2157 => x"0598180c",
          2158 => x"7483ff06",
          2159 => x"16b4059c",
          2160 => x"180c8058",
          2161 => x"778293c8",
          2162 => x"0c8a3d0d",
          2163 => x"04f93d0d",
          2164 => x"797b7108",
          2165 => x"901308a0",
          2166 => x"05595959",
          2167 => x"55f0800a",
          2168 => x"76278638",
          2169 => x"800b9816",
          2170 => x"0c845398",
          2171 => x"1508802e",
          2172 => x"81da3875",
          2173 => x"83ff0654",
          2174 => x"7381c138",
          2175 => x"98150881",
          2176 => x"0598160c",
          2177 => x"94150898",
          2178 => x"3875852a",
          2179 => x"88182259",
          2180 => x"53777326",
          2181 => x"81a63873",
          2182 => x"98160c84",
          2183 => x"5381ad39",
          2184 => x"8a1722ff",
          2185 => x"1177892a",
          2186 => x"06515372",
          2187 => x"818e3894",
          2188 => x"15085274",
          2189 => x"51f3b03f",
          2190 => x"8293c808",
          2191 => x"54825381",
          2192 => x"0b8293c8",
          2193 => x"08278184",
          2194 => x"38815382",
          2195 => x"93c808ff",
          2196 => x"2e80f938",
          2197 => x"98170882",
          2198 => x"93c80826",
          2199 => x"80cc3877",
          2200 => x"8a387798",
          2201 => x"160c8453",
          2202 => x"80e23994",
          2203 => x"15085274",
          2204 => x"51f8eb3f",
          2205 => x"8293c808",
          2206 => x"54875382",
          2207 => x"93c80880",
          2208 => x"2e80c938",
          2209 => x"82538293",
          2210 => x"c808812e",
          2211 => x"bf388153",
          2212 => x"8293c808",
          2213 => x"ff2eb538",
          2214 => x"8293c808",
          2215 => x"527651fb",
          2216 => x"e13f8153",
          2217 => x"8293c808",
          2218 => x"a3387394",
          2219 => x"160c7352",
          2220 => x"7651f289",
          2221 => x"3f8293c8",
          2222 => x"0898160c",
          2223 => x"7590160c",
          2224 => x"7583ff06",
          2225 => x"17b4059c",
          2226 => x"160c8053",
          2227 => x"728293c8",
          2228 => x"0c893d0d",
          2229 => x"04f83d0d",
          2230 => x"7a7c7108",
          2231 => x"5a5a5680",
          2232 => x"527551fc",
          2233 => x"933f8293",
          2234 => x"c8085482",
          2235 => x"93c80880",
          2236 => x"e1388293",
          2237 => x"c8085798",
          2238 => x"16085277",
          2239 => x"51efc83f",
          2240 => x"8293c808",
          2241 => x"548293c8",
          2242 => x"0880c738",
          2243 => x"8293c808",
          2244 => x"9c170870",
          2245 => x"33515455",
          2246 => x"7281e52e",
          2247 => x"09810683",
          2248 => x"38815572",
          2249 => x"30708025",
          2250 => x"76075153",
          2251 => x"72802e8b",
          2252 => x"38811757",
          2253 => x"76792e9a",
          2254 => x"38833980",
          2255 => x"57815275",
          2256 => x"51fd8a3f",
          2257 => x"8293c808",
          2258 => x"548293c8",
          2259 => x"08802eff",
          2260 => x"a6387384",
          2261 => x"2e098106",
          2262 => x"83388754",
          2263 => x"738293c8",
          2264 => x"0c8a3d0d",
          2265 => x"04fd3d0d",
          2266 => x"769a1152",
          2267 => x"54ebaa3f",
          2268 => x"8293c808",
          2269 => x"83ffff06",
          2270 => x"76703351",
          2271 => x"53537183",
          2272 => x"2e098106",
          2273 => x"90389414",
          2274 => x"51eb8e3f",
          2275 => x"8293c808",
          2276 => x"902b7307",
          2277 => x"53728293",
          2278 => x"c80c853d",
          2279 => x"0d04fc3d",
          2280 => x"0d777970",
          2281 => x"83ffff06",
          2282 => x"549a1253",
          2283 => x"5555ebab",
          2284 => x"3f767033",
          2285 => x"51537283",
          2286 => x"2e098106",
          2287 => x"8b387390",
          2288 => x"2a529415",
          2289 => x"51eb943f",
          2290 => x"863d0d04",
          2291 => x"f73d0d7b",
          2292 => x"7d5b5684",
          2293 => x"76085a58",
          2294 => x"98160880",
          2295 => x"2e818638",
          2296 => x"98160852",
          2297 => x"7851eddf",
          2298 => x"3f8293c8",
          2299 => x"08588293",
          2300 => x"c80880f1",
          2301 => x"389c1608",
          2302 => x"70335653",
          2303 => x"74863884",
          2304 => x"5880e239",
          2305 => x"9c16088b",
          2306 => x"113370bf",
          2307 => x"067081ff",
          2308 => x"065a5151",
          2309 => x"53728617",
          2310 => x"347481e5",
          2311 => x"32703076",
          2312 => x"ae327030",
          2313 => x"7073069f",
          2314 => x"2a535155",
          2315 => x"51547380",
          2316 => x"2e9b3876",
          2317 => x"8f2e9638",
          2318 => x"8077df06",
          2319 => x"54547288",
          2320 => x"2e098106",
          2321 => x"83388154",
          2322 => x"737a2e99",
          2323 => x"38805275",
          2324 => x"51fafa3f",
          2325 => x"8293c808",
          2326 => x"588293c8",
          2327 => x"08873898",
          2328 => x"1608fefc",
          2329 => x"3877802e",
          2330 => x"8638800b",
          2331 => x"98170c77",
          2332 => x"8293c80c",
          2333 => x"8b3d0d04",
          2334 => x"f83d0d7a",
          2335 => x"70085956",
          2336 => x"80527551",
          2337 => x"f8f23f82",
          2338 => x"93c80854",
          2339 => x"8293c808",
          2340 => x"80ef3886",
          2341 => x"39845780",
          2342 => x"e6399816",
          2343 => x"08527751",
          2344 => x"eca53f82",
          2345 => x"93c80857",
          2346 => x"8293c808",
          2347 => x"80d1389c",
          2348 => x"16087033",
          2349 => x"51547380",
          2350 => x"2edb389c",
          2351 => x"16088b11",
          2352 => x"33bf0655",
          2353 => x"55738617",
          2354 => x"348b1533",
          2355 => x"70832a70",
          2356 => x"81065155",
          2357 => x"59739338",
          2358 => x"8b53a016",
          2359 => x"527451ea",
          2360 => x"853f8293",
          2361 => x"c808802e",
          2362 => x"96388052",
          2363 => x"7551f9dd",
          2364 => x"3f8293c8",
          2365 => x"08578293",
          2366 => x"c808802e",
          2367 => x"ff9c3876",
          2368 => x"54738293",
          2369 => x"c80c8a3d",
          2370 => x"0d04fb3d",
          2371 => x"0d777008",
          2372 => x"57548152",
          2373 => x"7351fbbd",
          2374 => x"3f8293c8",
          2375 => x"08558293",
          2376 => x"c808b438",
          2377 => x"98140852",
          2378 => x"7551eb9b",
          2379 => x"3f8293c8",
          2380 => x"08558293",
          2381 => x"c808a038",
          2382 => x"a0538293",
          2383 => x"c808529c",
          2384 => x"140851e9",
          2385 => x"873f8b53",
          2386 => x"a014529c",
          2387 => x"140851e8",
          2388 => x"d73f810b",
          2389 => x"83173474",
          2390 => x"8293c80c",
          2391 => x"873d0d04",
          2392 => x"fc3d0d76",
          2393 => x"70089812",
          2394 => x"08547053",
          2395 => x"5653ead7",
          2396 => x"3f8293c8",
          2397 => x"08548293",
          2398 => x"c8088d38",
          2399 => x"9c130853",
          2400 => x"e5733481",
          2401 => x"0b831634",
          2402 => x"738293c8",
          2403 => x"0c863d0d",
          2404 => x"04fa3d0d",
          2405 => x"787a5757",
          2406 => x"800b8917",
          2407 => x"34981708",
          2408 => x"802e8189",
          2409 => x"38807055",
          2410 => x"559c1708",
          2411 => x"14703381",
          2412 => x"16565452",
          2413 => x"72a02ead",
          2414 => x"3872852e",
          2415 => x"09810684",
          2416 => x"3881e553",
          2417 => x"73892e09",
          2418 => x"81068e38",
          2419 => x"75158805",
          2420 => x"52ae0b81",
          2421 => x"13348115",
          2422 => x"55751588",
          2423 => x"05527281",
          2424 => x"13348115",
          2425 => x"558a7427",
          2426 => x"c0387515",
          2427 => x"88055280",
          2428 => x"0b811334",
          2429 => x"9c170852",
          2430 => x"8b123388",
          2431 => x"17349c17",
          2432 => x"089c0551",
          2433 => x"e6ac3f82",
          2434 => x"93c80876",
          2435 => x"0c9c1708",
          2436 => x"960551e6",
          2437 => x"843f8293",
          2438 => x"c8088617",
          2439 => x"239c1708",
          2440 => x"980551e5",
          2441 => x"f43f8293",
          2442 => x"c8088417",
          2443 => x"23883d0d",
          2444 => x"04f53d0d",
          2445 => x"7e70087f",
          2446 => x"a0055d5a",
          2447 => x"5c8b53a0",
          2448 => x"527a51e7",
          2449 => x"873f8070",
          2450 => x"58588879",
          2451 => x"33555a73",
          2452 => x"ae2e0981",
          2453 => x"0680df38",
          2454 => x"78177033",
          2455 => x"811971ae",
          2456 => x"32703070",
          2457 => x"9f2a7382",
          2458 => x"26075151",
          2459 => x"53595754",
          2460 => x"738c387a",
          2461 => x"18547574",
          2462 => x"34811858",
          2463 => x"db3975af",
          2464 => x"32703077",
          2465 => x"80dc3270",
          2466 => x"30707306",
          2467 => x"9f2a5351",
          2468 => x"56515574",
          2469 => x"802e8938",
          2470 => x"865475a0",
          2471 => x"2682e438",
          2472 => x"76197c0c",
          2473 => x"a454a076",
          2474 => x"278338a0",
          2475 => x"54738b1c",
          2476 => x"34805482",
          2477 => x"ce397817",
          2478 => x"70338119",
          2479 => x"595754a0",
          2480 => x"7627828c",
          2481 => x"3875af32",
          2482 => x"70307780",
          2483 => x"dc327030",
          2484 => x"72802571",
          2485 => x"80250753",
          2486 => x"51565155",
          2487 => x"74802eb5",
          2488 => x"38843981",
          2489 => x"17578077",
          2490 => x"1a703351",
          2491 => x"555a73af",
          2492 => x"2e098106",
          2493 => x"8338815a",
          2494 => x"80771a70",
          2495 => x"33515555",
          2496 => x"7380dc2e",
          2497 => x"09810683",
          2498 => x"38815579",
          2499 => x"75075473",
          2500 => x"d23881bc",
          2501 => x"3975ae32",
          2502 => x"70307080",
          2503 => x"257a7d27",
          2504 => x"07515154",
          2505 => x"73802ea2",
          2506 => x"38798b32",
          2507 => x"703077ae",
          2508 => x"32703072",
          2509 => x"8025719f",
          2510 => x"2a075351",
          2511 => x"56515574",
          2512 => x"81b13888",
          2513 => x"588b5afe",
          2514 => x"ed397598",
          2515 => x"2b547380",
          2516 => x"258c3875",
          2517 => x"80ff0681",
          2518 => x"fbf81133",
          2519 => x"57547551",
          2520 => x"e5e63f82",
          2521 => x"93c80880",
          2522 => x"2eb93878",
          2523 => x"17703381",
          2524 => x"19715459",
          2525 => x"5654e5d7",
          2526 => x"3f8293c8",
          2527 => x"08802e89",
          2528 => x"38ff1a54",
          2529 => x"73782686",
          2530 => x"38865480",
          2531 => x"f6397a18",
          2532 => x"54757434",
          2533 => x"81187b11",
          2534 => x"55587474",
          2535 => x"34811858",
          2536 => x"fe943975",
          2537 => x"5281faf0",
          2538 => x"51e4ec3f",
          2539 => x"8293c808",
          2540 => x"80c538ff",
          2541 => x"9f165473",
          2542 => x"99268938",
          2543 => x"e0167081",
          2544 => x"ff065754",
          2545 => x"7a185475",
          2546 => x"74348118",
          2547 => x"58fde739",
          2548 => x"76197c0c",
          2549 => x"86547780",
          2550 => x"2ea9387a",
          2551 => x"33547381",
          2552 => x"e52e0981",
          2553 => x"06843885",
          2554 => x"7b348454",
          2555 => x"a076278d",
          2556 => x"38893986",
          2557 => x"548d3986",
          2558 => x"54893980",
          2559 => x"54738b1c",
          2560 => x"34805473",
          2561 => x"8293c80c",
          2562 => x"8d3d0d04",
          2563 => x"fa3d0d78",
          2564 => x"70085856",
          2565 => x"807a7033",
          2566 => x"51545572",
          2567 => x"af2e8338",
          2568 => x"8155807a",
          2569 => x"70335154",
          2570 => x"547280dc",
          2571 => x"2e833881",
          2572 => x"54747406",
          2573 => x"5372802e",
          2574 => x"8c389417",
          2575 => x"0888170c",
          2576 => x"b339811a",
          2577 => x"5a807a70",
          2578 => x"33515455",
          2579 => x"72af2e09",
          2580 => x"81068338",
          2581 => x"8155807a",
          2582 => x"70335154",
          2583 => x"547280dc",
          2584 => x"2e098106",
          2585 => x"83388154",
          2586 => x"74740753",
          2587 => x"72d43880",
          2588 => x"0b88170c",
          2589 => x"79703351",
          2590 => x"53729f26",
          2591 => x"9b38ff80",
          2592 => x"0bab1734",
          2593 => x"80527551",
          2594 => x"f0ee3f82",
          2595 => x"93c80855",
          2596 => x"81aa3985",
          2597 => x"5581a539",
          2598 => x"893d8405",
          2599 => x"527551fb",
          2600 => x"903f8293",
          2601 => x"c8085582",
          2602 => x"93c80881",
          2603 => x"8f387551",
          2604 => x"f7c63f82",
          2605 => x"93c808ab",
          2606 => x"17335555",
          2607 => x"8293c808",
          2608 => x"802e80c2",
          2609 => x"388293c8",
          2610 => x"08842e09",
          2611 => x"810680ec",
          2612 => x"3873852a",
          2613 => x"70810651",
          2614 => x"5372802e",
          2615 => x"9a387382",
          2616 => x"2a708106",
          2617 => x"51537280",
          2618 => x"2effad38",
          2619 => x"ff800bab",
          2620 => x"17348055",
          2621 => x"80c63973",
          2622 => x"822a7081",
          2623 => x"06515372",
          2624 => x"bb388555",
          2625 => x"b7397382",
          2626 => x"2a708106",
          2627 => x"515372ac",
          2628 => x"38861633",
          2629 => x"70842a70",
          2630 => x"81065154",
          2631 => x"5472802e",
          2632 => x"fef13890",
          2633 => x"160883ff",
          2634 => x"0617b405",
          2635 => x"527651f4",
          2636 => x"b43f8293",
          2637 => x"c8088817",
          2638 => x"0cfedd39",
          2639 => x"748293c8",
          2640 => x"0c883d0d",
          2641 => x"04f63d0d",
          2642 => x"7c59ff79",
          2643 => x"08707254",
          2644 => x"59565a74",
          2645 => x"802e81d0",
          2646 => x"38767081",
          2647 => x"05583370",
          2648 => x"ba327030",
          2649 => x"72a02671",
          2650 => x"9f2a0651",
          2651 => x"51525370",
          2652 => x"e83872ba",
          2653 => x"2e098106",
          2654 => x"81a93874",
          2655 => x"33d01152",
          2656 => x"52708926",
          2657 => x"92388215",
          2658 => x"7281ff06",
          2659 => x"d0115159",
          2660 => x"5170772e",
          2661 => x"80ff3880",
          2662 => x"0b81fbe8",
          2663 => x"5c587710",
          2664 => x"101b7008",
          2665 => x"7a085757",
          2666 => x"51757081",
          2667 => x"05573375",
          2668 => x"70810557",
          2669 => x"33ff9f12",
          2670 => x"53545470",
          2671 => x"99268938",
          2672 => x"e0147081",
          2673 => x"ff065551",
          2674 => x"ff9f1351",
          2675 => x"70992689",
          2676 => x"38e01370",
          2677 => x"81ff0654",
          2678 => x"51733074",
          2679 => x"74327030",
          2680 => x"70720780",
          2681 => x"25739f2a",
          2682 => x"06535553",
          2683 => x"5170ffb9",
          2684 => x"38733075",
          2685 => x"78327030",
          2686 => x"7072079f",
          2687 => x"2a739f2a",
          2688 => x"07535553",
          2689 => x"5170802e",
          2690 => x"8c388118",
          2691 => x"58837825",
          2692 => x"ff8c388b",
          2693 => x"39778324",
          2694 => x"86387777",
          2695 => x"7a0c5a79",
          2696 => x"51863982",
          2697 => x"93f83351",
          2698 => x"708293c8",
          2699 => x"0c8c3d0d",
          2700 => x"04fb3d0d",
          2701 => x"7756800b",
          2702 => x"831734ff",
          2703 => x"0bb0170c",
          2704 => x"78527551",
          2705 => x"e1813f84",
          2706 => x"558293c8",
          2707 => x"08818438",
          2708 => x"84b21651",
          2709 => x"ddc33f82",
          2710 => x"93c80883",
          2711 => x"ffff0654",
          2712 => x"83557382",
          2713 => x"d4d52e09",
          2714 => x"810680e7",
          2715 => x"38800bb4",
          2716 => x"17335555",
          2717 => x"7381e92e",
          2718 => x"09810683",
          2719 => x"38815573",
          2720 => x"81eb3270",
          2721 => x"30708025",
          2722 => x"77075151",
          2723 => x"54738e38",
          2724 => x"b4163354",
          2725 => x"7381e82e",
          2726 => x"098106b5",
          2727 => x"38835381",
          2728 => x"fb805280",
          2729 => x"ea1651de",
          2730 => x"bd3f8293",
          2731 => x"c8085582",
          2732 => x"93c80880",
          2733 => x"2e9d3885",
          2734 => x"5381fb84",
          2735 => x"52818616",
          2736 => x"51dea33f",
          2737 => x"8293c808",
          2738 => x"558293c8",
          2739 => x"08802e83",
          2740 => x"38825574",
          2741 => x"8293c80c",
          2742 => x"873d0d04",
          2743 => x"f33d0d60",
          2744 => x"02840580",
          2745 => x"c7053358",
          2746 => x"5480740c",
          2747 => x"7f51fcd5",
          2748 => x"3f8293c8",
          2749 => x"08588b56",
          2750 => x"800b8293",
          2751 => x"c8082487",
          2752 => x"9e388293",
          2753 => x"c8081010",
          2754 => x"8293e405",
          2755 => x"70085653",
          2756 => x"8c567480",
          2757 => x"2e878838",
          2758 => x"74740c76",
          2759 => x"81fe0675",
          2760 => x"33545772",
          2761 => x"802eaf38",
          2762 => x"81153351",
          2763 => x"d6a63f82",
          2764 => x"93c80881",
          2765 => x"ff067081",
          2766 => x"06545472",
          2767 => x"99387680",
          2768 => x"2e8f3873",
          2769 => x"822a7081",
          2770 => x"0651538a",
          2771 => x"567286cf",
          2772 => x"38805686",
          2773 => x"ca398075",
          2774 => x"34778116",
          2775 => x"34815281",
          2776 => x"153351d6",
          2777 => x"8d3f8293",
          2778 => x"c80881ff",
          2779 => x"06708106",
          2780 => x"54548356",
          2781 => x"7286a838",
          2782 => x"76802e8f",
          2783 => x"3873822a",
          2784 => x"70810651",
          2785 => x"538a5672",
          2786 => x"86953880",
          2787 => x"70537552",
          2788 => x"5afd9e3f",
          2789 => x"8293c808",
          2790 => x"81ff0657",
          2791 => x"76822e09",
          2792 => x"810680e4",
          2793 => x"38795473",
          2794 => x"90291590",
          2795 => x"3d751010",
          2796 => x"05f00583",
          2797 => x"f6123355",
          2798 => x"59568057",
          2799 => x"72772e8d",
          2800 => x"3883fa16",
          2801 => x"51daeb3f",
          2802 => x"8293c808",
          2803 => x"5776780c",
          2804 => x"81145483",
          2805 => x"7427d038",
          2806 => x"80548f3d",
          2807 => x"74101005",
          2808 => x"f011085b",
          2809 => x"53835779",
          2810 => x"802e9038",
          2811 => x"79527451",
          2812 => x"fcbf3f82",
          2813 => x"93c80881",
          2814 => x"ff065781",
          2815 => x"77278938",
          2816 => x"81145483",
          2817 => x"7427d338",
          2818 => x"81567684",
          2819 => x"2e859038",
          2820 => x"8d567681",
          2821 => x"26858838",
          2822 => x"bf1551d9",
          2823 => x"fc3f8293",
          2824 => x"c80883ff",
          2825 => x"ff06538d",
          2826 => x"56728480",
          2827 => x"2e098106",
          2828 => x"84ed3880",
          2829 => x"ca1551d9",
          2830 => x"e03f8293",
          2831 => x"c80883ff",
          2832 => x"ff065473",
          2833 => x"8d3880d8",
          2834 => x"1551d9e6",
          2835 => x"3f8293c8",
          2836 => x"0854739c",
          2837 => x"160c80c4",
          2838 => x"15338216",
          2839 => x"3480c415",
          2840 => x"33ff0553",
          2841 => x"8d567281",
          2842 => x"2684b438",
          2843 => x"82153374",
          2844 => x"712980c1",
          2845 => x"17335255",
          2846 => x"53728a16",
          2847 => x"237283ff",
          2848 => x"ff065372",
          2849 => x"802e8b38",
          2850 => x"ff137306",
          2851 => x"5372802e",
          2852 => x"86388d56",
          2853 => x"84893980",
          2854 => x"c51551d8",
          2855 => x"fc3f8293",
          2856 => x"c8088816",
          2857 => x"238293c8",
          2858 => x"0883ffff",
          2859 => x"068f0653",
          2860 => x"8d567283",
          2861 => x"ea3880c7",
          2862 => x"1551d8dd",
          2863 => x"3f8293c8",
          2864 => x"0883ffff",
          2865 => x"0653728d",
          2866 => x"3880d415",
          2867 => x"51d8e33f",
          2868 => x"8293c808",
          2869 => x"5380c215",
          2870 => x"51d8be3f",
          2871 => x"8293c808",
          2872 => x"83ffff06",
          2873 => x"598d5678",
          2874 => x"802e83b3",
          2875 => x"38881522",
          2876 => x"741a7184",
          2877 => x"2a055956",
          2878 => x"8d567773",
          2879 => x"2683a038",
          2880 => x"8a152252",
          2881 => x"72783151",
          2882 => x"ffb0ab3f",
          2883 => x"8293c808",
          2884 => x"538d5682",
          2885 => x"93c80880",
          2886 => x"2e838438",
          2887 => x"80578293",
          2888 => x"c80880ff",
          2889 => x"fffff526",
          2890 => x"83388357",
          2891 => x"7283fff5",
          2892 => x"26833882",
          2893 => x"57729ff5",
          2894 => x"26833881",
          2895 => x"578d5676",
          2896 => x"802e82db",
          2897 => x"38821398",
          2898 => x"160c79a0",
          2899 => x"160c7919",
          2900 => x"a4160c77",
          2901 => x"1aac160c",
          2902 => x"76832e09",
          2903 => x"8106b738",
          2904 => x"80de1551",
          2905 => x"d7b33f82",
          2906 => x"93c80883",
          2907 => x"ffff0653",
          2908 => x"8d567282",
          2909 => x"aa388815",
          2910 => x"22538d56",
          2911 => x"7282a038",
          2912 => x"80e01551",
          2913 => x"d7ac3f82",
          2914 => x"93c808a8",
          2915 => x"160c9815",
          2916 => x"08822b53",
          2917 => x"b6398815",
          2918 => x"22538d56",
          2919 => x"72802e81",
          2920 => x"fe38a415",
          2921 => x"0814a816",
          2922 => x"0c76822e",
          2923 => x"09810688",
          2924 => x"38981508",
          2925 => x"10539439",
          2926 => x"98150810",
          2927 => x"98160805",
          2928 => x"70812a98",
          2929 => x"17088106",
          2930 => x"05515383",
          2931 => x"ff13892a",
          2932 => x"538d5672",
          2933 => x"9c160826",
          2934 => x"81c538ff",
          2935 => x"0b90160c",
          2936 => x"ff0b8c16",
          2937 => x"0cff800b",
          2938 => x"84163476",
          2939 => x"832e0981",
          2940 => x"06819238",
          2941 => x"80e41551",
          2942 => x"d69f3f82",
          2943 => x"93c80883",
          2944 => x"ffff0653",
          2945 => x"72812e09",
          2946 => x"810680f9",
          2947 => x"38811a52",
          2948 => x"7451d9b3",
          2949 => x"3f8293c8",
          2950 => x"0880ea38",
          2951 => x"8293c808",
          2952 => x"84163484",
          2953 => x"b21551d5",
          2954 => x"f03f8293",
          2955 => x"c80883ff",
          2956 => x"ff065372",
          2957 => x"82d4d52e",
          2958 => x"09810680",
          2959 => x"c838b415",
          2960 => x"51d5ef3f",
          2961 => x"8293c808",
          2962 => x"848b85a4",
          2963 => x"d22e0981",
          2964 => x"06b33884",
          2965 => x"981551d5",
          2966 => x"d93f8293",
          2967 => x"c808868a",
          2968 => x"85e4f22e",
          2969 => x"0981069d",
          2970 => x"38849c15",
          2971 => x"51d5c33f",
          2972 => x"8293c808",
          2973 => x"90160c84",
          2974 => x"a01551d5",
          2975 => x"b53f8293",
          2976 => x"c8088c16",
          2977 => x"0c767534",
          2978 => x"8293f422",
          2979 => x"81055372",
          2980 => x"8293f423",
          2981 => x"72861623",
          2982 => x"800b9416",
          2983 => x"0c805675",
          2984 => x"8293c80c",
          2985 => x"8f3d0d04",
          2986 => x"fb3d0d77",
          2987 => x"54895573",
          2988 => x"802eb538",
          2989 => x"7308802e",
          2990 => x"af387308",
          2991 => x"70335353",
          2992 => x"71802ea4",
          2993 => x"38841422",
          2994 => x"86142257",
          2995 => x"5271762e",
          2996 => x"09810694",
          2997 => x"38811333",
          2998 => x"51cef93f",
          2999 => x"8293c808",
          3000 => x"81065271",
          3001 => x"83387155",
          3002 => x"80537473",
          3003 => x"2e098106",
          3004 => x"84387308",
          3005 => x"53787371",
          3006 => x"0c527482",
          3007 => x"93c80c87",
          3008 => x"3d0d04fa",
          3009 => x"3d0d02ab",
          3010 => x"05337a58",
          3011 => x"893dfc05",
          3012 => x"5256f4b1",
          3013 => x"3f8293c8",
          3014 => x"08558b54",
          3015 => x"800b8293",
          3016 => x"c8082480",
          3017 => x"c4388293",
          3018 => x"c8081010",
          3019 => x"8293e405",
          3020 => x"70085154",
          3021 => x"73802e84",
          3022 => x"38807434",
          3023 => x"78802e86",
          3024 => x"38785480",
          3025 => x"74347410",
          3026 => x"108293e4",
          3027 => x"0579710c",
          3028 => x"54755475",
          3029 => x"802e9238",
          3030 => x"8053893d",
          3031 => x"70538405",
          3032 => x"51f6f93f",
          3033 => x"8293c808",
          3034 => x"54738293",
          3035 => x"c80c883d",
          3036 => x"0d04eb3d",
          3037 => x"0d670284",
          3038 => x"0580e705",
          3039 => x"33585889",
          3040 => x"5577802e",
          3041 => x"84e93876",
          3042 => x"bf067054",
          3043 => x"983dd005",
          3044 => x"53993d84",
          3045 => x"055257f6",
          3046 => x"c33f8293",
          3047 => x"c8085682",
          3048 => x"93c80884",
          3049 => x"c5387a5c",
          3050 => x"6852973d",
          3051 => x"d40551f0",
          3052 => x"db3f8293",
          3053 => x"c8085682",
          3054 => x"93c80892",
          3055 => x"380280d7",
          3056 => x"05337098",
          3057 => x"2b565974",
          3058 => x"80258338",
          3059 => x"8656769c",
          3060 => x"06557480",
          3061 => x"2e81c338",
          3062 => x"75802e9c",
          3063 => x"3875842e",
          3064 => x"0981068e",
          3065 => x"38973dd4",
          3066 => x"0551ea9e",
          3067 => x"3f8293c8",
          3068 => x"08567688",
          3069 => x"0757a039",
          3070 => x"02b20533",
          3071 => x"91065574",
          3072 => x"802e8538",
          3073 => x"87569039",
          3074 => x"76822a70",
          3075 => x"81065155",
          3076 => x"74802e83",
          3077 => x"38885675",
          3078 => x"83d03876",
          3079 => x"832a7081",
          3080 => x"06515574",
          3081 => x"802e81a7",
          3082 => x"3862527a",
          3083 => x"51e6b63f",
          3084 => x"8293c808",
          3085 => x"598288b2",
          3086 => x"0a52628e",
          3087 => x"0551d2b9",
          3088 => x"3f6255a0",
          3089 => x"0b8b1634",
          3090 => x"75536252",
          3091 => x"7a51e6ce",
          3092 => x"3f755262",
          3093 => x"9c0551d2",
          3094 => x"a03f7a55",
          3095 => x"810b8316",
          3096 => x"3478802e",
          3097 => x"80e9387a",
          3098 => x"b0110877",
          3099 => x"557a5499",
          3100 => x"3dd40553",
          3101 => x"5155dbb3",
          3102 => x"3f8293c8",
          3103 => x"08568293",
          3104 => x"c80882e6",
          3105 => x"3874527a",
          3106 => x"51d4bc3f",
          3107 => x"8293c808",
          3108 => x"7bff1b8c",
          3109 => x"120c5656",
          3110 => x"b6397582",
          3111 => x"cd3802b2",
          3112 => x"05337084",
          3113 => x"2a708106",
          3114 => x"51565974",
          3115 => x"802e8538",
          3116 => x"84569c39",
          3117 => x"76812a70",
          3118 => x"81065155",
          3119 => x"74802e8f",
          3120 => x"3802b205",
          3121 => x"33810655",
          3122 => x"74802e83",
          3123 => x"38875675",
          3124 => x"82983876",
          3125 => x"832a7081",
          3126 => x"06515574",
          3127 => x"802e8638",
          3128 => x"7680c007",
          3129 => x"577ab011",
          3130 => x"08a01a0c",
          3131 => x"63a41a0c",
          3132 => x"557581f6",
          3133 => x"38625274",
          3134 => x"51e4ea3f",
          3135 => x"8293c808",
          3136 => x"88190c62",
          3137 => x"9c0551d0",
          3138 => x"a93f8293",
          3139 => x"c8088c19",
          3140 => x"0c74780c",
          3141 => x"86152284",
          3142 => x"19237690",
          3143 => x"19347591",
          3144 => x"1934759c",
          3145 => x"190c7594",
          3146 => x"190c8480",
          3147 => x"537552a8",
          3148 => x"1851d198",
          3149 => x"3f76852a",
          3150 => x"70810651",
          3151 => x"5574802e",
          3152 => x"81a3388c",
          3153 => x"1808802e",
          3154 => x"819b388c",
          3155 => x"18089419",
          3156 => x"0c7a8a11",
          3157 => x"2270892b",
          3158 => x"881b088c",
          3159 => x"1c085d5a",
          3160 => x"5c5155a5",
          3161 => x"39765277",
          3162 => x"51d4fc3f",
          3163 => x"8293c808",
          3164 => x"578293c8",
          3165 => x"08812683",
          3166 => x"38825676",
          3167 => x"ff2e0981",
          3168 => x"06833881",
          3169 => x"56787a31",
          3170 => x"59753070",
          3171 => x"77078025",
          3172 => x"707b7d26",
          3173 => x"06515155",
          3174 => x"74cb3876",
          3175 => x"98190c75",
          3176 => x"80c83878",
          3177 => x"83ff0655",
          3178 => x"74802eb9",
          3179 => x"3876527a",
          3180 => x"51d48a3f",
          3181 => x"8293c808",
          3182 => x"85388256",
          3183 => x"a8397889",
          3184 => x"2a8293c8",
          3185 => x"0805709c",
          3186 => x"1a0c5581",
          3187 => x"547453a8",
          3188 => x"18527a81",
          3189 => x"11335255",
          3190 => x"caa43f82",
          3191 => x"93c80880",
          3192 => x"2e833881",
          3193 => x"5675802e",
          3194 => x"84388078",
          3195 => x"0c755574",
          3196 => x"8293c80c",
          3197 => x"973d0d04",
          3198 => x"f33d0d7f",
          3199 => x"6264635f",
          3200 => x"5f5a5780",
          3201 => x"7d0c8f3d",
          3202 => x"fc055276",
          3203 => x"51f9993f",
          3204 => x"8293c808",
          3205 => x"558293c8",
          3206 => x"088a3891",
          3207 => x"17335574",
          3208 => x"802e8638",
          3209 => x"745683ae",
          3210 => x"39901733",
          3211 => x"81065587",
          3212 => x"5674802e",
          3213 => x"83a038bd",
          3214 => x"39820b91",
          3215 => x"18348256",
          3216 => x"83943981",
          3217 => x"0b911834",
          3218 => x"8156838a",
          3219 => x"39820b91",
          3220 => x"18348256",
          3221 => x"83803981",
          3222 => x"0b911834",
          3223 => x"815682f6",
          3224 => x"39810b91",
          3225 => x"18348156",
          3226 => x"82ec3981",
          3227 => x"0b911834",
          3228 => x"815682e2",
          3229 => x"398c1708",
          3230 => x"94180831",
          3231 => x"55747927",
          3232 => x"83387459",
          3233 => x"78802e82",
          3234 => x"cb389417",
          3235 => x"087083ff",
          3236 => x"06565674",
          3237 => x"8283387d",
          3238 => x"8a1122ff",
          3239 => x"0577892a",
          3240 => x"065c557a",
          3241 => x"a8387587",
          3242 => x"38881708",
          3243 => x"558f3998",
          3244 => x"17085276",
          3245 => x"51d2b03f",
          3246 => x"8293c808",
          3247 => x"55817527",
          3248 => x"fef73874",
          3249 => x"ff2efefb",
          3250 => x"38749818",
          3251 => x"0c981708",
          3252 => x"527d51d1",
          3253 => x"e83f8293",
          3254 => x"c808802e",
          3255 => x"feef3882",
          3256 => x"93c8081b",
          3257 => x"79892a5b",
          3258 => x"5879802e",
          3259 => x"80d73879",
          3260 => x"1b7e8a11",
          3261 => x"22515656",
          3262 => x"74762785",
          3263 => x"38747b31",
          3264 => x"5a795477",
          3265 => x"537b527d",
          3266 => x"81113352",
          3267 => x"55c7ef3f",
          3268 => x"8293c808",
          3269 => x"fec13890",
          3270 => x"17337098",
          3271 => x"2b565674",
          3272 => x"80259b38",
          3273 => x"9c170878",
          3274 => x"3155747a",
          3275 => x"27903884",
          3276 => x"8053a817",
          3277 => x"52748480",
          3278 => x"291c51cc",
          3279 => x"eb3f7989",
          3280 => x"2b5680f9",
          3281 => x"399c1708",
          3282 => x"782e80c9",
          3283 => x"38901733",
          3284 => x"70982b56",
          3285 => x"56748025",
          3286 => x"a5388154",
          3287 => x"9c170853",
          3288 => x"a817527d",
          3289 => x"81113352",
          3290 => x"55c8ec3f",
          3291 => x"8293c808",
          3292 => x"fdef3890",
          3293 => x"173380ff",
          3294 => x"06557490",
          3295 => x"18348154",
          3296 => x"7753a817",
          3297 => x"527d8111",
          3298 => x"335255c6",
          3299 => x"f13f8293",
          3300 => x"c808fdd7",
          3301 => x"38779c18",
          3302 => x"0c941708",
          3303 => x"83ff0684",
          3304 => x"80713157",
          3305 => x"55787627",
          3306 => x"83387856",
          3307 => x"75539417",
          3308 => x"0883ff06",
          3309 => x"17a80552",
          3310 => x"7b51cbec",
          3311 => x"3f787631",
          3312 => x"7d08177e",
          3313 => x"0c761d94",
          3314 => x"19081894",
          3315 => x"1a0c5d59",
          3316 => x"78fdb738",
          3317 => x"80567582",
          3318 => x"93c80c8f",
          3319 => x"3d0d04f3",
          3320 => x"3d0d7f62",
          3321 => x"64635f5f",
          3322 => x"5a57807d",
          3323 => x"0c8f3dfc",
          3324 => x"05527651",
          3325 => x"f5b23f82",
          3326 => x"93c80855",
          3327 => x"8293c808",
          3328 => x"8a389117",
          3329 => x"33557480",
          3330 => x"2e863874",
          3331 => x"56848239",
          3332 => x"90173370",
          3333 => x"812a7081",
          3334 => x"06515656",
          3335 => x"87567480",
          3336 => x"2e83ee38",
          3337 => x"bd39820b",
          3338 => x"91183482",
          3339 => x"5683e239",
          3340 => x"810b9118",
          3341 => x"34815683",
          3342 => x"d839810b",
          3343 => x"91183481",
          3344 => x"5683ce39",
          3345 => x"820b9118",
          3346 => x"34825683",
          3347 => x"c439810b",
          3348 => x"91183481",
          3349 => x"5683ba39",
          3350 => x"810b9118",
          3351 => x"34815683",
          3352 => x"b0399417",
          3353 => x"08195574",
          3354 => x"94180827",
          3355 => x"86389417",
          3356 => x"08095978",
          3357 => x"802e838c",
          3358 => x"38941708",
          3359 => x"7083ff06",
          3360 => x"56567482",
          3361 => x"a8387d8a",
          3362 => x"1122ff05",
          3363 => x"77892a06",
          3364 => x"5c557a80",
          3365 => x"c6387596",
          3366 => x"38881708",
          3367 => x"5574a338",
          3368 => x"7a527651",
          3369 => x"d4b83f82",
          3370 => x"93c80855",
          3371 => x"8f399817",
          3372 => x"08527651",
          3373 => x"d4a83f82",
          3374 => x"93c80855",
          3375 => x"74802e82",
          3376 => x"c3387481",
          3377 => x"2efedf38",
          3378 => x"74ff2efe",
          3379 => x"e3387498",
          3380 => x"180c8817",
          3381 => x"08853874",
          3382 => x"88180c90",
          3383 => x"17337098",
          3384 => x"2b565874",
          3385 => x"8025a538",
          3386 => x"81549c17",
          3387 => x"0853a817",
          3388 => x"527d8111",
          3389 => x"335255c5",
          3390 => x"de3f8293",
          3391 => x"c808feba",
          3392 => x"38901733",
          3393 => x"80ff0655",
          3394 => x"74901834",
          3395 => x"98170852",
          3396 => x"7d51cda9",
          3397 => x"3f8293c8",
          3398 => x"08802efe",
          3399 => x"a7388293",
          3400 => x"c8081b79",
          3401 => x"892a5b58",
          3402 => x"79802e80",
          3403 => x"d538791b",
          3404 => x"7e8a1122",
          3405 => x"51565674",
          3406 => x"76278538",
          3407 => x"747b315a",
          3408 => x"79547753",
          3409 => x"7b527d81",
          3410 => x"11335255",
          3411 => x"c5893f82",
          3412 => x"93c808fd",
          3413 => x"f9389c17",
          3414 => x"08783155",
          3415 => x"747a279b",
          3416 => x"38848053",
          3417 => x"74848029",
          3418 => x"1c52a817",
          3419 => x"51c8b93f",
          3420 => x"90173380",
          3421 => x"ff065574",
          3422 => x"90183479",
          3423 => x"892b5680",
          3424 => x"db399c17",
          3425 => x"08782ea1",
          3426 => x"38941708",
          3427 => x"8c180827",
          3428 => x"98388154",
          3429 => x"7753a817",
          3430 => x"527d8111",
          3431 => x"335255c2",
          3432 => x"dd3f8293",
          3433 => x"c808fdb0",
          3434 => x"38779c18",
          3435 => x"0c941708",
          3436 => x"83ff0684",
          3437 => x"80713157",
          3438 => x"55787627",
          3439 => x"83387856",
          3440 => x"75537b52",
          3441 => x"94170883",
          3442 => x"ff0617a8",
          3443 => x"0551c7d8",
          3444 => x"3f901733",
          3445 => x"ff800755",
          3446 => x"74901834",
          3447 => x"7876317d",
          3448 => x"08177e0c",
          3449 => x"761d9419",
          3450 => x"08187094",
          3451 => x"1b0c8c1a",
          3452 => x"0858585d",
          3453 => x"59747627",
          3454 => x"83387555",
          3455 => x"748c180c",
          3456 => x"78fcf638",
          3457 => x"90173380",
          3458 => x"c0075574",
          3459 => x"90183480",
          3460 => x"56758293",
          3461 => x"c80c8f3d",
          3462 => x"0d04f73d",
          3463 => x"0d7b8c3d",
          3464 => x"fc055370",
          3465 => x"5258f180",
          3466 => x"3f8293c8",
          3467 => x"08578293",
          3468 => x"c80881aa",
          3469 => x"38901833",
          3470 => x"70862a70",
          3471 => x"81065156",
          3472 => x"5674802e",
          3473 => x"81983875",
          3474 => x"982b5574",
          3475 => x"8025a738",
          3476 => x"81549c18",
          3477 => x"0853a818",
          3478 => x"52798111",
          3479 => x"335255c2",
          3480 => x"f63f8155",
          3481 => x"8293c808",
          3482 => x"80f63890",
          3483 => x"183380ff",
          3484 => x"06557490",
          3485 => x"1934a018",
          3486 => x"08527951",
          3487 => x"c8c93f82",
          3488 => x"93c80857",
          3489 => x"8293c808",
          3490 => x"80d438a4",
          3491 => x"18088b11",
          3492 => x"33a00756",
          3493 => x"56748b17",
          3494 => x"34881808",
          3495 => x"53755277",
          3496 => x"0851d9fa",
          3497 => x"3f8c1808",
          3498 => x"529c1651",
          3499 => x"c5cb3f82",
          3500 => x"88b20a52",
          3501 => x"961651c5",
          3502 => x"c03f7652",
          3503 => x"921651c5",
          3504 => x"9a3f7955",
          3505 => x"810b8316",
          3506 => x"347951c8",
          3507 => x"c13f8293",
          3508 => x"c8089019",
          3509 => x"3381bf06",
          3510 => x"56577490",
          3511 => x"19347655",
          3512 => x"748293c8",
          3513 => x"0c8b3d0d",
          3514 => x"04fc3d0d",
          3515 => x"76705254",
          3516 => x"fea83f82",
          3517 => x"93c80853",
          3518 => x"8293c808",
          3519 => x"9c38863d",
          3520 => x"fc055273",
          3521 => x"51efa13f",
          3522 => x"8293c808",
          3523 => x"538293c8",
          3524 => x"08873882",
          3525 => x"93c80874",
          3526 => x"0c728293",
          3527 => x"c80c863d",
          3528 => x"0d04fe3d",
          3529 => x"0d853d51",
          3530 => x"e49b3f8b",
          3531 => x"53800b82",
          3532 => x"93c80824",
          3533 => x"8b388293",
          3534 => x"c8088293",
          3535 => x"f8348053",
          3536 => x"728293c8",
          3537 => x"0c843d0d",
          3538 => x"04ef3d0d",
          3539 => x"8053933d",
          3540 => x"d0055294",
          3541 => x"3d51e784",
          3542 => x"3f8293c8",
          3543 => x"08558293",
          3544 => x"c80880df",
          3545 => x"38765863",
          3546 => x"52933dd4",
          3547 => x"0551e19c",
          3548 => x"3f8293c8",
          3549 => x"08558293",
          3550 => x"c808be38",
          3551 => x"0280c705",
          3552 => x"3370982b",
          3553 => x"55567380",
          3554 => x"25893876",
          3555 => x"7a94120c",
          3556 => x"54a73902",
          3557 => x"a2053370",
          3558 => x"842a7081",
          3559 => x"06515556",
          3560 => x"73802e93",
          3561 => x"38767f53",
          3562 => x"705254d7",
          3563 => x"b83f8293",
          3564 => x"c8089415",
          3565 => x"0c833985",
          3566 => x"5574842e",
          3567 => x"09810683",
          3568 => x"38855574",
          3569 => x"8293c80c",
          3570 => x"933d0d04",
          3571 => x"e13d0da3",
          3572 => x"3d08a33d",
          3573 => x"085b5c80",
          3574 => x"7a348053",
          3575 => x"a13dffb8",
          3576 => x"0552a23d",
          3577 => x"51e5f53f",
          3578 => x"8293c808",
          3579 => x"578293c8",
          3580 => x"08839338",
          3581 => x"7e467b7f",
          3582 => x"9411084a",
          3583 => x"55685659",
          3584 => x"74802e81",
          3585 => x"f938963d",
          3586 => x"70943d40",
          3587 => x"5e5ba052",
          3588 => x"7a51d1e4",
          3589 => x"3f8293c8",
          3590 => x"08578293",
          3591 => x"c80881de",
          3592 => x"386b527e",
          3593 => x"51c5a03f",
          3594 => x"8293c808",
          3595 => x"578293c8",
          3596 => x"0881cb38",
          3597 => x"6c527e51",
          3598 => x"d6ab3f82",
          3599 => x"93c80848",
          3600 => x"76527a51",
          3601 => x"d1b23f82",
          3602 => x"93c80857",
          3603 => x"8293c808",
          3604 => x"81ac387c",
          3605 => x"54805273",
          3606 => x"51d6f13f",
          3607 => x"8293c808",
          3608 => x"578293c8",
          3609 => x"08a4386c",
          3610 => x"527e51d5",
          3611 => x"f83f8293",
          3612 => x"c808752e",
          3613 => x"95387652",
          3614 => x"7351d2d1",
          3615 => x"3f8293c8",
          3616 => x"08578293",
          3617 => x"c808802e",
          3618 => x"cc387684",
          3619 => x"2e098106",
          3620 => x"83388257",
          3621 => x"7681ef38",
          3622 => x"a13dffbc",
          3623 => x"1153d405",
          3624 => x"51d9ee3f",
          3625 => x"76933d70",
          3626 => x"79128111",
          3627 => x"33515257",
          3628 => x"55567380",
          3629 => x"2e8e3881",
          3630 => x"16701681",
          3631 => x"11335155",
          3632 => x"5673f438",
          3633 => x"81165478",
          3634 => x"74278538",
          3635 => x"9157af39",
          3636 => x"75802e99",
          3637 => x"387d58ff",
          3638 => x"19a33d08",
          3639 => x"11ff1870",
          3640 => x"1b575856",
          3641 => x"59811433",
          3642 => x"753475eb",
          3643 => x"38ff19a3",
          3644 => x"3d081155",
          3645 => x"59af7434",
          3646 => x"675574fe",
          3647 => x"91387681",
          3648 => x"8538787c",
          3649 => x"2e098106",
          3650 => x"8c38ff19",
          3651 => x"a33d0811",
          3652 => x"5559af74",
          3653 => x"34807082",
          3654 => x"93f83370",
          3655 => x"101081fb",
          3656 => x"e8057008",
          3657 => x"70335252",
          3658 => x"57575758",
          3659 => x"73782e8d",
          3660 => x"38811670",
          3661 => x"16703351",
          3662 => x"555673f5",
          3663 => x"38821654",
          3664 => x"737926a5",
          3665 => x"38805877",
          3666 => x"76279438",
          3667 => x"77155473",
          3668 => x"337a7081",
          3669 => x"055c3481",
          3670 => x"18587578",
          3671 => x"26ee38ba",
          3672 => x"7a708105",
          3673 => x"5c348118",
          3674 => x"58778338",
          3675 => x"91577696",
          3676 => x"38a23d08",
          3677 => x"19811a5a",
          3678 => x"5473337a",
          3679 => x"7081055c",
          3680 => x"347b7926",
          3681 => x"ec38807a",
          3682 => x"34768293",
          3683 => x"c80ca13d",
          3684 => x"0d04f43d",
          3685 => x"0d7e6090",
          3686 => x"3dfc0554",
          3687 => x"71535957",
          3688 => x"ea863f82",
          3689 => x"93c8085a",
          3690 => x"8293c808",
          3691 => x"8a389117",
          3692 => x"335a7980",
          3693 => x"2e863879",
          3694 => x"5583f939",
          3695 => x"8c170878",
          3696 => x"27943890",
          3697 => x"17337081",
          3698 => x"2a708106",
          3699 => x"51565674",
          3700 => x"85388c17",
          3701 => x"08589417",
          3702 => x"08568070",
          3703 => x"94190c5b",
          3704 => x"777b2e82",
          3705 => x"b3387c8a",
          3706 => x"11227089",
          3707 => x"2b5b5155",
          3708 => x"757b2eb6",
          3709 => x"387852ff",
          3710 => x"1851ff96",
          3711 => x"b93f8293",
          3712 => x"c808ff17",
          3713 => x"7a547053",
          3714 => x"5755ff96",
          3715 => x"a93f8293",
          3716 => x"c8087526",
          3717 => x"95387830",
          3718 => x"76069418",
          3719 => x"0c779418",
          3720 => x"08319818",
          3721 => x"08575880",
          3722 => x"c9398817",
          3723 => x"085675be",
          3724 => x"38755276",
          3725 => x"51c9a73f",
          3726 => x"8293c808",
          3727 => x"568293c8",
          3728 => x"08812e09",
          3729 => x"81068b38",
          3730 => x"820b9118",
          3731 => x"34825582",
          3732 => x"e3398293",
          3733 => x"c808ff2e",
          3734 => x"0981068b",
          3735 => x"38810b91",
          3736 => x"18348155",
          3737 => x"82ce3982",
          3738 => x"93c80888",
          3739 => x"180c7598",
          3740 => x"180c7580",
          3741 => x"2e81a138",
          3742 => x"78782780",
          3743 => x"ea387779",
          3744 => x"31941808",
          3745 => x"1a94190c",
          3746 => x"90183370",
          3747 => x"812a7081",
          3748 => x"0651575d",
          3749 => x"5874802e",
          3750 => x"9a387552",
          3751 => x"7651c8be",
          3752 => x"3f8293c8",
          3753 => x"08568293",
          3754 => x"c8089438",
          3755 => x"8293c808",
          3756 => x"58b53975",
          3757 => x"527651c2",
          3758 => x"ae3f8293",
          3759 => x"c8085675",
          3760 => x"ff2e81e1",
          3761 => x"38817627",
          3762 => x"8a387c55",
          3763 => x"98150876",
          3764 => x"268b3882",
          3765 => x"0b911834",
          3766 => x"825581d8",
          3767 => x"39759818",
          3768 => x"0c777926",
          3769 => x"ff983894",
          3770 => x"17081894",
          3771 => x"180c7783",
          3772 => x"ff065574",
          3773 => x"802ea138",
          3774 => x"75527c51",
          3775 => x"c1bf3f82",
          3776 => x"93c8088b",
          3777 => x"38820b91",
          3778 => x"18348255",
          3779 => x"81a63977",
          3780 => x"892a8293",
          3781 => x"c808055b",
          3782 => x"8c170894",
          3783 => x"18082792",
          3784 => x"38941708",
          3785 => x"8c180c90",
          3786 => x"173380c0",
          3787 => x"07557490",
          3788 => x"18349417",
          3789 => x"0883ff06",
          3790 => x"5574802e",
          3791 => x"80f4389c",
          3792 => x"17087b2e",
          3793 => x"80ec3890",
          3794 => x"17337098",
          3795 => x"2b565c74",
          3796 => x"8025b038",
          3797 => x"81549c17",
          3798 => x"0853a817",
          3799 => x"527c8111",
          3800 => x"335255ff",
          3801 => x"b8f13f82",
          3802 => x"93c80880",
          3803 => x"2e8a3881",
          3804 => x"0b911834",
          3805 => x"8155bd39",
          3806 => x"90173380",
          3807 => x"ff065574",
          3808 => x"90183481",
          3809 => x"547a53a8",
          3810 => x"17527c81",
          3811 => x"11335255",
          3812 => x"ffb6eb3f",
          3813 => x"8293c808",
          3814 => x"802e9338",
          3815 => x"810b9118",
          3816 => x"34815590",
          3817 => x"39810b91",
          3818 => x"18348155",
          3819 => x"87397a9c",
          3820 => x"180c7955",
          3821 => x"748293c8",
          3822 => x"0c8e3d0d",
          3823 => x"04f93d0d",
          3824 => x"79568954",
          3825 => x"75802e81",
          3826 => x"8f388053",
          3827 => x"893dfc05",
          3828 => x"528a3d84",
          3829 => x"0551de84",
          3830 => x"3f8293c8",
          3831 => x"08558293",
          3832 => x"c80880ef",
          3833 => x"3877760c",
          3834 => x"7a527551",
          3835 => x"d89e3f82",
          3836 => x"93c80855",
          3837 => x"8293c808",
          3838 => x"80ca38ab",
          3839 => x"16337098",
          3840 => x"2b555780",
          3841 => x"7424a638",
          3842 => x"86163370",
          3843 => x"842a7081",
          3844 => x"06515557",
          3845 => x"73802e93",
          3846 => x"389c1608",
          3847 => x"527751ce",
          3848 => x"c43f8293",
          3849 => x"c8088817",
          3850 => x"0c833985",
          3851 => x"55749538",
          3852 => x"77548614",
          3853 => x"22841723",
          3854 => x"74527551",
          3855 => x"c9ba3f82",
          3856 => x"93c80855",
          3857 => x"74842e09",
          3858 => x"81068338",
          3859 => x"85557480",
          3860 => x"2e843880",
          3861 => x"760c7454",
          3862 => x"738293c8",
          3863 => x"0c893d0d",
          3864 => x"04fc3d0d",
          3865 => x"76873dfc",
          3866 => x"05537052",
          3867 => x"54e4b93f",
          3868 => x"8293c808",
          3869 => x"538293c8",
          3870 => x"08873882",
          3871 => x"93c80874",
          3872 => x"0c728293",
          3873 => x"c80c863d",
          3874 => x"0d04fb3d",
          3875 => x"0d777989",
          3876 => x"3dfc0554",
          3877 => x"71535654",
          3878 => x"e48e3f82",
          3879 => x"93c80853",
          3880 => x"8293c808",
          3881 => x"80d13874",
          3882 => x"92388293",
          3883 => x"c8085273",
          3884 => x"51c8c53f",
          3885 => x"8293c808",
          3886 => x"53bd3980",
          3887 => x"527351ce",
          3888 => x"8b3f8293",
          3889 => x"c8085382",
          3890 => x"93c80884",
          3891 => x"2e098106",
          3892 => x"83388053",
          3893 => x"72a13874",
          3894 => x"527351d1",
          3895 => x"b43f7252",
          3896 => x"7351c9e9",
          3897 => x"3f8293c8",
          3898 => x"08538293",
          3899 => x"c808842e",
          3900 => x"09810683",
          3901 => x"38805372",
          3902 => x"8293c80c",
          3903 => x"873d0d04",
          3904 => x"ef3d0d64",
          3905 => x"56805388",
          3906 => x"3d705395",
          3907 => x"3d5254db",
          3908 => x"cb3f8293",
          3909 => x"c8085582",
          3910 => x"93c808b5",
          3911 => x"38635273",
          3912 => x"51d5e93f",
          3913 => x"8293c808",
          3914 => x"558293c8",
          3915 => x"08a33802",
          3916 => x"80c70533",
          3917 => x"70982b55",
          3918 => x"57738025",
          3919 => x"85388655",
          3920 => x"90397580",
          3921 => x"2e8b3875",
          3922 => x"52933dd4",
          3923 => x"0551d0c1",
          3924 => x"3f748293",
          3925 => x"c80c933d",
          3926 => x"0d04f23d",
          3927 => x"0d616355",
          3928 => x"5a805390",
          3929 => x"3dec0552",
          3930 => x"913d51da",
          3931 => x"ef3f8293",
          3932 => x"c8085982",
          3933 => x"93c80882",
          3934 => x"84387a74",
          3935 => x"0c730898",
          3936 => x"1108fe05",
          3937 => x"55559015",
          3938 => x"08742693",
          3939 => x"38901508",
          3940 => x"7a0c81e9",
          3941 => x"39815981",
          3942 => x"cf398259",
          3943 => x"81ca3980",
          3944 => x"7b703356",
          3945 => x"56577381",
          3946 => x"2e098106",
          3947 => x"80c03882",
          3948 => x"755d5675",
          3949 => x"52903df0",
          3950 => x"0551ffbc",
          3951 => x"aa3f8293",
          3952 => x"c808ff2e",
          3953 => x"d0388293",
          3954 => x"c808812e",
          3955 => x"cd388293",
          3956 => x"c8083070",
          3957 => x"8293c808",
          3958 => x"07802578",
          3959 => x"0581187d",
          3960 => x"53585854",
          3961 => x"98140876",
          3962 => x"26c93880",
          3963 => x"fb397a98",
          3964 => x"1108a412",
          3965 => x"085a5754",
          3966 => x"80557498",
          3967 => x"38775281",
          3968 => x"187b5258",
          3969 => x"ffb9c03f",
          3970 => x"8293c808",
          3971 => x"598293c8",
          3972 => x"0880d538",
          3973 => x"7a703351",
          3974 => x"5473822e",
          3975 => x"098106a0",
          3976 => x"387a15b4",
          3977 => x"0551ffb5",
          3978 => x"f03f8293",
          3979 => x"c80883ff",
          3980 => x"ff067030",
          3981 => x"70802519",
          3982 => x"82185859",
          3983 => x"51549d39",
          3984 => x"7a15b405",
          3985 => x"51ffb5ea",
          3986 => x"3f8293c8",
          3987 => x"08f00a06",
          3988 => x"70307080",
          3989 => x"25198418",
          3990 => x"58595154",
          3991 => x"7483ff06",
          3992 => x"ff175755",
          3993 => x"75ff9338",
          3994 => x"767a0c7a",
          3995 => x"7790120c",
          3996 => x"547a8411",
          3997 => x"33810755",
          3998 => x"55738416",
          3999 => x"34788293",
          4000 => x"c80c903d",
          4001 => x"0d04f83d",
          4002 => x"0d7a8b3d",
          4003 => x"fc055370",
          4004 => x"5258e094",
          4005 => x"3f8293c8",
          4006 => x"08578293",
          4007 => x"c8088a38",
          4008 => x"91183357",
          4009 => x"76802e86",
          4010 => x"38765681",
          4011 => x"dc399018",
          4012 => x"3370812a",
          4013 => x"70810651",
          4014 => x"56568756",
          4015 => x"74802e81",
          4016 => x"c8389418",
          4017 => x"088c1908",
          4018 => x"2781bc38",
          4019 => x"9418089a",
          4020 => x"38805388",
          4021 => x"18085277",
          4022 => x"51ffbecf",
          4023 => x"3f8293c8",
          4024 => x"0857800b",
          4025 => x"88190c80",
          4026 => x"ca399818",
          4027 => x"08527751",
          4028 => x"ffb9f43f",
          4029 => x"8293c808",
          4030 => x"8293c808",
          4031 => x"ff327030",
          4032 => x"70720780",
          4033 => x"25525758",
          4034 => x"568293c8",
          4035 => x"08812e09",
          4036 => x"81068338",
          4037 => x"8257769b",
          4038 => x"38785575",
          4039 => x"98160827",
          4040 => x"92389818",
          4041 => x"08537552",
          4042 => x"7751ffbd",
          4043 => x"fe3f8293",
          4044 => x"c8085794",
          4045 => x"18088c19",
          4046 => x"0c901833",
          4047 => x"80c00755",
          4048 => x"74901934",
          4049 => x"76b93874",
          4050 => x"982b5574",
          4051 => x"8025ab38",
          4052 => x"81549c18",
          4053 => x"0853a818",
          4054 => x"52788111",
          4055 => x"335255ff",
          4056 => x"b0f53f82",
          4057 => x"93c80880",
          4058 => x"2e853881",
          4059 => x"578c3990",
          4060 => x"183380ff",
          4061 => x"06557490",
          4062 => x"19347680",
          4063 => x"2e893876",
          4064 => x"91193476",
          4065 => x"56833976",
          4066 => x"56758293",
          4067 => x"c80c8a3d",
          4068 => x"0d04e33d",
          4069 => x"0d81fb8c",
          4070 => x"51ff96d5",
          4071 => x"3f82539f",
          4072 => x"3dffa405",
          4073 => x"52a03d51",
          4074 => x"d6b23f82",
          4075 => x"93c80856",
          4076 => x"8293c808",
          4077 => x"82d33881",
          4078 => x"fb9051ff",
          4079 => x"96b33f77",
          4080 => x"446f529f",
          4081 => x"3dd40551",
          4082 => x"d0c23f82",
          4083 => x"93c80881",
          4084 => x"fb945256",
          4085 => x"ff969a3f",
          4086 => x"7582ae38",
          4087 => x"0280f705",
          4088 => x"3370852a",
          4089 => x"70810651",
          4090 => x"55557380",
          4091 => x"2e833886",
          4092 => x"56758295",
          4093 => x"3881fb98",
          4094 => x"51ff95f5",
          4095 => x"3f0280f7",
          4096 => x"05337098",
          4097 => x"2b555573",
          4098 => x"80258538",
          4099 => x"86569039",
          4100 => x"0280d205",
          4101 => x"33810654",
          4102 => x"73802e83",
          4103 => x"38875675",
          4104 => x"81e7386a",
          4105 => x"527751c6",
          4106 => x"bc3f8293",
          4107 => x"c8080284",
          4108 => x"0580d205",
          4109 => x"3370842a",
          4110 => x"70810651",
          4111 => x"56565773",
          4112 => x"802e80e5",
          4113 => x"3881fb9c",
          4114 => x"51ff95a5",
          4115 => x"3f877855",
          4116 => x"56941408",
          4117 => x"772e80d1",
          4118 => x"3881fba0",
          4119 => x"51ff9591",
          4120 => x"3f775976",
          4121 => x"5b81fba4",
          4122 => x"51ff9585",
          4123 => x"3f805289",
          4124 => x"3d705254",
          4125 => x"c1823f82",
          4126 => x"93c80856",
          4127 => x"8293c808",
          4128 => x"81873882",
          4129 => x"93c80852",
          4130 => x"7351c6c0",
          4131 => x"3f8293c8",
          4132 => x"08568293",
          4133 => x"c8088338",
          4134 => x"87567584",
          4135 => x"32703070",
          4136 => x"72079f2c",
          4137 => x"78065856",
          4138 => x"547580dd",
          4139 => x"3881fba8",
          4140 => x"51ff94bd",
          4141 => x"3f9f3dd4",
          4142 => x"0551c9a4",
          4143 => x"3f8293c8",
          4144 => x"088293c8",
          4145 => x"08307082",
          4146 => x"93c80807",
          4147 => x"80257930",
          4148 => x"707b079f",
          4149 => x"2a720652",
          4150 => x"57515656",
          4151 => x"74802e9b",
          4152 => x"3881fbac",
          4153 => x"51ff9489",
          4154 => x"3f805376",
          4155 => x"529f3dd4",
          4156 => x"0551ffba",
          4157 => x"b63f8293",
          4158 => x"c8085675",
          4159 => x"8c387751",
          4160 => x"ffb48b3f",
          4161 => x"8293c808",
          4162 => x"5681fbb0",
          4163 => x"51ff93e1",
          4164 => x"3f758293",
          4165 => x"c80c9f3d",
          4166 => x"0d04ea3d",
          4167 => x"0d825398",
          4168 => x"3dc00552",
          4169 => x"993d51d3",
          4170 => x"b33f8293",
          4171 => x"c8085582",
          4172 => x"93c80882",
          4173 => x"b538775d",
          4174 => x"6852983d",
          4175 => x"d40551cd",
          4176 => x"cb3f8293",
          4177 => x"c8085582",
          4178 => x"93c80883",
          4179 => x"38885574",
          4180 => x"842e0981",
          4181 => x"06829338",
          4182 => x"0280db05",
          4183 => x"3370852a",
          4184 => x"70810651",
          4185 => x"55567380",
          4186 => x"2e833886",
          4187 => x"5574842e",
          4188 => x"09810681",
          4189 => x"f5387759",
          4190 => x"8052983d",
          4191 => x"c40551ff",
          4192 => x"badc3f82",
          4193 => x"93c80856",
          4194 => x"80558293",
          4195 => x"c808752e",
          4196 => x"09810683",
          4197 => x"38875575",
          4198 => x"812e0981",
          4199 => x"06833882",
          4200 => x"5575ff2e",
          4201 => x"09810683",
          4202 => x"38815582",
          4203 => x"88b20a57",
          4204 => x"7481aa38",
          4205 => x"75527751",
          4206 => x"ffbdc73f",
          4207 => x"8293c808",
          4208 => x"558293c8",
          4209 => x"08819638",
          4210 => x"8b53a052",
          4211 => x"b41851ff",
          4212 => x"affa3f77",
          4213 => x"54ae0bb4",
          4214 => x"15347754",
          4215 => x"900bbf15",
          4216 => x"34765280",
          4217 => x"ca1851ff",
          4218 => x"af8f3f75",
          4219 => x"53b41852",
          4220 => x"7751c3aa",
          4221 => x"3fa053b4",
          4222 => x"185280d4",
          4223 => x"1851ffaf",
          4224 => x"a73f7754",
          4225 => x"ae0b80d5",
          4226 => x"15347e53",
          4227 => x"80d41852",
          4228 => x"7751c38a",
          4229 => x"3f775481",
          4230 => x"0b831534",
          4231 => x"983dd405",
          4232 => x"51c5e73f",
          4233 => x"8293c808",
          4234 => x"558293c8",
          4235 => x"08af3876",
          4236 => x"52639605",
          4237 => x"51ffaec1",
          4238 => x"3f755363",
          4239 => x"527751c2",
          4240 => x"dd3f6354",
          4241 => x"900b8b15",
          4242 => x"34775481",
          4243 => x"0b831534",
          4244 => x"7751ffb1",
          4245 => x"b93f8293",
          4246 => x"c808558e",
          4247 => x"39805375",
          4248 => x"52983dc4",
          4249 => x"0551ffb7",
          4250 => x"c23f7482",
          4251 => x"93c80c98",
          4252 => x"3d0d04db",
          4253 => x"3d0da83d",
          4254 => x"840551cd",
          4255 => x"c83f8253",
          4256 => x"a73dff84",
          4257 => x"0552a83d",
          4258 => x"51d0d13f",
          4259 => x"8293c808",
          4260 => x"558293c8",
          4261 => x"0882d738",
          4262 => x"774ca83d",
          4263 => x"0852a73d",
          4264 => x"d40551ca",
          4265 => x"e73f8293",
          4266 => x"c8085582",
          4267 => x"93c80882",
          4268 => x"bd380281",
          4269 => x"97053381",
          4270 => x"a0065473",
          4271 => x"802e8338",
          4272 => x"86557482",
          4273 => x"a938a053",
          4274 => x"a33d0852",
          4275 => x"a73dff88",
          4276 => x"0551ffad",
          4277 => x"d33fac53",
          4278 => x"a73dd405",
          4279 => x"52913d70",
          4280 => x"5254ffad",
          4281 => x"c33fa93d",
          4282 => x"08527351",
          4283 => x"ca9e3f82",
          4284 => x"93c80855",
          4285 => x"8293c808",
          4286 => x"9438626e",
          4287 => x"2e098106",
          4288 => x"8a388455",
          4289 => x"64a13d08",
          4290 => x"2e833888",
          4291 => x"5574842e",
          4292 => x"09810681",
          4293 => x"b838a73d",
          4294 => x"ffa80551",
          4295 => x"c3ec3f82",
          4296 => x"93c80855",
          4297 => x"8293c808",
          4298 => x"81c43867",
          4299 => x"569353a7",
          4300 => x"3dff9505",
          4301 => x"528d1651",
          4302 => x"ffaced3f",
          4303 => x"02ab0533",
          4304 => x"8b17348b",
          4305 => x"16337084",
          4306 => x"2a708106",
          4307 => x"51555773",
          4308 => x"893876a0",
          4309 => x"0754738b",
          4310 => x"17347754",
          4311 => x"810b8315",
          4312 => x"348b1633",
          4313 => x"70842a70",
          4314 => x"81065155",
          4315 => x"5773802e",
          4316 => x"80db386d",
          4317 => x"632e80d5",
          4318 => x"38755277",
          4319 => x"51ffbfe5",
          4320 => x"3f8293c8",
          4321 => x"08527751",
          4322 => x"ffb0b23f",
          4323 => x"82558293",
          4324 => x"c808802e",
          4325 => x"b8388293",
          4326 => x"c8085277",
          4327 => x"51ffaea7",
          4328 => x"3f8293c8",
          4329 => x"0880d419",
          4330 => x"57558293",
          4331 => x"c808bf38",
          4332 => x"81163354",
          4333 => x"73ae2e09",
          4334 => x"81069238",
          4335 => x"62537552",
          4336 => x"7751ffbf",
          4337 => x"d93f7754",
          4338 => x"810b8315",
          4339 => x"34749f38",
          4340 => x"a73dd405",
          4341 => x"51c3893f",
          4342 => x"8293c808",
          4343 => x"558293c8",
          4344 => x"088c3877",
          4345 => x"51ffaea6",
          4346 => x"3f8293c8",
          4347 => x"08557482",
          4348 => x"93c80ca7",
          4349 => x"3d0d04ed",
          4350 => x"3d0d0280",
          4351 => x"db053302",
          4352 => x"840580df",
          4353 => x"05335757",
          4354 => x"8253953d",
          4355 => x"d0055296",
          4356 => x"3d51cdc8",
          4357 => x"3f8293c8",
          4358 => x"08558293",
          4359 => x"c80880d4",
          4360 => x"38785a65",
          4361 => x"52953dd4",
          4362 => x"0551c7e0",
          4363 => x"3f8293c8",
          4364 => x"08558293",
          4365 => x"c808bd38",
          4366 => x"0280cf05",
          4367 => x"3381a006",
          4368 => x"5473802e",
          4369 => x"83388655",
          4370 => x"74aa3875",
          4371 => x"a7066171",
          4372 => x"098b1233",
          4373 => x"71067a74",
          4374 => x"06075157",
          4375 => x"5556748b",
          4376 => x"15347854",
          4377 => x"810b8315",
          4378 => x"347851ff",
          4379 => x"ada03f82",
          4380 => x"93c80855",
          4381 => x"748293c8",
          4382 => x"0c953d0d",
          4383 => x"04ee3d0d",
          4384 => x"65568253",
          4385 => x"943dd005",
          4386 => x"52953d51",
          4387 => x"ccce3f82",
          4388 => x"93c80855",
          4389 => x"8293c808",
          4390 => x"80d33877",
          4391 => x"59645294",
          4392 => x"3dd40551",
          4393 => x"c6e63f82",
          4394 => x"93c80855",
          4395 => x"8293c808",
          4396 => x"bc380280",
          4397 => x"cb053381",
          4398 => x"a0065473",
          4399 => x"802e8338",
          4400 => x"865574a9",
          4401 => x"38861622",
          4402 => x"84172270",
          4403 => x"902b7207",
          4404 => x"5457547f",
          4405 => x"960551ff",
          4406 => x"a99f3f77",
          4407 => x"54810b83",
          4408 => x"15347751",
          4409 => x"ffaca73f",
          4410 => x"8293c808",
          4411 => x"55748293",
          4412 => x"c80c943d",
          4413 => x"0d04ea3d",
          4414 => x"0d696b5c",
          4415 => x"59805398",
          4416 => x"3dd00552",
          4417 => x"993d51cb",
          4418 => x"d33f8293",
          4419 => x"c8088293",
          4420 => x"c8083070",
          4421 => x"8293c808",
          4422 => x"0780257b",
          4423 => x"30707d07",
          4424 => x"9f2a7206",
          4425 => x"52575156",
          4426 => x"5674802e",
          4427 => x"80f6387b",
          4428 => x"5d805f80",
          4429 => x"528d3d70",
          4430 => x"5254ffb7",
          4431 => x"bb3f8293",
          4432 => x"c8085682",
          4433 => x"93c80880",
          4434 => x"ce388152",
          4435 => x"7351ffbc",
          4436 => x"fb3f8293",
          4437 => x"c8085682",
          4438 => x"93c808bb",
          4439 => x"388293c8",
          4440 => x"088293c8",
          4441 => x"08655c58",
          4442 => x"58791781",
          4443 => x"187a1a56",
          4444 => x"58557433",
          4445 => x"74348118",
          4446 => x"588a7727",
          4447 => x"ec387719",
          4448 => x"54807434",
          4449 => x"77802e8f",
          4450 => x"38ff1879",
          4451 => x"11703351",
          4452 => x"555873a0",
          4453 => x"2ee83875",
          4454 => x"842e0981",
          4455 => x"06863880",
          4456 => x"79348056",
          4457 => x"75307077",
          4458 => x"0780257c",
          4459 => x"30707e07",
          4460 => x"9f2a7206",
          4461 => x"52565155",
          4462 => x"74802ebc",
          4463 => x"387ba011",
          4464 => x"085351ff",
          4465 => x"aa813f82",
          4466 => x"93c80856",
          4467 => x"8293c808",
          4468 => x"a7387b70",
          4469 => x"33515480",
          4470 => x"c3587383",
          4471 => x"2e8b3880",
          4472 => x"e4587384",
          4473 => x"2e8338a7",
          4474 => x"587b18b4",
          4475 => x"0551ffa6",
          4476 => x"c13f8293",
          4477 => x"c8087b0c",
          4478 => x"758293c8",
          4479 => x"0c983d0d",
          4480 => x"04e83d0d",
          4481 => x"82539a3d",
          4482 => x"ffb80552",
          4483 => x"9b3d51c9",
          4484 => x"cb3f8293",
          4485 => x"c8085582",
          4486 => x"93c80883",
          4487 => x"c8388b53",
          4488 => x"a0529a3d",
          4489 => x"ffbc0551",
          4490 => x"ffa7a13f",
          4491 => x"806b7071",
          4492 => x"33525755",
          4493 => x"579f7427",
          4494 => x"81b53874",
          4495 => x"336b8105",
          4496 => x"4c7081ff",
          4497 => x"065256ff",
          4498 => x"a7fe3f82",
          4499 => x"93c80880",
          4500 => x"2ea2386a",
          4501 => x"70337053",
          4502 => x"5154ffa7",
          4503 => x"f23f8293",
          4504 => x"c808802e",
          4505 => x"8d387588",
          4506 => x"2b74076b",
          4507 => x"81054c56",
          4508 => x"83398056",
          4509 => x"ff9f1654",
          4510 => x"7399268a",
          4511 => x"38e01670",
          4512 => x"83ffff06",
          4513 => x"575480ff",
          4514 => x"76278738",
          4515 => x"81faf816",
          4516 => x"33567580",
          4517 => x"2ea33875",
          4518 => x"5281fcf8",
          4519 => x"51ffa6f7",
          4520 => x"3f8293c8",
          4521 => x"08933881",
          4522 => x"ff762788",
          4523 => x"38768926",
          4524 => x"88388b39",
          4525 => x"8a772786",
          4526 => x"38865582",
          4527 => x"a83981ff",
          4528 => x"76279338",
          4529 => x"9a3d7705",
          4530 => x"ffbc0576",
          4531 => x"882a5555",
          4532 => x"73753481",
          4533 => x"17579a3d",
          4534 => x"7705ffbc",
          4535 => x"05547574",
          4536 => x"3481176b",
          4537 => x"70335656",
          4538 => x"57739f26",
          4539 => x"fecd3889",
          4540 => x"3d335486",
          4541 => x"557381e5",
          4542 => x"2e81ea38",
          4543 => x"76802ea8",
          4544 => x"38029f05",
          4545 => x"70781270",
          4546 => x"33515256",
          4547 => x"5473a02e",
          4548 => x"09810694",
          4549 => x"38ff1757",
          4550 => x"76802e8c",
          4551 => x"38761570",
          4552 => x"33515473",
          4553 => x"a02eee38",
          4554 => x"775f8041",
          4555 => x"80528f3d",
          4556 => x"705255ff",
          4557 => x"b3c23f82",
          4558 => x"93c80854",
          4559 => x"8293c808",
          4560 => x"81a13881",
          4561 => x"527451ff",
          4562 => x"b9823f82",
          4563 => x"93c80854",
          4564 => x"8293c808",
          4565 => x"b0387680",
          4566 => x"2e91388b",
          4567 => x"539a3dff",
          4568 => x"bc055265",
          4569 => x"51ffa4c0",
          4570 => x"3f863965",
          4571 => x"54e57434",
          4572 => x"7754810b",
          4573 => x"83153477",
          4574 => x"51ffa792",
          4575 => x"3f8293c8",
          4576 => x"085480df",
          4577 => x"398293c8",
          4578 => x"08842e09",
          4579 => x"810680d3",
          4580 => x"38805476",
          4581 => x"742e80cb",
          4582 => x"3881529a",
          4583 => x"3dd40551",
          4584 => x"ffb6b23f",
          4585 => x"8293c808",
          4586 => x"548293c8",
          4587 => x"08b538a0",
          4588 => x"538293c8",
          4589 => x"08526551",
          4590 => x"ffa4913f",
          4591 => x"6554880b",
          4592 => x"8b15348b",
          4593 => x"539a3dff",
          4594 => x"bc055265",
          4595 => x"51ffa3d8",
          4596 => x"3f775481",
          4597 => x"0b831534",
          4598 => x"7751ffa6",
          4599 => x"b13f8293",
          4600 => x"c8085473",
          4601 => x"55748293",
          4602 => x"c80c9a3d",
          4603 => x"0d04f13d",
          4604 => x"0d616302",
          4605 => x"880580cf",
          4606 => x"0533943d",
          4607 => x"fc055572",
          4608 => x"545e5c58",
          4609 => x"cda23f82",
          4610 => x"93c80857",
          4611 => x"8293c808",
          4612 => x"8a389118",
          4613 => x"33577680",
          4614 => x"2e863876",
          4615 => x"5482b739",
          4616 => x"7a802e95",
          4617 => x"388c1808",
          4618 => x"90389018",
          4619 => x"3370812a",
          4620 => x"70810651",
          4621 => x"55557390",
          4622 => x"38875482",
          4623 => x"99398257",
          4624 => x"81893981",
          4625 => x"57818439",
          4626 => x"7f8a1122",
          4627 => x"70892b70",
          4628 => x"557d5458",
          4629 => x"5154fef9",
          4630 => x"dd3fff16",
          4631 => x"7b067030",
          4632 => x"7072079f",
          4633 => x"2a8293c8",
          4634 => x"0805628c",
          4635 => x"11085d52",
          4636 => x"40555580",
          4637 => x"5f817927",
          4638 => x"88389814",
          4639 => x"08792683",
          4640 => x"38825978",
          4641 => x"79565d80",
          4642 => x"5a745277",
          4643 => x"51ffa6d7",
          4644 => x"3f8293c8",
          4645 => x"08811661",
          4646 => x"56565698",
          4647 => x"14087526",
          4648 => x"83388255",
          4649 => x"75812eff",
          4650 => x"953875ff",
          4651 => x"2eff9438",
          4652 => x"758b3881",
          4653 => x"1a5a797e",
          4654 => x"2e913885",
          4655 => x"39745d80",
          4656 => x"5a74792e",
          4657 => x"098106c1",
          4658 => x"38875776",
          4659 => x"8186387b",
          4660 => x"802eb938",
          4661 => x"7c7e5755",
          4662 => x"7d802eb3",
          4663 => x"38811554",
          4664 => x"75812e09",
          4665 => x"81068338",
          4666 => x"ff547353",
          4667 => x"74527f51",
          4668 => x"ffa7f03f",
          4669 => x"8293c808",
          4670 => x"578293c8",
          4671 => x"08913874",
          4672 => x"8116ff18",
          4673 => x"58565f75",
          4674 => x"d4388439",
          4675 => x"ff1d5f76",
          4676 => x"80c2387f",
          4677 => x"7f8c120c",
          4678 => x"547b802e",
          4679 => x"b7387c88",
          4680 => x"190c7a8c",
          4681 => x"190c9018",
          4682 => x"3380c007",
          4683 => x"54739019",
          4684 => x"347f9811",
          4685 => x"08fe0555",
          4686 => x"55901508",
          4687 => x"74269538",
          4688 => x"9015087e",
          4689 => x"3190160c",
          4690 => x"7f841133",
          4691 => x"81075555",
          4692 => x"73841634",
          4693 => x"76547382",
          4694 => x"93c80c91",
          4695 => x"3d0d04ea",
          4696 => x"3d0d6a02",
          4697 => x"840580e7",
          4698 => x"05339b3d",
          4699 => x"535e58ff",
          4700 => x"bfd33f82",
          4701 => x"93c80856",
          4702 => x"8b57800b",
          4703 => x"8293c808",
          4704 => x"248cd138",
          4705 => x"8293c808",
          4706 => x"10108293",
          4707 => x"e4055574",
          4708 => x"08802e87",
          4709 => x"38740855",
          4710 => x"80753475",
          4711 => x"81ff065a",
          4712 => x"81527951",
          4713 => x"ff99cb3f",
          4714 => x"8293c808",
          4715 => x"81ff0670",
          4716 => x"81065656",
          4717 => x"8357748c",
          4718 => x"9b387582",
          4719 => x"2a708106",
          4720 => x"51558a57",
          4721 => x"748c8d38",
          4722 => x"983dfc05",
          4723 => x"53835279",
          4724 => x"51ff9ddd",
          4725 => x"3f8293c8",
          4726 => x"08983866",
          4727 => x"802e9338",
          4728 => x"66828080",
          4729 => x"268c3866",
          4730 => x"ff056706",
          4731 => x"5574802e",
          4732 => x"83388147",
          4733 => x"84805e77",
          4734 => x"802e8638",
          4735 => x"7d782692",
          4736 => x"38778180",
          4737 => x"0a268b38",
          4738 => x"ff187806",
          4739 => x"5574802e",
          4740 => x"86389357",
          4741 => x"8bbe397d",
          4742 => x"527751fe",
          4743 => x"f6983f82",
          4744 => x"93c8086c",
          4745 => x"7f546e53",
          4746 => x"4058fef6",
          4747 => x"893f8293",
          4748 => x"c8087e82",
          4749 => x"93c80829",
          4750 => x"60307062",
          4751 => x"07802582",
          4752 => x"93c80830",
          4753 => x"708293c8",
          4754 => x"08078025",
          4755 => x"72075259",
          4756 => x"51584641",
          4757 => x"9157758a",
          4758 => x"fb38983d",
          4759 => x"f8055381",
          4760 => x"527951ff",
          4761 => x"9ccb3f81",
          4762 => x"578293c8",
          4763 => x"088ae538",
          4764 => x"7c832a70",
          4765 => x"81065155",
          4766 => x"80447464",
          4767 => x"2e098106",
          4768 => x"8338bf44",
          4769 => x"8e576366",
          4770 => x"268ac938",
          4771 => x"65643146",
          4772 => x"8e5780ff",
          4773 => x"66278abc",
          4774 => x"38935777",
          4775 => x"8180268a",
          4776 => x"b3387c81",
          4777 => x"2a708106",
          4778 => x"51557480",
          4779 => x"2e95387c",
          4780 => x"87065574",
          4781 => x"822e8838",
          4782 => x"7c810655",
          4783 => x"74853883",
          4784 => x"428f397c",
          4785 => x"81065593",
          4786 => x"57824274",
          4787 => x"802e8a84",
          4788 => x"38775961",
          4789 => x"832e0981",
          4790 => x"0680f138",
          4791 => x"77b43865",
          4792 => x"912a785c",
          4793 => x"57810b81",
          4794 => x"fd9c7071",
          4795 => x"22525856",
          4796 => x"5974802e",
          4797 => x"9d387477",
          4798 => x"26983881",
          4799 => x"1b791071",
          4800 => x"10187022",
          4801 => x"51575a5b",
          4802 => x"74802e86",
          4803 => x"38767527",
          4804 => x"ea387852",
          4805 => x"6551fef4",
          4806 => x"9d3f8293",
          4807 => x"c8088293",
          4808 => x"c8081010",
          4809 => x"1f7f5487",
          4810 => x"055256fe",
          4811 => x"f4883f82",
          4812 => x"93c8085c",
          4813 => x"a05b800b",
          4814 => x"fc808a17",
          4815 => x"5643fdff",
          4816 => x"f00a7527",
          4817 => x"818b388e",
          4818 => x"57898939",
          4819 => x"77b43865",
          4820 => x"8c2a785c",
          4821 => x"57810b81",
          4822 => x"fd8c7071",
          4823 => x"22525856",
          4824 => x"5974802e",
          4825 => x"9d387477",
          4826 => x"26983881",
          4827 => x"1b791071",
          4828 => x"10187022",
          4829 => x"51575a5b",
          4830 => x"74802e86",
          4831 => x"38767527",
          4832 => x"ea387852",
          4833 => x"6551fef3",
          4834 => x"ad3f8293",
          4835 => x"c8081084",
          4836 => x"05578293",
          4837 => x"c8089ff5",
          4838 => x"26923881",
          4839 => x"0b8293c8",
          4840 => x"08832911",
          4841 => x"70722a83",
          4842 => x"05515842",
          4843 => x"7d52761e",
          4844 => x"ff0551fe",
          4845 => x"f3803f82",
          4846 => x"93c8085c",
          4847 => x"817e535b",
          4848 => x"81808051",
          4849 => x"fef2ef3f",
          4850 => x"8293c808",
          4851 => x"83ffff06",
          4852 => x"43631b7c",
          4853 => x"11640568",
          4854 => x"11ff0569",
          4855 => x"30707206",
          4856 => x"73315258",
          4857 => x"59574061",
          4858 => x"832e0981",
          4859 => x"06893876",
          4860 => x"1b601841",
          4861 => x"5b843976",
          4862 => x"1c5c7890",
          4863 => x"29167065",
          4864 => x"31515574",
          4865 => x"662687be",
          4866 => x"38657b31",
          4867 => x"7c317953",
          4868 => x"70643152",
          4869 => x"56fef29e",
          4870 => x"3f8293c8",
          4871 => x"08566183",
          4872 => x"2e098106",
          4873 => x"9b388293",
          4874 => x"c80883ff",
          4875 => x"f5269138",
          4876 => x"77893878",
          4877 => x"812a5877",
          4878 => x"fd97388e",
          4879 => x"57879539",
          4880 => x"61822e09",
          4881 => x"810680d3",
          4882 => x"3883fff5",
          4883 => x"7627b438",
          4884 => x"778f3878",
          4885 => x"19557480",
          4886 => x"c0268638",
          4887 => x"7458fcf1",
          4888 => x"397c812a",
          4889 => x"81065574",
          4890 => x"802e8638",
          4891 => x"8342fce1",
          4892 => x"39778b38",
          4893 => x"78195881",
          4894 => x"807827fc",
          4895 => x"d4388e57",
          4896 => x"86d23975",
          4897 => x"9ff52693",
          4898 => x"38778b38",
          4899 => x"78195881",
          4900 => x"807827fc",
          4901 => x"bc388e57",
          4902 => x"86ba3980",
          4903 => x"5561812e",
          4904 => x"09810683",
          4905 => x"38615575",
          4906 => x"9ff52675",
          4907 => x"06558e57",
          4908 => x"7486a138",
          4909 => x"7d538052",
          4910 => x"7e51ff9a",
          4911 => x"8f3f8b53",
          4912 => x"81fbb452",
          4913 => x"7e51ff99",
          4914 => x"df3f7d52",
          4915 => x"8b1f51ff",
          4916 => x"99893f78",
          4917 => x"7f8d0534",
          4918 => x"7a83ffff",
          4919 => x"06528e1f",
          4920 => x"51ff98f7",
          4921 => x"3f817f90",
          4922 => x"05346183",
          4923 => x"32703070",
          4924 => x"962a8480",
          4925 => x"06545155",
          4926 => x"911f51ff",
          4927 => x"98dd3f65",
          4928 => x"83ffff26",
          4929 => x"90380280",
          4930 => x"d6052252",
          4931 => x"931f51ff",
          4932 => x"98c93f8a",
          4933 => x"396552a0",
          4934 => x"1f51ff98",
          4935 => x"dc3ff87f",
          4936 => x"950534bf",
          4937 => x"52981f51",
          4938 => x"ff98b03f",
          4939 => x"81ff529a",
          4940 => x"1f51ff98",
          4941 => x"a63f6352",
          4942 => x"9c1f51ff",
          4943 => x"98bb3f61",
          4944 => x"832e0981",
          4945 => x"0680cf38",
          4946 => x"8288b20a",
          4947 => x"5280c31f",
          4948 => x"51ff98a5",
          4949 => x"3f7b52a4",
          4950 => x"1f51ff98",
          4951 => x"9c3f8252",
          4952 => x"ac1f51ff",
          4953 => x"98933f81",
          4954 => x"52b01f51",
          4955 => x"ff97ec3f",
          4956 => x"8652b21f",
          4957 => x"51ff97e3",
          4958 => x"3fff807f",
          4959 => x"80c00534",
          4960 => x"a97f80c2",
          4961 => x"05349353",
          4962 => x"81fbc052",
          4963 => x"80c71f51",
          4964 => x"ff98953f",
          4965 => x"b2398288",
          4966 => x"b20a52a7",
          4967 => x"1f51ff97",
          4968 => x"d83f7b83",
          4969 => x"ffff0652",
          4970 => x"961f51ff",
          4971 => x"97ad3fff",
          4972 => x"807fa405",
          4973 => x"34a97fa6",
          4974 => x"05349353",
          4975 => x"81fbd452",
          4976 => x"ab1f51ff",
          4977 => x"97e23f82",
          4978 => x"d4d55283",
          4979 => x"fe1f51ff",
          4980 => x"97893f81",
          4981 => x"5463537e",
          4982 => x"527951ff",
          4983 => x"93f93f81",
          4984 => x"578293c8",
          4985 => x"0883ed38",
          4986 => x"61832e09",
          4987 => x"810680f0",
          4988 => x"38815463",
          4989 => x"8605537e",
          4990 => x"527951ff",
          4991 => x"93d93f7d",
          4992 => x"5380527e",
          4993 => x"51ff97c4",
          4994 => x"3f848b85",
          4995 => x"a4d2527e",
          4996 => x"51ff96e5",
          4997 => x"3f868a85",
          4998 => x"e4f25283",
          4999 => x"e41f51ff",
          5000 => x"96d73fff",
          5001 => x"165283e8",
          5002 => x"1f51ff96",
          5003 => x"cc3f8252",
          5004 => x"83ec1f51",
          5005 => x"ff96c23f",
          5006 => x"82d4d552",
          5007 => x"83fe1f51",
          5008 => x"ff96983f",
          5009 => x"81546387",
          5010 => x"05537e52",
          5011 => x"7951ff93",
          5012 => x"863f8154",
          5013 => x"63810553",
          5014 => x"7e527951",
          5015 => x"ff92f83f",
          5016 => x"64538052",
          5017 => x"7e51ff96",
          5018 => x"e33f7f56",
          5019 => x"805b6183",
          5020 => x"2e098106",
          5021 => x"9e38f852",
          5022 => x"7e51ff95",
          5023 => x"fc3fff52",
          5024 => x"841f51ff",
          5025 => x"95f33ff0",
          5026 => x"0a52881f",
          5027 => x"51ff95e9",
          5028 => x"3f953987",
          5029 => x"fffff855",
          5030 => x"61812e83",
          5031 => x"38f85574",
          5032 => x"527e51ff",
          5033 => x"95d33f7b",
          5034 => x"55605774",
          5035 => x"61268338",
          5036 => x"74577654",
          5037 => x"75537e52",
          5038 => x"7951ff92",
          5039 => x"9a3f8293",
          5040 => x"c8088286",
          5041 => x"387d5380",
          5042 => x"527e51ff",
          5043 => x"95fe3f76",
          5044 => x"16757831",
          5045 => x"565674d1",
          5046 => x"38811b5b",
          5047 => x"7a802eff",
          5048 => x"8d387855",
          5049 => x"61832e83",
          5050 => x"38625560",
          5051 => x"57746126",
          5052 => x"83387457",
          5053 => x"76547553",
          5054 => x"7e527951",
          5055 => x"ff91d83f",
          5056 => x"8293c808",
          5057 => x"81c83876",
          5058 => x"16757831",
          5059 => x"565674db",
          5060 => x"388c5761",
          5061 => x"832e9338",
          5062 => x"86576583",
          5063 => x"ffff268a",
          5064 => x"38845761",
          5065 => x"822e8338",
          5066 => x"81577c83",
          5067 => x"2a810658",
          5068 => x"7780ff38",
          5069 => x"7d537752",
          5070 => x"7e51ff95",
          5071 => x"8f3f82d4",
          5072 => x"d55283fe",
          5073 => x"1f51ff94",
          5074 => x"923f83be",
          5075 => x"1f567776",
          5076 => x"34810b81",
          5077 => x"1734810b",
          5078 => x"82173477",
          5079 => x"83173476",
          5080 => x"84173463",
          5081 => x"66055780",
          5082 => x"fdc15276",
          5083 => x"51feebc6",
          5084 => x"3ffe0b85",
          5085 => x"17348293",
          5086 => x"c808822a",
          5087 => x"bf075574",
          5088 => x"86173482",
          5089 => x"93c80887",
          5090 => x"17346352",
          5091 => x"83c61f51",
          5092 => x"ff93e63f",
          5093 => x"655283ca",
          5094 => x"1f51ff93",
          5095 => x"dc3f8154",
          5096 => x"77537e52",
          5097 => x"7951ff90",
          5098 => x"ae3f8157",
          5099 => x"8293c808",
          5100 => x"a3388053",
          5101 => x"80527951",
          5102 => x"ff91f63f",
          5103 => x"81578293",
          5104 => x"c8089138",
          5105 => x"8d398e57",
          5106 => x"8b398157",
          5107 => x"87398157",
          5108 => x"83398057",
          5109 => x"768293c8",
          5110 => x"0c983d0d",
          5111 => x"04ff3d0d",
          5112 => x"73527193",
          5113 => x"2681e238",
          5114 => x"71101081",
          5115 => x"f1b80552",
          5116 => x"71080482",
          5117 => x"81f851ff",
          5118 => x"80a93f81",
          5119 => x"d4398282",
          5120 => x"8451ff80",
          5121 => x"9e3f81c9",
          5122 => x"39828298",
          5123 => x"51ff8093",
          5124 => x"3f81be39",
          5125 => x"8282ac51",
          5126 => x"ff80883f",
          5127 => x"81b33982",
          5128 => x"82bc51fe",
          5129 => x"fffd3f81",
          5130 => x"a8398282",
          5131 => x"cc51feff",
          5132 => x"f23f819d",
          5133 => x"398282e0",
          5134 => x"51feffe7",
          5135 => x"3f819239",
          5136 => x"8282f051",
          5137 => x"feffdc3f",
          5138 => x"81873982",
          5139 => x"838851fe",
          5140 => x"ffd13f80",
          5141 => x"fc398283",
          5142 => x"a051feff",
          5143 => x"c63f80f1",
          5144 => x"398283b8",
          5145 => x"51feffbb",
          5146 => x"3f80e639",
          5147 => x"8283d451",
          5148 => x"feffb03f",
          5149 => x"80db3982",
          5150 => x"83e851fe",
          5151 => x"ffa53f80",
          5152 => x"d0398284",
          5153 => x"9451feff",
          5154 => x"9a3f80c5",
          5155 => x"398284a8",
          5156 => x"51feff8f",
          5157 => x"3fbb3982",
          5158 => x"84c851fe",
          5159 => x"ff853fb1",
          5160 => x"398284dc",
          5161 => x"51fefefb",
          5162 => x"3fa73982",
          5163 => x"84f451fe",
          5164 => x"fef13f9d",
          5165 => x"3982858c",
          5166 => x"51fefee7",
          5167 => x"3f933982",
          5168 => x"85a451fe",
          5169 => x"fedd3f89",
          5170 => x"398285b0",
          5171 => x"51fefed3",
          5172 => x"3f833d0d",
          5173 => x"04fb3d0d",
          5174 => x"77795656",
          5175 => x"7487e726",
          5176 => x"93387452",
          5177 => x"7587e829",
          5178 => x"51fee8ca",
          5179 => x"3f8293c8",
          5180 => x"08559a39",
          5181 => x"87e85274",
          5182 => x"51fee8ba",
          5183 => x"3f8293c8",
          5184 => x"08527551",
          5185 => x"fee8af3f",
          5186 => x"8293c808",
          5187 => x"55745479",
          5188 => x"53755282",
          5189 => x"85c051ff",
          5190 => x"84833f87",
          5191 => x"3d0d04fe",
          5192 => x"ec3d0d81",
          5193 => x"973d0881",
          5194 => x"993d0802",
          5195 => x"880584e3",
          5196 => x"05337173",
          5197 => x"30707507",
          5198 => x"802587ff",
          5199 => x"75270754",
          5200 => x"595a5c57",
          5201 => x"58935575",
          5202 => x"81873881",
          5203 => x"53775281",
          5204 => x"963dfbd8",
          5205 => x"0551ffbc",
          5206 => x"993f8293",
          5207 => x"c8085882",
          5208 => x"93c808bb",
          5209 => x"388293c8",
          5210 => x"0887c098",
          5211 => x"880c8293",
          5212 => x"c8085981",
          5213 => x"963dfbd4",
          5214 => x"11555584",
          5215 => x"80537652",
          5216 => x"fbd81551",
          5217 => x"c0f23f82",
          5218 => x"93c80858",
          5219 => x"8293c808",
          5220 => x"8e387a80",
          5221 => x"2e89387a",
          5222 => x"197b1858",
          5223 => x"59d53981",
          5224 => x"963dfbd8",
          5225 => x"0551cac1",
          5226 => x"3f773070",
          5227 => x"79078025",
          5228 => x"7b30709f",
          5229 => x"2a720651",
          5230 => x"57515674",
          5231 => x"802e9038",
          5232 => x"8285e453",
          5233 => x"87c09888",
          5234 => x"08527851",
          5235 => x"fe873f77",
          5236 => x"55748293",
          5237 => x"c80c8196",
          5238 => x"3d0d04f8",
          5239 => x"3d0d02b7",
          5240 => x"053357ff",
          5241 => x"7d575980",
          5242 => x"537b527a",
          5243 => x"51feb03f",
          5244 => x"8293c808",
          5245 => x"a4387680",
          5246 => x"2e883876",
          5247 => x"812e9838",
          5248 => x"98396155",
          5249 => x"60548293",
          5250 => x"c8537f52",
          5251 => x"7e51752d",
          5252 => x"8293c808",
          5253 => x"59833975",
          5254 => x"04788293",
          5255 => x"c80c8a3d",
          5256 => x"0d04fb3d",
          5257 => x"0d029f05",
          5258 => x"338285ec",
          5259 => x"538285f4",
          5260 => x"5256ff81",
          5261 => x"e83f828b",
          5262 => x"e8702252",
          5263 => x"55fef9d6",
          5264 => x"3f828680",
          5265 => x"5482868c",
          5266 => x"53811533",
          5267 => x"52828694",
          5268 => x"51ff81c9",
          5269 => x"3f75802e",
          5270 => x"8538fef6",
          5271 => x"ff3f873d",
          5272 => x"0d04fe3d",
          5273 => x"0d87c096",
          5274 => x"800853fe",
          5275 => x"f9ff3f81",
          5276 => x"51feeeff",
          5277 => x"3f8286b0",
          5278 => x"51fef0f5",
          5279 => x"3f8051fe",
          5280 => x"eef13f72",
          5281 => x"812a7081",
          5282 => x"06515271",
          5283 => x"802e9538",
          5284 => x"8151feee",
          5285 => x"de3f8286",
          5286 => x"cc51fef0",
          5287 => x"d43f8051",
          5288 => x"feeed03f",
          5289 => x"72822a70",
          5290 => x"81065152",
          5291 => x"71802e95",
          5292 => x"388151fe",
          5293 => x"eebd3f82",
          5294 => x"86e051fe",
          5295 => x"f0b33f80",
          5296 => x"51feeeaf",
          5297 => x"3f72832a",
          5298 => x"70810651",
          5299 => x"5271802e",
          5300 => x"95388151",
          5301 => x"feee9c3f",
          5302 => x"8286f051",
          5303 => x"fef0923f",
          5304 => x"8051feee",
          5305 => x"8e3f7284",
          5306 => x"2a708106",
          5307 => x"51527180",
          5308 => x"2e953881",
          5309 => x"51feedfb",
          5310 => x"3f828784",
          5311 => x"51feeff1",
          5312 => x"3f8051fe",
          5313 => x"eded3f72",
          5314 => x"852a7081",
          5315 => x"06515271",
          5316 => x"802e9538",
          5317 => x"8151feed",
          5318 => x"da3f8287",
          5319 => x"9851feef",
          5320 => x"d03f8051",
          5321 => x"feedcc3f",
          5322 => x"72862a70",
          5323 => x"81065152",
          5324 => x"71802e95",
          5325 => x"388151fe",
          5326 => x"edb93f82",
          5327 => x"87ac51fe",
          5328 => x"efaf3f80",
          5329 => x"51feedab",
          5330 => x"3f72872a",
          5331 => x"70810651",
          5332 => x"5271802e",
          5333 => x"95388151",
          5334 => x"feed983f",
          5335 => x"8287c051",
          5336 => x"feef8e3f",
          5337 => x"8051feed",
          5338 => x"8a3f7288",
          5339 => x"2a708106",
          5340 => x"51527180",
          5341 => x"2e953881",
          5342 => x"51feecf7",
          5343 => x"3f8287d4",
          5344 => x"51feeeed",
          5345 => x"3f8051fe",
          5346 => x"ece93ffe",
          5347 => x"f8a83f84",
          5348 => x"3d0d04fa",
          5349 => x"3d0d7870",
          5350 => x"08705556",
          5351 => x"5774802e",
          5352 => x"80ed388e",
          5353 => x"3974770c",
          5354 => x"85143353",
          5355 => x"80e13981",
          5356 => x"15558075",
          5357 => x"33545472",
          5358 => x"a02e8338",
          5359 => x"81547230",
          5360 => x"709f2a75",
          5361 => x"06515372",
          5362 => x"e6387433",
          5363 => x"5372a02e",
          5364 => x"09810688",
          5365 => x"38807570",
          5366 => x"81055734",
          5367 => x"80567590",
          5368 => x"29828c88",
          5369 => x"05770853",
          5370 => x"70085254",
          5371 => x"fee6d03f",
          5372 => x"8293c808",
          5373 => x"8b388414",
          5374 => x"33537281",
          5375 => x"2effa638",
          5376 => x"81167081",
          5377 => x"ff065753",
          5378 => x"bb7627d2",
          5379 => x"38ff5372",
          5380 => x"8293c80c",
          5381 => x"883d0d04",
          5382 => x"ce3d0d80",
          5383 => x"7082b6c8",
          5384 => x"72710c5d",
          5385 => x"5e5c8c5a",
          5386 => x"81527b51",
          5387 => x"ff84c33f",
          5388 => x"8293c808",
          5389 => x"81ff0659",
          5390 => x"787c2e09",
          5391 => x"81069f38",
          5392 => x"82889452",
          5393 => x"963d7052",
          5394 => x"59fefde7",
          5395 => x"3f7b5378",
          5396 => x"52eab01b",
          5397 => x"51ffb5ab",
          5398 => x"3f8293c8",
          5399 => x"085a7980",
          5400 => x"2e8b3882",
          5401 => x"889851fe",
          5402 => x"fdb33f85",
          5403 => x"3981705e",
          5404 => x"5c8288d0",
          5405 => x"51fef7ab",
          5406 => x"3f963d70",
          5407 => x"435980f8",
          5408 => x"70545a80",
          5409 => x"527851fe",
          5410 => x"e4a43f79",
          5411 => x"526151fe",
          5412 => x"fde53fb4",
          5413 => x"3dfef805",
          5414 => x"51fdf83f",
          5415 => x"8293c808",
          5416 => x"902b7090",
          5417 => x"2c515978",
          5418 => x"81872685",
          5419 => x"af387810",
          5420 => x"1081f288",
          5421 => x"05597808",
          5422 => x"04b43dfe",
          5423 => x"f41153fe",
          5424 => x"f80551fe",
          5425 => x"fee23f82",
          5426 => x"93c8088c",
          5427 => x"388288d4",
          5428 => x"51fefcc9",
          5429 => x"3fff9a39",
          5430 => x"b43dfef0",
          5431 => x"1153fef8",
          5432 => x"0551fefe",
          5433 => x"c33f8293",
          5434 => x"c808802e",
          5435 => x"88388160",
          5436 => x"25833880",
          5437 => x"4002bf05",
          5438 => x"33520280",
          5439 => x"c3053351",
          5440 => x"ff82ef3f",
          5441 => x"8293c808",
          5442 => x"81ff0659",
          5443 => x"788e3882",
          5444 => x"88e451fe",
          5445 => x"f68d3f81",
          5446 => x"5dfed639",
          5447 => x"8288f451",
          5448 => x"fef6803f",
          5449 => x"fecb39b4",
          5450 => x"3dfef411",
          5451 => x"53fef805",
          5452 => x"51fefdf4",
          5453 => x"3f8293c8",
          5454 => x"08802efe",
          5455 => x"b4388053",
          5456 => x"80520280",
          5457 => x"c3053351",
          5458 => x"ff86e63f",
          5459 => x"8293c808",
          5460 => x"5282898c",
          5461 => x"51fefbc5",
          5462 => x"3ffe9639",
          5463 => x"b43dfef4",
          5464 => x"1153fef8",
          5465 => x"0551fefd",
          5466 => x"bf3f8293",
          5467 => x"c808802e",
          5468 => x"87386089",
          5469 => x"26fdfa38",
          5470 => x"b43dfef0",
          5471 => x"1153fef8",
          5472 => x"0551fefd",
          5473 => x"a33f8293",
          5474 => x"c8088638",
          5475 => x"8293c808",
          5476 => x"40605382",
          5477 => x"89945296",
          5478 => x"3d705259",
          5479 => x"fefb943f",
          5480 => x"02bf0533",
          5481 => x"53785260",
          5482 => x"84b42982",
          5483 => x"a0f80551",
          5484 => x"ffb2d03f",
          5485 => x"8293c808",
          5486 => x"802e8c38",
          5487 => x"8293c808",
          5488 => x"51f49a3f",
          5489 => x"fdab3982",
          5490 => x"88e451fe",
          5491 => x"f4d53f81",
          5492 => x"5cfd9e39",
          5493 => x"b43dfef8",
          5494 => x"0551fee4",
          5495 => x"a43f8293",
          5496 => x"c808b53d",
          5497 => x"fef80552",
          5498 => x"5bfee4fa",
          5499 => x"3f815382",
          5500 => x"93c80852",
          5501 => x"7a51f6a7",
          5502 => x"3f8293c8",
          5503 => x"08802efc",
          5504 => x"f0388293",
          5505 => x"c80851f3",
          5506 => x"d43ffce5",
          5507 => x"39b43dfe",
          5508 => x"f80551fe",
          5509 => x"e3eb3f82",
          5510 => x"93c808b5",
          5511 => x"3dfef805",
          5512 => x"525bfee4",
          5513 => x"c13f8293",
          5514 => x"c808b53d",
          5515 => x"fef80552",
          5516 => x"5afee4b2",
          5517 => x"3f8293c8",
          5518 => x"08b53dfe",
          5519 => x"f8055259",
          5520 => x"fee4a33f",
          5521 => x"828bc458",
          5522 => x"8293fc57",
          5523 => x"80568055",
          5524 => x"8293c808",
          5525 => x"81ff0654",
          5526 => x"78537952",
          5527 => x"7a51f6fb",
          5528 => x"3f8293c8",
          5529 => x"08802efc",
          5530 => x"88388293",
          5531 => x"c80851f2",
          5532 => x"ec3ffbfd",
          5533 => x"39828998",
          5534 => x"51fef3a7",
          5535 => x"3f8251fe",
          5536 => x"f28f3ffb",
          5537 => x"ec398289",
          5538 => x"b051fef3",
          5539 => x"963fa251",
          5540 => x"fef1e23f",
          5541 => x"fbdb3984",
          5542 => x"80810b87",
          5543 => x"c094840c",
          5544 => x"8480810b",
          5545 => x"87c09494",
          5546 => x"0c8289c8",
          5547 => x"51fef2f3",
          5548 => x"3ffbbe39",
          5549 => x"8289dc51",
          5550 => x"fef2e83f",
          5551 => x"8c80830b",
          5552 => x"87c09484",
          5553 => x"0c8c8083",
          5554 => x"0b87c094",
          5555 => x"940cfba1",
          5556 => x"39b43dfe",
          5557 => x"f41153fe",
          5558 => x"f80551fe",
          5559 => x"faca3f82",
          5560 => x"93c80880",
          5561 => x"2efb8a38",
          5562 => x"60528289",
          5563 => x"f051fef8",
          5564 => x"ac3f6059",
          5565 => x"7804b43d",
          5566 => x"fef41153",
          5567 => x"fef80551",
          5568 => x"fefaa53f",
          5569 => x"8293c808",
          5570 => x"802efae5",
          5571 => x"38605282",
          5572 => x"8a8c51fe",
          5573 => x"f8873f60",
          5574 => x"59782d82",
          5575 => x"93c8085e",
          5576 => x"8293c808",
          5577 => x"802efac9",
          5578 => x"388293c8",
          5579 => x"0852828a",
          5580 => x"a851fef7",
          5581 => x"e83ffab9",
          5582 => x"39828ac4",
          5583 => x"51fef1e3",
          5584 => x"3ffed1bc",
          5585 => x"3ffaaa39",
          5586 => x"828ae051",
          5587 => x"fef1d43f",
          5588 => x"8059ffa0",
          5589 => x"39feed84",
          5590 => x"3ffa9639",
          5591 => x"61703351",
          5592 => x"5978802e",
          5593 => x"fa8b387c",
          5594 => x"7c065978",
          5595 => x"802e80cb",
          5596 => x"38b43dfe",
          5597 => x"f80551fe",
          5598 => x"e1873f82",
          5599 => x"8af45682",
          5600 => x"93c80855",
          5601 => x"828af854",
          5602 => x"8053828a",
          5603 => x"fc52a03d",
          5604 => x"705259fe",
          5605 => x"f79d3f82",
          5606 => x"8bc45882",
          5607 => x"93fc5780",
          5608 => x"56618105",
          5609 => x"42615580",
          5610 => x"54838080",
          5611 => x"53838080",
          5612 => x"527851f4",
          5613 => x"a63f8293",
          5614 => x"c8085e7c",
          5615 => x"81327c81",
          5616 => x"32075978",
          5617 => x"8a387dff",
          5618 => x"2e098106",
          5619 => x"f9a33882",
          5620 => x"8b8c51fe",
          5621 => x"f6c73ff9",
          5622 => x"9839803d",
          5623 => x"0d800b82",
          5624 => x"93fc349b",
          5625 => x"9086e40b",
          5626 => x"87c0948c",
          5627 => x"0c9b9086",
          5628 => x"e40b87c0",
          5629 => x"949c0c8c",
          5630 => x"80830b87",
          5631 => x"c094840c",
          5632 => x"8c80830b",
          5633 => x"87c09494",
          5634 => x"0c80d48d",
          5635 => x"0b8293d8",
          5636 => x"0c80d780",
          5637 => x"0b8293dc",
          5638 => x"0cfee887",
          5639 => x"3ffeeecd",
          5640 => x"3f828b9c",
          5641 => x"51fee5c9",
          5642 => x"3f828ba8",
          5643 => x"51feeff3",
          5644 => x"3f81e4e2",
          5645 => x"51feeeb0",
          5646 => x"3f8151f3",
          5647 => x"e53ff7d8",
          5648 => x"3f800400",
          5649 => x"00002f5d",
          5650 => x"00002f30",
          5651 => x"00002f39",
          5652 => x"00002f42",
          5653 => x"00002f4b",
          5654 => x"00002f54",
          5655 => x"000031cf",
          5656 => x"000031c0",
          5657 => x"000031d7",
          5658 => x"000031df",
          5659 => x"000031df",
          5660 => x"000031df",
          5661 => x"000031df",
          5662 => x"000031df",
          5663 => x"000031df",
          5664 => x"000031df",
          5665 => x"000031df",
          5666 => x"000031df",
          5667 => x"000031df",
          5668 => x"000031d3",
          5669 => x"000031df",
          5670 => x"000031df",
          5671 => x"000031df",
          5672 => x"00003153",
          5673 => x"000031df",
          5674 => x"000031d7",
          5675 => x"000031df",
          5676 => x"000031df",
          5677 => x"000031db",
          5678 => x"000070bf",
          5679 => x"00006ff3",
          5680 => x"00006ffe",
          5681 => x"00007009",
          5682 => x"00007014",
          5683 => x"0000701f",
          5684 => x"0000702a",
          5685 => x"00007035",
          5686 => x"00007040",
          5687 => x"0000704b",
          5688 => x"00007056",
          5689 => x"00007061",
          5690 => x"0000706c",
          5691 => x"00007077",
          5692 => x"00007082",
          5693 => x"0000708d",
          5694 => x"00007097",
          5695 => x"000070a1",
          5696 => x"000070ab",
          5697 => x"000070b5",
          5698 => x"00007471",
          5699 => x"0000775c",
          5700 => x"000074b9",
          5701 => x"0000775c",
          5702 => x"00007527",
          5703 => x"0000775c",
          5704 => x"0000775c",
          5705 => x"0000775c",
          5706 => x"0000775c",
          5707 => x"0000775c",
          5708 => x"0000775c",
          5709 => x"0000775c",
          5710 => x"0000775c",
          5711 => x"0000775c",
          5712 => x"0000775c",
          5713 => x"0000775c",
          5714 => x"0000775c",
          5715 => x"0000775c",
          5716 => x"0000775c",
          5717 => x"0000775c",
          5718 => x"0000755c",
          5719 => x"0000775c",
          5720 => x"0000775c",
          5721 => x"0000775c",
          5722 => x"0000775c",
          5723 => x"0000775c",
          5724 => x"0000775c",
          5725 => x"0000775c",
          5726 => x"0000775c",
          5727 => x"0000775c",
          5728 => x"0000775c",
          5729 => x"0000775c",
          5730 => x"0000775c",
          5731 => x"0000775c",
          5732 => x"0000775c",
          5733 => x"0000775c",
          5734 => x"0000775c",
          5735 => x"0000775c",
          5736 => x"0000775c",
          5737 => x"0000775c",
          5738 => x"0000775c",
          5739 => x"0000775c",
          5740 => x"0000775c",
          5741 => x"000075d4",
          5742 => x"0000775c",
          5743 => x"0000775c",
          5744 => x"0000775c",
          5745 => x"0000775c",
          5746 => x"0000760d",
          5747 => x"0000775c",
          5748 => x"0000775c",
          5749 => x"0000775c",
          5750 => x"0000775c",
          5751 => x"0000775c",
          5752 => x"0000775c",
          5753 => x"0000775c",
          5754 => x"0000775c",
          5755 => x"0000775c",
          5756 => x"0000775c",
          5757 => x"0000775c",
          5758 => x"0000775c",
          5759 => x"0000775c",
          5760 => x"0000775c",
          5761 => x"0000775c",
          5762 => x"0000775c",
          5763 => x"0000775c",
          5764 => x"0000775c",
          5765 => x"0000775c",
          5766 => x"0000775c",
          5767 => x"0000775c",
          5768 => x"0000775c",
          5769 => x"0000775c",
          5770 => x"0000775c",
          5771 => x"0000775c",
          5772 => x"0000775c",
          5773 => x"0000775c",
          5774 => x"0000775c",
          5775 => x"0000775c",
          5776 => x"0000775c",
          5777 => x"0000775c",
          5778 => x"00007675",
          5779 => x"00007686",
          5780 => x"0000775c",
          5781 => x"0000775c",
          5782 => x"00007697",
          5783 => x"000076b4",
          5784 => x"0000775c",
          5785 => x"0000775c",
          5786 => x"0000775c",
          5787 => x"0000775c",
          5788 => x"0000775c",
          5789 => x"0000775c",
          5790 => x"0000775c",
          5791 => x"0000775c",
          5792 => x"0000775c",
          5793 => x"0000775c",
          5794 => x"0000775c",
          5795 => x"0000775c",
          5796 => x"0000775c",
          5797 => x"0000775c",
          5798 => x"0000775c",
          5799 => x"0000775c",
          5800 => x"0000775c",
          5801 => x"0000775c",
          5802 => x"0000775c",
          5803 => x"0000775c",
          5804 => x"0000775c",
          5805 => x"0000775c",
          5806 => x"0000775c",
          5807 => x"0000775c",
          5808 => x"0000775c",
          5809 => x"0000775c",
          5810 => x"0000775c",
          5811 => x"0000775c",
          5812 => x"0000775c",
          5813 => x"0000775c",
          5814 => x"0000775c",
          5815 => x"0000775c",
          5816 => x"0000775c",
          5817 => x"0000775c",
          5818 => x"000076d1",
          5819 => x"000076f6",
          5820 => x"0000775c",
          5821 => x"0000775c",
          5822 => x"0000775c",
          5823 => x"0000775c",
          5824 => x"0000775c",
          5825 => x"0000775c",
          5826 => x"0000775c",
          5827 => x"0000775c",
          5828 => x"00007739",
          5829 => x"00007748",
          5830 => x"0000775c",
          5831 => x"00007755",
          5832 => x"0000775c",
          5833 => x"00007471",
          5834 => x"25642f25",
          5835 => x"642f2564",
          5836 => x"2025643a",
          5837 => x"25643a25",
          5838 => x"642e2564",
          5839 => x"25640a00",
          5840 => x"536f4320",
          5841 => x"436f6e66",
          5842 => x"69677572",
          5843 => x"6174696f",
          5844 => x"6e000000",
          5845 => x"20286672",
          5846 => x"6f6d2053",
          5847 => x"6f432063",
          5848 => x"6f6e6669",
          5849 => x"67290000",
          5850 => x"3a0a4465",
          5851 => x"76696365",
          5852 => x"7320696d",
          5853 => x"706c656d",
          5854 => x"656e7465",
          5855 => x"643a0a00",
          5856 => x"20202020",
          5857 => x"494e534e",
          5858 => x"20425241",
          5859 => x"4d202853",
          5860 => x"74617274",
          5861 => x"3d253038",
          5862 => x"582c2053",
          5863 => x"697a653d",
          5864 => x"25303858",
          5865 => x"292e0a00",
          5866 => x"20202020",
          5867 => x"4252414d",
          5868 => x"20285374",
          5869 => x"6172743d",
          5870 => x"25303858",
          5871 => x"2c205369",
          5872 => x"7a653d25",
          5873 => x"30385829",
          5874 => x"2e0a0000",
          5875 => x"20202020",
          5876 => x"52414d20",
          5877 => x"28537461",
          5878 => x"72743d25",
          5879 => x"3038582c",
          5880 => x"2053697a",
          5881 => x"653d2530",
          5882 => x"3858292e",
          5883 => x"0a000000",
          5884 => x"20202020",
          5885 => x"494f4354",
          5886 => x"4c0a0000",
          5887 => x"20202020",
          5888 => x"5053320a",
          5889 => x"00000000",
          5890 => x"20202020",
          5891 => x"5350490a",
          5892 => x"00000000",
          5893 => x"20202020",
          5894 => x"53442043",
          5895 => x"61726420",
          5896 => x"28446576",
          5897 => x"69636573",
          5898 => x"3d253032",
          5899 => x"58292e0a",
          5900 => x"00000000",
          5901 => x"20202020",
          5902 => x"494e5445",
          5903 => x"52525550",
          5904 => x"5420434f",
          5905 => x"4e54524f",
          5906 => x"4c4c4552",
          5907 => x"0a000000",
          5908 => x"20202020",
          5909 => x"54494d45",
          5910 => x"52312028",
          5911 => x"54696d65",
          5912 => x"72733d25",
          5913 => x"30315829",
          5914 => x"2e0a0000",
          5915 => x"41646472",
          5916 => x"65737365",
          5917 => x"733a0a00",
          5918 => x"20202020",
          5919 => x"43505520",
          5920 => x"52657365",
          5921 => x"74205665",
          5922 => x"63746f72",
          5923 => x"20416464",
          5924 => x"72657373",
          5925 => x"203d2025",
          5926 => x"3038580a",
          5927 => x"00000000",
          5928 => x"20202020",
          5929 => x"43505520",
          5930 => x"4d656d6f",
          5931 => x"72792053",
          5932 => x"74617274",
          5933 => x"20416464",
          5934 => x"72657373",
          5935 => x"203d2025",
          5936 => x"3038580a",
          5937 => x"00000000",
          5938 => x"20202020",
          5939 => x"53746163",
          5940 => x"6b205374",
          5941 => x"61727420",
          5942 => x"41646472",
          5943 => x"65737320",
          5944 => x"20202020",
          5945 => x"203d2025",
          5946 => x"3038580a",
          5947 => x"00000000",
          5948 => x"20202020",
          5949 => x"5a505520",
          5950 => x"49642020",
          5951 => x"20202020",
          5952 => x"20202020",
          5953 => x"20202020",
          5954 => x"20202020",
          5955 => x"203d2025",
          5956 => x"3038580a",
          5957 => x"00000000",
          5958 => x"20202020",
          5959 => x"53797374",
          5960 => x"656d2043",
          5961 => x"6c6f636b",
          5962 => x"20467265",
          5963 => x"71202020",
          5964 => x"20202020",
          5965 => x"203d2025",
          5966 => x"3038580a",
          5967 => x"00000000",
          5968 => x"536d616c",
          5969 => x"6c000000",
          5970 => x"4d656469",
          5971 => x"756d0000",
          5972 => x"466c6578",
          5973 => x"00000000",
          5974 => x"45564f00",
          5975 => x"45564f6d",
          5976 => x"696e0000",
          5977 => x"556e6b6e",
          5978 => x"6f776e00",
          5979 => x"53440000",
          5980 => x"222a2b2c",
          5981 => x"3a3b3c3d",
          5982 => x"3e3f5b5d",
          5983 => x"7c7f0000",
          5984 => x"46415400",
          5985 => x"46415433",
          5986 => x"32000000",
          5987 => x"300a0000",
          5988 => x"310a0000",
          5989 => x"320a0000",
          5990 => x"330a0000",
          5991 => x"350a0000",
          5992 => x"360a0000",
          5993 => x"370a0000",
          5994 => x"380a0000",
          5995 => x"390a0000",
          5996 => x"31300a00",
          5997 => x"ebfe904d",
          5998 => x"53444f53",
          5999 => x"352e3000",
          6000 => x"4e4f204e",
          6001 => x"414d4520",
          6002 => x"20202046",
          6003 => x"41543332",
          6004 => x"20202000",
          6005 => x"4e4f204e",
          6006 => x"414d4520",
          6007 => x"20202046",
          6008 => x"41542020",
          6009 => x"20202000",
          6010 => x"00007d6c",
          6011 => x"00000000",
          6012 => x"00000000",
          6013 => x"00000000",
          6014 => x"809a4541",
          6015 => x"8e418f80",
          6016 => x"45454549",
          6017 => x"49498e8f",
          6018 => x"9092924f",
          6019 => x"994f5555",
          6020 => x"59999a9b",
          6021 => x"9c9d9e9f",
          6022 => x"41494f55",
          6023 => x"a5a5a6a7",
          6024 => x"a8a9aaab",
          6025 => x"acadaeaf",
          6026 => x"b0b1b2b3",
          6027 => x"b4b5b6b7",
          6028 => x"b8b9babb",
          6029 => x"bcbdbebf",
          6030 => x"c0c1c2c3",
          6031 => x"c4c5c6c7",
          6032 => x"c8c9cacb",
          6033 => x"cccdcecf",
          6034 => x"d0d1d2d3",
          6035 => x"d4d5d6d7",
          6036 => x"d8d9dadb",
          6037 => x"dcdddedf",
          6038 => x"e0e1e2e3",
          6039 => x"e4e5e6e7",
          6040 => x"e8e9eaeb",
          6041 => x"ecedeeef",
          6042 => x"f0f1f2f3",
          6043 => x"f4f5f6f7",
          6044 => x"f8f9fafb",
          6045 => x"fcfdfeff",
          6046 => x"2b2e2c3b",
          6047 => x"3d5b5d2f",
          6048 => x"5c222a3a",
          6049 => x"3c3e3f7c",
          6050 => x"7f000000",
          6051 => x"00010004",
          6052 => x"00100040",
          6053 => x"01000200",
          6054 => x"00000000",
          6055 => x"00010002",
          6056 => x"00040008",
          6057 => x"00100020",
          6058 => x"00000000",
          6059 => x"46415431",
          6060 => x"32000000",
          6061 => x"46415431",
          6062 => x"36000000",
          6063 => x"65784641",
          6064 => x"54000000",
          6065 => x"4449534b",
          6066 => x"20494f20",
          6067 => x"434f4e54",
          6068 => x"524f4c53",
          6069 => x"00000000",
          6070 => x"4449534b",
          6071 => x"20425546",
          6072 => x"46455220",
          6073 => x"434f4e54",
          6074 => x"524f4c53",
          6075 => x"00000000",
          6076 => x"46494c45",
          6077 => x"53595354",
          6078 => x"454d2043",
          6079 => x"4f4e5452",
          6080 => x"4f4c5300",
          6081 => x"4d454d4f",
          6082 => x"52590000",
          6083 => x"48415244",
          6084 => x"57415245",
          6085 => x"00000000",
          6086 => x"54455354",
          6087 => x"494e4700",
          6088 => x"45584543",
          6089 => x"5554494f",
          6090 => x"4e000000",
          6091 => x"4d495343",
          6092 => x"20434f4d",
          6093 => x"4d414e44",
          6094 => x"53000000",
          6095 => x"6464756d",
          6096 => x"70000000",
          6097 => x"64696e69",
          6098 => x"74000000",
          6099 => x"64737461",
          6100 => x"74000000",
          6101 => x"64696f63",
          6102 => x"746c0000",
          6103 => x"6264756d",
          6104 => x"70000000",
          6105 => x"62656469",
          6106 => x"74000000",
          6107 => x"62726561",
          6108 => x"64000000",
          6109 => x"62777269",
          6110 => x"74650000",
          6111 => x"6266696c",
          6112 => x"6c000000",
          6113 => x"626c656e",
          6114 => x"00000000",
          6115 => x"66696e69",
          6116 => x"74000000",
          6117 => x"666f7065",
          6118 => x"6e000000",
          6119 => x"66636c6f",
          6120 => x"73650000",
          6121 => x"66736565",
          6122 => x"6b000000",
          6123 => x"66726561",
          6124 => x"64000000",
          6125 => x"66696e73",
          6126 => x"70656374",
          6127 => x"00000000",
          6128 => x"66777269",
          6129 => x"74650000",
          6130 => x"66747275",
          6131 => x"6e630000",
          6132 => x"66616c6c",
          6133 => x"6f630000",
          6134 => x"66617474",
          6135 => x"72000000",
          6136 => x"6674696d",
          6137 => x"65000000",
          6138 => x"6672656e",
          6139 => x"616d6500",
          6140 => x"6664656c",
          6141 => x"00000000",
          6142 => x"666d6b64",
          6143 => x"69720000",
          6144 => x"66737461",
          6145 => x"74000000",
          6146 => x"66646972",
          6147 => x"00000000",
          6148 => x"66636174",
          6149 => x"00000000",
          6150 => x"66637000",
          6151 => x"66636f6e",
          6152 => x"63617400",
          6153 => x"66787472",
          6154 => x"61637400",
          6155 => x"666c6f61",
          6156 => x"64000000",
          6157 => x"66657865",
          6158 => x"63000000",
          6159 => x"66736176",
          6160 => x"65000000",
          6161 => x"6664756d",
          6162 => x"70000000",
          6163 => x"66636400",
          6164 => x"66647269",
          6165 => x"76650000",
          6166 => x"6673686f",
          6167 => x"77646972",
          6168 => x"00000000",
          6169 => x"666c6162",
          6170 => x"656c0000",
          6171 => x"666d6b66",
          6172 => x"73000000",
          6173 => x"6d636c72",
          6174 => x"00000000",
          6175 => x"6d64756d",
          6176 => x"70000000",
          6177 => x"6d656200",
          6178 => x"6d656800",
          6179 => x"6d657700",
          6180 => x"68696400",
          6181 => x"68696500",
          6182 => x"68720000",
          6183 => x"68740000",
          6184 => x"68666400",
          6185 => x"68666500",
          6186 => x"64687279",
          6187 => x"00000000",
          6188 => x"636f7265",
          6189 => x"6d61726b",
          6190 => x"00000000",
          6191 => x"63616c6c",
          6192 => x"00000000",
          6193 => x"6a6d7000",
          6194 => x"72657374",
          6195 => x"61727400",
          6196 => x"72657365",
          6197 => x"74000000",
          6198 => x"68656c70",
          6199 => x"00000000",
          6200 => x"696e666f",
          6201 => x"00000000",
          6202 => x"74696d65",
          6203 => x"00000000",
          6204 => x"74657374",
          6205 => x"00000000",
          6206 => x"4469736b",
          6207 => x"20457272",
          6208 => x"6f720a00",
          6209 => x"496e7465",
          6210 => x"726e616c",
          6211 => x"20657272",
          6212 => x"6f722e0a",
          6213 => x"00000000",
          6214 => x"4469736b",
          6215 => x"206e6f74",
          6216 => x"20726561",
          6217 => x"64792e0a",
          6218 => x"00000000",
          6219 => x"4e6f2066",
          6220 => x"696c6520",
          6221 => x"666f756e",
          6222 => x"642e0a00",
          6223 => x"4e6f2070",
          6224 => x"61746820",
          6225 => x"666f756e",
          6226 => x"642e0a00",
          6227 => x"496e7661",
          6228 => x"6c696420",
          6229 => x"66696c65",
          6230 => x"6e616d65",
          6231 => x"2e0a0000",
          6232 => x"41636365",
          6233 => x"73732064",
          6234 => x"656e6965",
          6235 => x"642e0a00",
          6236 => x"46696c65",
          6237 => x"20616c72",
          6238 => x"65616479",
          6239 => x"20657869",
          6240 => x"7374732e",
          6241 => x"0a000000",
          6242 => x"46696c65",
          6243 => x"2068616e",
          6244 => x"646c6520",
          6245 => x"696e7661",
          6246 => x"6c69642e",
          6247 => x"0a000000",
          6248 => x"53442069",
          6249 => x"73207772",
          6250 => x"69746520",
          6251 => x"70726f74",
          6252 => x"65637465",
          6253 => x"642e0a00",
          6254 => x"44726976",
          6255 => x"65206e75",
          6256 => x"6d626572",
          6257 => x"20697320",
          6258 => x"696e7661",
          6259 => x"6c69642e",
          6260 => x"0a000000",
          6261 => x"4469736b",
          6262 => x"206e6f74",
          6263 => x"20656e61",
          6264 => x"626c6564",
          6265 => x"2e0a0000",
          6266 => x"4e6f2063",
          6267 => x"6f6d7061",
          6268 => x"7469626c",
          6269 => x"65206669",
          6270 => x"6c657379",
          6271 => x"7374656d",
          6272 => x"20666f75",
          6273 => x"6e64206f",
          6274 => x"6e206469",
          6275 => x"736b2e0a",
          6276 => x"00000000",
          6277 => x"466f726d",
          6278 => x"61742061",
          6279 => x"626f7274",
          6280 => x"65642e0a",
          6281 => x"00000000",
          6282 => x"54696d65",
          6283 => x"6f75742c",
          6284 => x"206f7065",
          6285 => x"72617469",
          6286 => x"6f6e2063",
          6287 => x"616e6365",
          6288 => x"6c6c6564",
          6289 => x"2e0a0000",
          6290 => x"46696c65",
          6291 => x"20697320",
          6292 => x"6c6f636b",
          6293 => x"65642e0a",
          6294 => x"00000000",
          6295 => x"496e7375",
          6296 => x"66666963",
          6297 => x"69656e74",
          6298 => x"206d656d",
          6299 => x"6f72792e",
          6300 => x"0a000000",
          6301 => x"546f6f20",
          6302 => x"6d616e79",
          6303 => x"206f7065",
          6304 => x"6e206669",
          6305 => x"6c65732e",
          6306 => x"0a000000",
          6307 => x"50617261",
          6308 => x"6d657465",
          6309 => x"72732069",
          6310 => x"6e636f72",
          6311 => x"72656374",
          6312 => x"2e0a0000",
          6313 => x"53756363",
          6314 => x"6573732e",
          6315 => x"0a000000",
          6316 => x"556e6b6e",
          6317 => x"6f776e20",
          6318 => x"6572726f",
          6319 => x"722e0a00",
          6320 => x"0a256c75",
          6321 => x"20627974",
          6322 => x"65732025",
          6323 => x"73206174",
          6324 => x"20256c75",
          6325 => x"20627974",
          6326 => x"65732f73",
          6327 => x"65632e0a",
          6328 => x"00000000",
          6329 => x"72656164",
          6330 => x"00000000",
          6331 => x"5a505554",
          6332 => x"41000000",
          6333 => x"0a2a2a20",
          6334 => x"25732028",
          6335 => x"00000000",
          6336 => x"31382f30",
          6337 => x"372f3230",
          6338 => x"31390000",
          6339 => x"76312e33",
          6340 => x"00000000",
          6341 => x"205a5055",
          6342 => x"2c207265",
          6343 => x"76202530",
          6344 => x"32782920",
          6345 => x"25732025",
          6346 => x"73202a2a",
          6347 => x"0a0a0000",
          6348 => x"5a505554",
          6349 => x"4120496e",
          6350 => x"74657272",
          6351 => x"75707420",
          6352 => x"48616e64",
          6353 => x"6c65720a",
          6354 => x"00000000",
          6355 => x"54696d65",
          6356 => x"7220696e",
          6357 => x"74657272",
          6358 => x"7570740a",
          6359 => x"00000000",
          6360 => x"50533220",
          6361 => x"696e7465",
          6362 => x"72727570",
          6363 => x"740a0000",
          6364 => x"494f4354",
          6365 => x"4c205244",
          6366 => x"20696e74",
          6367 => x"65727275",
          6368 => x"70740a00",
          6369 => x"494f4354",
          6370 => x"4c205752",
          6371 => x"20696e74",
          6372 => x"65727275",
          6373 => x"70740a00",
          6374 => x"55415254",
          6375 => x"30205258",
          6376 => x"20696e74",
          6377 => x"65727275",
          6378 => x"70740a00",
          6379 => x"55415254",
          6380 => x"30205458",
          6381 => x"20696e74",
          6382 => x"65727275",
          6383 => x"70740a00",
          6384 => x"55415254",
          6385 => x"31205258",
          6386 => x"20696e74",
          6387 => x"65727275",
          6388 => x"70740a00",
          6389 => x"55415254",
          6390 => x"31205458",
          6391 => x"20696e74",
          6392 => x"65727275",
          6393 => x"70740a00",
          6394 => x"53657474",
          6395 => x"696e6720",
          6396 => x"75702074",
          6397 => x"696d6572",
          6398 => x"2e2e2e0a",
          6399 => x"00000000",
          6400 => x"456e6162",
          6401 => x"6c696e67",
          6402 => x"2074696d",
          6403 => x"65722e2e",
          6404 => x"2e0a0000",
          6405 => x"303a0000",
          6406 => x"4661696c",
          6407 => x"65642074",
          6408 => x"6f20696e",
          6409 => x"69746961",
          6410 => x"6c697365",
          6411 => x"20736420",
          6412 => x"63617264",
          6413 => x"20302c20",
          6414 => x"706c6561",
          6415 => x"73652069",
          6416 => x"6e697420",
          6417 => x"6d616e75",
          6418 => x"616c6c79",
          6419 => x"2e0a0000",
          6420 => x"2a200000",
          6421 => x"42616420",
          6422 => x"6469736b",
          6423 => x"20696421",
          6424 => x"0a000000",
          6425 => x"496e6974",
          6426 => x"69616c69",
          6427 => x"7365642e",
          6428 => x"0a000000",
          6429 => x"4661696c",
          6430 => x"65642074",
          6431 => x"6f20696e",
          6432 => x"69746961",
          6433 => x"6c697365",
          6434 => x"2e0a0000",
          6435 => x"72633d25",
          6436 => x"640a0000",
          6437 => x"25753a00",
          6438 => x"44697361",
          6439 => x"626c696e",
          6440 => x"6720696e",
          6441 => x"74657272",
          6442 => x"75707473",
          6443 => x"0a000000",
          6444 => x"456e6162",
          6445 => x"6c696e67",
          6446 => x"20696e74",
          6447 => x"65727275",
          6448 => x"7074730a",
          6449 => x"00000000",
          6450 => x"44697361",
          6451 => x"626c6564",
          6452 => x"20756172",
          6453 => x"74206669",
          6454 => x"666f0a00",
          6455 => x"456e6162",
          6456 => x"6c696e67",
          6457 => x"20756172",
          6458 => x"74206669",
          6459 => x"666f0a00",
          6460 => x"45786563",
          6461 => x"7574696e",
          6462 => x"6720636f",
          6463 => x"64652040",
          6464 => x"20253038",
          6465 => x"78202e2e",
          6466 => x"2e0a0000",
          6467 => x"43616c6c",
          6468 => x"696e6720",
          6469 => x"636f6465",
          6470 => x"20402025",
          6471 => x"30387820",
          6472 => x"2e2e2e0a",
          6473 => x"00000000",
          6474 => x"43616c6c",
          6475 => x"20726574",
          6476 => x"75726e65",
          6477 => x"6420636f",
          6478 => x"64652028",
          6479 => x"2564292e",
          6480 => x"0a000000",
          6481 => x"52657374",
          6482 => x"61727469",
          6483 => x"6e672061",
          6484 => x"70706c69",
          6485 => x"63617469",
          6486 => x"6f6e2e2e",
          6487 => x"2e0a0000",
          6488 => x"436f6c64",
          6489 => x"20726562",
          6490 => x"6f6f7469",
          6491 => x"6e672e2e",
          6492 => x"2e0a0000",
          6493 => x"5a505500",
          6494 => x"62696e00",
          6495 => x"25643a5c",
          6496 => x"25735c25",
          6497 => x"732e2573",
          6498 => x"00000000",
          6499 => x"42616420",
          6500 => x"636f6d6d",
          6501 => x"616e642e",
          6502 => x"0a000000",
          6503 => x"52756e6e",
          6504 => x"696e672e",
          6505 => x"2e2e0a00",
          6506 => x"456e6162",
          6507 => x"6c696e67",
          6508 => x"20696e74",
          6509 => x"65727275",
          6510 => x"7074732e",
          6511 => x"2e2e0a00",
          6512 => x"00000000",
          6513 => x"00000000",
          6514 => x"00007fff",
          6515 => x"00000000",
          6516 => x"00007fff",
          6517 => x"00010000",
          6518 => x"00007fff",
          6519 => x"00000000",
          6520 => x"00000000",
          6521 => x"00007800",
          6522 => x"00000000",
          6523 => x"05f5e100",
          6524 => x"00010101",
          6525 => x"01010101",
          6526 => x"80010101",
          6527 => x"01000000",
          6528 => x"00000000",
          6529 => x"01000000",
          6530 => x"00007f3c",
          6531 => x"00010100",
          6532 => x"00000000",
          6533 => x"00000000",
          6534 => x"00007f44",
          6535 => x"01020100",
          6536 => x"00000000",
          6537 => x"00000000",
          6538 => x"00007f4c",
          6539 => x"00030100",
          6540 => x"00000000",
          6541 => x"00000000",
          6542 => x"00007f54",
          6543 => x"01040100",
          6544 => x"00000000",
          6545 => x"00000000",
          6546 => x"00007f5c",
          6547 => x"000a0200",
          6548 => x"00000000",
          6549 => x"00000000",
          6550 => x"00007f64",
          6551 => x"000b0200",
          6552 => x"00000000",
          6553 => x"00000000",
          6554 => x"00007f6c",
          6555 => x"000c0200",
          6556 => x"00000000",
          6557 => x"00000000",
          6558 => x"00007f74",
          6559 => x"000d0200",
          6560 => x"00000000",
          6561 => x"00000000",
          6562 => x"00007f7c",
          6563 => x"000e0200",
          6564 => x"00000000",
          6565 => x"00000000",
          6566 => x"00007f84",
          6567 => x"000f0200",
          6568 => x"00000000",
          6569 => x"00000000",
          6570 => x"00007f8c",
          6571 => x"01140300",
          6572 => x"00000000",
          6573 => x"00000000",
          6574 => x"00007f94",
          6575 => x"00170300",
          6576 => x"00000000",
          6577 => x"00000000",
          6578 => x"00007f9c",
          6579 => x"00180300",
          6580 => x"00000000",
          6581 => x"00000000",
          6582 => x"00007fa4",
          6583 => x"00190300",
          6584 => x"00000000",
          6585 => x"00000000",
          6586 => x"00007fac",
          6587 => x"001a0300",
          6588 => x"00000000",
          6589 => x"00000000",
          6590 => x"00007fb4",
          6591 => x"001c0300",
          6592 => x"00000000",
          6593 => x"00000000",
          6594 => x"00007fc0",
          6595 => x"001d0300",
          6596 => x"00000000",
          6597 => x"00000000",
          6598 => x"00007fc8",
          6599 => x"001e0300",
          6600 => x"00000000",
          6601 => x"00000000",
          6602 => x"00007fd0",
          6603 => x"00220300",
          6604 => x"00000000",
          6605 => x"00000000",
          6606 => x"00007fd8",
          6607 => x"00230300",
          6608 => x"00000000",
          6609 => x"00000000",
          6610 => x"00007fe0",
          6611 => x"00240300",
          6612 => x"00000000",
          6613 => x"00000000",
          6614 => x"00007fe8",
          6615 => x"001f0300",
          6616 => x"00000000",
          6617 => x"00000000",
          6618 => x"00007ff0",
          6619 => x"00200300",
          6620 => x"00000000",
          6621 => x"00000000",
          6622 => x"00007ff8",
          6623 => x"00210300",
          6624 => x"00000000",
          6625 => x"00000000",
          6626 => x"00008000",
          6627 => x"00150300",
          6628 => x"00000000",
          6629 => x"00000000",
          6630 => x"00008008",
          6631 => x"00160300",
          6632 => x"00000000",
          6633 => x"00000000",
          6634 => x"00008010",
          6635 => x"001b0300",
          6636 => x"00000000",
          6637 => x"00000000",
          6638 => x"00008018",
          6639 => x"00250300",
          6640 => x"00000000",
          6641 => x"00000000",
          6642 => x"0000801c",
          6643 => x"002d0300",
          6644 => x"00000000",
          6645 => x"00000000",
          6646 => x"00008024",
          6647 => x"002e0300",
          6648 => x"00000000",
          6649 => x"00000000",
          6650 => x"0000802c",
          6651 => x"012b0300",
          6652 => x"00000000",
          6653 => x"00000000",
          6654 => x"00008034",
          6655 => x"01300300",
          6656 => x"00000000",
          6657 => x"00000000",
          6658 => x"0000803c",
          6659 => x"002f0300",
          6660 => x"00000000",
          6661 => x"00000000",
          6662 => x"00008044",
          6663 => x"002c0300",
          6664 => x"00000000",
          6665 => x"00000000",
          6666 => x"0000804c",
          6667 => x"00260300",
          6668 => x"00000000",
          6669 => x"00000000",
          6670 => x"00008050",
          6671 => x"00270300",
          6672 => x"00000000",
          6673 => x"00000000",
          6674 => x"00008058",
          6675 => x"00280300",
          6676 => x"00000000",
          6677 => x"00000000",
          6678 => x"00008064",
          6679 => x"00290300",
          6680 => x"00000000",
          6681 => x"00000000",
          6682 => x"0000806c",
          6683 => x"002a0300",
          6684 => x"00000000",
          6685 => x"00000000",
          6686 => x"00008074",
          6687 => x"003c0400",
          6688 => x"00000000",
          6689 => x"00000000",
          6690 => x"0000807c",
          6691 => x"003d0400",
          6692 => x"00000000",
          6693 => x"00000000",
          6694 => x"00008084",
          6695 => x"003e0400",
          6696 => x"00000000",
          6697 => x"00000000",
          6698 => x"00008088",
          6699 => x"003f0400",
          6700 => x"00000000",
          6701 => x"00000000",
          6702 => x"0000808c",
          6703 => x"00400400",
          6704 => x"00000000",
          6705 => x"00000000",
          6706 => x"00008090",
          6707 => x"01500500",
          6708 => x"00000000",
          6709 => x"00000000",
          6710 => x"00008094",
          6711 => x"01510500",
          6712 => x"00000000",
          6713 => x"00000000",
          6714 => x"00008098",
          6715 => x"00520500",
          6716 => x"00000000",
          6717 => x"00000000",
          6718 => x"0000809c",
          6719 => x"00530500",
          6720 => x"00000000",
          6721 => x"00000000",
          6722 => x"000080a0",
          6723 => x"01540500",
          6724 => x"00000000",
          6725 => x"00000000",
          6726 => x"000080a4",
          6727 => x"01550500",
          6728 => x"00000000",
          6729 => x"00000000",
          6730 => x"000080a8",
          6731 => x"00640600",
          6732 => x"00000000",
          6733 => x"00000000",
          6734 => x"000080b0",
          6735 => x"00650600",
          6736 => x"00000000",
          6737 => x"00000000",
          6738 => x"000080bc",
          6739 => x"01790700",
          6740 => x"00000000",
          6741 => x"00000000",
          6742 => x"000080c4",
          6743 => x"01780700",
          6744 => x"00000000",
          6745 => x"00000000",
          6746 => x"000080c8",
          6747 => x"01820800",
          6748 => x"00000000",
          6749 => x"00000000",
          6750 => x"000080d0",
          6751 => x"01830800",
          6752 => x"00000000",
          6753 => x"00000000",
          6754 => x"000080d8",
          6755 => x"00840800",
          6756 => x"00000000",
          6757 => x"00000000",
          6758 => x"000080e0",
          6759 => x"01850800",
          6760 => x"00000000",
          6761 => x"00000000",
          6762 => x"000080e8",
          6763 => x"00860800",
          6764 => x"00000000",
          6765 => x"00000000",
          6766 => x"000080f0",
          6767 => x"01870800",
          6768 => x"00000000",
          6769 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

