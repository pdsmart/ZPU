IOCP_SinglePortBRAM.vhd