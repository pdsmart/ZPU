SinglePortBRAM.vhd.uninitialized