IOCP_DualPortBootBRAM.vhd