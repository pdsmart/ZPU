-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"92",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"92",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"9f",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"bc",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"93",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"95",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"90",
           386 => x"2d",
           387 => x"08",
           388 => x"04",
           389 => x"0c",
           390 => x"81",
           391 => x"82",
           392 => x"81",
           393 => x"ab",
           394 => x"d3",
           395 => x"a0",
           396 => x"d3",
           397 => x"b9",
           398 => x"90",
           399 => x"90",
           400 => x"90",
           401 => x"2d",
           402 => x"08",
           403 => x"04",
           404 => x"0c",
           405 => x"81",
           406 => x"82",
           407 => x"81",
           408 => x"ab",
           409 => x"d3",
           410 => x"a0",
           411 => x"d3",
           412 => x"92",
           413 => x"90",
           414 => x"90",
           415 => x"90",
           416 => x"2d",
           417 => x"08",
           418 => x"04",
           419 => x"0c",
           420 => x"81",
           421 => x"82",
           422 => x"81",
           423 => x"b1",
           424 => x"d3",
           425 => x"a0",
           426 => x"d3",
           427 => x"d7",
           428 => x"90",
           429 => x"90",
           430 => x"90",
           431 => x"2d",
           432 => x"08",
           433 => x"04",
           434 => x"0c",
           435 => x"81",
           436 => x"82",
           437 => x"81",
           438 => x"9b",
           439 => x"d3",
           440 => x"a0",
           441 => x"d3",
           442 => x"dd",
           443 => x"90",
           444 => x"90",
           445 => x"90",
           446 => x"2d",
           447 => x"08",
           448 => x"04",
           449 => x"0c",
           450 => x"2d",
           451 => x"08",
           452 => x"04",
           453 => x"0c",
           454 => x"2d",
           455 => x"08",
           456 => x"04",
           457 => x"0c",
           458 => x"2d",
           459 => x"08",
           460 => x"04",
           461 => x"0c",
           462 => x"2d",
           463 => x"08",
           464 => x"04",
           465 => x"0c",
           466 => x"2d",
           467 => x"08",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"04",
           485 => x"0c",
           486 => x"2d",
           487 => x"08",
           488 => x"04",
           489 => x"0c",
           490 => x"2d",
           491 => x"08",
           492 => x"04",
           493 => x"0c",
           494 => x"2d",
           495 => x"08",
           496 => x"04",
           497 => x"0c",
           498 => x"2d",
           499 => x"08",
           500 => x"04",
           501 => x"0c",
           502 => x"2d",
           503 => x"08",
           504 => x"04",
           505 => x"0c",
           506 => x"2d",
           507 => x"08",
           508 => x"04",
           509 => x"0c",
           510 => x"2d",
           511 => x"08",
           512 => x"04",
           513 => x"0c",
           514 => x"2d",
           515 => x"08",
           516 => x"04",
           517 => x"0c",
           518 => x"2d",
           519 => x"08",
           520 => x"04",
           521 => x"0c",
           522 => x"2d",
           523 => x"08",
           524 => x"04",
           525 => x"0c",
           526 => x"2d",
           527 => x"08",
           528 => x"04",
           529 => x"0c",
           530 => x"2d",
           531 => x"08",
           532 => x"04",
           533 => x"0c",
           534 => x"2d",
           535 => x"08",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"04",
           549 => x"0c",
           550 => x"81",
           551 => x"82",
           552 => x"81",
           553 => x"b9",
           554 => x"d3",
           555 => x"a0",
           556 => x"d3",
           557 => x"e1",
           558 => x"90",
           559 => x"90",
           560 => x"90",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"81",
           566 => x"82",
           567 => x"81",
           568 => x"9f",
           569 => x"d3",
           570 => x"a0",
           571 => x"d3",
           572 => x"a2",
           573 => x"d3",
           574 => x"a0",
           575 => x"04",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"53",
           584 => x"00",
           585 => x"06",
           586 => x"09",
           587 => x"05",
           588 => x"2b",
           589 => x"06",
           590 => x"04",
           591 => x"72",
           592 => x"05",
           593 => x"05",
           594 => x"72",
           595 => x"53",
           596 => x"51",
           597 => x"04",
           598 => x"70",
           599 => x"27",
           600 => x"71",
           601 => x"53",
           602 => x"0b",
           603 => x"8c",
           604 => x"bb",
           605 => x"81",
           606 => x"02",
           607 => x"0c",
           608 => x"80",
           609 => x"90",
           610 => x"08",
           611 => x"90",
           612 => x"08",
           613 => x"3f",
           614 => x"08",
           615 => x"84",
           616 => x"3d",
           617 => x"90",
           618 => x"d3",
           619 => x"81",
           620 => x"fd",
           621 => x"53",
           622 => x"08",
           623 => x"52",
           624 => x"08",
           625 => x"51",
           626 => x"81",
           627 => x"70",
           628 => x"0c",
           629 => x"0d",
           630 => x"0c",
           631 => x"90",
           632 => x"d3",
           633 => x"3d",
           634 => x"81",
           635 => x"fc",
           636 => x"d3",
           637 => x"05",
           638 => x"b9",
           639 => x"90",
           640 => x"08",
           641 => x"90",
           642 => x"0c",
           643 => x"d3",
           644 => x"05",
           645 => x"90",
           646 => x"08",
           647 => x"0b",
           648 => x"08",
           649 => x"81",
           650 => x"f4",
           651 => x"d3",
           652 => x"05",
           653 => x"90",
           654 => x"08",
           655 => x"38",
           656 => x"08",
           657 => x"30",
           658 => x"08",
           659 => x"80",
           660 => x"90",
           661 => x"0c",
           662 => x"08",
           663 => x"8a",
           664 => x"81",
           665 => x"f0",
           666 => x"d3",
           667 => x"05",
           668 => x"90",
           669 => x"0c",
           670 => x"d3",
           671 => x"05",
           672 => x"d3",
           673 => x"05",
           674 => x"df",
           675 => x"84",
           676 => x"d3",
           677 => x"05",
           678 => x"d3",
           679 => x"05",
           680 => x"90",
           681 => x"90",
           682 => x"08",
           683 => x"90",
           684 => x"0c",
           685 => x"08",
           686 => x"70",
           687 => x"0c",
           688 => x"0d",
           689 => x"0c",
           690 => x"90",
           691 => x"d3",
           692 => x"3d",
           693 => x"81",
           694 => x"fc",
           695 => x"d3",
           696 => x"05",
           697 => x"99",
           698 => x"90",
           699 => x"08",
           700 => x"90",
           701 => x"0c",
           702 => x"d3",
           703 => x"05",
           704 => x"90",
           705 => x"08",
           706 => x"38",
           707 => x"08",
           708 => x"30",
           709 => x"08",
           710 => x"81",
           711 => x"90",
           712 => x"08",
           713 => x"90",
           714 => x"08",
           715 => x"81",
           716 => x"70",
           717 => x"08",
           718 => x"54",
           719 => x"08",
           720 => x"80",
           721 => x"81",
           722 => x"f8",
           723 => x"81",
           724 => x"f8",
           725 => x"d3",
           726 => x"05",
           727 => x"d3",
           728 => x"87",
           729 => x"d3",
           730 => x"81",
           731 => x"02",
           732 => x"0c",
           733 => x"81",
           734 => x"90",
           735 => x"0c",
           736 => x"d3",
           737 => x"05",
           738 => x"90",
           739 => x"08",
           740 => x"08",
           741 => x"27",
           742 => x"d3",
           743 => x"05",
           744 => x"ae",
           745 => x"81",
           746 => x"8c",
           747 => x"a2",
           748 => x"90",
           749 => x"08",
           750 => x"90",
           751 => x"0c",
           752 => x"08",
           753 => x"10",
           754 => x"08",
           755 => x"ff",
           756 => x"d3",
           757 => x"05",
           758 => x"80",
           759 => x"d3",
           760 => x"05",
           761 => x"90",
           762 => x"08",
           763 => x"81",
           764 => x"88",
           765 => x"d3",
           766 => x"05",
           767 => x"d3",
           768 => x"05",
           769 => x"90",
           770 => x"08",
           771 => x"08",
           772 => x"07",
           773 => x"08",
           774 => x"81",
           775 => x"fc",
           776 => x"2a",
           777 => x"08",
           778 => x"81",
           779 => x"8c",
           780 => x"2a",
           781 => x"08",
           782 => x"ff",
           783 => x"d3",
           784 => x"05",
           785 => x"93",
           786 => x"90",
           787 => x"08",
           788 => x"90",
           789 => x"0c",
           790 => x"81",
           791 => x"f8",
           792 => x"81",
           793 => x"f4",
           794 => x"81",
           795 => x"f4",
           796 => x"d3",
           797 => x"3d",
           798 => x"90",
           799 => x"3d",
           800 => x"71",
           801 => x"9f",
           802 => x"55",
           803 => x"72",
           804 => x"74",
           805 => x"70",
           806 => x"38",
           807 => x"71",
           808 => x"38",
           809 => x"81",
           810 => x"ff",
           811 => x"ff",
           812 => x"06",
           813 => x"81",
           814 => x"86",
           815 => x"74",
           816 => x"75",
           817 => x"90",
           818 => x"54",
           819 => x"27",
           820 => x"71",
           821 => x"53",
           822 => x"70",
           823 => x"0c",
           824 => x"84",
           825 => x"72",
           826 => x"05",
           827 => x"12",
           828 => x"26",
           829 => x"72",
           830 => x"72",
           831 => x"05",
           832 => x"12",
           833 => x"26",
           834 => x"53",
           835 => x"fb",
           836 => x"79",
           837 => x"83",
           838 => x"52",
           839 => x"71",
           840 => x"54",
           841 => x"73",
           842 => x"c6",
           843 => x"54",
           844 => x"70",
           845 => x"52",
           846 => x"2e",
           847 => x"33",
           848 => x"2e",
           849 => x"95",
           850 => x"81",
           851 => x"70",
           852 => x"54",
           853 => x"70",
           854 => x"33",
           855 => x"ff",
           856 => x"ff",
           857 => x"31",
           858 => x"0c",
           859 => x"3d",
           860 => x"09",
           861 => x"fd",
           862 => x"70",
           863 => x"81",
           864 => x"51",
           865 => x"38",
           866 => x"16",
           867 => x"56",
           868 => x"08",
           869 => x"73",
           870 => x"ff",
           871 => x"0b",
           872 => x"0c",
           873 => x"04",
           874 => x"80",
           875 => x"71",
           876 => x"87",
           877 => x"d3",
           878 => x"ff",
           879 => x"ff",
           880 => x"72",
           881 => x"38",
           882 => x"84",
           883 => x"0d",
           884 => x"0d",
           885 => x"70",
           886 => x"71",
           887 => x"ca",
           888 => x"51",
           889 => x"09",
           890 => x"38",
           891 => x"f1",
           892 => x"84",
           893 => x"53",
           894 => x"70",
           895 => x"53",
           896 => x"a0",
           897 => x"81",
           898 => x"2e",
           899 => x"e5",
           900 => x"ff",
           901 => x"a0",
           902 => x"06",
           903 => x"73",
           904 => x"55",
           905 => x"0c",
           906 => x"81",
           907 => x"87",
           908 => x"fc",
           909 => x"53",
           910 => x"2e",
           911 => x"3d",
           912 => x"72",
           913 => x"3f",
           914 => x"08",
           915 => x"53",
           916 => x"53",
           917 => x"84",
           918 => x"0d",
           919 => x"0d",
           920 => x"33",
           921 => x"53",
           922 => x"8b",
           923 => x"38",
           924 => x"ff",
           925 => x"52",
           926 => x"81",
           927 => x"13",
           928 => x"52",
           929 => x"80",
           930 => x"13",
           931 => x"52",
           932 => x"80",
           933 => x"13",
           934 => x"52",
           935 => x"80",
           936 => x"13",
           937 => x"52",
           938 => x"26",
           939 => x"8a",
           940 => x"87",
           941 => x"e7",
           942 => x"38",
           943 => x"c0",
           944 => x"72",
           945 => x"98",
           946 => x"13",
           947 => x"98",
           948 => x"13",
           949 => x"98",
           950 => x"13",
           951 => x"98",
           952 => x"13",
           953 => x"98",
           954 => x"13",
           955 => x"98",
           956 => x"87",
           957 => x"0c",
           958 => x"98",
           959 => x"0b",
           960 => x"9c",
           961 => x"71",
           962 => x"0c",
           963 => x"04",
           964 => x"7f",
           965 => x"98",
           966 => x"7d",
           967 => x"98",
           968 => x"7d",
           969 => x"c0",
           970 => x"5a",
           971 => x"34",
           972 => x"b4",
           973 => x"83",
           974 => x"c0",
           975 => x"5a",
           976 => x"34",
           977 => x"ac",
           978 => x"85",
           979 => x"c0",
           980 => x"5a",
           981 => x"34",
           982 => x"a4",
           983 => x"88",
           984 => x"c0",
           985 => x"5a",
           986 => x"23",
           987 => x"79",
           988 => x"06",
           989 => x"ff",
           990 => x"86",
           991 => x"85",
           992 => x"84",
           993 => x"83",
           994 => x"82",
           995 => x"7d",
           996 => x"06",
           997 => x"d0",
           998 => x"3f",
           999 => x"04",
          1000 => x"02",
          1001 => x"70",
          1002 => x"2a",
          1003 => x"70",
          1004 => x"cf",
          1005 => x"3d",
          1006 => x"3d",
          1007 => x"0b",
          1008 => x"33",
          1009 => x"06",
          1010 => x"87",
          1011 => x"51",
          1012 => x"86",
          1013 => x"94",
          1014 => x"08",
          1015 => x"70",
          1016 => x"54",
          1017 => x"2e",
          1018 => x"91",
          1019 => x"06",
          1020 => x"d7",
          1021 => x"32",
          1022 => x"51",
          1023 => x"2e",
          1024 => x"93",
          1025 => x"06",
          1026 => x"ff",
          1027 => x"81",
          1028 => x"87",
          1029 => x"52",
          1030 => x"86",
          1031 => x"94",
          1032 => x"72",
          1033 => x"d3",
          1034 => x"3d",
          1035 => x"3d",
          1036 => x"05",
          1037 => x"81",
          1038 => x"70",
          1039 => x"57",
          1040 => x"c0",
          1041 => x"74",
          1042 => x"38",
          1043 => x"94",
          1044 => x"70",
          1045 => x"81",
          1046 => x"52",
          1047 => x"8c",
          1048 => x"2a",
          1049 => x"51",
          1050 => x"38",
          1051 => x"70",
          1052 => x"51",
          1053 => x"8d",
          1054 => x"2a",
          1055 => x"51",
          1056 => x"be",
          1057 => x"ff",
          1058 => x"c0",
          1059 => x"70",
          1060 => x"38",
          1061 => x"90",
          1062 => x"0c",
          1063 => x"04",
          1064 => x"79",
          1065 => x"33",
          1066 => x"06",
          1067 => x"70",
          1068 => x"fe",
          1069 => x"ff",
          1070 => x"0b",
          1071 => x"fc",
          1072 => x"ff",
          1073 => x"55",
          1074 => x"94",
          1075 => x"80",
          1076 => x"87",
          1077 => x"51",
          1078 => x"96",
          1079 => x"06",
          1080 => x"70",
          1081 => x"38",
          1082 => x"70",
          1083 => x"51",
          1084 => x"72",
          1085 => x"81",
          1086 => x"70",
          1087 => x"38",
          1088 => x"70",
          1089 => x"51",
          1090 => x"38",
          1091 => x"06",
          1092 => x"94",
          1093 => x"80",
          1094 => x"87",
          1095 => x"52",
          1096 => x"81",
          1097 => x"70",
          1098 => x"53",
          1099 => x"ff",
          1100 => x"81",
          1101 => x"89",
          1102 => x"fe",
          1103 => x"0b",
          1104 => x"33",
          1105 => x"06",
          1106 => x"c0",
          1107 => x"72",
          1108 => x"38",
          1109 => x"94",
          1110 => x"70",
          1111 => x"81",
          1112 => x"51",
          1113 => x"e2",
          1114 => x"ff",
          1115 => x"c0",
          1116 => x"70",
          1117 => x"38",
          1118 => x"90",
          1119 => x"70",
          1120 => x"81",
          1121 => x"51",
          1122 => x"04",
          1123 => x"0b",
          1124 => x"fc",
          1125 => x"ff",
          1126 => x"87",
          1127 => x"52",
          1128 => x"86",
          1129 => x"94",
          1130 => x"08",
          1131 => x"70",
          1132 => x"51",
          1133 => x"70",
          1134 => x"38",
          1135 => x"06",
          1136 => x"94",
          1137 => x"80",
          1138 => x"87",
          1139 => x"52",
          1140 => x"98",
          1141 => x"2c",
          1142 => x"71",
          1143 => x"0c",
          1144 => x"04",
          1145 => x"87",
          1146 => x"08",
          1147 => x"8a",
          1148 => x"70",
          1149 => x"93",
          1150 => x"9e",
          1151 => x"d0",
          1152 => x"c0",
          1153 => x"81",
          1154 => x"87",
          1155 => x"08",
          1156 => x"0c",
          1157 => x"90",
          1158 => x"8c",
          1159 => x"9e",
          1160 => x"d0",
          1161 => x"c0",
          1162 => x"81",
          1163 => x"87",
          1164 => x"08",
          1165 => x"0c",
          1166 => x"a8",
          1167 => x"9c",
          1168 => x"9e",
          1169 => x"d0",
          1170 => x"c0",
          1171 => x"51",
          1172 => x"a4",
          1173 => x"9e",
          1174 => x"d0",
          1175 => x"0b",
          1176 => x"34",
          1177 => x"c0",
          1178 => x"70",
          1179 => x"51",
          1180 => x"80",
          1181 => x"81",
          1182 => x"d0",
          1183 => x"0b",
          1184 => x"88",
          1185 => x"80",
          1186 => x"52",
          1187 => x"2e",
          1188 => x"52",
          1189 => x"ae",
          1190 => x"87",
          1191 => x"08",
          1192 => x"80",
          1193 => x"52",
          1194 => x"83",
          1195 => x"71",
          1196 => x"34",
          1197 => x"c0",
          1198 => x"70",
          1199 => x"51",
          1200 => x"80",
          1201 => x"81",
          1202 => x"d0",
          1203 => x"0b",
          1204 => x"88",
          1205 => x"80",
          1206 => x"52",
          1207 => x"83",
          1208 => x"71",
          1209 => x"34",
          1210 => x"c0",
          1211 => x"70",
          1212 => x"51",
          1213 => x"80",
          1214 => x"81",
          1215 => x"d0",
          1216 => x"0b",
          1217 => x"88",
          1218 => x"80",
          1219 => x"52",
          1220 => x"83",
          1221 => x"71",
          1222 => x"34",
          1223 => x"c0",
          1224 => x"70",
          1225 => x"51",
          1226 => x"80",
          1227 => x"81",
          1228 => x"d0",
          1229 => x"c0",
          1230 => x"70",
          1231 => x"70",
          1232 => x"51",
          1233 => x"d0",
          1234 => x"0b",
          1235 => x"88",
          1236 => x"06",
          1237 => x"70",
          1238 => x"38",
          1239 => x"81",
          1240 => x"80",
          1241 => x"9e",
          1242 => x"88",
          1243 => x"52",
          1244 => x"83",
          1245 => x"71",
          1246 => x"34",
          1247 => x"88",
          1248 => x"06",
          1249 => x"81",
          1250 => x"83",
          1251 => x"fd",
          1252 => x"bd",
          1253 => x"a1",
          1254 => x"ac",
          1255 => x"80",
          1256 => x"81",
          1257 => x"84",
          1258 => x"be",
          1259 => x"89",
          1260 => x"ad",
          1261 => x"80",
          1262 => x"81",
          1263 => x"53",
          1264 => x"08",
          1265 => x"a8",
          1266 => x"3f",
          1267 => x"33",
          1268 => x"2e",
          1269 => x"d0",
          1270 => x"81",
          1271 => x"52",
          1272 => x"51",
          1273 => x"81",
          1274 => x"54",
          1275 => x"81",
          1276 => x"54",
          1277 => x"92",
          1278 => x"94",
          1279 => x"d0",
          1280 => x"81",
          1281 => x"89",
          1282 => x"d0",
          1283 => x"73",
          1284 => x"38",
          1285 => x"51",
          1286 => x"81",
          1287 => x"54",
          1288 => x"88",
          1289 => x"a4",
          1290 => x"3f",
          1291 => x"33",
          1292 => x"2e",
          1293 => x"bf",
          1294 => x"fd",
          1295 => x"b4",
          1296 => x"80",
          1297 => x"81",
          1298 => x"52",
          1299 => x"51",
          1300 => x"81",
          1301 => x"54",
          1302 => x"88",
          1303 => x"dc",
          1304 => x"3f",
          1305 => x"33",
          1306 => x"2e",
          1307 => x"d0",
          1308 => x"81",
          1309 => x"88",
          1310 => x"c0",
          1311 => x"b9",
          1312 => x"98",
          1313 => x"c0",
          1314 => x"91",
          1315 => x"9c",
          1316 => x"c0",
          1317 => x"85",
          1318 => x"a0",
          1319 => x"c0",
          1320 => x"f9",
          1321 => x"a4",
          1322 => x"c1",
          1323 => x"ed",
          1324 => x"a8",
          1325 => x"c1",
          1326 => x"e1",
          1327 => x"0d",
          1328 => x"0d",
          1329 => x"33",
          1330 => x"71",
          1331 => x"38",
          1332 => x"81",
          1333 => x"52",
          1334 => x"81",
          1335 => x"9d",
          1336 => x"f0",
          1337 => x"81",
          1338 => x"91",
          1339 => x"80",
          1340 => x"81",
          1341 => x"85",
          1342 => x"8c",
          1343 => x"3f",
          1344 => x"04",
          1345 => x"0c",
          1346 => x"87",
          1347 => x"0c",
          1348 => x"0d",
          1349 => x"84",
          1350 => x"52",
          1351 => x"70",
          1352 => x"81",
          1353 => x"72",
          1354 => x"0d",
          1355 => x"0d",
          1356 => x"84",
          1357 => x"d0",
          1358 => x"80",
          1359 => x"09",
          1360 => x"bc",
          1361 => x"81",
          1362 => x"73",
          1363 => x"3d",
          1364 => x"d0",
          1365 => x"c0",
          1366 => x"04",
          1367 => x"02",
          1368 => x"53",
          1369 => x"09",
          1370 => x"38",
          1371 => x"3f",
          1372 => x"08",
          1373 => x"2e",
          1374 => x"72",
          1375 => x"9c",
          1376 => x"81",
          1377 => x"8f",
          1378 => x"94",
          1379 => x"80",
          1380 => x"72",
          1381 => x"84",
          1382 => x"fe",
          1383 => x"97",
          1384 => x"d3",
          1385 => x"81",
          1386 => x"54",
          1387 => x"3f",
          1388 => x"94",
          1389 => x"0d",
          1390 => x"0d",
          1391 => x"33",
          1392 => x"06",
          1393 => x"80",
          1394 => x"72",
          1395 => x"51",
          1396 => x"ff",
          1397 => x"39",
          1398 => x"04",
          1399 => x"77",
          1400 => x"08",
          1401 => x"94",
          1402 => x"73",
          1403 => x"ff",
          1404 => x"71",
          1405 => x"38",
          1406 => x"06",
          1407 => x"54",
          1408 => x"e7",
          1409 => x"d3",
          1410 => x"3d",
          1411 => x"3d",
          1412 => x"59",
          1413 => x"81",
          1414 => x"56",
          1415 => x"84",
          1416 => x"a5",
          1417 => x"06",
          1418 => x"80",
          1419 => x"81",
          1420 => x"58",
          1421 => x"b0",
          1422 => x"06",
          1423 => x"5a",
          1424 => x"ad",
          1425 => x"06",
          1426 => x"5a",
          1427 => x"05",
          1428 => x"75",
          1429 => x"81",
          1430 => x"77",
          1431 => x"08",
          1432 => x"05",
          1433 => x"5d",
          1434 => x"39",
          1435 => x"72",
          1436 => x"38",
          1437 => x"7b",
          1438 => x"05",
          1439 => x"70",
          1440 => x"33",
          1441 => x"39",
          1442 => x"32",
          1443 => x"72",
          1444 => x"78",
          1445 => x"70",
          1446 => x"07",
          1447 => x"07",
          1448 => x"51",
          1449 => x"80",
          1450 => x"79",
          1451 => x"70",
          1452 => x"33",
          1453 => x"80",
          1454 => x"38",
          1455 => x"e0",
          1456 => x"38",
          1457 => x"81",
          1458 => x"53",
          1459 => x"2e",
          1460 => x"73",
          1461 => x"a2",
          1462 => x"c3",
          1463 => x"38",
          1464 => x"24",
          1465 => x"80",
          1466 => x"8c",
          1467 => x"39",
          1468 => x"2e",
          1469 => x"81",
          1470 => x"80",
          1471 => x"80",
          1472 => x"d5",
          1473 => x"73",
          1474 => x"8e",
          1475 => x"39",
          1476 => x"2e",
          1477 => x"80",
          1478 => x"84",
          1479 => x"56",
          1480 => x"74",
          1481 => x"72",
          1482 => x"38",
          1483 => x"15",
          1484 => x"54",
          1485 => x"38",
          1486 => x"56",
          1487 => x"81",
          1488 => x"72",
          1489 => x"38",
          1490 => x"90",
          1491 => x"06",
          1492 => x"2e",
          1493 => x"51",
          1494 => x"74",
          1495 => x"53",
          1496 => x"fd",
          1497 => x"51",
          1498 => x"ef",
          1499 => x"19",
          1500 => x"53",
          1501 => x"39",
          1502 => x"39",
          1503 => x"39",
          1504 => x"39",
          1505 => x"39",
          1506 => x"d0",
          1507 => x"39",
          1508 => x"70",
          1509 => x"53",
          1510 => x"88",
          1511 => x"19",
          1512 => x"39",
          1513 => x"54",
          1514 => x"74",
          1515 => x"70",
          1516 => x"07",
          1517 => x"55",
          1518 => x"80",
          1519 => x"72",
          1520 => x"38",
          1521 => x"90",
          1522 => x"80",
          1523 => x"5e",
          1524 => x"74",
          1525 => x"3f",
          1526 => x"08",
          1527 => x"7c",
          1528 => x"54",
          1529 => x"81",
          1530 => x"55",
          1531 => x"92",
          1532 => x"53",
          1533 => x"2e",
          1534 => x"14",
          1535 => x"ff",
          1536 => x"14",
          1537 => x"70",
          1538 => x"34",
          1539 => x"30",
          1540 => x"9f",
          1541 => x"57",
          1542 => x"85",
          1543 => x"b1",
          1544 => x"2a",
          1545 => x"51",
          1546 => x"2e",
          1547 => x"3d",
          1548 => x"05",
          1549 => x"34",
          1550 => x"76",
          1551 => x"54",
          1552 => x"72",
          1553 => x"54",
          1554 => x"70",
          1555 => x"56",
          1556 => x"81",
          1557 => x"7b",
          1558 => x"73",
          1559 => x"3f",
          1560 => x"53",
          1561 => x"74",
          1562 => x"53",
          1563 => x"eb",
          1564 => x"77",
          1565 => x"53",
          1566 => x"14",
          1567 => x"54",
          1568 => x"3f",
          1569 => x"74",
          1570 => x"53",
          1571 => x"fb",
          1572 => x"51",
          1573 => x"ef",
          1574 => x"0d",
          1575 => x"0d",
          1576 => x"70",
          1577 => x"08",
          1578 => x"51",
          1579 => x"85",
          1580 => x"fe",
          1581 => x"81",
          1582 => x"85",
          1583 => x"52",
          1584 => x"ca",
          1585 => x"9c",
          1586 => x"73",
          1587 => x"81",
          1588 => x"84",
          1589 => x"fd",
          1590 => x"d3",
          1591 => x"81",
          1592 => x"87",
          1593 => x"53",
          1594 => x"fa",
          1595 => x"81",
          1596 => x"85",
          1597 => x"fb",
          1598 => x"79",
          1599 => x"08",
          1600 => x"57",
          1601 => x"71",
          1602 => x"e0",
          1603 => x"98",
          1604 => x"2d",
          1605 => x"08",
          1606 => x"53",
          1607 => x"80",
          1608 => x"8d",
          1609 => x"72",
          1610 => x"30",
          1611 => x"51",
          1612 => x"80",
          1613 => x"71",
          1614 => x"38",
          1615 => x"97",
          1616 => x"25",
          1617 => x"16",
          1618 => x"25",
          1619 => x"14",
          1620 => x"34",
          1621 => x"72",
          1622 => x"3f",
          1623 => x"73",
          1624 => x"72",
          1625 => x"f7",
          1626 => x"53",
          1627 => x"84",
          1628 => x"0d",
          1629 => x"0d",
          1630 => x"08",
          1631 => x"98",
          1632 => x"76",
          1633 => x"ef",
          1634 => x"d3",
          1635 => x"3d",
          1636 => x"3d",
          1637 => x"5a",
          1638 => x"7a",
          1639 => x"08",
          1640 => x"53",
          1641 => x"09",
          1642 => x"38",
          1643 => x"0c",
          1644 => x"ad",
          1645 => x"06",
          1646 => x"76",
          1647 => x"0c",
          1648 => x"33",
          1649 => x"73",
          1650 => x"81",
          1651 => x"38",
          1652 => x"05",
          1653 => x"08",
          1654 => x"53",
          1655 => x"2e",
          1656 => x"57",
          1657 => x"2e",
          1658 => x"39",
          1659 => x"13",
          1660 => x"08",
          1661 => x"53",
          1662 => x"55",
          1663 => x"80",
          1664 => x"14",
          1665 => x"88",
          1666 => x"27",
          1667 => x"eb",
          1668 => x"53",
          1669 => x"89",
          1670 => x"38",
          1671 => x"55",
          1672 => x"8a",
          1673 => x"a0",
          1674 => x"c2",
          1675 => x"74",
          1676 => x"e0",
          1677 => x"ff",
          1678 => x"d0",
          1679 => x"ff",
          1680 => x"90",
          1681 => x"38",
          1682 => x"81",
          1683 => x"53",
          1684 => x"ca",
          1685 => x"27",
          1686 => x"77",
          1687 => x"08",
          1688 => x"0c",
          1689 => x"33",
          1690 => x"ff",
          1691 => x"80",
          1692 => x"74",
          1693 => x"79",
          1694 => x"74",
          1695 => x"0c",
          1696 => x"04",
          1697 => x"7a",
          1698 => x"80",
          1699 => x"58",
          1700 => x"33",
          1701 => x"a0",
          1702 => x"06",
          1703 => x"13",
          1704 => x"39",
          1705 => x"09",
          1706 => x"38",
          1707 => x"11",
          1708 => x"08",
          1709 => x"54",
          1710 => x"2e",
          1711 => x"80",
          1712 => x"08",
          1713 => x"0c",
          1714 => x"33",
          1715 => x"80",
          1716 => x"38",
          1717 => x"80",
          1718 => x"38",
          1719 => x"57",
          1720 => x"0c",
          1721 => x"33",
          1722 => x"39",
          1723 => x"74",
          1724 => x"38",
          1725 => x"80",
          1726 => x"89",
          1727 => x"38",
          1728 => x"d0",
          1729 => x"55",
          1730 => x"80",
          1731 => x"39",
          1732 => x"d9",
          1733 => x"80",
          1734 => x"27",
          1735 => x"80",
          1736 => x"89",
          1737 => x"70",
          1738 => x"55",
          1739 => x"70",
          1740 => x"55",
          1741 => x"27",
          1742 => x"14",
          1743 => x"06",
          1744 => x"74",
          1745 => x"73",
          1746 => x"38",
          1747 => x"14",
          1748 => x"05",
          1749 => x"08",
          1750 => x"54",
          1751 => x"39",
          1752 => x"84",
          1753 => x"55",
          1754 => x"81",
          1755 => x"d3",
          1756 => x"3d",
          1757 => x"3d",
          1758 => x"05",
          1759 => x"52",
          1760 => x"87",
          1761 => x"c0",
          1762 => x"71",
          1763 => x"0c",
          1764 => x"04",
          1765 => x"02",
          1766 => x"02",
          1767 => x"05",
          1768 => x"83",
          1769 => x"26",
          1770 => x"72",
          1771 => x"c0",
          1772 => x"53",
          1773 => x"74",
          1774 => x"38",
          1775 => x"73",
          1776 => x"c0",
          1777 => x"51",
          1778 => x"85",
          1779 => x"98",
          1780 => x"52",
          1781 => x"82",
          1782 => x"70",
          1783 => x"38",
          1784 => x"8c",
          1785 => x"ec",
          1786 => x"fc",
          1787 => x"52",
          1788 => x"87",
          1789 => x"08",
          1790 => x"2e",
          1791 => x"81",
          1792 => x"34",
          1793 => x"13",
          1794 => x"81",
          1795 => x"86",
          1796 => x"f3",
          1797 => x"62",
          1798 => x"05",
          1799 => x"57",
          1800 => x"83",
          1801 => x"fe",
          1802 => x"d3",
          1803 => x"06",
          1804 => x"71",
          1805 => x"71",
          1806 => x"2b",
          1807 => x"80",
          1808 => x"92",
          1809 => x"c0",
          1810 => x"41",
          1811 => x"5a",
          1812 => x"87",
          1813 => x"0c",
          1814 => x"84",
          1815 => x"08",
          1816 => x"70",
          1817 => x"53",
          1818 => x"2e",
          1819 => x"08",
          1820 => x"70",
          1821 => x"34",
          1822 => x"80",
          1823 => x"53",
          1824 => x"2e",
          1825 => x"53",
          1826 => x"26",
          1827 => x"80",
          1828 => x"87",
          1829 => x"08",
          1830 => x"38",
          1831 => x"8c",
          1832 => x"80",
          1833 => x"78",
          1834 => x"99",
          1835 => x"0c",
          1836 => x"8c",
          1837 => x"08",
          1838 => x"51",
          1839 => x"38",
          1840 => x"8d",
          1841 => x"17",
          1842 => x"81",
          1843 => x"53",
          1844 => x"2e",
          1845 => x"fc",
          1846 => x"52",
          1847 => x"7d",
          1848 => x"ed",
          1849 => x"80",
          1850 => x"71",
          1851 => x"38",
          1852 => x"53",
          1853 => x"84",
          1854 => x"0d",
          1855 => x"0d",
          1856 => x"02",
          1857 => x"05",
          1858 => x"58",
          1859 => x"80",
          1860 => x"fc",
          1861 => x"d3",
          1862 => x"06",
          1863 => x"71",
          1864 => x"81",
          1865 => x"38",
          1866 => x"2b",
          1867 => x"80",
          1868 => x"92",
          1869 => x"c0",
          1870 => x"40",
          1871 => x"5a",
          1872 => x"c0",
          1873 => x"76",
          1874 => x"76",
          1875 => x"75",
          1876 => x"2a",
          1877 => x"51",
          1878 => x"80",
          1879 => x"7a",
          1880 => x"5c",
          1881 => x"81",
          1882 => x"81",
          1883 => x"06",
          1884 => x"80",
          1885 => x"87",
          1886 => x"08",
          1887 => x"38",
          1888 => x"8c",
          1889 => x"80",
          1890 => x"77",
          1891 => x"99",
          1892 => x"0c",
          1893 => x"8c",
          1894 => x"08",
          1895 => x"51",
          1896 => x"38",
          1897 => x"8d",
          1898 => x"70",
          1899 => x"84",
          1900 => x"5b",
          1901 => x"2e",
          1902 => x"fc",
          1903 => x"52",
          1904 => x"7d",
          1905 => x"f8",
          1906 => x"80",
          1907 => x"71",
          1908 => x"38",
          1909 => x"53",
          1910 => x"84",
          1911 => x"0d",
          1912 => x"0d",
          1913 => x"05",
          1914 => x"02",
          1915 => x"05",
          1916 => x"54",
          1917 => x"fe",
          1918 => x"84",
          1919 => x"53",
          1920 => x"80",
          1921 => x"0b",
          1922 => x"8c",
          1923 => x"71",
          1924 => x"dc",
          1925 => x"24",
          1926 => x"84",
          1927 => x"92",
          1928 => x"54",
          1929 => x"8d",
          1930 => x"39",
          1931 => x"80",
          1932 => x"cb",
          1933 => x"70",
          1934 => x"81",
          1935 => x"52",
          1936 => x"8a",
          1937 => x"98",
          1938 => x"71",
          1939 => x"c0",
          1940 => x"52",
          1941 => x"81",
          1942 => x"c0",
          1943 => x"53",
          1944 => x"82",
          1945 => x"71",
          1946 => x"39",
          1947 => x"39",
          1948 => x"77",
          1949 => x"81",
          1950 => x"72",
          1951 => x"84",
          1952 => x"73",
          1953 => x"0c",
          1954 => x"04",
          1955 => x"74",
          1956 => x"71",
          1957 => x"2b",
          1958 => x"84",
          1959 => x"84",
          1960 => x"fd",
          1961 => x"83",
          1962 => x"12",
          1963 => x"2b",
          1964 => x"07",
          1965 => x"70",
          1966 => x"2b",
          1967 => x"07",
          1968 => x"0c",
          1969 => x"56",
          1970 => x"3d",
          1971 => x"3d",
          1972 => x"84",
          1973 => x"22",
          1974 => x"72",
          1975 => x"54",
          1976 => x"2a",
          1977 => x"34",
          1978 => x"04",
          1979 => x"73",
          1980 => x"70",
          1981 => x"05",
          1982 => x"88",
          1983 => x"72",
          1984 => x"54",
          1985 => x"2a",
          1986 => x"70",
          1987 => x"34",
          1988 => x"51",
          1989 => x"83",
          1990 => x"fe",
          1991 => x"75",
          1992 => x"51",
          1993 => x"92",
          1994 => x"81",
          1995 => x"73",
          1996 => x"55",
          1997 => x"51",
          1998 => x"3d",
          1999 => x"3d",
          2000 => x"76",
          2001 => x"72",
          2002 => x"05",
          2003 => x"11",
          2004 => x"38",
          2005 => x"04",
          2006 => x"78",
          2007 => x"56",
          2008 => x"81",
          2009 => x"74",
          2010 => x"56",
          2011 => x"31",
          2012 => x"52",
          2013 => x"80",
          2014 => x"71",
          2015 => x"38",
          2016 => x"84",
          2017 => x"0d",
          2018 => x"0d",
          2019 => x"51",
          2020 => x"73",
          2021 => x"81",
          2022 => x"33",
          2023 => x"38",
          2024 => x"d3",
          2025 => x"3d",
          2026 => x"0b",
          2027 => x"0c",
          2028 => x"81",
          2029 => x"04",
          2030 => x"7b",
          2031 => x"83",
          2032 => x"5a",
          2033 => x"80",
          2034 => x"54",
          2035 => x"53",
          2036 => x"53",
          2037 => x"52",
          2038 => x"3f",
          2039 => x"08",
          2040 => x"81",
          2041 => x"81",
          2042 => x"83",
          2043 => x"16",
          2044 => x"18",
          2045 => x"18",
          2046 => x"58",
          2047 => x"9f",
          2048 => x"33",
          2049 => x"2e",
          2050 => x"93",
          2051 => x"76",
          2052 => x"52",
          2053 => x"51",
          2054 => x"83",
          2055 => x"79",
          2056 => x"0c",
          2057 => x"04",
          2058 => x"78",
          2059 => x"80",
          2060 => x"17",
          2061 => x"38",
          2062 => x"fc",
          2063 => x"84",
          2064 => x"d3",
          2065 => x"38",
          2066 => x"53",
          2067 => x"81",
          2068 => x"f7",
          2069 => x"d3",
          2070 => x"2e",
          2071 => x"55",
          2072 => x"b0",
          2073 => x"81",
          2074 => x"88",
          2075 => x"f8",
          2076 => x"70",
          2077 => x"c0",
          2078 => x"84",
          2079 => x"d3",
          2080 => x"91",
          2081 => x"55",
          2082 => x"09",
          2083 => x"f0",
          2084 => x"33",
          2085 => x"2e",
          2086 => x"80",
          2087 => x"80",
          2088 => x"84",
          2089 => x"17",
          2090 => x"fd",
          2091 => x"d4",
          2092 => x"b2",
          2093 => x"96",
          2094 => x"85",
          2095 => x"75",
          2096 => x"3f",
          2097 => x"e4",
          2098 => x"98",
          2099 => x"9c",
          2100 => x"08",
          2101 => x"17",
          2102 => x"3f",
          2103 => x"52",
          2104 => x"51",
          2105 => x"a0",
          2106 => x"05",
          2107 => x"0c",
          2108 => x"75",
          2109 => x"33",
          2110 => x"3f",
          2111 => x"34",
          2112 => x"52",
          2113 => x"51",
          2114 => x"81",
          2115 => x"80",
          2116 => x"81",
          2117 => x"d3",
          2118 => x"3d",
          2119 => x"3d",
          2120 => x"1a",
          2121 => x"fe",
          2122 => x"54",
          2123 => x"73",
          2124 => x"8a",
          2125 => x"71",
          2126 => x"08",
          2127 => x"75",
          2128 => x"0c",
          2129 => x"04",
          2130 => x"7a",
          2131 => x"56",
          2132 => x"77",
          2133 => x"38",
          2134 => x"08",
          2135 => x"38",
          2136 => x"54",
          2137 => x"2e",
          2138 => x"72",
          2139 => x"38",
          2140 => x"8d",
          2141 => x"39",
          2142 => x"81",
          2143 => x"b6",
          2144 => x"2a",
          2145 => x"2a",
          2146 => x"05",
          2147 => x"55",
          2148 => x"81",
          2149 => x"81",
          2150 => x"83",
          2151 => x"b4",
          2152 => x"17",
          2153 => x"a4",
          2154 => x"55",
          2155 => x"57",
          2156 => x"3f",
          2157 => x"08",
          2158 => x"74",
          2159 => x"14",
          2160 => x"70",
          2161 => x"07",
          2162 => x"71",
          2163 => x"52",
          2164 => x"72",
          2165 => x"75",
          2166 => x"58",
          2167 => x"76",
          2168 => x"15",
          2169 => x"73",
          2170 => x"3f",
          2171 => x"08",
          2172 => x"76",
          2173 => x"06",
          2174 => x"05",
          2175 => x"3f",
          2176 => x"08",
          2177 => x"06",
          2178 => x"76",
          2179 => x"15",
          2180 => x"73",
          2181 => x"3f",
          2182 => x"08",
          2183 => x"82",
          2184 => x"06",
          2185 => x"05",
          2186 => x"3f",
          2187 => x"08",
          2188 => x"58",
          2189 => x"58",
          2190 => x"84",
          2191 => x"0d",
          2192 => x"0d",
          2193 => x"5a",
          2194 => x"59",
          2195 => x"82",
          2196 => x"98",
          2197 => x"82",
          2198 => x"33",
          2199 => x"2e",
          2200 => x"72",
          2201 => x"38",
          2202 => x"8d",
          2203 => x"39",
          2204 => x"81",
          2205 => x"f7",
          2206 => x"2a",
          2207 => x"2a",
          2208 => x"05",
          2209 => x"55",
          2210 => x"81",
          2211 => x"59",
          2212 => x"08",
          2213 => x"74",
          2214 => x"16",
          2215 => x"16",
          2216 => x"59",
          2217 => x"53",
          2218 => x"8f",
          2219 => x"2b",
          2220 => x"74",
          2221 => x"71",
          2222 => x"72",
          2223 => x"0b",
          2224 => x"74",
          2225 => x"17",
          2226 => x"75",
          2227 => x"3f",
          2228 => x"08",
          2229 => x"84",
          2230 => x"38",
          2231 => x"06",
          2232 => x"78",
          2233 => x"54",
          2234 => x"77",
          2235 => x"33",
          2236 => x"71",
          2237 => x"51",
          2238 => x"34",
          2239 => x"76",
          2240 => x"17",
          2241 => x"75",
          2242 => x"3f",
          2243 => x"08",
          2244 => x"84",
          2245 => x"38",
          2246 => x"ff",
          2247 => x"10",
          2248 => x"76",
          2249 => x"51",
          2250 => x"be",
          2251 => x"2a",
          2252 => x"05",
          2253 => x"f9",
          2254 => x"d3",
          2255 => x"81",
          2256 => x"ab",
          2257 => x"0a",
          2258 => x"2b",
          2259 => x"70",
          2260 => x"70",
          2261 => x"54",
          2262 => x"81",
          2263 => x"8f",
          2264 => x"07",
          2265 => x"f7",
          2266 => x"0b",
          2267 => x"78",
          2268 => x"0c",
          2269 => x"04",
          2270 => x"7a",
          2271 => x"08",
          2272 => x"59",
          2273 => x"a4",
          2274 => x"17",
          2275 => x"38",
          2276 => x"aa",
          2277 => x"73",
          2278 => x"fd",
          2279 => x"d3",
          2280 => x"81",
          2281 => x"80",
          2282 => x"39",
          2283 => x"eb",
          2284 => x"80",
          2285 => x"d3",
          2286 => x"80",
          2287 => x"52",
          2288 => x"84",
          2289 => x"84",
          2290 => x"d3",
          2291 => x"2e",
          2292 => x"81",
          2293 => x"81",
          2294 => x"81",
          2295 => x"ff",
          2296 => x"80",
          2297 => x"75",
          2298 => x"3f",
          2299 => x"08",
          2300 => x"16",
          2301 => x"90",
          2302 => x"55",
          2303 => x"27",
          2304 => x"15",
          2305 => x"84",
          2306 => x"07",
          2307 => x"17",
          2308 => x"76",
          2309 => x"a6",
          2310 => x"73",
          2311 => x"0c",
          2312 => x"04",
          2313 => x"7c",
          2314 => x"59",
          2315 => x"95",
          2316 => x"08",
          2317 => x"2e",
          2318 => x"17",
          2319 => x"b2",
          2320 => x"ae",
          2321 => x"7a",
          2322 => x"3f",
          2323 => x"81",
          2324 => x"27",
          2325 => x"81",
          2326 => x"55",
          2327 => x"08",
          2328 => x"d2",
          2329 => x"08",
          2330 => x"08",
          2331 => x"38",
          2332 => x"17",
          2333 => x"54",
          2334 => x"82",
          2335 => x"7a",
          2336 => x"06",
          2337 => x"81",
          2338 => x"17",
          2339 => x"83",
          2340 => x"75",
          2341 => x"f9",
          2342 => x"59",
          2343 => x"08",
          2344 => x"81",
          2345 => x"81",
          2346 => x"59",
          2347 => x"08",
          2348 => x"70",
          2349 => x"25",
          2350 => x"81",
          2351 => x"54",
          2352 => x"55",
          2353 => x"38",
          2354 => x"08",
          2355 => x"38",
          2356 => x"54",
          2357 => x"90",
          2358 => x"18",
          2359 => x"38",
          2360 => x"39",
          2361 => x"38",
          2362 => x"16",
          2363 => x"08",
          2364 => x"38",
          2365 => x"78",
          2366 => x"38",
          2367 => x"51",
          2368 => x"81",
          2369 => x"80",
          2370 => x"80",
          2371 => x"84",
          2372 => x"09",
          2373 => x"38",
          2374 => x"08",
          2375 => x"84",
          2376 => x"30",
          2377 => x"80",
          2378 => x"07",
          2379 => x"55",
          2380 => x"38",
          2381 => x"09",
          2382 => x"ae",
          2383 => x"80",
          2384 => x"53",
          2385 => x"51",
          2386 => x"81",
          2387 => x"81",
          2388 => x"30",
          2389 => x"84",
          2390 => x"25",
          2391 => x"79",
          2392 => x"38",
          2393 => x"8f",
          2394 => x"79",
          2395 => x"f9",
          2396 => x"d3",
          2397 => x"74",
          2398 => x"8c",
          2399 => x"17",
          2400 => x"90",
          2401 => x"54",
          2402 => x"86",
          2403 => x"90",
          2404 => x"17",
          2405 => x"54",
          2406 => x"34",
          2407 => x"56",
          2408 => x"90",
          2409 => x"80",
          2410 => x"81",
          2411 => x"55",
          2412 => x"56",
          2413 => x"81",
          2414 => x"8c",
          2415 => x"f8",
          2416 => x"70",
          2417 => x"f0",
          2418 => x"84",
          2419 => x"56",
          2420 => x"08",
          2421 => x"7b",
          2422 => x"f6",
          2423 => x"d3",
          2424 => x"d3",
          2425 => x"17",
          2426 => x"80",
          2427 => x"b4",
          2428 => x"57",
          2429 => x"77",
          2430 => x"81",
          2431 => x"15",
          2432 => x"78",
          2433 => x"81",
          2434 => x"53",
          2435 => x"15",
          2436 => x"e9",
          2437 => x"84",
          2438 => x"df",
          2439 => x"22",
          2440 => x"30",
          2441 => x"70",
          2442 => x"51",
          2443 => x"81",
          2444 => x"8a",
          2445 => x"f8",
          2446 => x"7c",
          2447 => x"56",
          2448 => x"80",
          2449 => x"f1",
          2450 => x"06",
          2451 => x"e9",
          2452 => x"18",
          2453 => x"08",
          2454 => x"38",
          2455 => x"82",
          2456 => x"38",
          2457 => x"54",
          2458 => x"74",
          2459 => x"82",
          2460 => x"22",
          2461 => x"79",
          2462 => x"38",
          2463 => x"98",
          2464 => x"cd",
          2465 => x"22",
          2466 => x"54",
          2467 => x"26",
          2468 => x"52",
          2469 => x"b0",
          2470 => x"84",
          2471 => x"d3",
          2472 => x"2e",
          2473 => x"0b",
          2474 => x"08",
          2475 => x"98",
          2476 => x"d3",
          2477 => x"85",
          2478 => x"bd",
          2479 => x"31",
          2480 => x"73",
          2481 => x"f4",
          2482 => x"d3",
          2483 => x"18",
          2484 => x"18",
          2485 => x"08",
          2486 => x"72",
          2487 => x"38",
          2488 => x"58",
          2489 => x"89",
          2490 => x"18",
          2491 => x"ff",
          2492 => x"05",
          2493 => x"80",
          2494 => x"d3",
          2495 => x"3d",
          2496 => x"3d",
          2497 => x"08",
          2498 => x"a0",
          2499 => x"54",
          2500 => x"77",
          2501 => x"80",
          2502 => x"0c",
          2503 => x"53",
          2504 => x"80",
          2505 => x"38",
          2506 => x"06",
          2507 => x"b5",
          2508 => x"98",
          2509 => x"14",
          2510 => x"92",
          2511 => x"2a",
          2512 => x"56",
          2513 => x"26",
          2514 => x"80",
          2515 => x"16",
          2516 => x"77",
          2517 => x"53",
          2518 => x"38",
          2519 => x"51",
          2520 => x"81",
          2521 => x"53",
          2522 => x"0b",
          2523 => x"08",
          2524 => x"38",
          2525 => x"d3",
          2526 => x"2e",
          2527 => x"98",
          2528 => x"d3",
          2529 => x"80",
          2530 => x"8a",
          2531 => x"15",
          2532 => x"80",
          2533 => x"14",
          2534 => x"51",
          2535 => x"81",
          2536 => x"53",
          2537 => x"d3",
          2538 => x"2e",
          2539 => x"82",
          2540 => x"84",
          2541 => x"ba",
          2542 => x"81",
          2543 => x"ff",
          2544 => x"81",
          2545 => x"52",
          2546 => x"f3",
          2547 => x"84",
          2548 => x"72",
          2549 => x"72",
          2550 => x"f2",
          2551 => x"d3",
          2552 => x"15",
          2553 => x"15",
          2554 => x"b4",
          2555 => x"0c",
          2556 => x"81",
          2557 => x"8a",
          2558 => x"f7",
          2559 => x"7d",
          2560 => x"5b",
          2561 => x"76",
          2562 => x"3f",
          2563 => x"08",
          2564 => x"84",
          2565 => x"38",
          2566 => x"08",
          2567 => x"08",
          2568 => x"f0",
          2569 => x"d3",
          2570 => x"81",
          2571 => x"80",
          2572 => x"d3",
          2573 => x"18",
          2574 => x"51",
          2575 => x"81",
          2576 => x"81",
          2577 => x"81",
          2578 => x"84",
          2579 => x"83",
          2580 => x"77",
          2581 => x"72",
          2582 => x"38",
          2583 => x"75",
          2584 => x"81",
          2585 => x"a5",
          2586 => x"84",
          2587 => x"52",
          2588 => x"8e",
          2589 => x"84",
          2590 => x"d3",
          2591 => x"2e",
          2592 => x"73",
          2593 => x"81",
          2594 => x"87",
          2595 => x"d3",
          2596 => x"3d",
          2597 => x"3d",
          2598 => x"11",
          2599 => x"ec",
          2600 => x"84",
          2601 => x"ff",
          2602 => x"33",
          2603 => x"71",
          2604 => x"81",
          2605 => x"94",
          2606 => x"d0",
          2607 => x"84",
          2608 => x"73",
          2609 => x"81",
          2610 => x"85",
          2611 => x"fc",
          2612 => x"79",
          2613 => x"ff",
          2614 => x"12",
          2615 => x"eb",
          2616 => x"70",
          2617 => x"72",
          2618 => x"81",
          2619 => x"73",
          2620 => x"94",
          2621 => x"d6",
          2622 => x"0d",
          2623 => x"0d",
          2624 => x"55",
          2625 => x"5a",
          2626 => x"08",
          2627 => x"8a",
          2628 => x"08",
          2629 => x"ee",
          2630 => x"d3",
          2631 => x"81",
          2632 => x"80",
          2633 => x"15",
          2634 => x"55",
          2635 => x"38",
          2636 => x"e6",
          2637 => x"33",
          2638 => x"70",
          2639 => x"58",
          2640 => x"86",
          2641 => x"d3",
          2642 => x"73",
          2643 => x"83",
          2644 => x"73",
          2645 => x"38",
          2646 => x"06",
          2647 => x"80",
          2648 => x"75",
          2649 => x"38",
          2650 => x"08",
          2651 => x"54",
          2652 => x"2e",
          2653 => x"83",
          2654 => x"73",
          2655 => x"38",
          2656 => x"51",
          2657 => x"81",
          2658 => x"58",
          2659 => x"08",
          2660 => x"15",
          2661 => x"38",
          2662 => x"0b",
          2663 => x"77",
          2664 => x"0c",
          2665 => x"04",
          2666 => x"77",
          2667 => x"54",
          2668 => x"51",
          2669 => x"81",
          2670 => x"55",
          2671 => x"08",
          2672 => x"14",
          2673 => x"51",
          2674 => x"81",
          2675 => x"55",
          2676 => x"08",
          2677 => x"53",
          2678 => x"08",
          2679 => x"08",
          2680 => x"3f",
          2681 => x"14",
          2682 => x"08",
          2683 => x"3f",
          2684 => x"17",
          2685 => x"d3",
          2686 => x"3d",
          2687 => x"3d",
          2688 => x"08",
          2689 => x"54",
          2690 => x"53",
          2691 => x"81",
          2692 => x"8d",
          2693 => x"08",
          2694 => x"34",
          2695 => x"15",
          2696 => x"0d",
          2697 => x"0d",
          2698 => x"57",
          2699 => x"17",
          2700 => x"08",
          2701 => x"82",
          2702 => x"89",
          2703 => x"55",
          2704 => x"14",
          2705 => x"16",
          2706 => x"71",
          2707 => x"38",
          2708 => x"09",
          2709 => x"38",
          2710 => x"73",
          2711 => x"81",
          2712 => x"ae",
          2713 => x"05",
          2714 => x"15",
          2715 => x"70",
          2716 => x"34",
          2717 => x"8a",
          2718 => x"38",
          2719 => x"05",
          2720 => x"81",
          2721 => x"17",
          2722 => x"12",
          2723 => x"34",
          2724 => x"9c",
          2725 => x"e8",
          2726 => x"d3",
          2727 => x"0c",
          2728 => x"e7",
          2729 => x"d3",
          2730 => x"17",
          2731 => x"51",
          2732 => x"81",
          2733 => x"84",
          2734 => x"3d",
          2735 => x"3d",
          2736 => x"08",
          2737 => x"61",
          2738 => x"55",
          2739 => x"2e",
          2740 => x"55",
          2741 => x"2e",
          2742 => x"80",
          2743 => x"94",
          2744 => x"1c",
          2745 => x"81",
          2746 => x"61",
          2747 => x"56",
          2748 => x"2e",
          2749 => x"83",
          2750 => x"73",
          2751 => x"70",
          2752 => x"25",
          2753 => x"51",
          2754 => x"38",
          2755 => x"0c",
          2756 => x"51",
          2757 => x"26",
          2758 => x"80",
          2759 => x"34",
          2760 => x"51",
          2761 => x"81",
          2762 => x"55",
          2763 => x"91",
          2764 => x"1d",
          2765 => x"8b",
          2766 => x"79",
          2767 => x"3f",
          2768 => x"57",
          2769 => x"55",
          2770 => x"2e",
          2771 => x"80",
          2772 => x"18",
          2773 => x"1a",
          2774 => x"70",
          2775 => x"2a",
          2776 => x"07",
          2777 => x"5a",
          2778 => x"8c",
          2779 => x"54",
          2780 => x"81",
          2781 => x"39",
          2782 => x"70",
          2783 => x"2a",
          2784 => x"75",
          2785 => x"8c",
          2786 => x"2e",
          2787 => x"a0",
          2788 => x"38",
          2789 => x"0c",
          2790 => x"76",
          2791 => x"38",
          2792 => x"b8",
          2793 => x"70",
          2794 => x"5a",
          2795 => x"76",
          2796 => x"38",
          2797 => x"70",
          2798 => x"dc",
          2799 => x"72",
          2800 => x"80",
          2801 => x"51",
          2802 => x"73",
          2803 => x"38",
          2804 => x"18",
          2805 => x"1a",
          2806 => x"55",
          2807 => x"2e",
          2808 => x"83",
          2809 => x"73",
          2810 => x"70",
          2811 => x"25",
          2812 => x"51",
          2813 => x"38",
          2814 => x"75",
          2815 => x"81",
          2816 => x"81",
          2817 => x"27",
          2818 => x"73",
          2819 => x"38",
          2820 => x"70",
          2821 => x"32",
          2822 => x"80",
          2823 => x"2a",
          2824 => x"56",
          2825 => x"81",
          2826 => x"57",
          2827 => x"f5",
          2828 => x"2b",
          2829 => x"25",
          2830 => x"80",
          2831 => x"c2",
          2832 => x"57",
          2833 => x"e6",
          2834 => x"d3",
          2835 => x"2e",
          2836 => x"18",
          2837 => x"1a",
          2838 => x"56",
          2839 => x"3f",
          2840 => x"08",
          2841 => x"e8",
          2842 => x"54",
          2843 => x"80",
          2844 => x"17",
          2845 => x"34",
          2846 => x"11",
          2847 => x"74",
          2848 => x"75",
          2849 => x"98",
          2850 => x"3f",
          2851 => x"08",
          2852 => x"9f",
          2853 => x"99",
          2854 => x"e0",
          2855 => x"ff",
          2856 => x"79",
          2857 => x"74",
          2858 => x"57",
          2859 => x"77",
          2860 => x"76",
          2861 => x"38",
          2862 => x"73",
          2863 => x"09",
          2864 => x"38",
          2865 => x"84",
          2866 => x"27",
          2867 => x"39",
          2868 => x"f2",
          2869 => x"80",
          2870 => x"54",
          2871 => x"34",
          2872 => x"58",
          2873 => x"f2",
          2874 => x"d3",
          2875 => x"81",
          2876 => x"80",
          2877 => x"1b",
          2878 => x"51",
          2879 => x"81",
          2880 => x"56",
          2881 => x"08",
          2882 => x"9c",
          2883 => x"33",
          2884 => x"80",
          2885 => x"38",
          2886 => x"bf",
          2887 => x"86",
          2888 => x"15",
          2889 => x"2a",
          2890 => x"51",
          2891 => x"92",
          2892 => x"79",
          2893 => x"e4",
          2894 => x"d3",
          2895 => x"2e",
          2896 => x"52",
          2897 => x"ba",
          2898 => x"39",
          2899 => x"33",
          2900 => x"80",
          2901 => x"74",
          2902 => x"81",
          2903 => x"38",
          2904 => x"70",
          2905 => x"82",
          2906 => x"54",
          2907 => x"96",
          2908 => x"06",
          2909 => x"2e",
          2910 => x"ff",
          2911 => x"1c",
          2912 => x"80",
          2913 => x"81",
          2914 => x"ba",
          2915 => x"b6",
          2916 => x"2a",
          2917 => x"51",
          2918 => x"38",
          2919 => x"70",
          2920 => x"81",
          2921 => x"55",
          2922 => x"e1",
          2923 => x"08",
          2924 => x"1d",
          2925 => x"7c",
          2926 => x"3f",
          2927 => x"08",
          2928 => x"fa",
          2929 => x"81",
          2930 => x"8f",
          2931 => x"f6",
          2932 => x"5b",
          2933 => x"70",
          2934 => x"59",
          2935 => x"73",
          2936 => x"c6",
          2937 => x"81",
          2938 => x"70",
          2939 => x"52",
          2940 => x"8d",
          2941 => x"38",
          2942 => x"09",
          2943 => x"a5",
          2944 => x"d0",
          2945 => x"ff",
          2946 => x"53",
          2947 => x"91",
          2948 => x"73",
          2949 => x"d0",
          2950 => x"71",
          2951 => x"f7",
          2952 => x"81",
          2953 => x"55",
          2954 => x"55",
          2955 => x"81",
          2956 => x"74",
          2957 => x"56",
          2958 => x"12",
          2959 => x"70",
          2960 => x"38",
          2961 => x"81",
          2962 => x"51",
          2963 => x"51",
          2964 => x"89",
          2965 => x"70",
          2966 => x"53",
          2967 => x"70",
          2968 => x"51",
          2969 => x"09",
          2970 => x"38",
          2971 => x"38",
          2972 => x"77",
          2973 => x"70",
          2974 => x"2a",
          2975 => x"07",
          2976 => x"51",
          2977 => x"8f",
          2978 => x"84",
          2979 => x"83",
          2980 => x"94",
          2981 => x"74",
          2982 => x"38",
          2983 => x"0c",
          2984 => x"86",
          2985 => x"b4",
          2986 => x"81",
          2987 => x"8c",
          2988 => x"fa",
          2989 => x"56",
          2990 => x"17",
          2991 => x"b0",
          2992 => x"52",
          2993 => x"e0",
          2994 => x"81",
          2995 => x"81",
          2996 => x"b2",
          2997 => x"b4",
          2998 => x"84",
          2999 => x"ff",
          3000 => x"55",
          3001 => x"d5",
          3002 => x"06",
          3003 => x"80",
          3004 => x"33",
          3005 => x"81",
          3006 => x"81",
          3007 => x"81",
          3008 => x"eb",
          3009 => x"70",
          3010 => x"07",
          3011 => x"73",
          3012 => x"81",
          3013 => x"81",
          3014 => x"83",
          3015 => x"a8",
          3016 => x"16",
          3017 => x"3f",
          3018 => x"08",
          3019 => x"84",
          3020 => x"9d",
          3021 => x"81",
          3022 => x"81",
          3023 => x"e0",
          3024 => x"d3",
          3025 => x"81",
          3026 => x"80",
          3027 => x"82",
          3028 => x"d3",
          3029 => x"3d",
          3030 => x"3d",
          3031 => x"84",
          3032 => x"05",
          3033 => x"80",
          3034 => x"51",
          3035 => x"81",
          3036 => x"58",
          3037 => x"0b",
          3038 => x"08",
          3039 => x"38",
          3040 => x"08",
          3041 => x"d3",
          3042 => x"08",
          3043 => x"56",
          3044 => x"86",
          3045 => x"75",
          3046 => x"fe",
          3047 => x"54",
          3048 => x"2e",
          3049 => x"14",
          3050 => x"ca",
          3051 => x"84",
          3052 => x"06",
          3053 => x"54",
          3054 => x"38",
          3055 => x"86",
          3056 => x"82",
          3057 => x"06",
          3058 => x"56",
          3059 => x"38",
          3060 => x"80",
          3061 => x"81",
          3062 => x"52",
          3063 => x"51",
          3064 => x"81",
          3065 => x"81",
          3066 => x"81",
          3067 => x"83",
          3068 => x"87",
          3069 => x"2e",
          3070 => x"82",
          3071 => x"06",
          3072 => x"56",
          3073 => x"38",
          3074 => x"74",
          3075 => x"a3",
          3076 => x"84",
          3077 => x"06",
          3078 => x"2e",
          3079 => x"80",
          3080 => x"3d",
          3081 => x"83",
          3082 => x"15",
          3083 => x"53",
          3084 => x"8d",
          3085 => x"15",
          3086 => x"3f",
          3087 => x"08",
          3088 => x"70",
          3089 => x"0c",
          3090 => x"16",
          3091 => x"80",
          3092 => x"80",
          3093 => x"54",
          3094 => x"84",
          3095 => x"5b",
          3096 => x"80",
          3097 => x"7a",
          3098 => x"fc",
          3099 => x"d3",
          3100 => x"ff",
          3101 => x"77",
          3102 => x"81",
          3103 => x"76",
          3104 => x"81",
          3105 => x"2e",
          3106 => x"8d",
          3107 => x"26",
          3108 => x"bf",
          3109 => x"f4",
          3110 => x"84",
          3111 => x"ff",
          3112 => x"84",
          3113 => x"81",
          3114 => x"38",
          3115 => x"51",
          3116 => x"81",
          3117 => x"83",
          3118 => x"58",
          3119 => x"80",
          3120 => x"db",
          3121 => x"d3",
          3122 => x"77",
          3123 => x"80",
          3124 => x"82",
          3125 => x"c4",
          3126 => x"11",
          3127 => x"06",
          3128 => x"8d",
          3129 => x"26",
          3130 => x"74",
          3131 => x"78",
          3132 => x"c1",
          3133 => x"59",
          3134 => x"15",
          3135 => x"2e",
          3136 => x"13",
          3137 => x"72",
          3138 => x"38",
          3139 => x"eb",
          3140 => x"14",
          3141 => x"3f",
          3142 => x"08",
          3143 => x"84",
          3144 => x"23",
          3145 => x"57",
          3146 => x"83",
          3147 => x"c7",
          3148 => x"d8",
          3149 => x"84",
          3150 => x"ff",
          3151 => x"8d",
          3152 => x"14",
          3153 => x"3f",
          3154 => x"08",
          3155 => x"14",
          3156 => x"3f",
          3157 => x"08",
          3158 => x"06",
          3159 => x"72",
          3160 => x"97",
          3161 => x"22",
          3162 => x"84",
          3163 => x"5a",
          3164 => x"83",
          3165 => x"14",
          3166 => x"79",
          3167 => x"af",
          3168 => x"d3",
          3169 => x"81",
          3170 => x"80",
          3171 => x"38",
          3172 => x"08",
          3173 => x"ff",
          3174 => x"38",
          3175 => x"83",
          3176 => x"83",
          3177 => x"74",
          3178 => x"85",
          3179 => x"89",
          3180 => x"76",
          3181 => x"c3",
          3182 => x"70",
          3183 => x"7b",
          3184 => x"73",
          3185 => x"17",
          3186 => x"ac",
          3187 => x"55",
          3188 => x"09",
          3189 => x"38",
          3190 => x"51",
          3191 => x"81",
          3192 => x"83",
          3193 => x"53",
          3194 => x"82",
          3195 => x"82",
          3196 => x"e0",
          3197 => x"ab",
          3198 => x"84",
          3199 => x"0c",
          3200 => x"53",
          3201 => x"56",
          3202 => x"81",
          3203 => x"13",
          3204 => x"74",
          3205 => x"82",
          3206 => x"74",
          3207 => x"81",
          3208 => x"06",
          3209 => x"83",
          3210 => x"2a",
          3211 => x"72",
          3212 => x"26",
          3213 => x"ff",
          3214 => x"0c",
          3215 => x"15",
          3216 => x"0b",
          3217 => x"76",
          3218 => x"81",
          3219 => x"38",
          3220 => x"51",
          3221 => x"81",
          3222 => x"83",
          3223 => x"53",
          3224 => x"09",
          3225 => x"f9",
          3226 => x"52",
          3227 => x"b8",
          3228 => x"84",
          3229 => x"38",
          3230 => x"08",
          3231 => x"84",
          3232 => x"d8",
          3233 => x"d3",
          3234 => x"ff",
          3235 => x"72",
          3236 => x"2e",
          3237 => x"80",
          3238 => x"14",
          3239 => x"3f",
          3240 => x"08",
          3241 => x"a4",
          3242 => x"81",
          3243 => x"84",
          3244 => x"d7",
          3245 => x"d3",
          3246 => x"8a",
          3247 => x"2e",
          3248 => x"9d",
          3249 => x"14",
          3250 => x"3f",
          3251 => x"08",
          3252 => x"84",
          3253 => x"d7",
          3254 => x"d3",
          3255 => x"15",
          3256 => x"34",
          3257 => x"22",
          3258 => x"72",
          3259 => x"23",
          3260 => x"23",
          3261 => x"15",
          3262 => x"75",
          3263 => x"0c",
          3264 => x"04",
          3265 => x"77",
          3266 => x"73",
          3267 => x"38",
          3268 => x"72",
          3269 => x"38",
          3270 => x"71",
          3271 => x"38",
          3272 => x"84",
          3273 => x"52",
          3274 => x"09",
          3275 => x"38",
          3276 => x"51",
          3277 => x"81",
          3278 => x"81",
          3279 => x"88",
          3280 => x"08",
          3281 => x"39",
          3282 => x"73",
          3283 => x"74",
          3284 => x"0c",
          3285 => x"04",
          3286 => x"02",
          3287 => x"7a",
          3288 => x"fc",
          3289 => x"f4",
          3290 => x"54",
          3291 => x"d3",
          3292 => x"bc",
          3293 => x"84",
          3294 => x"81",
          3295 => x"70",
          3296 => x"73",
          3297 => x"38",
          3298 => x"78",
          3299 => x"2e",
          3300 => x"74",
          3301 => x"0c",
          3302 => x"80",
          3303 => x"80",
          3304 => x"70",
          3305 => x"51",
          3306 => x"81",
          3307 => x"54",
          3308 => x"84",
          3309 => x"0d",
          3310 => x"0d",
          3311 => x"05",
          3312 => x"33",
          3313 => x"54",
          3314 => x"84",
          3315 => x"bf",
          3316 => x"98",
          3317 => x"53",
          3318 => x"05",
          3319 => x"fa",
          3320 => x"84",
          3321 => x"d3",
          3322 => x"a4",
          3323 => x"68",
          3324 => x"70",
          3325 => x"c6",
          3326 => x"84",
          3327 => x"d3",
          3328 => x"38",
          3329 => x"05",
          3330 => x"2b",
          3331 => x"80",
          3332 => x"86",
          3333 => x"06",
          3334 => x"2e",
          3335 => x"74",
          3336 => x"38",
          3337 => x"09",
          3338 => x"38",
          3339 => x"f8",
          3340 => x"84",
          3341 => x"39",
          3342 => x"33",
          3343 => x"73",
          3344 => x"77",
          3345 => x"81",
          3346 => x"73",
          3347 => x"38",
          3348 => x"bc",
          3349 => x"07",
          3350 => x"b4",
          3351 => x"2a",
          3352 => x"51",
          3353 => x"2e",
          3354 => x"62",
          3355 => x"e8",
          3356 => x"d3",
          3357 => x"82",
          3358 => x"52",
          3359 => x"51",
          3360 => x"62",
          3361 => x"8b",
          3362 => x"53",
          3363 => x"51",
          3364 => x"80",
          3365 => x"05",
          3366 => x"3f",
          3367 => x"0b",
          3368 => x"75",
          3369 => x"f1",
          3370 => x"11",
          3371 => x"80",
          3372 => x"97",
          3373 => x"51",
          3374 => x"81",
          3375 => x"55",
          3376 => x"08",
          3377 => x"b7",
          3378 => x"c4",
          3379 => x"05",
          3380 => x"2a",
          3381 => x"51",
          3382 => x"80",
          3383 => x"84",
          3384 => x"39",
          3385 => x"70",
          3386 => x"54",
          3387 => x"a9",
          3388 => x"06",
          3389 => x"2e",
          3390 => x"55",
          3391 => x"73",
          3392 => x"d6",
          3393 => x"d3",
          3394 => x"ff",
          3395 => x"0c",
          3396 => x"d3",
          3397 => x"f8",
          3398 => x"2a",
          3399 => x"51",
          3400 => x"2e",
          3401 => x"80",
          3402 => x"7a",
          3403 => x"a0",
          3404 => x"a4",
          3405 => x"53",
          3406 => x"e6",
          3407 => x"d3",
          3408 => x"d3",
          3409 => x"1b",
          3410 => x"05",
          3411 => x"d3",
          3412 => x"84",
          3413 => x"84",
          3414 => x"0c",
          3415 => x"56",
          3416 => x"84",
          3417 => x"90",
          3418 => x"0b",
          3419 => x"80",
          3420 => x"0c",
          3421 => x"1a",
          3422 => x"2a",
          3423 => x"51",
          3424 => x"2e",
          3425 => x"81",
          3426 => x"80",
          3427 => x"38",
          3428 => x"08",
          3429 => x"8a",
          3430 => x"89",
          3431 => x"59",
          3432 => x"76",
          3433 => x"d7",
          3434 => x"d3",
          3435 => x"81",
          3436 => x"81",
          3437 => x"82",
          3438 => x"84",
          3439 => x"09",
          3440 => x"38",
          3441 => x"78",
          3442 => x"30",
          3443 => x"80",
          3444 => x"77",
          3445 => x"38",
          3446 => x"06",
          3447 => x"c3",
          3448 => x"1a",
          3449 => x"38",
          3450 => x"06",
          3451 => x"2e",
          3452 => x"52",
          3453 => x"a6",
          3454 => x"84",
          3455 => x"82",
          3456 => x"75",
          3457 => x"d3",
          3458 => x"9c",
          3459 => x"39",
          3460 => x"74",
          3461 => x"d3",
          3462 => x"3d",
          3463 => x"3d",
          3464 => x"65",
          3465 => x"5d",
          3466 => x"0c",
          3467 => x"05",
          3468 => x"f9",
          3469 => x"d3",
          3470 => x"81",
          3471 => x"8a",
          3472 => x"33",
          3473 => x"2e",
          3474 => x"56",
          3475 => x"90",
          3476 => x"06",
          3477 => x"74",
          3478 => x"b6",
          3479 => x"82",
          3480 => x"34",
          3481 => x"aa",
          3482 => x"91",
          3483 => x"56",
          3484 => x"8c",
          3485 => x"1a",
          3486 => x"74",
          3487 => x"38",
          3488 => x"80",
          3489 => x"38",
          3490 => x"70",
          3491 => x"56",
          3492 => x"b2",
          3493 => x"11",
          3494 => x"77",
          3495 => x"5b",
          3496 => x"38",
          3497 => x"88",
          3498 => x"8f",
          3499 => x"08",
          3500 => x"d5",
          3501 => x"d3",
          3502 => x"81",
          3503 => x"9f",
          3504 => x"2e",
          3505 => x"74",
          3506 => x"98",
          3507 => x"7e",
          3508 => x"3f",
          3509 => x"08",
          3510 => x"83",
          3511 => x"84",
          3512 => x"89",
          3513 => x"77",
          3514 => x"d6",
          3515 => x"7f",
          3516 => x"58",
          3517 => x"75",
          3518 => x"75",
          3519 => x"77",
          3520 => x"7c",
          3521 => x"33",
          3522 => x"3f",
          3523 => x"08",
          3524 => x"7e",
          3525 => x"56",
          3526 => x"2e",
          3527 => x"16",
          3528 => x"55",
          3529 => x"94",
          3530 => x"53",
          3531 => x"b0",
          3532 => x"31",
          3533 => x"05",
          3534 => x"3f",
          3535 => x"56",
          3536 => x"9c",
          3537 => x"19",
          3538 => x"06",
          3539 => x"31",
          3540 => x"76",
          3541 => x"7b",
          3542 => x"08",
          3543 => x"d1",
          3544 => x"d3",
          3545 => x"81",
          3546 => x"94",
          3547 => x"ff",
          3548 => x"05",
          3549 => x"cf",
          3550 => x"76",
          3551 => x"17",
          3552 => x"1e",
          3553 => x"18",
          3554 => x"5e",
          3555 => x"39",
          3556 => x"81",
          3557 => x"90",
          3558 => x"f2",
          3559 => x"63",
          3560 => x"40",
          3561 => x"7e",
          3562 => x"fc",
          3563 => x"51",
          3564 => x"81",
          3565 => x"55",
          3566 => x"08",
          3567 => x"18",
          3568 => x"80",
          3569 => x"74",
          3570 => x"39",
          3571 => x"70",
          3572 => x"81",
          3573 => x"56",
          3574 => x"80",
          3575 => x"38",
          3576 => x"0b",
          3577 => x"82",
          3578 => x"39",
          3579 => x"19",
          3580 => x"83",
          3581 => x"18",
          3582 => x"56",
          3583 => x"27",
          3584 => x"09",
          3585 => x"2e",
          3586 => x"94",
          3587 => x"83",
          3588 => x"56",
          3589 => x"38",
          3590 => x"22",
          3591 => x"89",
          3592 => x"55",
          3593 => x"75",
          3594 => x"18",
          3595 => x"9c",
          3596 => x"85",
          3597 => x"08",
          3598 => x"d7",
          3599 => x"d3",
          3600 => x"81",
          3601 => x"80",
          3602 => x"38",
          3603 => x"ff",
          3604 => x"ff",
          3605 => x"38",
          3606 => x"0c",
          3607 => x"85",
          3608 => x"19",
          3609 => x"b0",
          3610 => x"19",
          3611 => x"81",
          3612 => x"74",
          3613 => x"3f",
          3614 => x"08",
          3615 => x"98",
          3616 => x"7e",
          3617 => x"3f",
          3618 => x"08",
          3619 => x"d2",
          3620 => x"84",
          3621 => x"89",
          3622 => x"78",
          3623 => x"d5",
          3624 => x"7f",
          3625 => x"58",
          3626 => x"75",
          3627 => x"75",
          3628 => x"78",
          3629 => x"7c",
          3630 => x"33",
          3631 => x"3f",
          3632 => x"08",
          3633 => x"7e",
          3634 => x"78",
          3635 => x"74",
          3636 => x"38",
          3637 => x"b0",
          3638 => x"31",
          3639 => x"05",
          3640 => x"51",
          3641 => x"7e",
          3642 => x"83",
          3643 => x"89",
          3644 => x"db",
          3645 => x"08",
          3646 => x"26",
          3647 => x"51",
          3648 => x"81",
          3649 => x"fd",
          3650 => x"77",
          3651 => x"55",
          3652 => x"0c",
          3653 => x"83",
          3654 => x"80",
          3655 => x"55",
          3656 => x"83",
          3657 => x"9c",
          3658 => x"7e",
          3659 => x"3f",
          3660 => x"08",
          3661 => x"75",
          3662 => x"94",
          3663 => x"ff",
          3664 => x"05",
          3665 => x"3f",
          3666 => x"0b",
          3667 => x"7b",
          3668 => x"08",
          3669 => x"76",
          3670 => x"08",
          3671 => x"1c",
          3672 => x"08",
          3673 => x"5c",
          3674 => x"83",
          3675 => x"74",
          3676 => x"fd",
          3677 => x"18",
          3678 => x"07",
          3679 => x"19",
          3680 => x"75",
          3681 => x"0c",
          3682 => x"04",
          3683 => x"7a",
          3684 => x"05",
          3685 => x"56",
          3686 => x"81",
          3687 => x"57",
          3688 => x"08",
          3689 => x"90",
          3690 => x"86",
          3691 => x"06",
          3692 => x"73",
          3693 => x"e9",
          3694 => x"08",
          3695 => x"cc",
          3696 => x"d3",
          3697 => x"81",
          3698 => x"80",
          3699 => x"16",
          3700 => x"33",
          3701 => x"55",
          3702 => x"34",
          3703 => x"53",
          3704 => x"08",
          3705 => x"3f",
          3706 => x"52",
          3707 => x"c9",
          3708 => x"88",
          3709 => x"96",
          3710 => x"f0",
          3711 => x"92",
          3712 => x"ca",
          3713 => x"81",
          3714 => x"34",
          3715 => x"df",
          3716 => x"84",
          3717 => x"33",
          3718 => x"55",
          3719 => x"17",
          3720 => x"d3",
          3721 => x"3d",
          3722 => x"3d",
          3723 => x"52",
          3724 => x"3f",
          3725 => x"08",
          3726 => x"84",
          3727 => x"86",
          3728 => x"52",
          3729 => x"bc",
          3730 => x"84",
          3731 => x"d3",
          3732 => x"38",
          3733 => x"08",
          3734 => x"81",
          3735 => x"86",
          3736 => x"ff",
          3737 => x"3d",
          3738 => x"3f",
          3739 => x"0b",
          3740 => x"08",
          3741 => x"81",
          3742 => x"81",
          3743 => x"80",
          3744 => x"d3",
          3745 => x"3d",
          3746 => x"3d",
          3747 => x"93",
          3748 => x"52",
          3749 => x"e9",
          3750 => x"d3",
          3751 => x"81",
          3752 => x"80",
          3753 => x"58",
          3754 => x"3d",
          3755 => x"e0",
          3756 => x"d3",
          3757 => x"81",
          3758 => x"bc",
          3759 => x"c7",
          3760 => x"98",
          3761 => x"73",
          3762 => x"38",
          3763 => x"12",
          3764 => x"39",
          3765 => x"33",
          3766 => x"70",
          3767 => x"55",
          3768 => x"2e",
          3769 => x"7f",
          3770 => x"54",
          3771 => x"81",
          3772 => x"94",
          3773 => x"39",
          3774 => x"08",
          3775 => x"81",
          3776 => x"85",
          3777 => x"d3",
          3778 => x"3d",
          3779 => x"3d",
          3780 => x"5b",
          3781 => x"34",
          3782 => x"3d",
          3783 => x"52",
          3784 => x"e8",
          3785 => x"d3",
          3786 => x"81",
          3787 => x"82",
          3788 => x"43",
          3789 => x"11",
          3790 => x"58",
          3791 => x"80",
          3792 => x"38",
          3793 => x"3d",
          3794 => x"d5",
          3795 => x"d3",
          3796 => x"81",
          3797 => x"82",
          3798 => x"52",
          3799 => x"c8",
          3800 => x"84",
          3801 => x"d3",
          3802 => x"c1",
          3803 => x"7b",
          3804 => x"3f",
          3805 => x"08",
          3806 => x"74",
          3807 => x"3f",
          3808 => x"08",
          3809 => x"84",
          3810 => x"38",
          3811 => x"51",
          3812 => x"81",
          3813 => x"57",
          3814 => x"08",
          3815 => x"52",
          3816 => x"f2",
          3817 => x"d3",
          3818 => x"a6",
          3819 => x"74",
          3820 => x"3f",
          3821 => x"08",
          3822 => x"84",
          3823 => x"cc",
          3824 => x"2e",
          3825 => x"86",
          3826 => x"81",
          3827 => x"81",
          3828 => x"3d",
          3829 => x"52",
          3830 => x"c9",
          3831 => x"3d",
          3832 => x"11",
          3833 => x"5a",
          3834 => x"2e",
          3835 => x"b9",
          3836 => x"16",
          3837 => x"33",
          3838 => x"73",
          3839 => x"16",
          3840 => x"26",
          3841 => x"75",
          3842 => x"38",
          3843 => x"05",
          3844 => x"6f",
          3845 => x"ff",
          3846 => x"55",
          3847 => x"74",
          3848 => x"38",
          3849 => x"11",
          3850 => x"74",
          3851 => x"39",
          3852 => x"09",
          3853 => x"38",
          3854 => x"11",
          3855 => x"74",
          3856 => x"81",
          3857 => x"70",
          3858 => x"c2",
          3859 => x"08",
          3860 => x"5c",
          3861 => x"73",
          3862 => x"38",
          3863 => x"1a",
          3864 => x"55",
          3865 => x"38",
          3866 => x"73",
          3867 => x"38",
          3868 => x"76",
          3869 => x"74",
          3870 => x"33",
          3871 => x"05",
          3872 => x"15",
          3873 => x"ba",
          3874 => x"05",
          3875 => x"ff",
          3876 => x"06",
          3877 => x"57",
          3878 => x"18",
          3879 => x"54",
          3880 => x"70",
          3881 => x"34",
          3882 => x"ee",
          3883 => x"34",
          3884 => x"84",
          3885 => x"0d",
          3886 => x"0d",
          3887 => x"3d",
          3888 => x"71",
          3889 => x"ec",
          3890 => x"d3",
          3891 => x"81",
          3892 => x"82",
          3893 => x"15",
          3894 => x"82",
          3895 => x"15",
          3896 => x"76",
          3897 => x"90",
          3898 => x"81",
          3899 => x"06",
          3900 => x"72",
          3901 => x"56",
          3902 => x"54",
          3903 => x"17",
          3904 => x"78",
          3905 => x"38",
          3906 => x"22",
          3907 => x"59",
          3908 => x"78",
          3909 => x"76",
          3910 => x"51",
          3911 => x"3f",
          3912 => x"08",
          3913 => x"54",
          3914 => x"53",
          3915 => x"3f",
          3916 => x"08",
          3917 => x"38",
          3918 => x"75",
          3919 => x"18",
          3920 => x"31",
          3921 => x"57",
          3922 => x"b1",
          3923 => x"08",
          3924 => x"38",
          3925 => x"51",
          3926 => x"81",
          3927 => x"54",
          3928 => x"08",
          3929 => x"9a",
          3930 => x"84",
          3931 => x"81",
          3932 => x"d3",
          3933 => x"16",
          3934 => x"16",
          3935 => x"2e",
          3936 => x"76",
          3937 => x"dc",
          3938 => x"31",
          3939 => x"18",
          3940 => x"90",
          3941 => x"81",
          3942 => x"06",
          3943 => x"56",
          3944 => x"9a",
          3945 => x"74",
          3946 => x"3f",
          3947 => x"08",
          3948 => x"84",
          3949 => x"81",
          3950 => x"56",
          3951 => x"52",
          3952 => x"84",
          3953 => x"84",
          3954 => x"ff",
          3955 => x"81",
          3956 => x"38",
          3957 => x"98",
          3958 => x"a6",
          3959 => x"16",
          3960 => x"39",
          3961 => x"16",
          3962 => x"75",
          3963 => x"53",
          3964 => x"aa",
          3965 => x"79",
          3966 => x"3f",
          3967 => x"08",
          3968 => x"0b",
          3969 => x"82",
          3970 => x"39",
          3971 => x"16",
          3972 => x"bb",
          3973 => x"2a",
          3974 => x"08",
          3975 => x"15",
          3976 => x"15",
          3977 => x"90",
          3978 => x"16",
          3979 => x"33",
          3980 => x"53",
          3981 => x"34",
          3982 => x"06",
          3983 => x"2e",
          3984 => x"9c",
          3985 => x"85",
          3986 => x"16",
          3987 => x"72",
          3988 => x"0c",
          3989 => x"04",
          3990 => x"79",
          3991 => x"75",
          3992 => x"8a",
          3993 => x"89",
          3994 => x"52",
          3995 => x"05",
          3996 => x"3f",
          3997 => x"08",
          3998 => x"84",
          3999 => x"38",
          4000 => x"7a",
          4001 => x"d8",
          4002 => x"d3",
          4003 => x"81",
          4004 => x"80",
          4005 => x"16",
          4006 => x"2b",
          4007 => x"74",
          4008 => x"86",
          4009 => x"84",
          4010 => x"06",
          4011 => x"73",
          4012 => x"38",
          4013 => x"52",
          4014 => x"da",
          4015 => x"84",
          4016 => x"0c",
          4017 => x"14",
          4018 => x"23",
          4019 => x"51",
          4020 => x"81",
          4021 => x"55",
          4022 => x"09",
          4023 => x"38",
          4024 => x"39",
          4025 => x"84",
          4026 => x"0c",
          4027 => x"81",
          4028 => x"89",
          4029 => x"fc",
          4030 => x"87",
          4031 => x"53",
          4032 => x"e7",
          4033 => x"d3",
          4034 => x"38",
          4035 => x"08",
          4036 => x"3d",
          4037 => x"3d",
          4038 => x"89",
          4039 => x"54",
          4040 => x"54",
          4041 => x"81",
          4042 => x"53",
          4043 => x"08",
          4044 => x"74",
          4045 => x"d3",
          4046 => x"73",
          4047 => x"3f",
          4048 => x"08",
          4049 => x"39",
          4050 => x"08",
          4051 => x"d3",
          4052 => x"d3",
          4053 => x"81",
          4054 => x"84",
          4055 => x"06",
          4056 => x"53",
          4057 => x"d3",
          4058 => x"38",
          4059 => x"51",
          4060 => x"72",
          4061 => x"cf",
          4062 => x"d3",
          4063 => x"32",
          4064 => x"72",
          4065 => x"70",
          4066 => x"08",
          4067 => x"54",
          4068 => x"d3",
          4069 => x"3d",
          4070 => x"3d",
          4071 => x"80",
          4072 => x"70",
          4073 => x"52",
          4074 => x"3f",
          4075 => x"08",
          4076 => x"84",
          4077 => x"64",
          4078 => x"d6",
          4079 => x"d3",
          4080 => x"81",
          4081 => x"a0",
          4082 => x"cb",
          4083 => x"98",
          4084 => x"73",
          4085 => x"38",
          4086 => x"39",
          4087 => x"88",
          4088 => x"75",
          4089 => x"3f",
          4090 => x"84",
          4091 => x"0d",
          4092 => x"0d",
          4093 => x"5c",
          4094 => x"3d",
          4095 => x"93",
          4096 => x"d6",
          4097 => x"84",
          4098 => x"d3",
          4099 => x"80",
          4100 => x"0c",
          4101 => x"11",
          4102 => x"90",
          4103 => x"56",
          4104 => x"74",
          4105 => x"75",
          4106 => x"e4",
          4107 => x"81",
          4108 => x"5b",
          4109 => x"81",
          4110 => x"75",
          4111 => x"73",
          4112 => x"81",
          4113 => x"82",
          4114 => x"76",
          4115 => x"f0",
          4116 => x"f4",
          4117 => x"84",
          4118 => x"d1",
          4119 => x"84",
          4120 => x"ce",
          4121 => x"84",
          4122 => x"81",
          4123 => x"07",
          4124 => x"05",
          4125 => x"53",
          4126 => x"98",
          4127 => x"26",
          4128 => x"f9",
          4129 => x"08",
          4130 => x"08",
          4131 => x"98",
          4132 => x"81",
          4133 => x"58",
          4134 => x"3f",
          4135 => x"08",
          4136 => x"84",
          4137 => x"38",
          4138 => x"77",
          4139 => x"5d",
          4140 => x"74",
          4141 => x"81",
          4142 => x"b4",
          4143 => x"bb",
          4144 => x"d3",
          4145 => x"ff",
          4146 => x"30",
          4147 => x"1b",
          4148 => x"5b",
          4149 => x"39",
          4150 => x"ff",
          4151 => x"81",
          4152 => x"f0",
          4153 => x"30",
          4154 => x"1b",
          4155 => x"5b",
          4156 => x"83",
          4157 => x"58",
          4158 => x"92",
          4159 => x"0c",
          4160 => x"12",
          4161 => x"33",
          4162 => x"54",
          4163 => x"34",
          4164 => x"84",
          4165 => x"0d",
          4166 => x"0d",
          4167 => x"fc",
          4168 => x"52",
          4169 => x"3f",
          4170 => x"08",
          4171 => x"84",
          4172 => x"38",
          4173 => x"56",
          4174 => x"38",
          4175 => x"70",
          4176 => x"81",
          4177 => x"55",
          4178 => x"80",
          4179 => x"38",
          4180 => x"54",
          4181 => x"08",
          4182 => x"38",
          4183 => x"81",
          4184 => x"53",
          4185 => x"52",
          4186 => x"8c",
          4187 => x"84",
          4188 => x"19",
          4189 => x"c9",
          4190 => x"08",
          4191 => x"ff",
          4192 => x"81",
          4193 => x"ff",
          4194 => x"06",
          4195 => x"56",
          4196 => x"08",
          4197 => x"81",
          4198 => x"82",
          4199 => x"75",
          4200 => x"54",
          4201 => x"08",
          4202 => x"27",
          4203 => x"17",
          4204 => x"d3",
          4205 => x"76",
          4206 => x"3f",
          4207 => x"08",
          4208 => x"08",
          4209 => x"90",
          4210 => x"c0",
          4211 => x"90",
          4212 => x"80",
          4213 => x"75",
          4214 => x"75",
          4215 => x"d3",
          4216 => x"3d",
          4217 => x"3d",
          4218 => x"a0",
          4219 => x"05",
          4220 => x"51",
          4221 => x"81",
          4222 => x"55",
          4223 => x"08",
          4224 => x"78",
          4225 => x"08",
          4226 => x"70",
          4227 => x"ae",
          4228 => x"84",
          4229 => x"d3",
          4230 => x"db",
          4231 => x"fb",
          4232 => x"85",
          4233 => x"06",
          4234 => x"86",
          4235 => x"c7",
          4236 => x"2b",
          4237 => x"24",
          4238 => x"02",
          4239 => x"33",
          4240 => x"58",
          4241 => x"76",
          4242 => x"6b",
          4243 => x"cc",
          4244 => x"d3",
          4245 => x"84",
          4246 => x"06",
          4247 => x"73",
          4248 => x"d4",
          4249 => x"81",
          4250 => x"94",
          4251 => x"81",
          4252 => x"5a",
          4253 => x"08",
          4254 => x"8a",
          4255 => x"54",
          4256 => x"81",
          4257 => x"55",
          4258 => x"08",
          4259 => x"81",
          4260 => x"52",
          4261 => x"e5",
          4262 => x"84",
          4263 => x"d3",
          4264 => x"38",
          4265 => x"cf",
          4266 => x"84",
          4267 => x"88",
          4268 => x"84",
          4269 => x"38",
          4270 => x"c2",
          4271 => x"84",
          4272 => x"84",
          4273 => x"81",
          4274 => x"07",
          4275 => x"55",
          4276 => x"2e",
          4277 => x"80",
          4278 => x"80",
          4279 => x"77",
          4280 => x"3f",
          4281 => x"08",
          4282 => x"38",
          4283 => x"ba",
          4284 => x"d3",
          4285 => x"74",
          4286 => x"0c",
          4287 => x"04",
          4288 => x"82",
          4289 => x"c0",
          4290 => x"3d",
          4291 => x"3f",
          4292 => x"08",
          4293 => x"84",
          4294 => x"38",
          4295 => x"52",
          4296 => x"52",
          4297 => x"3f",
          4298 => x"08",
          4299 => x"84",
          4300 => x"88",
          4301 => x"39",
          4302 => x"08",
          4303 => x"81",
          4304 => x"38",
          4305 => x"05",
          4306 => x"2a",
          4307 => x"55",
          4308 => x"81",
          4309 => x"5a",
          4310 => x"3d",
          4311 => x"c1",
          4312 => x"d3",
          4313 => x"55",
          4314 => x"84",
          4315 => x"87",
          4316 => x"84",
          4317 => x"09",
          4318 => x"38",
          4319 => x"d3",
          4320 => x"2e",
          4321 => x"86",
          4322 => x"81",
          4323 => x"81",
          4324 => x"d3",
          4325 => x"78",
          4326 => x"3f",
          4327 => x"08",
          4328 => x"84",
          4329 => x"38",
          4330 => x"52",
          4331 => x"ff",
          4332 => x"78",
          4333 => x"b4",
          4334 => x"54",
          4335 => x"15",
          4336 => x"b2",
          4337 => x"ca",
          4338 => x"b6",
          4339 => x"53",
          4340 => x"53",
          4341 => x"3f",
          4342 => x"b4",
          4343 => x"d4",
          4344 => x"b6",
          4345 => x"54",
          4346 => x"d5",
          4347 => x"53",
          4348 => x"11",
          4349 => x"d7",
          4350 => x"81",
          4351 => x"34",
          4352 => x"a4",
          4353 => x"84",
          4354 => x"d3",
          4355 => x"38",
          4356 => x"0a",
          4357 => x"05",
          4358 => x"d0",
          4359 => x"64",
          4360 => x"c9",
          4361 => x"54",
          4362 => x"15",
          4363 => x"81",
          4364 => x"34",
          4365 => x"b8",
          4366 => x"d3",
          4367 => x"8b",
          4368 => x"75",
          4369 => x"ff",
          4370 => x"73",
          4371 => x"0c",
          4372 => x"04",
          4373 => x"a9",
          4374 => x"51",
          4375 => x"82",
          4376 => x"ff",
          4377 => x"a9",
          4378 => x"ee",
          4379 => x"84",
          4380 => x"d3",
          4381 => x"d3",
          4382 => x"a9",
          4383 => x"9d",
          4384 => x"58",
          4385 => x"81",
          4386 => x"55",
          4387 => x"08",
          4388 => x"02",
          4389 => x"33",
          4390 => x"54",
          4391 => x"82",
          4392 => x"53",
          4393 => x"52",
          4394 => x"88",
          4395 => x"b4",
          4396 => x"53",
          4397 => x"3d",
          4398 => x"ff",
          4399 => x"aa",
          4400 => x"73",
          4401 => x"3f",
          4402 => x"08",
          4403 => x"84",
          4404 => x"63",
          4405 => x"81",
          4406 => x"65",
          4407 => x"2e",
          4408 => x"55",
          4409 => x"81",
          4410 => x"84",
          4411 => x"06",
          4412 => x"73",
          4413 => x"3f",
          4414 => x"08",
          4415 => x"84",
          4416 => x"38",
          4417 => x"53",
          4418 => x"95",
          4419 => x"16",
          4420 => x"87",
          4421 => x"05",
          4422 => x"34",
          4423 => x"70",
          4424 => x"81",
          4425 => x"55",
          4426 => x"74",
          4427 => x"73",
          4428 => x"78",
          4429 => x"83",
          4430 => x"16",
          4431 => x"2a",
          4432 => x"51",
          4433 => x"80",
          4434 => x"38",
          4435 => x"80",
          4436 => x"52",
          4437 => x"be",
          4438 => x"84",
          4439 => x"51",
          4440 => x"3f",
          4441 => x"d3",
          4442 => x"2e",
          4443 => x"81",
          4444 => x"52",
          4445 => x"b5",
          4446 => x"d3",
          4447 => x"80",
          4448 => x"58",
          4449 => x"84",
          4450 => x"38",
          4451 => x"54",
          4452 => x"09",
          4453 => x"38",
          4454 => x"52",
          4455 => x"af",
          4456 => x"81",
          4457 => x"34",
          4458 => x"d3",
          4459 => x"38",
          4460 => x"ca",
          4461 => x"84",
          4462 => x"d3",
          4463 => x"38",
          4464 => x"b5",
          4465 => x"d3",
          4466 => x"74",
          4467 => x"0c",
          4468 => x"04",
          4469 => x"02",
          4470 => x"33",
          4471 => x"80",
          4472 => x"57",
          4473 => x"95",
          4474 => x"52",
          4475 => x"d2",
          4476 => x"d3",
          4477 => x"81",
          4478 => x"80",
          4479 => x"5a",
          4480 => x"3d",
          4481 => x"c9",
          4482 => x"d3",
          4483 => x"81",
          4484 => x"b8",
          4485 => x"cf",
          4486 => x"a0",
          4487 => x"55",
          4488 => x"75",
          4489 => x"71",
          4490 => x"33",
          4491 => x"74",
          4492 => x"57",
          4493 => x"8b",
          4494 => x"54",
          4495 => x"15",
          4496 => x"ff",
          4497 => x"81",
          4498 => x"55",
          4499 => x"84",
          4500 => x"0d",
          4501 => x"0d",
          4502 => x"53",
          4503 => x"05",
          4504 => x"51",
          4505 => x"81",
          4506 => x"55",
          4507 => x"08",
          4508 => x"76",
          4509 => x"93",
          4510 => x"51",
          4511 => x"81",
          4512 => x"55",
          4513 => x"08",
          4514 => x"80",
          4515 => x"81",
          4516 => x"86",
          4517 => x"38",
          4518 => x"86",
          4519 => x"90",
          4520 => x"54",
          4521 => x"ff",
          4522 => x"76",
          4523 => x"83",
          4524 => x"51",
          4525 => x"3f",
          4526 => x"08",
          4527 => x"d3",
          4528 => x"3d",
          4529 => x"3d",
          4530 => x"5c",
          4531 => x"98",
          4532 => x"52",
          4533 => x"d1",
          4534 => x"d3",
          4535 => x"d3",
          4536 => x"70",
          4537 => x"08",
          4538 => x"51",
          4539 => x"80",
          4540 => x"38",
          4541 => x"06",
          4542 => x"80",
          4543 => x"38",
          4544 => x"5f",
          4545 => x"3d",
          4546 => x"ff",
          4547 => x"81",
          4548 => x"57",
          4549 => x"08",
          4550 => x"74",
          4551 => x"c3",
          4552 => x"d3",
          4553 => x"81",
          4554 => x"bf",
          4555 => x"84",
          4556 => x"84",
          4557 => x"59",
          4558 => x"81",
          4559 => x"56",
          4560 => x"33",
          4561 => x"16",
          4562 => x"27",
          4563 => x"56",
          4564 => x"80",
          4565 => x"80",
          4566 => x"ff",
          4567 => x"70",
          4568 => x"56",
          4569 => x"e8",
          4570 => x"76",
          4571 => x"81",
          4572 => x"80",
          4573 => x"57",
          4574 => x"78",
          4575 => x"51",
          4576 => x"2e",
          4577 => x"73",
          4578 => x"38",
          4579 => x"08",
          4580 => x"b1",
          4581 => x"d3",
          4582 => x"81",
          4583 => x"a7",
          4584 => x"33",
          4585 => x"c3",
          4586 => x"2e",
          4587 => x"e4",
          4588 => x"2e",
          4589 => x"56",
          4590 => x"05",
          4591 => x"e3",
          4592 => x"84",
          4593 => x"76",
          4594 => x"0c",
          4595 => x"04",
          4596 => x"82",
          4597 => x"ff",
          4598 => x"9d",
          4599 => x"fa",
          4600 => x"84",
          4601 => x"84",
          4602 => x"81",
          4603 => x"83",
          4604 => x"53",
          4605 => x"3d",
          4606 => x"ff",
          4607 => x"73",
          4608 => x"70",
          4609 => x"52",
          4610 => x"9f",
          4611 => x"bc",
          4612 => x"74",
          4613 => x"6d",
          4614 => x"70",
          4615 => x"af",
          4616 => x"d3",
          4617 => x"2e",
          4618 => x"70",
          4619 => x"57",
          4620 => x"fd",
          4621 => x"84",
          4622 => x"8d",
          4623 => x"2b",
          4624 => x"81",
          4625 => x"86",
          4626 => x"84",
          4627 => x"9f",
          4628 => x"ff",
          4629 => x"54",
          4630 => x"8a",
          4631 => x"70",
          4632 => x"06",
          4633 => x"ff",
          4634 => x"38",
          4635 => x"15",
          4636 => x"80",
          4637 => x"74",
          4638 => x"f8",
          4639 => x"89",
          4640 => x"84",
          4641 => x"81",
          4642 => x"88",
          4643 => x"26",
          4644 => x"39",
          4645 => x"86",
          4646 => x"81",
          4647 => x"ff",
          4648 => x"38",
          4649 => x"54",
          4650 => x"81",
          4651 => x"81",
          4652 => x"78",
          4653 => x"5a",
          4654 => x"6d",
          4655 => x"81",
          4656 => x"57",
          4657 => x"9f",
          4658 => x"38",
          4659 => x"54",
          4660 => x"81",
          4661 => x"b1",
          4662 => x"2e",
          4663 => x"a7",
          4664 => x"15",
          4665 => x"54",
          4666 => x"09",
          4667 => x"38",
          4668 => x"76",
          4669 => x"41",
          4670 => x"52",
          4671 => x"52",
          4672 => x"b3",
          4673 => x"84",
          4674 => x"d3",
          4675 => x"f7",
          4676 => x"74",
          4677 => x"e5",
          4678 => x"84",
          4679 => x"d3",
          4680 => x"38",
          4681 => x"38",
          4682 => x"74",
          4683 => x"39",
          4684 => x"08",
          4685 => x"81",
          4686 => x"38",
          4687 => x"74",
          4688 => x"38",
          4689 => x"51",
          4690 => x"3f",
          4691 => x"08",
          4692 => x"84",
          4693 => x"a0",
          4694 => x"84",
          4695 => x"51",
          4696 => x"3f",
          4697 => x"0b",
          4698 => x"8b",
          4699 => x"67",
          4700 => x"a7",
          4701 => x"81",
          4702 => x"34",
          4703 => x"ad",
          4704 => x"d3",
          4705 => x"73",
          4706 => x"d3",
          4707 => x"3d",
          4708 => x"3d",
          4709 => x"02",
          4710 => x"cb",
          4711 => x"3d",
          4712 => x"72",
          4713 => x"5a",
          4714 => x"81",
          4715 => x"58",
          4716 => x"08",
          4717 => x"91",
          4718 => x"77",
          4719 => x"7c",
          4720 => x"38",
          4721 => x"59",
          4722 => x"90",
          4723 => x"81",
          4724 => x"06",
          4725 => x"73",
          4726 => x"54",
          4727 => x"82",
          4728 => x"39",
          4729 => x"8b",
          4730 => x"11",
          4731 => x"2b",
          4732 => x"54",
          4733 => x"fe",
          4734 => x"ff",
          4735 => x"70",
          4736 => x"07",
          4737 => x"d3",
          4738 => x"8c",
          4739 => x"40",
          4740 => x"55",
          4741 => x"88",
          4742 => x"08",
          4743 => x"38",
          4744 => x"77",
          4745 => x"56",
          4746 => x"51",
          4747 => x"3f",
          4748 => x"55",
          4749 => x"08",
          4750 => x"38",
          4751 => x"d3",
          4752 => x"2e",
          4753 => x"81",
          4754 => x"ff",
          4755 => x"38",
          4756 => x"08",
          4757 => x"16",
          4758 => x"2e",
          4759 => x"87",
          4760 => x"74",
          4761 => x"74",
          4762 => x"81",
          4763 => x"38",
          4764 => x"ff",
          4765 => x"2e",
          4766 => x"7b",
          4767 => x"80",
          4768 => x"81",
          4769 => x"81",
          4770 => x"06",
          4771 => x"56",
          4772 => x"52",
          4773 => x"af",
          4774 => x"d3",
          4775 => x"81",
          4776 => x"80",
          4777 => x"81",
          4778 => x"56",
          4779 => x"d3",
          4780 => x"ff",
          4781 => x"7c",
          4782 => x"55",
          4783 => x"b3",
          4784 => x"1b",
          4785 => x"1b",
          4786 => x"33",
          4787 => x"54",
          4788 => x"34",
          4789 => x"fe",
          4790 => x"08",
          4791 => x"74",
          4792 => x"75",
          4793 => x"16",
          4794 => x"33",
          4795 => x"73",
          4796 => x"77",
          4797 => x"d3",
          4798 => x"3d",
          4799 => x"3d",
          4800 => x"02",
          4801 => x"eb",
          4802 => x"3d",
          4803 => x"59",
          4804 => x"8b",
          4805 => x"81",
          4806 => x"24",
          4807 => x"81",
          4808 => x"84",
          4809 => x"a0",
          4810 => x"51",
          4811 => x"2e",
          4812 => x"75",
          4813 => x"84",
          4814 => x"06",
          4815 => x"7e",
          4816 => x"d0",
          4817 => x"84",
          4818 => x"06",
          4819 => x"56",
          4820 => x"74",
          4821 => x"76",
          4822 => x"81",
          4823 => x"8a",
          4824 => x"b2",
          4825 => x"fc",
          4826 => x"52",
          4827 => x"a4",
          4828 => x"d3",
          4829 => x"38",
          4830 => x"80",
          4831 => x"74",
          4832 => x"26",
          4833 => x"15",
          4834 => x"74",
          4835 => x"38",
          4836 => x"80",
          4837 => x"84",
          4838 => x"92",
          4839 => x"80",
          4840 => x"38",
          4841 => x"06",
          4842 => x"2e",
          4843 => x"56",
          4844 => x"78",
          4845 => x"89",
          4846 => x"2b",
          4847 => x"43",
          4848 => x"38",
          4849 => x"30",
          4850 => x"77",
          4851 => x"91",
          4852 => x"c2",
          4853 => x"f8",
          4854 => x"52",
          4855 => x"a4",
          4856 => x"56",
          4857 => x"08",
          4858 => x"77",
          4859 => x"77",
          4860 => x"84",
          4861 => x"45",
          4862 => x"bf",
          4863 => x"8e",
          4864 => x"26",
          4865 => x"74",
          4866 => x"48",
          4867 => x"75",
          4868 => x"38",
          4869 => x"81",
          4870 => x"fa",
          4871 => x"2a",
          4872 => x"56",
          4873 => x"2e",
          4874 => x"87",
          4875 => x"82",
          4876 => x"38",
          4877 => x"55",
          4878 => x"83",
          4879 => x"81",
          4880 => x"56",
          4881 => x"80",
          4882 => x"38",
          4883 => x"83",
          4884 => x"06",
          4885 => x"78",
          4886 => x"91",
          4887 => x"0b",
          4888 => x"22",
          4889 => x"80",
          4890 => x"74",
          4891 => x"38",
          4892 => x"56",
          4893 => x"17",
          4894 => x"57",
          4895 => x"2e",
          4896 => x"75",
          4897 => x"79",
          4898 => x"fe",
          4899 => x"81",
          4900 => x"84",
          4901 => x"05",
          4902 => x"5e",
          4903 => x"80",
          4904 => x"84",
          4905 => x"8a",
          4906 => x"fd",
          4907 => x"75",
          4908 => x"38",
          4909 => x"78",
          4910 => x"8c",
          4911 => x"0b",
          4912 => x"22",
          4913 => x"80",
          4914 => x"74",
          4915 => x"38",
          4916 => x"56",
          4917 => x"17",
          4918 => x"57",
          4919 => x"2e",
          4920 => x"75",
          4921 => x"79",
          4922 => x"fe",
          4923 => x"81",
          4924 => x"10",
          4925 => x"81",
          4926 => x"9f",
          4927 => x"38",
          4928 => x"d3",
          4929 => x"81",
          4930 => x"05",
          4931 => x"2a",
          4932 => x"56",
          4933 => x"17",
          4934 => x"81",
          4935 => x"60",
          4936 => x"65",
          4937 => x"12",
          4938 => x"30",
          4939 => x"74",
          4940 => x"59",
          4941 => x"7d",
          4942 => x"81",
          4943 => x"76",
          4944 => x"41",
          4945 => x"76",
          4946 => x"90",
          4947 => x"62",
          4948 => x"51",
          4949 => x"26",
          4950 => x"75",
          4951 => x"31",
          4952 => x"65",
          4953 => x"fe",
          4954 => x"81",
          4955 => x"58",
          4956 => x"09",
          4957 => x"38",
          4958 => x"08",
          4959 => x"26",
          4960 => x"78",
          4961 => x"79",
          4962 => x"78",
          4963 => x"86",
          4964 => x"82",
          4965 => x"06",
          4966 => x"83",
          4967 => x"81",
          4968 => x"27",
          4969 => x"8f",
          4970 => x"55",
          4971 => x"26",
          4972 => x"59",
          4973 => x"62",
          4974 => x"74",
          4975 => x"38",
          4976 => x"88",
          4977 => x"84",
          4978 => x"26",
          4979 => x"86",
          4980 => x"1a",
          4981 => x"79",
          4982 => x"38",
          4983 => x"80",
          4984 => x"2e",
          4985 => x"83",
          4986 => x"9f",
          4987 => x"8b",
          4988 => x"06",
          4989 => x"74",
          4990 => x"84",
          4991 => x"52",
          4992 => x"a2",
          4993 => x"53",
          4994 => x"52",
          4995 => x"a2",
          4996 => x"80",
          4997 => x"51",
          4998 => x"3f",
          4999 => x"34",
          5000 => x"ff",
          5001 => x"1b",
          5002 => x"a2",
          5003 => x"90",
          5004 => x"83",
          5005 => x"70",
          5006 => x"80",
          5007 => x"55",
          5008 => x"ff",
          5009 => x"66",
          5010 => x"ff",
          5011 => x"38",
          5012 => x"ff",
          5013 => x"1b",
          5014 => x"f2",
          5015 => x"74",
          5016 => x"51",
          5017 => x"3f",
          5018 => x"1c",
          5019 => x"98",
          5020 => x"a0",
          5021 => x"ff",
          5022 => x"51",
          5023 => x"3f",
          5024 => x"1b",
          5025 => x"e4",
          5026 => x"2e",
          5027 => x"80",
          5028 => x"88",
          5029 => x"80",
          5030 => x"ff",
          5031 => x"7c",
          5032 => x"51",
          5033 => x"3f",
          5034 => x"1b",
          5035 => x"bc",
          5036 => x"b0",
          5037 => x"a0",
          5038 => x"52",
          5039 => x"ff",
          5040 => x"ff",
          5041 => x"c0",
          5042 => x"0b",
          5043 => x"34",
          5044 => x"c2",
          5045 => x"c7",
          5046 => x"39",
          5047 => x"0a",
          5048 => x"51",
          5049 => x"3f",
          5050 => x"ff",
          5051 => x"1b",
          5052 => x"da",
          5053 => x"0b",
          5054 => x"a9",
          5055 => x"34",
          5056 => x"c2",
          5057 => x"1b",
          5058 => x"8f",
          5059 => x"d5",
          5060 => x"1b",
          5061 => x"ff",
          5062 => x"81",
          5063 => x"7a",
          5064 => x"ff",
          5065 => x"81",
          5066 => x"84",
          5067 => x"38",
          5068 => x"09",
          5069 => x"ee",
          5070 => x"60",
          5071 => x"7a",
          5072 => x"ff",
          5073 => x"84",
          5074 => x"52",
          5075 => x"9f",
          5076 => x"8b",
          5077 => x"52",
          5078 => x"9f",
          5079 => x"8a",
          5080 => x"52",
          5081 => x"51",
          5082 => x"3f",
          5083 => x"83",
          5084 => x"ff",
          5085 => x"82",
          5086 => x"1b",
          5087 => x"ec",
          5088 => x"d5",
          5089 => x"ff",
          5090 => x"75",
          5091 => x"05",
          5092 => x"7e",
          5093 => x"e5",
          5094 => x"60",
          5095 => x"52",
          5096 => x"9a",
          5097 => x"53",
          5098 => x"51",
          5099 => x"3f",
          5100 => x"58",
          5101 => x"09",
          5102 => x"38",
          5103 => x"51",
          5104 => x"3f",
          5105 => x"1b",
          5106 => x"a0",
          5107 => x"52",
          5108 => x"91",
          5109 => x"ff",
          5110 => x"81",
          5111 => x"f8",
          5112 => x"7a",
          5113 => x"84",
          5114 => x"61",
          5115 => x"26",
          5116 => x"57",
          5117 => x"53",
          5118 => x"51",
          5119 => x"3f",
          5120 => x"08",
          5121 => x"84",
          5122 => x"d3",
          5123 => x"7a",
          5124 => x"aa",
          5125 => x"75",
          5126 => x"56",
          5127 => x"81",
          5128 => x"80",
          5129 => x"38",
          5130 => x"83",
          5131 => x"63",
          5132 => x"74",
          5133 => x"38",
          5134 => x"54",
          5135 => x"52",
          5136 => x"99",
          5137 => x"d3",
          5138 => x"c1",
          5139 => x"75",
          5140 => x"56",
          5141 => x"8c",
          5142 => x"2e",
          5143 => x"56",
          5144 => x"ff",
          5145 => x"84",
          5146 => x"2e",
          5147 => x"56",
          5148 => x"58",
          5149 => x"38",
          5150 => x"77",
          5151 => x"ff",
          5152 => x"82",
          5153 => x"78",
          5154 => x"c2",
          5155 => x"1b",
          5156 => x"34",
          5157 => x"16",
          5158 => x"82",
          5159 => x"83",
          5160 => x"84",
          5161 => x"67",
          5162 => x"fd",
          5163 => x"51",
          5164 => x"3f",
          5165 => x"16",
          5166 => x"84",
          5167 => x"bf",
          5168 => x"86",
          5169 => x"d3",
          5170 => x"16",
          5171 => x"83",
          5172 => x"ff",
          5173 => x"66",
          5174 => x"1b",
          5175 => x"8c",
          5176 => x"77",
          5177 => x"7e",
          5178 => x"91",
          5179 => x"81",
          5180 => x"a2",
          5181 => x"80",
          5182 => x"ff",
          5183 => x"81",
          5184 => x"84",
          5185 => x"89",
          5186 => x"8a",
          5187 => x"86",
          5188 => x"84",
          5189 => x"81",
          5190 => x"99",
          5191 => x"ff",
          5192 => x"52",
          5193 => x"81",
          5194 => x"84",
          5195 => x"80",
          5196 => x"08",
          5197 => x"ac",
          5198 => x"39",
          5199 => x"51",
          5200 => x"81",
          5201 => x"80",
          5202 => x"c5",
          5203 => x"eb",
          5204 => x"f0",
          5205 => x"39",
          5206 => x"51",
          5207 => x"81",
          5208 => x"80",
          5209 => x"c6",
          5210 => x"cf",
          5211 => x"bc",
          5212 => x"39",
          5213 => x"51",
          5214 => x"81",
          5215 => x"bb",
          5216 => x"88",
          5217 => x"81",
          5218 => x"af",
          5219 => x"c8",
          5220 => x"81",
          5221 => x"a3",
          5222 => x"fc",
          5223 => x"81",
          5224 => x"97",
          5225 => x"a8",
          5226 => x"81",
          5227 => x"8b",
          5228 => x"d8",
          5229 => x"81",
          5230 => x"ff",
          5231 => x"83",
          5232 => x"fb",
          5233 => x"79",
          5234 => x"87",
          5235 => x"38",
          5236 => x"87",
          5237 => x"91",
          5238 => x"52",
          5239 => x"ef",
          5240 => x"d3",
          5241 => x"75",
          5242 => x"8b",
          5243 => x"84",
          5244 => x"53",
          5245 => x"c8",
          5246 => x"8d",
          5247 => x"3d",
          5248 => x"3d",
          5249 => x"61",
          5250 => x"80",
          5251 => x"73",
          5252 => x"5f",
          5253 => x"5c",
          5254 => x"52",
          5255 => x"51",
          5256 => x"3f",
          5257 => x"51",
          5258 => x"3f",
          5259 => x"77",
          5260 => x"38",
          5261 => x"89",
          5262 => x"2e",
          5263 => x"c6",
          5264 => x"53",
          5265 => x"8e",
          5266 => x"52",
          5267 => x"51",
          5268 => x"3f",
          5269 => x"c9",
          5270 => x"86",
          5271 => x"15",
          5272 => x"39",
          5273 => x"72",
          5274 => x"38",
          5275 => x"81",
          5276 => x"ff",
          5277 => x"89",
          5278 => x"ac",
          5279 => x"b9",
          5280 => x"55",
          5281 => x"16",
          5282 => x"27",
          5283 => x"33",
          5284 => x"b8",
          5285 => x"85",
          5286 => x"81",
          5287 => x"ff",
          5288 => x"81",
          5289 => x"51",
          5290 => x"3f",
          5291 => x"81",
          5292 => x"ff",
          5293 => x"80",
          5294 => x"27",
          5295 => x"16",
          5296 => x"72",
          5297 => x"53",
          5298 => x"90",
          5299 => x"2e",
          5300 => x"80",
          5301 => x"38",
          5302 => x"39",
          5303 => x"f9",
          5304 => x"15",
          5305 => x"81",
          5306 => x"ff",
          5307 => x"76",
          5308 => x"5a",
          5309 => x"94",
          5310 => x"84",
          5311 => x"70",
          5312 => x"55",
          5313 => x"09",
          5314 => x"38",
          5315 => x"3f",
          5316 => x"08",
          5317 => x"98",
          5318 => x"32",
          5319 => x"72",
          5320 => x"51",
          5321 => x"55",
          5322 => x"8c",
          5323 => x"38",
          5324 => x"09",
          5325 => x"38",
          5326 => x"39",
          5327 => x"72",
          5328 => x"d6",
          5329 => x"72",
          5330 => x"0c",
          5331 => x"04",
          5332 => x"66",
          5333 => x"80",
          5334 => x"69",
          5335 => x"74",
          5336 => x"70",
          5337 => x"27",
          5338 => x"58",
          5339 => x"93",
          5340 => x"fb",
          5341 => x"75",
          5342 => x"70",
          5343 => x"b9",
          5344 => x"84",
          5345 => x"d3",
          5346 => x"38",
          5347 => x"08",
          5348 => x"88",
          5349 => x"84",
          5350 => x"3d",
          5351 => x"84",
          5352 => x"52",
          5353 => x"f6",
          5354 => x"84",
          5355 => x"d3",
          5356 => x"38",
          5357 => x"80",
          5358 => x"74",
          5359 => x"59",
          5360 => x"96",
          5361 => x"51",
          5362 => x"75",
          5363 => x"07",
          5364 => x"55",
          5365 => x"95",
          5366 => x"2e",
          5367 => x"c9",
          5368 => x"c0",
          5369 => x"52",
          5370 => x"d7",
          5371 => x"76",
          5372 => x"0c",
          5373 => x"04",
          5374 => x"7b",
          5375 => x"b3",
          5376 => x"58",
          5377 => x"53",
          5378 => x"51",
          5379 => x"81",
          5380 => x"a4",
          5381 => x"2e",
          5382 => x"81",
          5383 => x"98",
          5384 => x"7f",
          5385 => x"84",
          5386 => x"7d",
          5387 => x"81",
          5388 => x"57",
          5389 => x"04",
          5390 => x"84",
          5391 => x"0d",
          5392 => x"0d",
          5393 => x"33",
          5394 => x"53",
          5395 => x"52",
          5396 => x"c9",
          5397 => x"a4",
          5398 => x"80",
          5399 => x"c9",
          5400 => x"c9",
          5401 => x"d0",
          5402 => x"81",
          5403 => x"ff",
          5404 => x"74",
          5405 => x"38",
          5406 => x"3f",
          5407 => x"04",
          5408 => x"87",
          5409 => x"08",
          5410 => x"fd",
          5411 => x"fe",
          5412 => x"81",
          5413 => x"fe",
          5414 => x"80",
          5415 => x"80",
          5416 => x"2a",
          5417 => x"51",
          5418 => x"2e",
          5419 => x"51",
          5420 => x"3f",
          5421 => x"51",
          5422 => x"3f",
          5423 => x"f5",
          5424 => x"82",
          5425 => x"06",
          5426 => x"80",
          5427 => x"81",
          5428 => x"cc",
          5429 => x"c8",
          5430 => x"c4",
          5431 => x"fe",
          5432 => x"72",
          5433 => x"81",
          5434 => x"71",
          5435 => x"38",
          5436 => x"f5",
          5437 => x"ca",
          5438 => x"f7",
          5439 => x"51",
          5440 => x"3f",
          5441 => x"70",
          5442 => x"52",
          5443 => x"95",
          5444 => x"fe",
          5445 => x"81",
          5446 => x"fe",
          5447 => x"80",
          5448 => x"fc",
          5449 => x"2a",
          5450 => x"51",
          5451 => x"2e",
          5452 => x"51",
          5453 => x"3f",
          5454 => x"51",
          5455 => x"3f",
          5456 => x"f4",
          5457 => x"86",
          5458 => x"06",
          5459 => x"80",
          5460 => x"81",
          5461 => x"c8",
          5462 => x"94",
          5463 => x"c0",
          5464 => x"fe",
          5465 => x"72",
          5466 => x"81",
          5467 => x"71",
          5468 => x"38",
          5469 => x"f4",
          5470 => x"cb",
          5471 => x"f6",
          5472 => x"51",
          5473 => x"3f",
          5474 => x"70",
          5475 => x"52",
          5476 => x"95",
          5477 => x"fe",
          5478 => x"81",
          5479 => x"fe",
          5480 => x"80",
          5481 => x"f8",
          5482 => x"a6",
          5483 => x"0d",
          5484 => x"0d",
          5485 => x"70",
          5486 => x"73",
          5487 => x"f0",
          5488 => x"73",
          5489 => x"15",
          5490 => x"e4",
          5491 => x"54",
          5492 => x"70",
          5493 => x"57",
          5494 => x"a0",
          5495 => x"81",
          5496 => x"2e",
          5497 => x"e5",
          5498 => x"ff",
          5499 => x"a0",
          5500 => x"06",
          5501 => x"74",
          5502 => x"56",
          5503 => x"75",
          5504 => x"d0",
          5505 => x"08",
          5506 => x"52",
          5507 => x"ff",
          5508 => x"84",
          5509 => x"84",
          5510 => x"72",
          5511 => x"a3",
          5512 => x"70",
          5513 => x"57",
          5514 => x"27",
          5515 => x"53",
          5516 => x"84",
          5517 => x"0d",
          5518 => x"0d",
          5519 => x"81",
          5520 => x"5e",
          5521 => x"7b",
          5522 => x"c8",
          5523 => x"84",
          5524 => x"06",
          5525 => x"2e",
          5526 => x"a2",
          5527 => x"fc",
          5528 => x"70",
          5529 => x"84",
          5530 => x"53",
          5531 => x"d4",
          5532 => x"b9",
          5533 => x"d3",
          5534 => x"2e",
          5535 => x"cc",
          5536 => x"e8",
          5537 => x"5e",
          5538 => x"b8",
          5539 => x"a9",
          5540 => x"70",
          5541 => x"f8",
          5542 => x"79",
          5543 => x"de",
          5544 => x"52",
          5545 => x"84",
          5546 => x"3d",
          5547 => x"51",
          5548 => x"81",
          5549 => x"90",
          5550 => x"2c",
          5551 => x"80",
          5552 => x"9b",
          5553 => x"c3",
          5554 => x"38",
          5555 => x"83",
          5556 => x"ab",
          5557 => x"78",
          5558 => x"af",
          5559 => x"24",
          5560 => x"80",
          5561 => x"38",
          5562 => x"78",
          5563 => x"82",
          5564 => x"2e",
          5565 => x"8c",
          5566 => x"80",
          5567 => x"8a",
          5568 => x"c0",
          5569 => x"78",
          5570 => x"a9",
          5571 => x"2e",
          5572 => x"8c",
          5573 => x"80",
          5574 => x"eb",
          5575 => x"c2",
          5576 => x"38",
          5577 => x"78",
          5578 => x"8b",
          5579 => x"80",
          5580 => x"38",
          5581 => x"2e",
          5582 => x"78",
          5583 => x"8b",
          5584 => x"d0",
          5585 => x"38",
          5586 => x"78",
          5587 => x"8a",
          5588 => x"80",
          5589 => x"f2",
          5590 => x"39",
          5591 => x"2e",
          5592 => x"78",
          5593 => x"92",
          5594 => x"f9",
          5595 => x"38",
          5596 => x"2e",
          5597 => x"8b",
          5598 => x"81",
          5599 => x"eb",
          5600 => x"87",
          5601 => x"38",
          5602 => x"b7",
          5603 => x"11",
          5604 => x"05",
          5605 => x"fa",
          5606 => x"84",
          5607 => x"81",
          5608 => x"8c",
          5609 => x"3d",
          5610 => x"53",
          5611 => x"51",
          5612 => x"3f",
          5613 => x"08",
          5614 => x"38",
          5615 => x"83",
          5616 => x"02",
          5617 => x"33",
          5618 => x"cf",
          5619 => x"ff",
          5620 => x"81",
          5621 => x"81",
          5622 => x"78",
          5623 => x"cc",
          5624 => x"fb",
          5625 => x"5d",
          5626 => x"81",
          5627 => x"89",
          5628 => x"3d",
          5629 => x"53",
          5630 => x"51",
          5631 => x"3f",
          5632 => x"08",
          5633 => x"81",
          5634 => x"80",
          5635 => x"cf",
          5636 => x"ff",
          5637 => x"81",
          5638 => x"52",
          5639 => x"51",
          5640 => x"b7",
          5641 => x"11",
          5642 => x"05",
          5643 => x"e2",
          5644 => x"84",
          5645 => x"87",
          5646 => x"26",
          5647 => x"b7",
          5648 => x"11",
          5649 => x"05",
          5650 => x"c6",
          5651 => x"84",
          5652 => x"81",
          5653 => x"43",
          5654 => x"cc",
          5655 => x"51",
          5656 => x"3f",
          5657 => x"05",
          5658 => x"52",
          5659 => x"29",
          5660 => x"05",
          5661 => x"e0",
          5662 => x"84",
          5663 => x"38",
          5664 => x"51",
          5665 => x"3f",
          5666 => x"fd",
          5667 => x"fe",
          5668 => x"fe",
          5669 => x"81",
          5670 => x"b8",
          5671 => x"05",
          5672 => x"eb",
          5673 => x"53",
          5674 => x"08",
          5675 => x"f5",
          5676 => x"d5",
          5677 => x"fe",
          5678 => x"fe",
          5679 => x"81",
          5680 => x"b8",
          5681 => x"05",
          5682 => x"ea",
          5683 => x"d3",
          5684 => x"3d",
          5685 => x"52",
          5686 => x"d7",
          5687 => x"84",
          5688 => x"fe",
          5689 => x"59",
          5690 => x"3f",
          5691 => x"58",
          5692 => x"57",
          5693 => x"55",
          5694 => x"08",
          5695 => x"54",
          5696 => x"52",
          5697 => x"f0",
          5698 => x"84",
          5699 => x"fa",
          5700 => x"d3",
          5701 => x"f0",
          5702 => x"ed",
          5703 => x"fe",
          5704 => x"fe",
          5705 => x"ff",
          5706 => x"81",
          5707 => x"80",
          5708 => x"38",
          5709 => x"f0",
          5710 => x"f8",
          5711 => x"80",
          5712 => x"d3",
          5713 => x"2e",
          5714 => x"b7",
          5715 => x"11",
          5716 => x"05",
          5717 => x"ba",
          5718 => x"84",
          5719 => x"81",
          5720 => x"42",
          5721 => x"51",
          5722 => x"3f",
          5723 => x"5a",
          5724 => x"8f",
          5725 => x"78",
          5726 => x"05",
          5727 => x"7a",
          5728 => x"81",
          5729 => x"86",
          5730 => x"3d",
          5731 => x"53",
          5732 => x"51",
          5733 => x"3f",
          5734 => x"08",
          5735 => x"81",
          5736 => x"59",
          5737 => x"88",
          5738 => x"80",
          5739 => x"39",
          5740 => x"33",
          5741 => x"2e",
          5742 => x"d0",
          5743 => x"a2",
          5744 => x"af",
          5745 => x"8b",
          5746 => x"b0",
          5747 => x"80",
          5748 => x"81",
          5749 => x"44",
          5750 => x"d0",
          5751 => x"80",
          5752 => x"3d",
          5753 => x"53",
          5754 => x"51",
          5755 => x"3f",
          5756 => x"08",
          5757 => x"81",
          5758 => x"59",
          5759 => x"88",
          5760 => x"84",
          5761 => x"39",
          5762 => x"33",
          5763 => x"2e",
          5764 => x"d0",
          5765 => x"a1",
          5766 => x"af",
          5767 => x"8b",
          5768 => x"b0",
          5769 => x"80",
          5770 => x"81",
          5771 => x"43",
          5772 => x"d0",
          5773 => x"05",
          5774 => x"fe",
          5775 => x"fe",
          5776 => x"fe",
          5777 => x"81",
          5778 => x"80",
          5779 => x"80",
          5780 => x"79",
          5781 => x"38",
          5782 => x"90",
          5783 => x"78",
          5784 => x"38",
          5785 => x"83",
          5786 => x"81",
          5787 => x"fe",
          5788 => x"a0",
          5789 => x"61",
          5790 => x"63",
          5791 => x"3f",
          5792 => x"51",
          5793 => x"b7",
          5794 => x"11",
          5795 => x"05",
          5796 => x"fe",
          5797 => x"84",
          5798 => x"f7",
          5799 => x"3d",
          5800 => x"53",
          5801 => x"51",
          5802 => x"3f",
          5803 => x"08",
          5804 => x"38",
          5805 => x"80",
          5806 => x"79",
          5807 => x"05",
          5808 => x"fe",
          5809 => x"fe",
          5810 => x"fe",
          5811 => x"81",
          5812 => x"e0",
          5813 => x"39",
          5814 => x"54",
          5815 => x"a8",
          5816 => x"b9",
          5817 => x"52",
          5818 => x"fc",
          5819 => x"45",
          5820 => x"78",
          5821 => x"91",
          5822 => x"27",
          5823 => x"3d",
          5824 => x"53",
          5825 => x"51",
          5826 => x"3f",
          5827 => x"08",
          5828 => x"38",
          5829 => x"80",
          5830 => x"79",
          5831 => x"05",
          5832 => x"39",
          5833 => x"51",
          5834 => x"3f",
          5835 => x"b7",
          5836 => x"11",
          5837 => x"05",
          5838 => x"c8",
          5839 => x"84",
          5840 => x"f6",
          5841 => x"3d",
          5842 => x"53",
          5843 => x"51",
          5844 => x"3f",
          5845 => x"08",
          5846 => x"38",
          5847 => x"be",
          5848 => x"70",
          5849 => x"23",
          5850 => x"3d",
          5851 => x"53",
          5852 => x"51",
          5853 => x"3f",
          5854 => x"08",
          5855 => x"89",
          5856 => x"22",
          5857 => x"cd",
          5858 => x"fa",
          5859 => x"f8",
          5860 => x"fe",
          5861 => x"79",
          5862 => x"59",
          5863 => x"f5",
          5864 => x"9f",
          5865 => x"60",
          5866 => x"d5",
          5867 => x"fe",
          5868 => x"fe",
          5869 => x"fe",
          5870 => x"81",
          5871 => x"80",
          5872 => x"60",
          5873 => x"05",
          5874 => x"82",
          5875 => x"78",
          5876 => x"39",
          5877 => x"51",
          5878 => x"3f",
          5879 => x"b7",
          5880 => x"11",
          5881 => x"05",
          5882 => x"98",
          5883 => x"84",
          5884 => x"f5",
          5885 => x"3d",
          5886 => x"53",
          5887 => x"51",
          5888 => x"3f",
          5889 => x"08",
          5890 => x"38",
          5891 => x"0c",
          5892 => x"05",
          5893 => x"fe",
          5894 => x"fe",
          5895 => x"fe",
          5896 => x"81",
          5897 => x"e4",
          5898 => x"39",
          5899 => x"54",
          5900 => x"c8",
          5901 => x"e5",
          5902 => x"52",
          5903 => x"f9",
          5904 => x"45",
          5905 => x"78",
          5906 => x"bd",
          5907 => x"27",
          5908 => x"3d",
          5909 => x"53",
          5910 => x"51",
          5911 => x"3f",
          5912 => x"08",
          5913 => x"38",
          5914 => x"52",
          5915 => x"51",
          5916 => x"3f",
          5917 => x"0c",
          5918 => x"05",
          5919 => x"39",
          5920 => x"51",
          5921 => x"3f",
          5922 => x"81",
          5923 => x"fe",
          5924 => x"82",
          5925 => x"95",
          5926 => x"39",
          5927 => x"51",
          5928 => x"3f",
          5929 => x"f0",
          5930 => x"dd",
          5931 => x"81",
          5932 => x"94",
          5933 => x"80",
          5934 => x"c0",
          5935 => x"81",
          5936 => x"fe",
          5937 => x"f3",
          5938 => x"ce",
          5939 => x"f1",
          5940 => x"80",
          5941 => x"c0",
          5942 => x"8c",
          5943 => x"87",
          5944 => x"0c",
          5945 => x"b7",
          5946 => x"11",
          5947 => x"05",
          5948 => x"9e",
          5949 => x"84",
          5950 => x"f3",
          5951 => x"52",
          5952 => x"51",
          5953 => x"3f",
          5954 => x"04",
          5955 => x"f4",
          5956 => x"f8",
          5957 => x"f8",
          5958 => x"d3",
          5959 => x"2e",
          5960 => x"63",
          5961 => x"c8",
          5962 => x"f1",
          5963 => x"78",
          5964 => x"84",
          5965 => x"d3",
          5966 => x"2e",
          5967 => x"81",
          5968 => x"52",
          5969 => x"51",
          5970 => x"3f",
          5971 => x"81",
          5972 => x"fe",
          5973 => x"fe",
          5974 => x"f2",
          5975 => x"cf",
          5976 => x"f0",
          5977 => x"59",
          5978 => x"fe",
          5979 => x"f2",
          5980 => x"70",
          5981 => x"78",
          5982 => x"8d",
          5983 => x"2e",
          5984 => x"7c",
          5985 => x"cc",
          5986 => x"fe",
          5987 => x"fe",
          5988 => x"81",
          5989 => x"81",
          5990 => x"55",
          5991 => x"54",
          5992 => x"cf",
          5993 => x"3d",
          5994 => x"fe",
          5995 => x"81",
          5996 => x"81",
          5997 => x"80",
          5998 => x"11",
          5999 => x"55",
          6000 => x"a0",
          6001 => x"a0",
          6002 => x"51",
          6003 => x"81",
          6004 => x"5e",
          6005 => x"7c",
          6006 => x"59",
          6007 => x"7d",
          6008 => x"81",
          6009 => x"38",
          6010 => x"51",
          6011 => x"3f",
          6012 => x"80",
          6013 => x"0b",
          6014 => x"34",
          6015 => x"e4",
          6016 => x"94",
          6017 => x"90",
          6018 => x"87",
          6019 => x"0c",
          6020 => x"0b",
          6021 => x"84",
          6022 => x"83",
          6023 => x"94",
          6024 => x"ba",
          6025 => x"94",
          6026 => x"0b",
          6027 => x"0c",
          6028 => x"3f",
          6029 => x"3f",
          6030 => x"51",
          6031 => x"3f",
          6032 => x"51",
          6033 => x"3f",
          6034 => x"51",
          6035 => x"3f",
          6036 => x"ed",
          6037 => x"3f",
          6038 => x"00",
          6039 => x"ff",
          6040 => x"ff",
          6041 => x"ff",
          6042 => x"00",
          6043 => x"db",
          6044 => x"e1",
          6045 => x"e7",
          6046 => x"ed",
          6047 => x"f3",
          6048 => x"b1",
          6049 => x"35",
          6050 => x"3c",
          6051 => x"43",
          6052 => x"4a",
          6053 => x"51",
          6054 => x"58",
          6055 => x"5f",
          6056 => x"66",
          6057 => x"6d",
          6058 => x"74",
          6059 => x"7b",
          6060 => x"81",
          6061 => x"87",
          6062 => x"8d",
          6063 => x"93",
          6064 => x"99",
          6065 => x"9f",
          6066 => x"a5",
          6067 => x"ab",
          6068 => x"25",
          6069 => x"64",
          6070 => x"3a",
          6071 => x"25",
          6072 => x"64",
          6073 => x"00",
          6074 => x"20",
          6075 => x"66",
          6076 => x"72",
          6077 => x"6f",
          6078 => x"00",
          6079 => x"72",
          6080 => x"53",
          6081 => x"63",
          6082 => x"69",
          6083 => x"00",
          6084 => x"65",
          6085 => x"65",
          6086 => x"6d",
          6087 => x"6d",
          6088 => x"65",
          6089 => x"00",
          6090 => x"20",
          6091 => x"4e",
          6092 => x"41",
          6093 => x"53",
          6094 => x"74",
          6095 => x"38",
          6096 => x"53",
          6097 => x"3d",
          6098 => x"58",
          6099 => x"00",
          6100 => x"20",
          6101 => x"4d",
          6102 => x"74",
          6103 => x"3d",
          6104 => x"58",
          6105 => x"69",
          6106 => x"25",
          6107 => x"29",
          6108 => x"00",
          6109 => x"20",
          6110 => x"20",
          6111 => x"61",
          6112 => x"25",
          6113 => x"2c",
          6114 => x"7a",
          6115 => x"30",
          6116 => x"2e",
          6117 => x"00",
          6118 => x"20",
          6119 => x"54",
          6120 => x"00",
          6121 => x"20",
          6122 => x"0a",
          6123 => x"00",
          6124 => x"20",
          6125 => x"0a",
          6126 => x"00",
          6127 => x"20",
          6128 => x"43",
          6129 => x"20",
          6130 => x"76",
          6131 => x"73",
          6132 => x"32",
          6133 => x"0a",
          6134 => x"00",
          6135 => x"20",
          6136 => x"45",
          6137 => x"50",
          6138 => x"4f",
          6139 => x"4f",
          6140 => x"52",
          6141 => x"00",
          6142 => x"20",
          6143 => x"45",
          6144 => x"28",
          6145 => x"65",
          6146 => x"25",
          6147 => x"29",
          6148 => x"00",
          6149 => x"72",
          6150 => x"65",
          6151 => x"00",
          6152 => x"20",
          6153 => x"20",
          6154 => x"65",
          6155 => x"65",
          6156 => x"72",
          6157 => x"64",
          6158 => x"73",
          6159 => x"25",
          6160 => x"0a",
          6161 => x"00",
          6162 => x"20",
          6163 => x"20",
          6164 => x"6f",
          6165 => x"53",
          6166 => x"74",
          6167 => x"64",
          6168 => x"73",
          6169 => x"25",
          6170 => x"0a",
          6171 => x"00",
          6172 => x"20",
          6173 => x"63",
          6174 => x"74",
          6175 => x"20",
          6176 => x"72",
          6177 => x"20",
          6178 => x"20",
          6179 => x"25",
          6180 => x"0a",
          6181 => x"00",
          6182 => x"20",
          6183 => x"20",
          6184 => x"20",
          6185 => x"20",
          6186 => x"20",
          6187 => x"20",
          6188 => x"20",
          6189 => x"25",
          6190 => x"0a",
          6191 => x"00",
          6192 => x"20",
          6193 => x"74",
          6194 => x"43",
          6195 => x"6b",
          6196 => x"65",
          6197 => x"20",
          6198 => x"20",
          6199 => x"25",
          6200 => x"0a",
          6201 => x"00",
          6202 => x"6c",
          6203 => x"00",
          6204 => x"69",
          6205 => x"00",
          6206 => x"78",
          6207 => x"00",
          6208 => x"00",
          6209 => x"6d",
          6210 => x"00",
          6211 => x"6e",
          6212 => x"00",
          6213 => x"00",
          6214 => x"2c",
          6215 => x"3d",
          6216 => x"5d",
          6217 => x"00",
          6218 => x"00",
          6219 => x"33",
          6220 => x"00",
          6221 => x"4d",
          6222 => x"53",
          6223 => x"00",
          6224 => x"4e",
          6225 => x"20",
          6226 => x"46",
          6227 => x"32",
          6228 => x"00",
          6229 => x"4e",
          6230 => x"20",
          6231 => x"46",
          6232 => x"20",
          6233 => x"00",
          6234 => x"14",
          6235 => x"00",
          6236 => x"00",
          6237 => x"00",
          6238 => x"41",
          6239 => x"80",
          6240 => x"49",
          6241 => x"8f",
          6242 => x"4f",
          6243 => x"55",
          6244 => x"9b",
          6245 => x"9f",
          6246 => x"55",
          6247 => x"a7",
          6248 => x"ab",
          6249 => x"af",
          6250 => x"b3",
          6251 => x"b7",
          6252 => x"bb",
          6253 => x"bf",
          6254 => x"c3",
          6255 => x"c7",
          6256 => x"cb",
          6257 => x"cf",
          6258 => x"d3",
          6259 => x"d7",
          6260 => x"db",
          6261 => x"df",
          6262 => x"e3",
          6263 => x"e7",
          6264 => x"eb",
          6265 => x"ef",
          6266 => x"f3",
          6267 => x"f7",
          6268 => x"fb",
          6269 => x"ff",
          6270 => x"3b",
          6271 => x"2f",
          6272 => x"3a",
          6273 => x"7c",
          6274 => x"00",
          6275 => x"04",
          6276 => x"40",
          6277 => x"00",
          6278 => x"00",
          6279 => x"02",
          6280 => x"08",
          6281 => x"20",
          6282 => x"00",
          6283 => x"69",
          6284 => x"00",
          6285 => x"63",
          6286 => x"00",
          6287 => x"69",
          6288 => x"00",
          6289 => x"61",
          6290 => x"00",
          6291 => x"65",
          6292 => x"00",
          6293 => x"65",
          6294 => x"00",
          6295 => x"6d",
          6296 => x"00",
          6297 => x"00",
          6298 => x"00",
          6299 => x"00",
          6300 => x"00",
          6301 => x"00",
          6302 => x"00",
          6303 => x"00",
          6304 => x"6c",
          6305 => x"00",
          6306 => x"00",
          6307 => x"74",
          6308 => x"00",
          6309 => x"65",
          6310 => x"00",
          6311 => x"6f",
          6312 => x"00",
          6313 => x"74",
          6314 => x"00",
          6315 => x"6b",
          6316 => x"72",
          6317 => x"00",
          6318 => x"65",
          6319 => x"6c",
          6320 => x"72",
          6321 => x"0a",
          6322 => x"00",
          6323 => x"6b",
          6324 => x"74",
          6325 => x"61",
          6326 => x"0a",
          6327 => x"00",
          6328 => x"66",
          6329 => x"20",
          6330 => x"6e",
          6331 => x"00",
          6332 => x"70",
          6333 => x"20",
          6334 => x"6e",
          6335 => x"00",
          6336 => x"61",
          6337 => x"20",
          6338 => x"65",
          6339 => x"65",
          6340 => x"00",
          6341 => x"65",
          6342 => x"64",
          6343 => x"65",
          6344 => x"00",
          6345 => x"65",
          6346 => x"72",
          6347 => x"79",
          6348 => x"69",
          6349 => x"2e",
          6350 => x"00",
          6351 => x"65",
          6352 => x"6e",
          6353 => x"20",
          6354 => x"61",
          6355 => x"2e",
          6356 => x"00",
          6357 => x"69",
          6358 => x"72",
          6359 => x"20",
          6360 => x"74",
          6361 => x"65",
          6362 => x"00",
          6363 => x"76",
          6364 => x"75",
          6365 => x"72",
          6366 => x"20",
          6367 => x"61",
          6368 => x"2e",
          6369 => x"00",
          6370 => x"6b",
          6371 => x"74",
          6372 => x"61",
          6373 => x"64",
          6374 => x"00",
          6375 => x"63",
          6376 => x"61",
          6377 => x"6c",
          6378 => x"69",
          6379 => x"79",
          6380 => x"6d",
          6381 => x"75",
          6382 => x"6f",
          6383 => x"69",
          6384 => x"0a",
          6385 => x"00",
          6386 => x"6d",
          6387 => x"61",
          6388 => x"74",
          6389 => x"0a",
          6390 => x"00",
          6391 => x"65",
          6392 => x"2c",
          6393 => x"65",
          6394 => x"69",
          6395 => x"63",
          6396 => x"65",
          6397 => x"64",
          6398 => x"00",
          6399 => x"65",
          6400 => x"20",
          6401 => x"6b",
          6402 => x"0a",
          6403 => x"00",
          6404 => x"75",
          6405 => x"63",
          6406 => x"74",
          6407 => x"6d",
          6408 => x"2e",
          6409 => x"00",
          6410 => x"20",
          6411 => x"79",
          6412 => x"65",
          6413 => x"69",
          6414 => x"2e",
          6415 => x"00",
          6416 => x"61",
          6417 => x"65",
          6418 => x"69",
          6419 => x"72",
          6420 => x"74",
          6421 => x"00",
          6422 => x"63",
          6423 => x"2e",
          6424 => x"00",
          6425 => x"6e",
          6426 => x"20",
          6427 => x"6f",
          6428 => x"00",
          6429 => x"75",
          6430 => x"74",
          6431 => x"25",
          6432 => x"74",
          6433 => x"75",
          6434 => x"74",
          6435 => x"73",
          6436 => x"0a",
          6437 => x"00",
          6438 => x"58",
          6439 => x"00",
          6440 => x"00",
          6441 => x"58",
          6442 => x"00",
          6443 => x"20",
          6444 => x"20",
          6445 => x"00",
          6446 => x"58",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"00",
          6451 => x"64",
          6452 => x"00",
          6453 => x"54",
          6454 => x"00",
          6455 => x"20",
          6456 => x"28",
          6457 => x"00",
          6458 => x"30",
          6459 => x"30",
          6460 => x"00",
          6461 => x"33",
          6462 => x"00",
          6463 => x"55",
          6464 => x"65",
          6465 => x"30",
          6466 => x"20",
          6467 => x"25",
          6468 => x"2a",
          6469 => x"00",
          6470 => x"54",
          6471 => x"6e",
          6472 => x"72",
          6473 => x"20",
          6474 => x"64",
          6475 => x"0a",
          6476 => x"00",
          6477 => x"65",
          6478 => x"6e",
          6479 => x"72",
          6480 => x"0a",
          6481 => x"00",
          6482 => x"20",
          6483 => x"65",
          6484 => x"70",
          6485 => x"00",
          6486 => x"54",
          6487 => x"44",
          6488 => x"74",
          6489 => x"75",
          6490 => x"00",
          6491 => x"54",
          6492 => x"52",
          6493 => x"74",
          6494 => x"75",
          6495 => x"00",
          6496 => x"54",
          6497 => x"58",
          6498 => x"74",
          6499 => x"75",
          6500 => x"00",
          6501 => x"54",
          6502 => x"58",
          6503 => x"74",
          6504 => x"75",
          6505 => x"00",
          6506 => x"54",
          6507 => x"58",
          6508 => x"74",
          6509 => x"75",
          6510 => x"00",
          6511 => x"54",
          6512 => x"58",
          6513 => x"74",
          6514 => x"75",
          6515 => x"00",
          6516 => x"74",
          6517 => x"20",
          6518 => x"74",
          6519 => x"72",
          6520 => x"0a",
          6521 => x"00",
          6522 => x"62",
          6523 => x"67",
          6524 => x"6d",
          6525 => x"2e",
          6526 => x"00",
          6527 => x"00",
          6528 => x"6c",
          6529 => x"74",
          6530 => x"6e",
          6531 => x"61",
          6532 => x"65",
          6533 => x"20",
          6534 => x"64",
          6535 => x"20",
          6536 => x"61",
          6537 => x"69",
          6538 => x"20",
          6539 => x"75",
          6540 => x"79",
          6541 => x"00",
          6542 => x"00",
          6543 => x"20",
          6544 => x"6b",
          6545 => x"21",
          6546 => x"00",
          6547 => x"74",
          6548 => x"69",
          6549 => x"2e",
          6550 => x"00",
          6551 => x"6c",
          6552 => x"74",
          6553 => x"6e",
          6554 => x"61",
          6555 => x"65",
          6556 => x"00",
          6557 => x"25",
          6558 => x"00",
          6559 => x"00",
          6560 => x"61",
          6561 => x"67",
          6562 => x"00",
          6563 => x"70",
          6564 => x"6d",
          6565 => x"0a",
          6566 => x"00",
          6567 => x"6d",
          6568 => x"74",
          6569 => x"00",
          6570 => x"58",
          6571 => x"32",
          6572 => x"00",
          6573 => x"0a",
          6574 => x"00",
          6575 => x"58",
          6576 => x"34",
          6577 => x"00",
          6578 => x"58",
          6579 => x"38",
          6580 => x"00",
          6581 => x"61",
          6582 => x"6e",
          6583 => x"6e",
          6584 => x"72",
          6585 => x"73",
          6586 => x"00",
          6587 => x"62",
          6588 => x"67",
          6589 => x"74",
          6590 => x"75",
          6591 => x"0a",
          6592 => x"00",
          6593 => x"61",
          6594 => x"64",
          6595 => x"72",
          6596 => x"69",
          6597 => x"00",
          6598 => x"62",
          6599 => x"67",
          6600 => x"72",
          6601 => x"69",
          6602 => x"00",
          6603 => x"63",
          6604 => x"6e",
          6605 => x"6f",
          6606 => x"40",
          6607 => x"38",
          6608 => x"2e",
          6609 => x"00",
          6610 => x"6c",
          6611 => x"20",
          6612 => x"65",
          6613 => x"25",
          6614 => x"20",
          6615 => x"0a",
          6616 => x"00",
          6617 => x"6c",
          6618 => x"74",
          6619 => x"65",
          6620 => x"6f",
          6621 => x"28",
          6622 => x"2e",
          6623 => x"00",
          6624 => x"74",
          6625 => x"69",
          6626 => x"61",
          6627 => x"69",
          6628 => x"69",
          6629 => x"2e",
          6630 => x"00",
          6631 => x"64",
          6632 => x"62",
          6633 => x"69",
          6634 => x"2e",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"5c",
          6639 => x"25",
          6640 => x"73",
          6641 => x"00",
          6642 => x"20",
          6643 => x"6d",
          6644 => x"2e",
          6645 => x"00",
          6646 => x"6e",
          6647 => x"2e",
          6648 => x"00",
          6649 => x"62",
          6650 => x"67",
          6651 => x"74",
          6652 => x"75",
          6653 => x"2e",
          6654 => x"00",
          6655 => x"00",
          6656 => x"00",
          6657 => x"ff",
          6658 => x"00",
          6659 => x"ff",
          6660 => x"00",
          6661 => x"ff",
          6662 => x"00",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"00",
          6667 => x"01",
          6668 => x"01",
          6669 => x"01",
          6670 => x"00",
          6671 => x"00",
          6672 => x"00",
          6673 => x"2c",
          6674 => x"00",
          6675 => x"00",
          6676 => x"00",
          6677 => x"34",
          6678 => x"00",
          6679 => x"00",
          6680 => x"00",
          6681 => x"3c",
          6682 => x"00",
          6683 => x"00",
          6684 => x"00",
          6685 => x"44",
          6686 => x"00",
          6687 => x"00",
          6688 => x"00",
          6689 => x"4c",
          6690 => x"00",
          6691 => x"00",
          6692 => x"00",
          6693 => x"54",
          6694 => x"00",
          6695 => x"00",
          6696 => x"00",
          6697 => x"5c",
          6698 => x"00",
          6699 => x"00",
          6700 => x"00",
          6701 => x"64",
          6702 => x"00",
          6703 => x"00",
          6704 => x"00",
          6705 => x"68",
          6706 => x"00",
          6707 => x"00",
          6708 => x"00",
          6709 => x"6c",
          6710 => x"00",
          6711 => x"00",
          6712 => x"00",
          6713 => x"70",
          6714 => x"00",
          6715 => x"00",
          6716 => x"00",
          6717 => x"74",
          6718 => x"00",
          6719 => x"00",
          6720 => x"00",
          6721 => x"78",
          6722 => x"00",
          6723 => x"00",
          6724 => x"00",
          6725 => x"7c",
          6726 => x"00",
          6727 => x"00",
          6728 => x"00",
          6729 => x"80",
          6730 => x"00",
          6731 => x"00",
          6732 => x"00",
          6733 => x"88",
          6734 => x"00",
          6735 => x"00",
          6736 => x"00",
          6737 => x"8c",
          6738 => x"00",
          6739 => x"00",
          6740 => x"00",
          6741 => x"94",
          6742 => x"00",
          6743 => x"00",
          6744 => x"00",
          6745 => x"9c",
          6746 => x"00",
          6747 => x"00",
          6748 => x"00",
          6749 => x"a4",
          6750 => x"00",
          6751 => x"00",
          6752 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"92",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"81",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a3",
           270 => x"0b",
           271 => x"0b",
           272 => x"c1",
           273 => x"0b",
           274 => x"0b",
           275 => x"df",
           276 => x"0b",
           277 => x"0b",
           278 => x"fd",
           279 => x"0b",
           280 => x"0b",
           281 => x"9b",
           282 => x"0b",
           283 => x"0b",
           284 => x"b9",
           285 => x"0b",
           286 => x"0b",
           287 => x"d7",
           288 => x"0b",
           289 => x"0b",
           290 => x"f5",
           291 => x"0b",
           292 => x"0b",
           293 => x"94",
           294 => x"0b",
           295 => x"0b",
           296 => x"b4",
           297 => x"0b",
           298 => x"0b",
           299 => x"d4",
           300 => x"0b",
           301 => x"0b",
           302 => x"f4",
           303 => x"0b",
           304 => x"0b",
           305 => x"94",
           306 => x"0b",
           307 => x"0b",
           308 => x"b4",
           309 => x"0b",
           310 => x"0b",
           311 => x"d4",
           312 => x"0b",
           313 => x"0b",
           314 => x"f4",
           315 => x"0b",
           316 => x"0b",
           317 => x"94",
           318 => x"0b",
           319 => x"0b",
           320 => x"b4",
           321 => x"0b",
           322 => x"0b",
           323 => x"d4",
           324 => x"0b",
           325 => x"0b",
           326 => x"f4",
           327 => x"0b",
           328 => x"0b",
           329 => x"94",
           330 => x"0b",
           331 => x"0b",
           332 => x"b2",
           333 => x"0b",
           334 => x"0b",
           335 => x"d0",
           336 => x"0b",
           337 => x"0b",
           338 => x"ee",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"d3",
           386 => x"ae",
           387 => x"90",
           388 => x"90",
           389 => x"90",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"81",
           395 => x"82",
           396 => x"81",
           397 => x"ab",
           398 => x"d3",
           399 => x"a0",
           400 => x"d3",
           401 => x"f7",
           402 => x"90",
           403 => x"90",
           404 => x"90",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"81",
           410 => x"82",
           411 => x"81",
           412 => x"b3",
           413 => x"d3",
           414 => x"a0",
           415 => x"d3",
           416 => x"84",
           417 => x"90",
           418 => x"90",
           419 => x"90",
           420 => x"2d",
           421 => x"08",
           422 => x"04",
           423 => x"0c",
           424 => x"81",
           425 => x"82",
           426 => x"81",
           427 => x"b1",
           428 => x"d3",
           429 => x"a0",
           430 => x"d3",
           431 => x"bb",
           432 => x"90",
           433 => x"90",
           434 => x"90",
           435 => x"2d",
           436 => x"08",
           437 => x"04",
           438 => x"0c",
           439 => x"81",
           440 => x"82",
           441 => x"81",
           442 => x"9c",
           443 => x"d3",
           444 => x"a0",
           445 => x"d3",
           446 => x"90",
           447 => x"90",
           448 => x"90",
           449 => x"90",
           450 => x"b9",
           451 => x"90",
           452 => x"90",
           453 => x"90",
           454 => x"aa",
           455 => x"90",
           456 => x"90",
           457 => x"90",
           458 => x"9e",
           459 => x"90",
           460 => x"90",
           461 => x"90",
           462 => x"9b",
           463 => x"90",
           464 => x"90",
           465 => x"90",
           466 => x"b9",
           467 => x"90",
           468 => x"90",
           469 => x"90",
           470 => x"99",
           471 => x"90",
           472 => x"90",
           473 => x"90",
           474 => x"8c",
           475 => x"90",
           476 => x"90",
           477 => x"90",
           478 => x"d8",
           479 => x"90",
           480 => x"90",
           481 => x"90",
           482 => x"f7",
           483 => x"90",
           484 => x"90",
           485 => x"90",
           486 => x"96",
           487 => x"90",
           488 => x"90",
           489 => x"90",
           490 => x"80",
           491 => x"90",
           492 => x"90",
           493 => x"90",
           494 => x"e6",
           495 => x"90",
           496 => x"90",
           497 => x"90",
           498 => x"d4",
           499 => x"90",
           500 => x"90",
           501 => x"90",
           502 => x"9a",
           503 => x"90",
           504 => x"90",
           505 => x"90",
           506 => x"d4",
           507 => x"90",
           508 => x"90",
           509 => x"90",
           510 => x"d5",
           511 => x"90",
           512 => x"90",
           513 => x"90",
           514 => x"8a",
           515 => x"90",
           516 => x"90",
           517 => x"90",
           518 => x"e3",
           519 => x"90",
           520 => x"90",
           521 => x"90",
           522 => x"8e",
           523 => x"90",
           524 => x"90",
           525 => x"90",
           526 => x"f1",
           527 => x"90",
           528 => x"90",
           529 => x"90",
           530 => x"c6",
           531 => x"90",
           532 => x"90",
           533 => x"90",
           534 => x"d0",
           535 => x"90",
           536 => x"90",
           537 => x"90",
           538 => x"92",
           539 => x"90",
           540 => x"90",
           541 => x"90",
           542 => x"d8",
           543 => x"90",
           544 => x"90",
           545 => x"90",
           546 => x"fe",
           547 => x"90",
           548 => x"90",
           549 => x"90",
           550 => x"2d",
           551 => x"08",
           552 => x"04",
           553 => x"0c",
           554 => x"81",
           555 => x"82",
           556 => x"81",
           557 => x"bb",
           558 => x"d3",
           559 => x"a0",
           560 => x"d3",
           561 => x"d1",
           562 => x"90",
           563 => x"90",
           564 => x"90",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"81",
           570 => x"82",
           571 => x"81",
           572 => x"81",
           573 => x"81",
           574 => x"82",
           575 => x"3c",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"00",
           585 => x"ff",
           586 => x"06",
           587 => x"83",
           588 => x"10",
           589 => x"fc",
           590 => x"51",
           591 => x"80",
           592 => x"ff",
           593 => x"06",
           594 => x"52",
           595 => x"0a",
           596 => x"38",
           597 => x"51",
           598 => x"84",
           599 => x"88",
           600 => x"80",
           601 => x"05",
           602 => x"0b",
           603 => x"04",
           604 => x"81",
           605 => x"00",
           606 => x"08",
           607 => x"90",
           608 => x"0d",
           609 => x"d3",
           610 => x"05",
           611 => x"d3",
           612 => x"05",
           613 => x"d4",
           614 => x"84",
           615 => x"d3",
           616 => x"85",
           617 => x"d3",
           618 => x"81",
           619 => x"02",
           620 => x"0c",
           621 => x"81",
           622 => x"90",
           623 => x"08",
           624 => x"90",
           625 => x"08",
           626 => x"3f",
           627 => x"08",
           628 => x"84",
           629 => x"3d",
           630 => x"90",
           631 => x"d3",
           632 => x"81",
           633 => x"f9",
           634 => x"0b",
           635 => x"08",
           636 => x"81",
           637 => x"88",
           638 => x"25",
           639 => x"d3",
           640 => x"05",
           641 => x"d3",
           642 => x"05",
           643 => x"81",
           644 => x"f4",
           645 => x"d3",
           646 => x"05",
           647 => x"81",
           648 => x"90",
           649 => x"0c",
           650 => x"08",
           651 => x"81",
           652 => x"fc",
           653 => x"d3",
           654 => x"05",
           655 => x"b9",
           656 => x"90",
           657 => x"08",
           658 => x"90",
           659 => x"0c",
           660 => x"d3",
           661 => x"05",
           662 => x"90",
           663 => x"08",
           664 => x"0b",
           665 => x"08",
           666 => x"81",
           667 => x"f0",
           668 => x"d3",
           669 => x"05",
           670 => x"81",
           671 => x"8c",
           672 => x"81",
           673 => x"88",
           674 => x"81",
           675 => x"d3",
           676 => x"81",
           677 => x"f8",
           678 => x"81",
           679 => x"fc",
           680 => x"2e",
           681 => x"d3",
           682 => x"05",
           683 => x"d3",
           684 => x"05",
           685 => x"90",
           686 => x"08",
           687 => x"84",
           688 => x"3d",
           689 => x"90",
           690 => x"d3",
           691 => x"81",
           692 => x"fb",
           693 => x"0b",
           694 => x"08",
           695 => x"81",
           696 => x"88",
           697 => x"25",
           698 => x"d3",
           699 => x"05",
           700 => x"d3",
           701 => x"05",
           702 => x"81",
           703 => x"fc",
           704 => x"d3",
           705 => x"05",
           706 => x"90",
           707 => x"90",
           708 => x"08",
           709 => x"90",
           710 => x"0c",
           711 => x"d3",
           712 => x"05",
           713 => x"d3",
           714 => x"05",
           715 => x"3f",
           716 => x"08",
           717 => x"90",
           718 => x"0c",
           719 => x"90",
           720 => x"08",
           721 => x"38",
           722 => x"08",
           723 => x"30",
           724 => x"08",
           725 => x"81",
           726 => x"f8",
           727 => x"81",
           728 => x"54",
           729 => x"81",
           730 => x"04",
           731 => x"08",
           732 => x"90",
           733 => x"0d",
           734 => x"d3",
           735 => x"05",
           736 => x"81",
           737 => x"f8",
           738 => x"d3",
           739 => x"05",
           740 => x"90",
           741 => x"08",
           742 => x"81",
           743 => x"fc",
           744 => x"2e",
           745 => x"0b",
           746 => x"08",
           747 => x"24",
           748 => x"d3",
           749 => x"05",
           750 => x"d3",
           751 => x"05",
           752 => x"90",
           753 => x"08",
           754 => x"90",
           755 => x"0c",
           756 => x"81",
           757 => x"fc",
           758 => x"2e",
           759 => x"81",
           760 => x"8c",
           761 => x"d3",
           762 => x"05",
           763 => x"38",
           764 => x"08",
           765 => x"81",
           766 => x"8c",
           767 => x"81",
           768 => x"88",
           769 => x"d3",
           770 => x"05",
           771 => x"90",
           772 => x"08",
           773 => x"90",
           774 => x"0c",
           775 => x"08",
           776 => x"81",
           777 => x"90",
           778 => x"0c",
           779 => x"08",
           780 => x"81",
           781 => x"90",
           782 => x"0c",
           783 => x"81",
           784 => x"90",
           785 => x"2e",
           786 => x"d3",
           787 => x"05",
           788 => x"d3",
           789 => x"05",
           790 => x"39",
           791 => x"08",
           792 => x"70",
           793 => x"08",
           794 => x"51",
           795 => x"08",
           796 => x"81",
           797 => x"85",
           798 => x"d3",
           799 => x"fc",
           800 => x"79",
           801 => x"05",
           802 => x"57",
           803 => x"83",
           804 => x"38",
           805 => x"51",
           806 => x"a4",
           807 => x"52",
           808 => x"93",
           809 => x"70",
           810 => x"34",
           811 => x"71",
           812 => x"81",
           813 => x"74",
           814 => x"0c",
           815 => x"04",
           816 => x"2b",
           817 => x"71",
           818 => x"51",
           819 => x"72",
           820 => x"72",
           821 => x"05",
           822 => x"71",
           823 => x"53",
           824 => x"70",
           825 => x"0c",
           826 => x"84",
           827 => x"f0",
           828 => x"8f",
           829 => x"83",
           830 => x"38",
           831 => x"84",
           832 => x"fc",
           833 => x"83",
           834 => x"70",
           835 => x"39",
           836 => x"77",
           837 => x"07",
           838 => x"54",
           839 => x"38",
           840 => x"08",
           841 => x"71",
           842 => x"80",
           843 => x"75",
           844 => x"33",
           845 => x"06",
           846 => x"80",
           847 => x"72",
           848 => x"75",
           849 => x"06",
           850 => x"12",
           851 => x"33",
           852 => x"06",
           853 => x"52",
           854 => x"72",
           855 => x"81",
           856 => x"81",
           857 => x"71",
           858 => x"84",
           859 => x"87",
           860 => x"71",
           861 => x"fb",
           862 => x"06",
           863 => x"82",
           864 => x"51",
           865 => x"97",
           866 => x"84",
           867 => x"54",
           868 => x"75",
           869 => x"38",
           870 => x"52",
           871 => x"80",
           872 => x"84",
           873 => x"0d",
           874 => x"0d",
           875 => x"53",
           876 => x"52",
           877 => x"81",
           878 => x"81",
           879 => x"07",
           880 => x"52",
           881 => x"e8",
           882 => x"d3",
           883 => x"3d",
           884 => x"3d",
           885 => x"08",
           886 => x"56",
           887 => x"80",
           888 => x"33",
           889 => x"2e",
           890 => x"86",
           891 => x"52",
           892 => x"53",
           893 => x"13",
           894 => x"33",
           895 => x"06",
           896 => x"70",
           897 => x"38",
           898 => x"80",
           899 => x"74",
           900 => x"81",
           901 => x"70",
           902 => x"81",
           903 => x"80",
           904 => x"05",
           905 => x"76",
           906 => x"70",
           907 => x"0c",
           908 => x"04",
           909 => x"76",
           910 => x"80",
           911 => x"86",
           912 => x"52",
           913 => x"bd",
           914 => x"84",
           915 => x"80",
           916 => x"74",
           917 => x"d3",
           918 => x"3d",
           919 => x"3d",
           920 => x"11",
           921 => x"52",
           922 => x"70",
           923 => x"98",
           924 => x"33",
           925 => x"82",
           926 => x"26",
           927 => x"84",
           928 => x"83",
           929 => x"26",
           930 => x"85",
           931 => x"84",
           932 => x"26",
           933 => x"86",
           934 => x"85",
           935 => x"26",
           936 => x"88",
           937 => x"86",
           938 => x"e7",
           939 => x"38",
           940 => x"54",
           941 => x"87",
           942 => x"cc",
           943 => x"87",
           944 => x"0c",
           945 => x"c0",
           946 => x"82",
           947 => x"c0",
           948 => x"83",
           949 => x"c0",
           950 => x"84",
           951 => x"c0",
           952 => x"85",
           953 => x"c0",
           954 => x"86",
           955 => x"c0",
           956 => x"74",
           957 => x"a4",
           958 => x"c0",
           959 => x"80",
           960 => x"98",
           961 => x"52",
           962 => x"84",
           963 => x"0d",
           964 => x"0d",
           965 => x"c0",
           966 => x"81",
           967 => x"c0",
           968 => x"5e",
           969 => x"87",
           970 => x"08",
           971 => x"1c",
           972 => x"98",
           973 => x"79",
           974 => x"87",
           975 => x"08",
           976 => x"1c",
           977 => x"98",
           978 => x"79",
           979 => x"87",
           980 => x"08",
           981 => x"1c",
           982 => x"98",
           983 => x"7b",
           984 => x"87",
           985 => x"08",
           986 => x"1c",
           987 => x"0c",
           988 => x"ff",
           989 => x"83",
           990 => x"58",
           991 => x"57",
           992 => x"56",
           993 => x"55",
           994 => x"54",
           995 => x"53",
           996 => x"ff",
           997 => x"bd",
           998 => x"82",
           999 => x"0d",
          1000 => x"0d",
          1001 => x"33",
          1002 => x"9f",
          1003 => x"52",
          1004 => x"81",
          1005 => x"83",
          1006 => x"fb",
          1007 => x"0b",
          1008 => x"fc",
          1009 => x"ff",
          1010 => x"56",
          1011 => x"84",
          1012 => x"2e",
          1013 => x"c0",
          1014 => x"70",
          1015 => x"2a",
          1016 => x"53",
          1017 => x"80",
          1018 => x"71",
          1019 => x"81",
          1020 => x"70",
          1021 => x"81",
          1022 => x"06",
          1023 => x"80",
          1024 => x"71",
          1025 => x"81",
          1026 => x"70",
          1027 => x"73",
          1028 => x"51",
          1029 => x"80",
          1030 => x"2e",
          1031 => x"c0",
          1032 => x"75",
          1033 => x"81",
          1034 => x"87",
          1035 => x"fb",
          1036 => x"9f",
          1037 => x"0b",
          1038 => x"33",
          1039 => x"06",
          1040 => x"87",
          1041 => x"51",
          1042 => x"86",
          1043 => x"94",
          1044 => x"08",
          1045 => x"70",
          1046 => x"54",
          1047 => x"2e",
          1048 => x"91",
          1049 => x"06",
          1050 => x"d7",
          1051 => x"32",
          1052 => x"51",
          1053 => x"2e",
          1054 => x"93",
          1055 => x"06",
          1056 => x"ff",
          1057 => x"81",
          1058 => x"87",
          1059 => x"52",
          1060 => x"86",
          1061 => x"94",
          1062 => x"72",
          1063 => x"0d",
          1064 => x"0d",
          1065 => x"74",
          1066 => x"ff",
          1067 => x"57",
          1068 => x"80",
          1069 => x"81",
          1070 => x"15",
          1071 => x"cf",
          1072 => x"81",
          1073 => x"57",
          1074 => x"c0",
          1075 => x"75",
          1076 => x"38",
          1077 => x"94",
          1078 => x"70",
          1079 => x"81",
          1080 => x"52",
          1081 => x"8c",
          1082 => x"2a",
          1083 => x"51",
          1084 => x"38",
          1085 => x"70",
          1086 => x"51",
          1087 => x"8d",
          1088 => x"2a",
          1089 => x"51",
          1090 => x"be",
          1091 => x"ff",
          1092 => x"c0",
          1093 => x"70",
          1094 => x"38",
          1095 => x"90",
          1096 => x"0c",
          1097 => x"33",
          1098 => x"06",
          1099 => x"70",
          1100 => x"76",
          1101 => x"0c",
          1102 => x"04",
          1103 => x"0b",
          1104 => x"fc",
          1105 => x"ff",
          1106 => x"87",
          1107 => x"51",
          1108 => x"86",
          1109 => x"94",
          1110 => x"08",
          1111 => x"70",
          1112 => x"51",
          1113 => x"2e",
          1114 => x"81",
          1115 => x"87",
          1116 => x"52",
          1117 => x"86",
          1118 => x"94",
          1119 => x"08",
          1120 => x"06",
          1121 => x"0c",
          1122 => x"0d",
          1123 => x"0d",
          1124 => x"cf",
          1125 => x"81",
          1126 => x"53",
          1127 => x"84",
          1128 => x"2e",
          1129 => x"c0",
          1130 => x"71",
          1131 => x"2a",
          1132 => x"51",
          1133 => x"52",
          1134 => x"a0",
          1135 => x"ff",
          1136 => x"c0",
          1137 => x"70",
          1138 => x"38",
          1139 => x"90",
          1140 => x"70",
          1141 => x"98",
          1142 => x"51",
          1143 => x"84",
          1144 => x"0d",
          1145 => x"0d",
          1146 => x"80",
          1147 => x"2a",
          1148 => x"51",
          1149 => x"83",
          1150 => x"c0",
          1151 => x"81",
          1152 => x"87",
          1153 => x"08",
          1154 => x"0c",
          1155 => x"8c",
          1156 => x"88",
          1157 => x"9e",
          1158 => x"d0",
          1159 => x"c0",
          1160 => x"81",
          1161 => x"87",
          1162 => x"08",
          1163 => x"0c",
          1164 => x"a4",
          1165 => x"98",
          1166 => x"9e",
          1167 => x"d0",
          1168 => x"c0",
          1169 => x"81",
          1170 => x"87",
          1171 => x"08",
          1172 => x"d0",
          1173 => x"c0",
          1174 => x"81",
          1175 => x"81",
          1176 => x"ac",
          1177 => x"87",
          1178 => x"08",
          1179 => x"06",
          1180 => x"70",
          1181 => x"38",
          1182 => x"81",
          1183 => x"80",
          1184 => x"9e",
          1185 => x"81",
          1186 => x"51",
          1187 => x"80",
          1188 => x"81",
          1189 => x"d0",
          1190 => x"0b",
          1191 => x"88",
          1192 => x"c0",
          1193 => x"52",
          1194 => x"2e",
          1195 => x"52",
          1196 => x"af",
          1197 => x"87",
          1198 => x"08",
          1199 => x"06",
          1200 => x"70",
          1201 => x"38",
          1202 => x"81",
          1203 => x"80",
          1204 => x"9e",
          1205 => x"88",
          1206 => x"52",
          1207 => x"2e",
          1208 => x"52",
          1209 => x"b1",
          1210 => x"87",
          1211 => x"08",
          1212 => x"06",
          1213 => x"70",
          1214 => x"38",
          1215 => x"81",
          1216 => x"80",
          1217 => x"9e",
          1218 => x"82",
          1219 => x"52",
          1220 => x"2e",
          1221 => x"52",
          1222 => x"b3",
          1223 => x"87",
          1224 => x"08",
          1225 => x"06",
          1226 => x"70",
          1227 => x"38",
          1228 => x"81",
          1229 => x"87",
          1230 => x"08",
          1231 => x"06",
          1232 => x"51",
          1233 => x"81",
          1234 => x"80",
          1235 => x"9e",
          1236 => x"90",
          1237 => x"52",
          1238 => x"83",
          1239 => x"71",
          1240 => x"34",
          1241 => x"c0",
          1242 => x"70",
          1243 => x"52",
          1244 => x"2e",
          1245 => x"52",
          1246 => x"b7",
          1247 => x"9e",
          1248 => x"87",
          1249 => x"70",
          1250 => x"34",
          1251 => x"04",
          1252 => x"81",
          1253 => x"84",
          1254 => x"d0",
          1255 => x"73",
          1256 => x"38",
          1257 => x"51",
          1258 => x"81",
          1259 => x"84",
          1260 => x"d0",
          1261 => x"73",
          1262 => x"38",
          1263 => x"08",
          1264 => x"80",
          1265 => x"be",
          1266 => x"d2",
          1267 => x"ae",
          1268 => x"80",
          1269 => x"81",
          1270 => x"53",
          1271 => x"08",
          1272 => x"d0",
          1273 => x"3f",
          1274 => x"33",
          1275 => x"38",
          1276 => x"33",
          1277 => x"2e",
          1278 => x"d0",
          1279 => x"81",
          1280 => x"52",
          1281 => x"51",
          1282 => x"81",
          1283 => x"54",
          1284 => x"88",
          1285 => x"98",
          1286 => x"3f",
          1287 => x"33",
          1288 => x"2e",
          1289 => x"bf",
          1290 => x"8e",
          1291 => x"b3",
          1292 => x"80",
          1293 => x"81",
          1294 => x"82",
          1295 => x"d0",
          1296 => x"73",
          1297 => x"38",
          1298 => x"33",
          1299 => x"bc",
          1300 => x"3f",
          1301 => x"33",
          1302 => x"2e",
          1303 => x"bf",
          1304 => x"d6",
          1305 => x"b7",
          1306 => x"80",
          1307 => x"81",
          1308 => x"52",
          1309 => x"51",
          1310 => x"81",
          1311 => x"82",
          1312 => x"d0",
          1313 => x"81",
          1314 => x"88",
          1315 => x"d0",
          1316 => x"81",
          1317 => x"88",
          1318 => x"d0",
          1319 => x"81",
          1320 => x"87",
          1321 => x"d0",
          1322 => x"81",
          1323 => x"87",
          1324 => x"d0",
          1325 => x"81",
          1326 => x"87",
          1327 => x"3d",
          1328 => x"3d",
          1329 => x"05",
          1330 => x"52",
          1331 => x"aa",
          1332 => x"29",
          1333 => x"05",
          1334 => x"04",
          1335 => x"51",
          1336 => x"c1",
          1337 => x"39",
          1338 => x"51",
          1339 => x"c2",
          1340 => x"39",
          1341 => x"51",
          1342 => x"c2",
          1343 => x"a1",
          1344 => x"0d",
          1345 => x"80",
          1346 => x"0b",
          1347 => x"84",
          1348 => x"3d",
          1349 => x"96",
          1350 => x"52",
          1351 => x"0c",
          1352 => x"70",
          1353 => x"0c",
          1354 => x"3d",
          1355 => x"3d",
          1356 => x"96",
          1357 => x"81",
          1358 => x"52",
          1359 => x"73",
          1360 => x"d0",
          1361 => x"70",
          1362 => x"0c",
          1363 => x"83",
          1364 => x"81",
          1365 => x"87",
          1366 => x"0c",
          1367 => x"0d",
          1368 => x"33",
          1369 => x"2e",
          1370 => x"85",
          1371 => x"ed",
          1372 => x"9c",
          1373 => x"80",
          1374 => x"72",
          1375 => x"d3",
          1376 => x"05",
          1377 => x"0c",
          1378 => x"d3",
          1379 => x"71",
          1380 => x"38",
          1381 => x"2d",
          1382 => x"04",
          1383 => x"02",
          1384 => x"81",
          1385 => x"76",
          1386 => x"0c",
          1387 => x"ad",
          1388 => x"d3",
          1389 => x"3d",
          1390 => x"3d",
          1391 => x"73",
          1392 => x"ff",
          1393 => x"71",
          1394 => x"38",
          1395 => x"06",
          1396 => x"54",
          1397 => x"e7",
          1398 => x"0d",
          1399 => x"0d",
          1400 => x"94",
          1401 => x"d3",
          1402 => x"54",
          1403 => x"81",
          1404 => x"53",
          1405 => x"8e",
          1406 => x"ff",
          1407 => x"14",
          1408 => x"3f",
          1409 => x"81",
          1410 => x"86",
          1411 => x"ec",
          1412 => x"68",
          1413 => x"70",
          1414 => x"33",
          1415 => x"2e",
          1416 => x"75",
          1417 => x"81",
          1418 => x"38",
          1419 => x"70",
          1420 => x"33",
          1421 => x"75",
          1422 => x"81",
          1423 => x"81",
          1424 => x"75",
          1425 => x"81",
          1426 => x"82",
          1427 => x"81",
          1428 => x"56",
          1429 => x"09",
          1430 => x"38",
          1431 => x"71",
          1432 => x"81",
          1433 => x"59",
          1434 => x"9d",
          1435 => x"53",
          1436 => x"95",
          1437 => x"29",
          1438 => x"76",
          1439 => x"79",
          1440 => x"5b",
          1441 => x"e5",
          1442 => x"ec",
          1443 => x"70",
          1444 => x"25",
          1445 => x"32",
          1446 => x"72",
          1447 => x"73",
          1448 => x"58",
          1449 => x"73",
          1450 => x"38",
          1451 => x"79",
          1452 => x"5b",
          1453 => x"75",
          1454 => x"de",
          1455 => x"80",
          1456 => x"89",
          1457 => x"70",
          1458 => x"55",
          1459 => x"cf",
          1460 => x"38",
          1461 => x"24",
          1462 => x"80",
          1463 => x"8e",
          1464 => x"c3",
          1465 => x"73",
          1466 => x"81",
          1467 => x"99",
          1468 => x"c4",
          1469 => x"38",
          1470 => x"73",
          1471 => x"81",
          1472 => x"80",
          1473 => x"38",
          1474 => x"2e",
          1475 => x"f9",
          1476 => x"d8",
          1477 => x"38",
          1478 => x"77",
          1479 => x"08",
          1480 => x"80",
          1481 => x"55",
          1482 => x"8d",
          1483 => x"70",
          1484 => x"51",
          1485 => x"f5",
          1486 => x"2a",
          1487 => x"74",
          1488 => x"53",
          1489 => x"8f",
          1490 => x"fc",
          1491 => x"81",
          1492 => x"80",
          1493 => x"73",
          1494 => x"3f",
          1495 => x"56",
          1496 => x"27",
          1497 => x"a0",
          1498 => x"3f",
          1499 => x"84",
          1500 => x"33",
          1501 => x"93",
          1502 => x"95",
          1503 => x"91",
          1504 => x"8d",
          1505 => x"89",
          1506 => x"fb",
          1507 => x"86",
          1508 => x"2a",
          1509 => x"51",
          1510 => x"2e",
          1511 => x"84",
          1512 => x"86",
          1513 => x"78",
          1514 => x"08",
          1515 => x"32",
          1516 => x"72",
          1517 => x"51",
          1518 => x"74",
          1519 => x"38",
          1520 => x"88",
          1521 => x"7a",
          1522 => x"55",
          1523 => x"3d",
          1524 => x"52",
          1525 => x"d3",
          1526 => x"84",
          1527 => x"06",
          1528 => x"52",
          1529 => x"3f",
          1530 => x"08",
          1531 => x"27",
          1532 => x"14",
          1533 => x"f8",
          1534 => x"87",
          1535 => x"81",
          1536 => x"b0",
          1537 => x"7d",
          1538 => x"5f",
          1539 => x"75",
          1540 => x"07",
          1541 => x"54",
          1542 => x"26",
          1543 => x"ff",
          1544 => x"84",
          1545 => x"06",
          1546 => x"80",
          1547 => x"96",
          1548 => x"e0",
          1549 => x"73",
          1550 => x"57",
          1551 => x"06",
          1552 => x"54",
          1553 => x"a0",
          1554 => x"2a",
          1555 => x"54",
          1556 => x"38",
          1557 => x"76",
          1558 => x"38",
          1559 => x"fd",
          1560 => x"06",
          1561 => x"38",
          1562 => x"56",
          1563 => x"26",
          1564 => x"3d",
          1565 => x"05",
          1566 => x"ff",
          1567 => x"53",
          1568 => x"d9",
          1569 => x"38",
          1570 => x"56",
          1571 => x"27",
          1572 => x"a0",
          1573 => x"3f",
          1574 => x"3d",
          1575 => x"3d",
          1576 => x"70",
          1577 => x"52",
          1578 => x"73",
          1579 => x"3f",
          1580 => x"04",
          1581 => x"74",
          1582 => x"0c",
          1583 => x"05",
          1584 => x"fa",
          1585 => x"d3",
          1586 => x"80",
          1587 => x"0b",
          1588 => x"0c",
          1589 => x"04",
          1590 => x"81",
          1591 => x"76",
          1592 => x"0c",
          1593 => x"05",
          1594 => x"53",
          1595 => x"72",
          1596 => x"0c",
          1597 => x"04",
          1598 => x"77",
          1599 => x"98",
          1600 => x"54",
          1601 => x"54",
          1602 => x"80",
          1603 => x"d3",
          1604 => x"71",
          1605 => x"84",
          1606 => x"06",
          1607 => x"2e",
          1608 => x"72",
          1609 => x"38",
          1610 => x"70",
          1611 => x"25",
          1612 => x"73",
          1613 => x"38",
          1614 => x"86",
          1615 => x"54",
          1616 => x"73",
          1617 => x"ff",
          1618 => x"72",
          1619 => x"74",
          1620 => x"72",
          1621 => x"54",
          1622 => x"81",
          1623 => x"39",
          1624 => x"80",
          1625 => x"51",
          1626 => x"81",
          1627 => x"d3",
          1628 => x"3d",
          1629 => x"3d",
          1630 => x"98",
          1631 => x"d3",
          1632 => x"53",
          1633 => x"fe",
          1634 => x"81",
          1635 => x"84",
          1636 => x"f8",
          1637 => x"7c",
          1638 => x"70",
          1639 => x"75",
          1640 => x"55",
          1641 => x"2e",
          1642 => x"87",
          1643 => x"76",
          1644 => x"73",
          1645 => x"81",
          1646 => x"81",
          1647 => x"77",
          1648 => x"70",
          1649 => x"58",
          1650 => x"09",
          1651 => x"c2",
          1652 => x"81",
          1653 => x"75",
          1654 => x"55",
          1655 => x"e2",
          1656 => x"90",
          1657 => x"f8",
          1658 => x"8f",
          1659 => x"81",
          1660 => x"75",
          1661 => x"55",
          1662 => x"81",
          1663 => x"27",
          1664 => x"d0",
          1665 => x"55",
          1666 => x"73",
          1667 => x"80",
          1668 => x"14",
          1669 => x"72",
          1670 => x"e0",
          1671 => x"80",
          1672 => x"39",
          1673 => x"55",
          1674 => x"80",
          1675 => x"e0",
          1676 => x"38",
          1677 => x"81",
          1678 => x"53",
          1679 => x"81",
          1680 => x"53",
          1681 => x"8e",
          1682 => x"70",
          1683 => x"55",
          1684 => x"27",
          1685 => x"77",
          1686 => x"74",
          1687 => x"76",
          1688 => x"77",
          1689 => x"70",
          1690 => x"55",
          1691 => x"77",
          1692 => x"38",
          1693 => x"74",
          1694 => x"55",
          1695 => x"84",
          1696 => x"0d",
          1697 => x"0d",
          1698 => x"56",
          1699 => x"0c",
          1700 => x"70",
          1701 => x"73",
          1702 => x"81",
          1703 => x"81",
          1704 => x"ed",
          1705 => x"2e",
          1706 => x"8e",
          1707 => x"08",
          1708 => x"76",
          1709 => x"56",
          1710 => x"b0",
          1711 => x"06",
          1712 => x"75",
          1713 => x"76",
          1714 => x"70",
          1715 => x"73",
          1716 => x"8b",
          1717 => x"73",
          1718 => x"85",
          1719 => x"82",
          1720 => x"76",
          1721 => x"70",
          1722 => x"ac",
          1723 => x"a0",
          1724 => x"fa",
          1725 => x"53",
          1726 => x"57",
          1727 => x"98",
          1728 => x"39",
          1729 => x"80",
          1730 => x"26",
          1731 => x"86",
          1732 => x"80",
          1733 => x"57",
          1734 => x"74",
          1735 => x"38",
          1736 => x"27",
          1737 => x"14",
          1738 => x"06",
          1739 => x"14",
          1740 => x"06",
          1741 => x"74",
          1742 => x"f9",
          1743 => x"ff",
          1744 => x"89",
          1745 => x"38",
          1746 => x"c5",
          1747 => x"29",
          1748 => x"81",
          1749 => x"76",
          1750 => x"56",
          1751 => x"ba",
          1752 => x"2e",
          1753 => x"30",
          1754 => x"0c",
          1755 => x"81",
          1756 => x"8a",
          1757 => x"ff",
          1758 => x"8f",
          1759 => x"81",
          1760 => x"26",
          1761 => x"d0",
          1762 => x"52",
          1763 => x"84",
          1764 => x"0d",
          1765 => x"0d",
          1766 => x"33",
          1767 => x"9f",
          1768 => x"53",
          1769 => x"81",
          1770 => x"38",
          1771 => x"87",
          1772 => x"11",
          1773 => x"54",
          1774 => x"84",
          1775 => x"54",
          1776 => x"87",
          1777 => x"11",
          1778 => x"0c",
          1779 => x"c0",
          1780 => x"70",
          1781 => x"70",
          1782 => x"51",
          1783 => x"8a",
          1784 => x"98",
          1785 => x"70",
          1786 => x"08",
          1787 => x"06",
          1788 => x"38",
          1789 => x"8c",
          1790 => x"80",
          1791 => x"71",
          1792 => x"14",
          1793 => x"c0",
          1794 => x"70",
          1795 => x"0c",
          1796 => x"04",
          1797 => x"60",
          1798 => x"8c",
          1799 => x"33",
          1800 => x"5b",
          1801 => x"5a",
          1802 => x"81",
          1803 => x"81",
          1804 => x"52",
          1805 => x"38",
          1806 => x"84",
          1807 => x"92",
          1808 => x"c0",
          1809 => x"87",
          1810 => x"13",
          1811 => x"57",
          1812 => x"0b",
          1813 => x"8c",
          1814 => x"0c",
          1815 => x"75",
          1816 => x"2a",
          1817 => x"51",
          1818 => x"80",
          1819 => x"7b",
          1820 => x"7b",
          1821 => x"5d",
          1822 => x"59",
          1823 => x"06",
          1824 => x"73",
          1825 => x"81",
          1826 => x"ff",
          1827 => x"72",
          1828 => x"38",
          1829 => x"8c",
          1830 => x"c3",
          1831 => x"98",
          1832 => x"71",
          1833 => x"38",
          1834 => x"2e",
          1835 => x"76",
          1836 => x"92",
          1837 => x"72",
          1838 => x"06",
          1839 => x"f7",
          1840 => x"5a",
          1841 => x"80",
          1842 => x"70",
          1843 => x"5a",
          1844 => x"80",
          1845 => x"73",
          1846 => x"06",
          1847 => x"38",
          1848 => x"fe",
          1849 => x"fc",
          1850 => x"52",
          1851 => x"83",
          1852 => x"71",
          1853 => x"d3",
          1854 => x"3d",
          1855 => x"3d",
          1856 => x"64",
          1857 => x"bf",
          1858 => x"40",
          1859 => x"59",
          1860 => x"58",
          1861 => x"81",
          1862 => x"81",
          1863 => x"52",
          1864 => x"09",
          1865 => x"b1",
          1866 => x"84",
          1867 => x"92",
          1868 => x"c0",
          1869 => x"87",
          1870 => x"13",
          1871 => x"56",
          1872 => x"87",
          1873 => x"0c",
          1874 => x"82",
          1875 => x"58",
          1876 => x"84",
          1877 => x"06",
          1878 => x"71",
          1879 => x"38",
          1880 => x"05",
          1881 => x"0c",
          1882 => x"73",
          1883 => x"81",
          1884 => x"71",
          1885 => x"38",
          1886 => x"8c",
          1887 => x"d0",
          1888 => x"98",
          1889 => x"71",
          1890 => x"38",
          1891 => x"2e",
          1892 => x"76",
          1893 => x"92",
          1894 => x"72",
          1895 => x"06",
          1896 => x"f7",
          1897 => x"59",
          1898 => x"1a",
          1899 => x"06",
          1900 => x"59",
          1901 => x"80",
          1902 => x"73",
          1903 => x"06",
          1904 => x"38",
          1905 => x"fe",
          1906 => x"fc",
          1907 => x"52",
          1908 => x"83",
          1909 => x"71",
          1910 => x"d3",
          1911 => x"3d",
          1912 => x"3d",
          1913 => x"84",
          1914 => x"33",
          1915 => x"b7",
          1916 => x"54",
          1917 => x"fa",
          1918 => x"d3",
          1919 => x"06",
          1920 => x"72",
          1921 => x"85",
          1922 => x"98",
          1923 => x"56",
          1924 => x"80",
          1925 => x"76",
          1926 => x"74",
          1927 => x"c0",
          1928 => x"54",
          1929 => x"2e",
          1930 => x"d4",
          1931 => x"2e",
          1932 => x"80",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"c0",
          1938 => x"52",
          1939 => x"87",
          1940 => x"08",
          1941 => x"38",
          1942 => x"87",
          1943 => x"14",
          1944 => x"70",
          1945 => x"52",
          1946 => x"96",
          1947 => x"92",
          1948 => x"0a",
          1949 => x"39",
          1950 => x"0c",
          1951 => x"39",
          1952 => x"54",
          1953 => x"84",
          1954 => x"0d",
          1955 => x"0d",
          1956 => x"33",
          1957 => x"88",
          1958 => x"d3",
          1959 => x"51",
          1960 => x"04",
          1961 => x"75",
          1962 => x"82",
          1963 => x"90",
          1964 => x"2b",
          1965 => x"33",
          1966 => x"88",
          1967 => x"71",
          1968 => x"84",
          1969 => x"54",
          1970 => x"85",
          1971 => x"ff",
          1972 => x"02",
          1973 => x"05",
          1974 => x"70",
          1975 => x"05",
          1976 => x"88",
          1977 => x"72",
          1978 => x"0d",
          1979 => x"0d",
          1980 => x"52",
          1981 => x"81",
          1982 => x"70",
          1983 => x"70",
          1984 => x"05",
          1985 => x"88",
          1986 => x"72",
          1987 => x"54",
          1988 => x"2a",
          1989 => x"34",
          1990 => x"04",
          1991 => x"76",
          1992 => x"54",
          1993 => x"2e",
          1994 => x"70",
          1995 => x"33",
          1996 => x"05",
          1997 => x"11",
          1998 => x"84",
          1999 => x"fe",
          2000 => x"77",
          2001 => x"53",
          2002 => x"81",
          2003 => x"ff",
          2004 => x"f4",
          2005 => x"0d",
          2006 => x"0d",
          2007 => x"56",
          2008 => x"70",
          2009 => x"33",
          2010 => x"05",
          2011 => x"71",
          2012 => x"56",
          2013 => x"72",
          2014 => x"38",
          2015 => x"e2",
          2016 => x"d3",
          2017 => x"3d",
          2018 => x"3d",
          2019 => x"54",
          2020 => x"71",
          2021 => x"38",
          2022 => x"70",
          2023 => x"f3",
          2024 => x"81",
          2025 => x"84",
          2026 => x"80",
          2027 => x"84",
          2028 => x"0b",
          2029 => x"0c",
          2030 => x"0d",
          2031 => x"0b",
          2032 => x"56",
          2033 => x"2e",
          2034 => x"81",
          2035 => x"08",
          2036 => x"70",
          2037 => x"33",
          2038 => x"a2",
          2039 => x"84",
          2040 => x"09",
          2041 => x"38",
          2042 => x"08",
          2043 => x"b0",
          2044 => x"a4",
          2045 => x"9c",
          2046 => x"56",
          2047 => x"27",
          2048 => x"16",
          2049 => x"82",
          2050 => x"06",
          2051 => x"54",
          2052 => x"78",
          2053 => x"33",
          2054 => x"3f",
          2055 => x"5a",
          2056 => x"84",
          2057 => x"0d",
          2058 => x"0d",
          2059 => x"56",
          2060 => x"b0",
          2061 => x"af",
          2062 => x"fe",
          2063 => x"d3",
          2064 => x"81",
          2065 => x"9f",
          2066 => x"74",
          2067 => x"52",
          2068 => x"51",
          2069 => x"81",
          2070 => x"80",
          2071 => x"ff",
          2072 => x"74",
          2073 => x"76",
          2074 => x"0c",
          2075 => x"04",
          2076 => x"7a",
          2077 => x"fe",
          2078 => x"d3",
          2079 => x"81",
          2080 => x"81",
          2081 => x"33",
          2082 => x"2e",
          2083 => x"80",
          2084 => x"17",
          2085 => x"81",
          2086 => x"06",
          2087 => x"84",
          2088 => x"d3",
          2089 => x"b4",
          2090 => x"56",
          2091 => x"82",
          2092 => x"84",
          2093 => x"fc",
          2094 => x"8b",
          2095 => x"52",
          2096 => x"a9",
          2097 => x"85",
          2098 => x"84",
          2099 => x"fc",
          2100 => x"17",
          2101 => x"9c",
          2102 => x"91",
          2103 => x"08",
          2104 => x"17",
          2105 => x"3f",
          2106 => x"81",
          2107 => x"19",
          2108 => x"53",
          2109 => x"17",
          2110 => x"82",
          2111 => x"18",
          2112 => x"80",
          2113 => x"33",
          2114 => x"3f",
          2115 => x"08",
          2116 => x"38",
          2117 => x"81",
          2118 => x"8a",
          2119 => x"fb",
          2120 => x"fe",
          2121 => x"08",
          2122 => x"56",
          2123 => x"74",
          2124 => x"38",
          2125 => x"75",
          2126 => x"16",
          2127 => x"53",
          2128 => x"84",
          2129 => x"0d",
          2130 => x"0d",
          2131 => x"08",
          2132 => x"81",
          2133 => x"df",
          2134 => x"15",
          2135 => x"d7",
          2136 => x"33",
          2137 => x"82",
          2138 => x"38",
          2139 => x"89",
          2140 => x"2e",
          2141 => x"bf",
          2142 => x"2e",
          2143 => x"81",
          2144 => x"81",
          2145 => x"89",
          2146 => x"08",
          2147 => x"52",
          2148 => x"3f",
          2149 => x"08",
          2150 => x"74",
          2151 => x"14",
          2152 => x"81",
          2153 => x"2a",
          2154 => x"05",
          2155 => x"57",
          2156 => x"f5",
          2157 => x"84",
          2158 => x"38",
          2159 => x"06",
          2160 => x"33",
          2161 => x"78",
          2162 => x"06",
          2163 => x"5c",
          2164 => x"53",
          2165 => x"38",
          2166 => x"06",
          2167 => x"39",
          2168 => x"a4",
          2169 => x"52",
          2170 => x"bd",
          2171 => x"84",
          2172 => x"38",
          2173 => x"fe",
          2174 => x"b4",
          2175 => x"8d",
          2176 => x"84",
          2177 => x"ff",
          2178 => x"39",
          2179 => x"a4",
          2180 => x"52",
          2181 => x"91",
          2182 => x"84",
          2183 => x"76",
          2184 => x"fc",
          2185 => x"b4",
          2186 => x"f8",
          2187 => x"84",
          2188 => x"06",
          2189 => x"81",
          2190 => x"d3",
          2191 => x"3d",
          2192 => x"3d",
          2193 => x"7e",
          2194 => x"82",
          2195 => x"27",
          2196 => x"76",
          2197 => x"27",
          2198 => x"75",
          2199 => x"79",
          2200 => x"38",
          2201 => x"89",
          2202 => x"2e",
          2203 => x"80",
          2204 => x"2e",
          2205 => x"81",
          2206 => x"81",
          2207 => x"89",
          2208 => x"08",
          2209 => x"52",
          2210 => x"3f",
          2211 => x"08",
          2212 => x"84",
          2213 => x"38",
          2214 => x"06",
          2215 => x"81",
          2216 => x"06",
          2217 => x"77",
          2218 => x"2e",
          2219 => x"84",
          2220 => x"06",
          2221 => x"06",
          2222 => x"53",
          2223 => x"81",
          2224 => x"34",
          2225 => x"a4",
          2226 => x"52",
          2227 => x"d9",
          2228 => x"84",
          2229 => x"d3",
          2230 => x"94",
          2231 => x"ff",
          2232 => x"05",
          2233 => x"54",
          2234 => x"38",
          2235 => x"74",
          2236 => x"06",
          2237 => x"07",
          2238 => x"74",
          2239 => x"39",
          2240 => x"a4",
          2241 => x"52",
          2242 => x"9d",
          2243 => x"84",
          2244 => x"d3",
          2245 => x"d8",
          2246 => x"ff",
          2247 => x"76",
          2248 => x"06",
          2249 => x"05",
          2250 => x"3f",
          2251 => x"87",
          2252 => x"08",
          2253 => x"51",
          2254 => x"81",
          2255 => x"59",
          2256 => x"08",
          2257 => x"f0",
          2258 => x"82",
          2259 => x"06",
          2260 => x"05",
          2261 => x"54",
          2262 => x"3f",
          2263 => x"08",
          2264 => x"74",
          2265 => x"51",
          2266 => x"81",
          2267 => x"34",
          2268 => x"84",
          2269 => x"0d",
          2270 => x"0d",
          2271 => x"72",
          2272 => x"56",
          2273 => x"27",
          2274 => x"98",
          2275 => x"9d",
          2276 => x"2e",
          2277 => x"53",
          2278 => x"51",
          2279 => x"81",
          2280 => x"54",
          2281 => x"08",
          2282 => x"93",
          2283 => x"80",
          2284 => x"54",
          2285 => x"81",
          2286 => x"54",
          2287 => x"74",
          2288 => x"fb",
          2289 => x"d3",
          2290 => x"81",
          2291 => x"80",
          2292 => x"38",
          2293 => x"08",
          2294 => x"38",
          2295 => x"08",
          2296 => x"38",
          2297 => x"52",
          2298 => x"d6",
          2299 => x"84",
          2300 => x"98",
          2301 => x"11",
          2302 => x"57",
          2303 => x"74",
          2304 => x"81",
          2305 => x"0c",
          2306 => x"81",
          2307 => x"84",
          2308 => x"55",
          2309 => x"ff",
          2310 => x"54",
          2311 => x"84",
          2312 => x"0d",
          2313 => x"0d",
          2314 => x"08",
          2315 => x"79",
          2316 => x"17",
          2317 => x"80",
          2318 => x"98",
          2319 => x"26",
          2320 => x"58",
          2321 => x"52",
          2322 => x"fd",
          2323 => x"74",
          2324 => x"08",
          2325 => x"38",
          2326 => x"08",
          2327 => x"84",
          2328 => x"82",
          2329 => x"17",
          2330 => x"84",
          2331 => x"c7",
          2332 => x"90",
          2333 => x"56",
          2334 => x"2e",
          2335 => x"77",
          2336 => x"81",
          2337 => x"38",
          2338 => x"98",
          2339 => x"26",
          2340 => x"56",
          2341 => x"51",
          2342 => x"80",
          2343 => x"84",
          2344 => x"09",
          2345 => x"38",
          2346 => x"08",
          2347 => x"84",
          2348 => x"30",
          2349 => x"80",
          2350 => x"07",
          2351 => x"08",
          2352 => x"55",
          2353 => x"ef",
          2354 => x"84",
          2355 => x"95",
          2356 => x"08",
          2357 => x"27",
          2358 => x"98",
          2359 => x"89",
          2360 => x"85",
          2361 => x"db",
          2362 => x"81",
          2363 => x"17",
          2364 => x"89",
          2365 => x"75",
          2366 => x"ac",
          2367 => x"7a",
          2368 => x"3f",
          2369 => x"08",
          2370 => x"38",
          2371 => x"d3",
          2372 => x"2e",
          2373 => x"86",
          2374 => x"84",
          2375 => x"d3",
          2376 => x"70",
          2377 => x"07",
          2378 => x"7c",
          2379 => x"55",
          2380 => x"f8",
          2381 => x"2e",
          2382 => x"ff",
          2383 => x"55",
          2384 => x"ff",
          2385 => x"76",
          2386 => x"3f",
          2387 => x"08",
          2388 => x"08",
          2389 => x"d3",
          2390 => x"80",
          2391 => x"55",
          2392 => x"94",
          2393 => x"2e",
          2394 => x"53",
          2395 => x"51",
          2396 => x"81",
          2397 => x"55",
          2398 => x"75",
          2399 => x"98",
          2400 => x"05",
          2401 => x"56",
          2402 => x"26",
          2403 => x"15",
          2404 => x"84",
          2405 => x"07",
          2406 => x"18",
          2407 => x"ff",
          2408 => x"2e",
          2409 => x"39",
          2410 => x"39",
          2411 => x"08",
          2412 => x"81",
          2413 => x"74",
          2414 => x"0c",
          2415 => x"04",
          2416 => x"7a",
          2417 => x"f3",
          2418 => x"d3",
          2419 => x"81",
          2420 => x"84",
          2421 => x"38",
          2422 => x"51",
          2423 => x"81",
          2424 => x"81",
          2425 => x"b0",
          2426 => x"84",
          2427 => x"52",
          2428 => x"52",
          2429 => x"3f",
          2430 => x"39",
          2431 => x"8a",
          2432 => x"75",
          2433 => x"38",
          2434 => x"19",
          2435 => x"81",
          2436 => x"ed",
          2437 => x"d3",
          2438 => x"2e",
          2439 => x"15",
          2440 => x"70",
          2441 => x"07",
          2442 => x"53",
          2443 => x"75",
          2444 => x"0c",
          2445 => x"04",
          2446 => x"7a",
          2447 => x"58",
          2448 => x"f0",
          2449 => x"80",
          2450 => x"9f",
          2451 => x"80",
          2452 => x"90",
          2453 => x"17",
          2454 => x"aa",
          2455 => x"53",
          2456 => x"88",
          2457 => x"08",
          2458 => x"38",
          2459 => x"53",
          2460 => x"17",
          2461 => x"72",
          2462 => x"fe",
          2463 => x"08",
          2464 => x"80",
          2465 => x"16",
          2466 => x"2b",
          2467 => x"75",
          2468 => x"73",
          2469 => x"f5",
          2470 => x"d3",
          2471 => x"81",
          2472 => x"ff",
          2473 => x"81",
          2474 => x"84",
          2475 => x"38",
          2476 => x"81",
          2477 => x"26",
          2478 => x"58",
          2479 => x"73",
          2480 => x"39",
          2481 => x"51",
          2482 => x"81",
          2483 => x"98",
          2484 => x"94",
          2485 => x"17",
          2486 => x"58",
          2487 => x"9a",
          2488 => x"81",
          2489 => x"74",
          2490 => x"98",
          2491 => x"83",
          2492 => x"b4",
          2493 => x"0c",
          2494 => x"81",
          2495 => x"8a",
          2496 => x"f8",
          2497 => x"70",
          2498 => x"08",
          2499 => x"57",
          2500 => x"0a",
          2501 => x"38",
          2502 => x"15",
          2503 => x"08",
          2504 => x"72",
          2505 => x"cb",
          2506 => x"ff",
          2507 => x"81",
          2508 => x"13",
          2509 => x"94",
          2510 => x"74",
          2511 => x"85",
          2512 => x"22",
          2513 => x"73",
          2514 => x"38",
          2515 => x"8a",
          2516 => x"05",
          2517 => x"06",
          2518 => x"8a",
          2519 => x"73",
          2520 => x"3f",
          2521 => x"08",
          2522 => x"81",
          2523 => x"84",
          2524 => x"ff",
          2525 => x"81",
          2526 => x"ff",
          2527 => x"38",
          2528 => x"81",
          2529 => x"26",
          2530 => x"7b",
          2531 => x"98",
          2532 => x"55",
          2533 => x"94",
          2534 => x"73",
          2535 => x"3f",
          2536 => x"08",
          2537 => x"81",
          2538 => x"80",
          2539 => x"38",
          2540 => x"d3",
          2541 => x"2e",
          2542 => x"55",
          2543 => x"08",
          2544 => x"38",
          2545 => x"08",
          2546 => x"fb",
          2547 => x"d3",
          2548 => x"38",
          2549 => x"0c",
          2550 => x"51",
          2551 => x"81",
          2552 => x"98",
          2553 => x"90",
          2554 => x"16",
          2555 => x"15",
          2556 => x"74",
          2557 => x"0c",
          2558 => x"04",
          2559 => x"7b",
          2560 => x"5b",
          2561 => x"52",
          2562 => x"ac",
          2563 => x"84",
          2564 => x"d3",
          2565 => x"ec",
          2566 => x"84",
          2567 => x"17",
          2568 => x"51",
          2569 => x"81",
          2570 => x"54",
          2571 => x"08",
          2572 => x"81",
          2573 => x"9c",
          2574 => x"33",
          2575 => x"72",
          2576 => x"09",
          2577 => x"38",
          2578 => x"d3",
          2579 => x"72",
          2580 => x"55",
          2581 => x"53",
          2582 => x"8e",
          2583 => x"56",
          2584 => x"09",
          2585 => x"38",
          2586 => x"d3",
          2587 => x"81",
          2588 => x"fd",
          2589 => x"d3",
          2590 => x"81",
          2591 => x"80",
          2592 => x"38",
          2593 => x"09",
          2594 => x"38",
          2595 => x"81",
          2596 => x"8b",
          2597 => x"fd",
          2598 => x"9a",
          2599 => x"eb",
          2600 => x"d3",
          2601 => x"ff",
          2602 => x"70",
          2603 => x"53",
          2604 => x"09",
          2605 => x"38",
          2606 => x"eb",
          2607 => x"d3",
          2608 => x"2b",
          2609 => x"72",
          2610 => x"0c",
          2611 => x"04",
          2612 => x"77",
          2613 => x"ff",
          2614 => x"9a",
          2615 => x"55",
          2616 => x"76",
          2617 => x"53",
          2618 => x"09",
          2619 => x"38",
          2620 => x"52",
          2621 => x"eb",
          2622 => x"3d",
          2623 => x"3d",
          2624 => x"5b",
          2625 => x"08",
          2626 => x"15",
          2627 => x"81",
          2628 => x"15",
          2629 => x"51",
          2630 => x"81",
          2631 => x"58",
          2632 => x"08",
          2633 => x"9c",
          2634 => x"33",
          2635 => x"86",
          2636 => x"80",
          2637 => x"13",
          2638 => x"06",
          2639 => x"06",
          2640 => x"72",
          2641 => x"81",
          2642 => x"53",
          2643 => x"2e",
          2644 => x"53",
          2645 => x"a9",
          2646 => x"74",
          2647 => x"72",
          2648 => x"38",
          2649 => x"99",
          2650 => x"84",
          2651 => x"06",
          2652 => x"88",
          2653 => x"06",
          2654 => x"54",
          2655 => x"a0",
          2656 => x"74",
          2657 => x"3f",
          2658 => x"08",
          2659 => x"84",
          2660 => x"98",
          2661 => x"fa",
          2662 => x"80",
          2663 => x"0c",
          2664 => x"84",
          2665 => x"0d",
          2666 => x"0d",
          2667 => x"57",
          2668 => x"73",
          2669 => x"3f",
          2670 => x"08",
          2671 => x"84",
          2672 => x"98",
          2673 => x"75",
          2674 => x"3f",
          2675 => x"08",
          2676 => x"84",
          2677 => x"a0",
          2678 => x"84",
          2679 => x"14",
          2680 => x"db",
          2681 => x"a0",
          2682 => x"14",
          2683 => x"ac",
          2684 => x"83",
          2685 => x"81",
          2686 => x"87",
          2687 => x"fd",
          2688 => x"70",
          2689 => x"08",
          2690 => x"55",
          2691 => x"3f",
          2692 => x"08",
          2693 => x"13",
          2694 => x"73",
          2695 => x"83",
          2696 => x"3d",
          2697 => x"3d",
          2698 => x"57",
          2699 => x"89",
          2700 => x"17",
          2701 => x"81",
          2702 => x"70",
          2703 => x"55",
          2704 => x"08",
          2705 => x"81",
          2706 => x"52",
          2707 => x"a8",
          2708 => x"2e",
          2709 => x"84",
          2710 => x"52",
          2711 => x"09",
          2712 => x"38",
          2713 => x"81",
          2714 => x"81",
          2715 => x"73",
          2716 => x"55",
          2717 => x"55",
          2718 => x"c5",
          2719 => x"88",
          2720 => x"0b",
          2721 => x"9c",
          2722 => x"8b",
          2723 => x"17",
          2724 => x"08",
          2725 => x"52",
          2726 => x"81",
          2727 => x"76",
          2728 => x"51",
          2729 => x"81",
          2730 => x"86",
          2731 => x"12",
          2732 => x"3f",
          2733 => x"08",
          2734 => x"88",
          2735 => x"f3",
          2736 => x"70",
          2737 => x"80",
          2738 => x"51",
          2739 => x"af",
          2740 => x"81",
          2741 => x"dc",
          2742 => x"74",
          2743 => x"38",
          2744 => x"88",
          2745 => x"39",
          2746 => x"80",
          2747 => x"56",
          2748 => x"af",
          2749 => x"06",
          2750 => x"56",
          2751 => x"32",
          2752 => x"80",
          2753 => x"51",
          2754 => x"dc",
          2755 => x"1c",
          2756 => x"33",
          2757 => x"9f",
          2758 => x"ff",
          2759 => x"1c",
          2760 => x"7a",
          2761 => x"3f",
          2762 => x"08",
          2763 => x"39",
          2764 => x"a0",
          2765 => x"5e",
          2766 => x"52",
          2767 => x"ff",
          2768 => x"59",
          2769 => x"33",
          2770 => x"ae",
          2771 => x"06",
          2772 => x"78",
          2773 => x"81",
          2774 => x"32",
          2775 => x"9f",
          2776 => x"26",
          2777 => x"53",
          2778 => x"73",
          2779 => x"17",
          2780 => x"34",
          2781 => x"db",
          2782 => x"32",
          2783 => x"9f",
          2784 => x"54",
          2785 => x"2e",
          2786 => x"80",
          2787 => x"75",
          2788 => x"bd",
          2789 => x"7e",
          2790 => x"a0",
          2791 => x"bd",
          2792 => x"82",
          2793 => x"18",
          2794 => x"1a",
          2795 => x"a0",
          2796 => x"fc",
          2797 => x"32",
          2798 => x"80",
          2799 => x"30",
          2800 => x"71",
          2801 => x"51",
          2802 => x"55",
          2803 => x"ac",
          2804 => x"81",
          2805 => x"78",
          2806 => x"51",
          2807 => x"af",
          2808 => x"06",
          2809 => x"55",
          2810 => x"32",
          2811 => x"80",
          2812 => x"51",
          2813 => x"db",
          2814 => x"39",
          2815 => x"09",
          2816 => x"38",
          2817 => x"7c",
          2818 => x"54",
          2819 => x"a2",
          2820 => x"32",
          2821 => x"ae",
          2822 => x"72",
          2823 => x"9f",
          2824 => x"51",
          2825 => x"74",
          2826 => x"88",
          2827 => x"fe",
          2828 => x"98",
          2829 => x"80",
          2830 => x"75",
          2831 => x"81",
          2832 => x"33",
          2833 => x"51",
          2834 => x"81",
          2835 => x"80",
          2836 => x"78",
          2837 => x"81",
          2838 => x"5a",
          2839 => x"d2",
          2840 => x"84",
          2841 => x"80",
          2842 => x"1c",
          2843 => x"27",
          2844 => x"79",
          2845 => x"74",
          2846 => x"7a",
          2847 => x"74",
          2848 => x"39",
          2849 => x"c2",
          2850 => x"fe",
          2851 => x"84",
          2852 => x"ff",
          2853 => x"73",
          2854 => x"38",
          2855 => x"81",
          2856 => x"54",
          2857 => x"75",
          2858 => x"17",
          2859 => x"39",
          2860 => x"0c",
          2861 => x"99",
          2862 => x"54",
          2863 => x"2e",
          2864 => x"84",
          2865 => x"34",
          2866 => x"76",
          2867 => x"8b",
          2868 => x"81",
          2869 => x"56",
          2870 => x"80",
          2871 => x"1b",
          2872 => x"08",
          2873 => x"51",
          2874 => x"81",
          2875 => x"56",
          2876 => x"08",
          2877 => x"98",
          2878 => x"76",
          2879 => x"3f",
          2880 => x"08",
          2881 => x"84",
          2882 => x"38",
          2883 => x"70",
          2884 => x"73",
          2885 => x"be",
          2886 => x"33",
          2887 => x"73",
          2888 => x"8b",
          2889 => x"83",
          2890 => x"06",
          2891 => x"73",
          2892 => x"53",
          2893 => x"51",
          2894 => x"81",
          2895 => x"80",
          2896 => x"75",
          2897 => x"f3",
          2898 => x"9f",
          2899 => x"1c",
          2900 => x"74",
          2901 => x"38",
          2902 => x"09",
          2903 => x"e7",
          2904 => x"2a",
          2905 => x"77",
          2906 => x"51",
          2907 => x"2e",
          2908 => x"81",
          2909 => x"80",
          2910 => x"38",
          2911 => x"ab",
          2912 => x"55",
          2913 => x"75",
          2914 => x"73",
          2915 => x"55",
          2916 => x"82",
          2917 => x"06",
          2918 => x"ab",
          2919 => x"33",
          2920 => x"70",
          2921 => x"55",
          2922 => x"2e",
          2923 => x"1b",
          2924 => x"06",
          2925 => x"52",
          2926 => x"db",
          2927 => x"84",
          2928 => x"0c",
          2929 => x"74",
          2930 => x"0c",
          2931 => x"04",
          2932 => x"7c",
          2933 => x"08",
          2934 => x"55",
          2935 => x"59",
          2936 => x"81",
          2937 => x"70",
          2938 => x"33",
          2939 => x"52",
          2940 => x"2e",
          2941 => x"ee",
          2942 => x"2e",
          2943 => x"81",
          2944 => x"33",
          2945 => x"81",
          2946 => x"52",
          2947 => x"26",
          2948 => x"14",
          2949 => x"06",
          2950 => x"52",
          2951 => x"80",
          2952 => x"0b",
          2953 => x"59",
          2954 => x"7a",
          2955 => x"70",
          2956 => x"33",
          2957 => x"05",
          2958 => x"9f",
          2959 => x"53",
          2960 => x"89",
          2961 => x"70",
          2962 => x"54",
          2963 => x"12",
          2964 => x"26",
          2965 => x"12",
          2966 => x"06",
          2967 => x"30",
          2968 => x"51",
          2969 => x"2e",
          2970 => x"85",
          2971 => x"be",
          2972 => x"74",
          2973 => x"30",
          2974 => x"9f",
          2975 => x"2a",
          2976 => x"54",
          2977 => x"2e",
          2978 => x"15",
          2979 => x"55",
          2980 => x"ff",
          2981 => x"39",
          2982 => x"86",
          2983 => x"7c",
          2984 => x"51",
          2985 => x"d3",
          2986 => x"70",
          2987 => x"0c",
          2988 => x"04",
          2989 => x"78",
          2990 => x"83",
          2991 => x"0b",
          2992 => x"79",
          2993 => x"e2",
          2994 => x"55",
          2995 => x"08",
          2996 => x"84",
          2997 => x"df",
          2998 => x"d3",
          2999 => x"ff",
          3000 => x"83",
          3001 => x"d4",
          3002 => x"81",
          3003 => x"38",
          3004 => x"17",
          3005 => x"74",
          3006 => x"09",
          3007 => x"38",
          3008 => x"81",
          3009 => x"30",
          3010 => x"79",
          3011 => x"54",
          3012 => x"74",
          3013 => x"09",
          3014 => x"38",
          3015 => x"c2",
          3016 => x"ea",
          3017 => x"b1",
          3018 => x"84",
          3019 => x"d3",
          3020 => x"2e",
          3021 => x"53",
          3022 => x"52",
          3023 => x"51",
          3024 => x"81",
          3025 => x"55",
          3026 => x"08",
          3027 => x"38",
          3028 => x"81",
          3029 => x"88",
          3030 => x"f2",
          3031 => x"02",
          3032 => x"cb",
          3033 => x"55",
          3034 => x"60",
          3035 => x"3f",
          3036 => x"08",
          3037 => x"80",
          3038 => x"84",
          3039 => x"fc",
          3040 => x"84",
          3041 => x"81",
          3042 => x"70",
          3043 => x"8c",
          3044 => x"2e",
          3045 => x"73",
          3046 => x"81",
          3047 => x"33",
          3048 => x"80",
          3049 => x"81",
          3050 => x"d7",
          3051 => x"d3",
          3052 => x"ff",
          3053 => x"06",
          3054 => x"98",
          3055 => x"2e",
          3056 => x"74",
          3057 => x"81",
          3058 => x"8a",
          3059 => x"ac",
          3060 => x"39",
          3061 => x"77",
          3062 => x"81",
          3063 => x"33",
          3064 => x"3f",
          3065 => x"08",
          3066 => x"70",
          3067 => x"55",
          3068 => x"86",
          3069 => x"80",
          3070 => x"74",
          3071 => x"81",
          3072 => x"8a",
          3073 => x"f4",
          3074 => x"53",
          3075 => x"fd",
          3076 => x"d3",
          3077 => x"ff",
          3078 => x"82",
          3079 => x"06",
          3080 => x"8c",
          3081 => x"58",
          3082 => x"f6",
          3083 => x"58",
          3084 => x"2e",
          3085 => x"fa",
          3086 => x"e8",
          3087 => x"84",
          3088 => x"78",
          3089 => x"5a",
          3090 => x"90",
          3091 => x"75",
          3092 => x"38",
          3093 => x"3d",
          3094 => x"70",
          3095 => x"08",
          3096 => x"7a",
          3097 => x"38",
          3098 => x"51",
          3099 => x"81",
          3100 => x"81",
          3101 => x"81",
          3102 => x"38",
          3103 => x"83",
          3104 => x"38",
          3105 => x"84",
          3106 => x"38",
          3107 => x"81",
          3108 => x"38",
          3109 => x"db",
          3110 => x"d3",
          3111 => x"ff",
          3112 => x"72",
          3113 => x"09",
          3114 => x"d0",
          3115 => x"14",
          3116 => x"3f",
          3117 => x"08",
          3118 => x"06",
          3119 => x"38",
          3120 => x"51",
          3121 => x"81",
          3122 => x"58",
          3123 => x"0c",
          3124 => x"33",
          3125 => x"80",
          3126 => x"ff",
          3127 => x"ff",
          3128 => x"55",
          3129 => x"81",
          3130 => x"38",
          3131 => x"06",
          3132 => x"80",
          3133 => x"52",
          3134 => x"8a",
          3135 => x"80",
          3136 => x"ff",
          3137 => x"53",
          3138 => x"86",
          3139 => x"83",
          3140 => x"c5",
          3141 => x"f5",
          3142 => x"84",
          3143 => x"d3",
          3144 => x"15",
          3145 => x"06",
          3146 => x"76",
          3147 => x"80",
          3148 => x"da",
          3149 => x"d3",
          3150 => x"ff",
          3151 => x"74",
          3152 => x"d4",
          3153 => x"dc",
          3154 => x"84",
          3155 => x"c2",
          3156 => x"b9",
          3157 => x"84",
          3158 => x"ff",
          3159 => x"56",
          3160 => x"83",
          3161 => x"14",
          3162 => x"71",
          3163 => x"5a",
          3164 => x"26",
          3165 => x"8a",
          3166 => x"74",
          3167 => x"ff",
          3168 => x"81",
          3169 => x"55",
          3170 => x"08",
          3171 => x"ec",
          3172 => x"84",
          3173 => x"ff",
          3174 => x"83",
          3175 => x"74",
          3176 => x"26",
          3177 => x"57",
          3178 => x"26",
          3179 => x"57",
          3180 => x"56",
          3181 => x"82",
          3182 => x"15",
          3183 => x"0c",
          3184 => x"0c",
          3185 => x"a4",
          3186 => x"1d",
          3187 => x"54",
          3188 => x"2e",
          3189 => x"af",
          3190 => x"14",
          3191 => x"3f",
          3192 => x"08",
          3193 => x"06",
          3194 => x"72",
          3195 => x"79",
          3196 => x"80",
          3197 => x"d9",
          3198 => x"d3",
          3199 => x"15",
          3200 => x"2b",
          3201 => x"8d",
          3202 => x"2e",
          3203 => x"77",
          3204 => x"0c",
          3205 => x"76",
          3206 => x"38",
          3207 => x"70",
          3208 => x"81",
          3209 => x"53",
          3210 => x"89",
          3211 => x"56",
          3212 => x"08",
          3213 => x"38",
          3214 => x"15",
          3215 => x"8c",
          3216 => x"80",
          3217 => x"34",
          3218 => x"09",
          3219 => x"92",
          3220 => x"14",
          3221 => x"3f",
          3222 => x"08",
          3223 => x"06",
          3224 => x"2e",
          3225 => x"80",
          3226 => x"1b",
          3227 => x"db",
          3228 => x"d3",
          3229 => x"ea",
          3230 => x"84",
          3231 => x"34",
          3232 => x"51",
          3233 => x"81",
          3234 => x"83",
          3235 => x"53",
          3236 => x"d5",
          3237 => x"06",
          3238 => x"b4",
          3239 => x"84",
          3240 => x"84",
          3241 => x"85",
          3242 => x"09",
          3243 => x"38",
          3244 => x"51",
          3245 => x"81",
          3246 => x"86",
          3247 => x"f2",
          3248 => x"06",
          3249 => x"9c",
          3250 => x"d8",
          3251 => x"84",
          3252 => x"0c",
          3253 => x"51",
          3254 => x"81",
          3255 => x"8c",
          3256 => x"74",
          3257 => x"b0",
          3258 => x"53",
          3259 => x"b0",
          3260 => x"15",
          3261 => x"94",
          3262 => x"56",
          3263 => x"84",
          3264 => x"0d",
          3265 => x"0d",
          3266 => x"55",
          3267 => x"b9",
          3268 => x"53",
          3269 => x"b1",
          3270 => x"52",
          3271 => x"a9",
          3272 => x"22",
          3273 => x"57",
          3274 => x"2e",
          3275 => x"99",
          3276 => x"33",
          3277 => x"3f",
          3278 => x"08",
          3279 => x"71",
          3280 => x"74",
          3281 => x"83",
          3282 => x"78",
          3283 => x"52",
          3284 => x"84",
          3285 => x"0d",
          3286 => x"0d",
          3287 => x"33",
          3288 => x"3d",
          3289 => x"56",
          3290 => x"8b",
          3291 => x"81",
          3292 => x"24",
          3293 => x"d3",
          3294 => x"29",
          3295 => x"05",
          3296 => x"55",
          3297 => x"84",
          3298 => x"34",
          3299 => x"80",
          3300 => x"80",
          3301 => x"75",
          3302 => x"75",
          3303 => x"38",
          3304 => x"3d",
          3305 => x"05",
          3306 => x"3f",
          3307 => x"08",
          3308 => x"d3",
          3309 => x"3d",
          3310 => x"3d",
          3311 => x"84",
          3312 => x"05",
          3313 => x"89",
          3314 => x"2e",
          3315 => x"77",
          3316 => x"54",
          3317 => x"05",
          3318 => x"84",
          3319 => x"f6",
          3320 => x"d3",
          3321 => x"81",
          3322 => x"84",
          3323 => x"5c",
          3324 => x"3d",
          3325 => x"ed",
          3326 => x"d3",
          3327 => x"81",
          3328 => x"92",
          3329 => x"d7",
          3330 => x"98",
          3331 => x"73",
          3332 => x"38",
          3333 => x"9c",
          3334 => x"80",
          3335 => x"38",
          3336 => x"95",
          3337 => x"2e",
          3338 => x"aa",
          3339 => x"ea",
          3340 => x"d3",
          3341 => x"9e",
          3342 => x"05",
          3343 => x"54",
          3344 => x"38",
          3345 => x"70",
          3346 => x"54",
          3347 => x"8e",
          3348 => x"83",
          3349 => x"88",
          3350 => x"83",
          3351 => x"83",
          3352 => x"06",
          3353 => x"80",
          3354 => x"38",
          3355 => x"51",
          3356 => x"81",
          3357 => x"56",
          3358 => x"0a",
          3359 => x"05",
          3360 => x"3f",
          3361 => x"0b",
          3362 => x"80",
          3363 => x"7a",
          3364 => x"3f",
          3365 => x"9c",
          3366 => x"d1",
          3367 => x"81",
          3368 => x"34",
          3369 => x"80",
          3370 => x"b0",
          3371 => x"54",
          3372 => x"52",
          3373 => x"05",
          3374 => x"3f",
          3375 => x"08",
          3376 => x"84",
          3377 => x"38",
          3378 => x"82",
          3379 => x"b2",
          3380 => x"84",
          3381 => x"06",
          3382 => x"73",
          3383 => x"38",
          3384 => x"ad",
          3385 => x"2a",
          3386 => x"51",
          3387 => x"2e",
          3388 => x"81",
          3389 => x"80",
          3390 => x"87",
          3391 => x"39",
          3392 => x"51",
          3393 => x"81",
          3394 => x"7b",
          3395 => x"12",
          3396 => x"81",
          3397 => x"81",
          3398 => x"83",
          3399 => x"06",
          3400 => x"80",
          3401 => x"77",
          3402 => x"58",
          3403 => x"08",
          3404 => x"63",
          3405 => x"63",
          3406 => x"57",
          3407 => x"81",
          3408 => x"81",
          3409 => x"88",
          3410 => x"9c",
          3411 => x"d2",
          3412 => x"d3",
          3413 => x"d3",
          3414 => x"1b",
          3415 => x"0c",
          3416 => x"22",
          3417 => x"77",
          3418 => x"80",
          3419 => x"34",
          3420 => x"1a",
          3421 => x"94",
          3422 => x"85",
          3423 => x"06",
          3424 => x"80",
          3425 => x"38",
          3426 => x"08",
          3427 => x"84",
          3428 => x"84",
          3429 => x"0c",
          3430 => x"70",
          3431 => x"52",
          3432 => x"39",
          3433 => x"51",
          3434 => x"81",
          3435 => x"57",
          3436 => x"08",
          3437 => x"38",
          3438 => x"d3",
          3439 => x"2e",
          3440 => x"83",
          3441 => x"75",
          3442 => x"74",
          3443 => x"07",
          3444 => x"54",
          3445 => x"8a",
          3446 => x"75",
          3447 => x"73",
          3448 => x"98",
          3449 => x"a9",
          3450 => x"ff",
          3451 => x"80",
          3452 => x"76",
          3453 => x"d6",
          3454 => x"d3",
          3455 => x"38",
          3456 => x"39",
          3457 => x"81",
          3458 => x"05",
          3459 => x"84",
          3460 => x"0c",
          3461 => x"81",
          3462 => x"97",
          3463 => x"f2",
          3464 => x"63",
          3465 => x"40",
          3466 => x"7e",
          3467 => x"fc",
          3468 => x"51",
          3469 => x"81",
          3470 => x"55",
          3471 => x"08",
          3472 => x"19",
          3473 => x"80",
          3474 => x"74",
          3475 => x"39",
          3476 => x"81",
          3477 => x"56",
          3478 => x"82",
          3479 => x"39",
          3480 => x"1a",
          3481 => x"82",
          3482 => x"0b",
          3483 => x"81",
          3484 => x"39",
          3485 => x"94",
          3486 => x"55",
          3487 => x"83",
          3488 => x"7b",
          3489 => x"89",
          3490 => x"08",
          3491 => x"06",
          3492 => x"81",
          3493 => x"8a",
          3494 => x"05",
          3495 => x"06",
          3496 => x"a8",
          3497 => x"38",
          3498 => x"55",
          3499 => x"19",
          3500 => x"51",
          3501 => x"81",
          3502 => x"55",
          3503 => x"ff",
          3504 => x"ff",
          3505 => x"38",
          3506 => x"0c",
          3507 => x"52",
          3508 => x"cb",
          3509 => x"84",
          3510 => x"ff",
          3511 => x"d3",
          3512 => x"7c",
          3513 => x"57",
          3514 => x"80",
          3515 => x"1a",
          3516 => x"22",
          3517 => x"75",
          3518 => x"38",
          3519 => x"58",
          3520 => x"53",
          3521 => x"1b",
          3522 => x"88",
          3523 => x"84",
          3524 => x"38",
          3525 => x"33",
          3526 => x"80",
          3527 => x"b0",
          3528 => x"31",
          3529 => x"27",
          3530 => x"80",
          3531 => x"52",
          3532 => x"77",
          3533 => x"7d",
          3534 => x"e0",
          3535 => x"2b",
          3536 => x"76",
          3537 => x"94",
          3538 => x"ff",
          3539 => x"71",
          3540 => x"7b",
          3541 => x"38",
          3542 => x"19",
          3543 => x"51",
          3544 => x"81",
          3545 => x"fe",
          3546 => x"53",
          3547 => x"83",
          3548 => x"b4",
          3549 => x"51",
          3550 => x"7b",
          3551 => x"08",
          3552 => x"76",
          3553 => x"08",
          3554 => x"0c",
          3555 => x"f3",
          3556 => x"75",
          3557 => x"0c",
          3558 => x"04",
          3559 => x"60",
          3560 => x"40",
          3561 => x"80",
          3562 => x"3d",
          3563 => x"77",
          3564 => x"3f",
          3565 => x"08",
          3566 => x"84",
          3567 => x"91",
          3568 => x"74",
          3569 => x"38",
          3570 => x"b8",
          3571 => x"33",
          3572 => x"70",
          3573 => x"56",
          3574 => x"74",
          3575 => x"a4",
          3576 => x"82",
          3577 => x"34",
          3578 => x"98",
          3579 => x"91",
          3580 => x"56",
          3581 => x"94",
          3582 => x"11",
          3583 => x"76",
          3584 => x"75",
          3585 => x"80",
          3586 => x"38",
          3587 => x"70",
          3588 => x"56",
          3589 => x"fd",
          3590 => x"11",
          3591 => x"77",
          3592 => x"5c",
          3593 => x"38",
          3594 => x"88",
          3595 => x"74",
          3596 => x"52",
          3597 => x"18",
          3598 => x"51",
          3599 => x"81",
          3600 => x"55",
          3601 => x"08",
          3602 => x"ab",
          3603 => x"2e",
          3604 => x"74",
          3605 => x"95",
          3606 => x"19",
          3607 => x"08",
          3608 => x"88",
          3609 => x"55",
          3610 => x"9c",
          3611 => x"09",
          3612 => x"38",
          3613 => x"c1",
          3614 => x"84",
          3615 => x"38",
          3616 => x"52",
          3617 => x"97",
          3618 => x"84",
          3619 => x"fe",
          3620 => x"d3",
          3621 => x"7c",
          3622 => x"57",
          3623 => x"80",
          3624 => x"1b",
          3625 => x"22",
          3626 => x"75",
          3627 => x"38",
          3628 => x"59",
          3629 => x"53",
          3630 => x"1a",
          3631 => x"be",
          3632 => x"84",
          3633 => x"38",
          3634 => x"08",
          3635 => x"56",
          3636 => x"9b",
          3637 => x"53",
          3638 => x"77",
          3639 => x"7d",
          3640 => x"16",
          3641 => x"3f",
          3642 => x"0b",
          3643 => x"78",
          3644 => x"80",
          3645 => x"18",
          3646 => x"08",
          3647 => x"7e",
          3648 => x"3f",
          3649 => x"08",
          3650 => x"7e",
          3651 => x"0c",
          3652 => x"19",
          3653 => x"08",
          3654 => x"84",
          3655 => x"57",
          3656 => x"27",
          3657 => x"56",
          3658 => x"52",
          3659 => x"f9",
          3660 => x"84",
          3661 => x"38",
          3662 => x"52",
          3663 => x"83",
          3664 => x"b4",
          3665 => x"d4",
          3666 => x"81",
          3667 => x"34",
          3668 => x"7e",
          3669 => x"0c",
          3670 => x"1a",
          3671 => x"94",
          3672 => x"1b",
          3673 => x"5e",
          3674 => x"27",
          3675 => x"55",
          3676 => x"0c",
          3677 => x"90",
          3678 => x"c0",
          3679 => x"90",
          3680 => x"56",
          3681 => x"84",
          3682 => x"0d",
          3683 => x"0d",
          3684 => x"fc",
          3685 => x"52",
          3686 => x"3f",
          3687 => x"08",
          3688 => x"84",
          3689 => x"38",
          3690 => x"70",
          3691 => x"81",
          3692 => x"55",
          3693 => x"80",
          3694 => x"16",
          3695 => x"51",
          3696 => x"81",
          3697 => x"57",
          3698 => x"08",
          3699 => x"a4",
          3700 => x"11",
          3701 => x"55",
          3702 => x"16",
          3703 => x"08",
          3704 => x"75",
          3705 => x"e8",
          3706 => x"08",
          3707 => x"51",
          3708 => x"82",
          3709 => x"52",
          3710 => x"c9",
          3711 => x"52",
          3712 => x"c9",
          3713 => x"54",
          3714 => x"15",
          3715 => x"cc",
          3716 => x"d3",
          3717 => x"17",
          3718 => x"06",
          3719 => x"90",
          3720 => x"81",
          3721 => x"8a",
          3722 => x"fc",
          3723 => x"70",
          3724 => x"d9",
          3725 => x"84",
          3726 => x"d3",
          3727 => x"38",
          3728 => x"05",
          3729 => x"f1",
          3730 => x"d3",
          3731 => x"81",
          3732 => x"87",
          3733 => x"84",
          3734 => x"72",
          3735 => x"0c",
          3736 => x"04",
          3737 => x"84",
          3738 => x"e4",
          3739 => x"80",
          3740 => x"84",
          3741 => x"38",
          3742 => x"08",
          3743 => x"34",
          3744 => x"81",
          3745 => x"83",
          3746 => x"ef",
          3747 => x"53",
          3748 => x"05",
          3749 => x"51",
          3750 => x"81",
          3751 => x"55",
          3752 => x"08",
          3753 => x"76",
          3754 => x"93",
          3755 => x"51",
          3756 => x"81",
          3757 => x"55",
          3758 => x"08",
          3759 => x"80",
          3760 => x"70",
          3761 => x"56",
          3762 => x"89",
          3763 => x"94",
          3764 => x"b2",
          3765 => x"05",
          3766 => x"2a",
          3767 => x"51",
          3768 => x"80",
          3769 => x"76",
          3770 => x"52",
          3771 => x"3f",
          3772 => x"08",
          3773 => x"8e",
          3774 => x"84",
          3775 => x"09",
          3776 => x"38",
          3777 => x"81",
          3778 => x"93",
          3779 => x"e4",
          3780 => x"6f",
          3781 => x"7a",
          3782 => x"9e",
          3783 => x"05",
          3784 => x"51",
          3785 => x"81",
          3786 => x"57",
          3787 => x"08",
          3788 => x"7b",
          3789 => x"94",
          3790 => x"55",
          3791 => x"73",
          3792 => x"ed",
          3793 => x"93",
          3794 => x"55",
          3795 => x"81",
          3796 => x"57",
          3797 => x"08",
          3798 => x"68",
          3799 => x"c9",
          3800 => x"d3",
          3801 => x"81",
          3802 => x"82",
          3803 => x"52",
          3804 => x"a3",
          3805 => x"84",
          3806 => x"52",
          3807 => x"b8",
          3808 => x"84",
          3809 => x"d3",
          3810 => x"a2",
          3811 => x"74",
          3812 => x"3f",
          3813 => x"08",
          3814 => x"84",
          3815 => x"69",
          3816 => x"d9",
          3817 => x"81",
          3818 => x"2e",
          3819 => x"52",
          3820 => x"cf",
          3821 => x"84",
          3822 => x"d3",
          3823 => x"2e",
          3824 => x"84",
          3825 => x"06",
          3826 => x"57",
          3827 => x"76",
          3828 => x"9e",
          3829 => x"05",
          3830 => x"dc",
          3831 => x"90",
          3832 => x"81",
          3833 => x"56",
          3834 => x"80",
          3835 => x"02",
          3836 => x"81",
          3837 => x"70",
          3838 => x"56",
          3839 => x"81",
          3840 => x"78",
          3841 => x"38",
          3842 => x"99",
          3843 => x"81",
          3844 => x"18",
          3845 => x"18",
          3846 => x"58",
          3847 => x"33",
          3848 => x"ee",
          3849 => x"6f",
          3850 => x"af",
          3851 => x"8d",
          3852 => x"2e",
          3853 => x"8a",
          3854 => x"6f",
          3855 => x"af",
          3856 => x"0b",
          3857 => x"33",
          3858 => x"81",
          3859 => x"70",
          3860 => x"52",
          3861 => x"56",
          3862 => x"8d",
          3863 => x"70",
          3864 => x"51",
          3865 => x"f5",
          3866 => x"54",
          3867 => x"a7",
          3868 => x"74",
          3869 => x"38",
          3870 => x"73",
          3871 => x"81",
          3872 => x"81",
          3873 => x"39",
          3874 => x"81",
          3875 => x"74",
          3876 => x"81",
          3877 => x"91",
          3878 => x"6e",
          3879 => x"59",
          3880 => x"7a",
          3881 => x"5c",
          3882 => x"26",
          3883 => x"7a",
          3884 => x"d3",
          3885 => x"3d",
          3886 => x"3d",
          3887 => x"8d",
          3888 => x"54",
          3889 => x"55",
          3890 => x"81",
          3891 => x"53",
          3892 => x"08",
          3893 => x"91",
          3894 => x"72",
          3895 => x"8c",
          3896 => x"73",
          3897 => x"38",
          3898 => x"70",
          3899 => x"81",
          3900 => x"57",
          3901 => x"73",
          3902 => x"08",
          3903 => x"94",
          3904 => x"75",
          3905 => x"97",
          3906 => x"11",
          3907 => x"2b",
          3908 => x"73",
          3909 => x"38",
          3910 => x"16",
          3911 => x"d8",
          3912 => x"84",
          3913 => x"78",
          3914 => x"55",
          3915 => x"c8",
          3916 => x"84",
          3917 => x"96",
          3918 => x"70",
          3919 => x"94",
          3920 => x"71",
          3921 => x"08",
          3922 => x"53",
          3923 => x"15",
          3924 => x"a6",
          3925 => x"74",
          3926 => x"3f",
          3927 => x"08",
          3928 => x"84",
          3929 => x"81",
          3930 => x"d3",
          3931 => x"2e",
          3932 => x"81",
          3933 => x"88",
          3934 => x"98",
          3935 => x"80",
          3936 => x"38",
          3937 => x"80",
          3938 => x"77",
          3939 => x"08",
          3940 => x"0c",
          3941 => x"70",
          3942 => x"81",
          3943 => x"5a",
          3944 => x"2e",
          3945 => x"52",
          3946 => x"f9",
          3947 => x"84",
          3948 => x"d3",
          3949 => x"38",
          3950 => x"08",
          3951 => x"73",
          3952 => x"c7",
          3953 => x"d3",
          3954 => x"73",
          3955 => x"38",
          3956 => x"af",
          3957 => x"73",
          3958 => x"27",
          3959 => x"98",
          3960 => x"a0",
          3961 => x"08",
          3962 => x"0c",
          3963 => x"06",
          3964 => x"2e",
          3965 => x"52",
          3966 => x"a3",
          3967 => x"84",
          3968 => x"82",
          3969 => x"34",
          3970 => x"c4",
          3971 => x"91",
          3972 => x"53",
          3973 => x"89",
          3974 => x"84",
          3975 => x"94",
          3976 => x"8c",
          3977 => x"27",
          3978 => x"8c",
          3979 => x"15",
          3980 => x"07",
          3981 => x"16",
          3982 => x"ff",
          3983 => x"80",
          3984 => x"77",
          3985 => x"2e",
          3986 => x"9c",
          3987 => x"53",
          3988 => x"84",
          3989 => x"0d",
          3990 => x"0d",
          3991 => x"54",
          3992 => x"81",
          3993 => x"53",
          3994 => x"05",
          3995 => x"84",
          3996 => x"e7",
          3997 => x"84",
          3998 => x"d3",
          3999 => x"ea",
          4000 => x"0c",
          4001 => x"51",
          4002 => x"81",
          4003 => x"55",
          4004 => x"08",
          4005 => x"ab",
          4006 => x"98",
          4007 => x"80",
          4008 => x"38",
          4009 => x"70",
          4010 => x"81",
          4011 => x"57",
          4012 => x"ad",
          4013 => x"08",
          4014 => x"d3",
          4015 => x"d3",
          4016 => x"17",
          4017 => x"86",
          4018 => x"17",
          4019 => x"75",
          4020 => x"3f",
          4021 => x"08",
          4022 => x"2e",
          4023 => x"85",
          4024 => x"86",
          4025 => x"2e",
          4026 => x"76",
          4027 => x"73",
          4028 => x"0c",
          4029 => x"04",
          4030 => x"76",
          4031 => x"05",
          4032 => x"53",
          4033 => x"81",
          4034 => x"87",
          4035 => x"84",
          4036 => x"86",
          4037 => x"fb",
          4038 => x"79",
          4039 => x"05",
          4040 => x"56",
          4041 => x"3f",
          4042 => x"08",
          4043 => x"84",
          4044 => x"38",
          4045 => x"81",
          4046 => x"52",
          4047 => x"f8",
          4048 => x"84",
          4049 => x"ca",
          4050 => x"84",
          4051 => x"51",
          4052 => x"81",
          4053 => x"53",
          4054 => x"08",
          4055 => x"81",
          4056 => x"80",
          4057 => x"81",
          4058 => x"a6",
          4059 => x"73",
          4060 => x"3f",
          4061 => x"51",
          4062 => x"81",
          4063 => x"84",
          4064 => x"70",
          4065 => x"2c",
          4066 => x"84",
          4067 => x"51",
          4068 => x"81",
          4069 => x"87",
          4070 => x"ee",
          4071 => x"57",
          4072 => x"3d",
          4073 => x"3d",
          4074 => x"af",
          4075 => x"84",
          4076 => x"d3",
          4077 => x"38",
          4078 => x"51",
          4079 => x"81",
          4080 => x"55",
          4081 => x"08",
          4082 => x"80",
          4083 => x"70",
          4084 => x"58",
          4085 => x"85",
          4086 => x"8d",
          4087 => x"2e",
          4088 => x"52",
          4089 => x"be",
          4090 => x"d3",
          4091 => x"3d",
          4092 => x"3d",
          4093 => x"55",
          4094 => x"92",
          4095 => x"52",
          4096 => x"de",
          4097 => x"d3",
          4098 => x"81",
          4099 => x"82",
          4100 => x"74",
          4101 => x"98",
          4102 => x"11",
          4103 => x"59",
          4104 => x"75",
          4105 => x"38",
          4106 => x"81",
          4107 => x"5b",
          4108 => x"82",
          4109 => x"39",
          4110 => x"08",
          4111 => x"59",
          4112 => x"09",
          4113 => x"38",
          4114 => x"57",
          4115 => x"3d",
          4116 => x"c1",
          4117 => x"d3",
          4118 => x"2e",
          4119 => x"d3",
          4120 => x"2e",
          4121 => x"d3",
          4122 => x"70",
          4123 => x"08",
          4124 => x"7a",
          4125 => x"7f",
          4126 => x"54",
          4127 => x"77",
          4128 => x"80",
          4129 => x"15",
          4130 => x"84",
          4131 => x"75",
          4132 => x"52",
          4133 => x"52",
          4134 => x"8d",
          4135 => x"84",
          4136 => x"d3",
          4137 => x"d6",
          4138 => x"33",
          4139 => x"1a",
          4140 => x"54",
          4141 => x"09",
          4142 => x"38",
          4143 => x"ff",
          4144 => x"81",
          4145 => x"83",
          4146 => x"70",
          4147 => x"25",
          4148 => x"59",
          4149 => x"9b",
          4150 => x"51",
          4151 => x"3f",
          4152 => x"08",
          4153 => x"70",
          4154 => x"25",
          4155 => x"59",
          4156 => x"75",
          4157 => x"7a",
          4158 => x"ff",
          4159 => x"7c",
          4160 => x"90",
          4161 => x"11",
          4162 => x"56",
          4163 => x"15",
          4164 => x"d3",
          4165 => x"3d",
          4166 => x"3d",
          4167 => x"3d",
          4168 => x"70",
          4169 => x"dd",
          4170 => x"84",
          4171 => x"d3",
          4172 => x"a8",
          4173 => x"33",
          4174 => x"a0",
          4175 => x"33",
          4176 => x"70",
          4177 => x"55",
          4178 => x"73",
          4179 => x"8e",
          4180 => x"08",
          4181 => x"18",
          4182 => x"80",
          4183 => x"38",
          4184 => x"08",
          4185 => x"08",
          4186 => x"c4",
          4187 => x"d3",
          4188 => x"88",
          4189 => x"80",
          4190 => x"17",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"08",
          4194 => x"81",
          4195 => x"81",
          4196 => x"84",
          4197 => x"09",
          4198 => x"38",
          4199 => x"39",
          4200 => x"77",
          4201 => x"84",
          4202 => x"08",
          4203 => x"98",
          4204 => x"81",
          4205 => x"52",
          4206 => x"bd",
          4207 => x"84",
          4208 => x"17",
          4209 => x"0c",
          4210 => x"80",
          4211 => x"73",
          4212 => x"75",
          4213 => x"38",
          4214 => x"34",
          4215 => x"81",
          4216 => x"89",
          4217 => x"e2",
          4218 => x"53",
          4219 => x"a4",
          4220 => x"3d",
          4221 => x"3f",
          4222 => x"08",
          4223 => x"84",
          4224 => x"38",
          4225 => x"3d",
          4226 => x"3d",
          4227 => x"d1",
          4228 => x"d3",
          4229 => x"81",
          4230 => x"81",
          4231 => x"80",
          4232 => x"70",
          4233 => x"81",
          4234 => x"56",
          4235 => x"81",
          4236 => x"98",
          4237 => x"74",
          4238 => x"38",
          4239 => x"05",
          4240 => x"06",
          4241 => x"55",
          4242 => x"38",
          4243 => x"51",
          4244 => x"81",
          4245 => x"74",
          4246 => x"81",
          4247 => x"56",
          4248 => x"80",
          4249 => x"54",
          4250 => x"08",
          4251 => x"2e",
          4252 => x"73",
          4253 => x"84",
          4254 => x"52",
          4255 => x"52",
          4256 => x"3f",
          4257 => x"08",
          4258 => x"84",
          4259 => x"38",
          4260 => x"08",
          4261 => x"cc",
          4262 => x"d3",
          4263 => x"81",
          4264 => x"86",
          4265 => x"80",
          4266 => x"d3",
          4267 => x"2e",
          4268 => x"d3",
          4269 => x"c0",
          4270 => x"ce",
          4271 => x"d3",
          4272 => x"d3",
          4273 => x"70",
          4274 => x"08",
          4275 => x"51",
          4276 => x"80",
          4277 => x"73",
          4278 => x"38",
          4279 => x"52",
          4280 => x"95",
          4281 => x"84",
          4282 => x"8c",
          4283 => x"ff",
          4284 => x"81",
          4285 => x"55",
          4286 => x"84",
          4287 => x"0d",
          4288 => x"0d",
          4289 => x"3d",
          4290 => x"9a",
          4291 => x"cb",
          4292 => x"84",
          4293 => x"d3",
          4294 => x"b0",
          4295 => x"69",
          4296 => x"70",
          4297 => x"97",
          4298 => x"84",
          4299 => x"d3",
          4300 => x"38",
          4301 => x"94",
          4302 => x"84",
          4303 => x"09",
          4304 => x"88",
          4305 => x"df",
          4306 => x"85",
          4307 => x"51",
          4308 => x"74",
          4309 => x"78",
          4310 => x"8a",
          4311 => x"57",
          4312 => x"81",
          4313 => x"75",
          4314 => x"d3",
          4315 => x"38",
          4316 => x"d3",
          4317 => x"2e",
          4318 => x"83",
          4319 => x"81",
          4320 => x"ff",
          4321 => x"06",
          4322 => x"54",
          4323 => x"73",
          4324 => x"81",
          4325 => x"52",
          4326 => x"a4",
          4327 => x"84",
          4328 => x"d3",
          4329 => x"9a",
          4330 => x"a0",
          4331 => x"51",
          4332 => x"3f",
          4333 => x"0b",
          4334 => x"78",
          4335 => x"bf",
          4336 => x"88",
          4337 => x"80",
          4338 => x"ff",
          4339 => x"75",
          4340 => x"11",
          4341 => x"f8",
          4342 => x"78",
          4343 => x"80",
          4344 => x"ff",
          4345 => x"78",
          4346 => x"80",
          4347 => x"7f",
          4348 => x"d4",
          4349 => x"c9",
          4350 => x"54",
          4351 => x"15",
          4352 => x"cb",
          4353 => x"d3",
          4354 => x"81",
          4355 => x"b2",
          4356 => x"b2",
          4357 => x"96",
          4358 => x"b5",
          4359 => x"53",
          4360 => x"51",
          4361 => x"64",
          4362 => x"8b",
          4363 => x"54",
          4364 => x"15",
          4365 => x"ff",
          4366 => x"81",
          4367 => x"54",
          4368 => x"53",
          4369 => x"51",
          4370 => x"3f",
          4371 => x"84",
          4372 => x"0d",
          4373 => x"0d",
          4374 => x"05",
          4375 => x"3f",
          4376 => x"3d",
          4377 => x"52",
          4378 => x"d5",
          4379 => x"d3",
          4380 => x"81",
          4381 => x"82",
          4382 => x"4d",
          4383 => x"52",
          4384 => x"52",
          4385 => x"3f",
          4386 => x"08",
          4387 => x"84",
          4388 => x"38",
          4389 => x"05",
          4390 => x"06",
          4391 => x"73",
          4392 => x"a0",
          4393 => x"08",
          4394 => x"ff",
          4395 => x"ff",
          4396 => x"ac",
          4397 => x"92",
          4398 => x"54",
          4399 => x"3f",
          4400 => x"52",
          4401 => x"f7",
          4402 => x"84",
          4403 => x"d3",
          4404 => x"38",
          4405 => x"09",
          4406 => x"38",
          4407 => x"08",
          4408 => x"88",
          4409 => x"39",
          4410 => x"08",
          4411 => x"81",
          4412 => x"38",
          4413 => x"b1",
          4414 => x"84",
          4415 => x"d3",
          4416 => x"c8",
          4417 => x"93",
          4418 => x"ff",
          4419 => x"8d",
          4420 => x"b4",
          4421 => x"af",
          4422 => x"17",
          4423 => x"33",
          4424 => x"70",
          4425 => x"55",
          4426 => x"38",
          4427 => x"54",
          4428 => x"34",
          4429 => x"0b",
          4430 => x"8b",
          4431 => x"84",
          4432 => x"06",
          4433 => x"73",
          4434 => x"e5",
          4435 => x"2e",
          4436 => x"75",
          4437 => x"c6",
          4438 => x"d3",
          4439 => x"78",
          4440 => x"bb",
          4441 => x"81",
          4442 => x"80",
          4443 => x"38",
          4444 => x"08",
          4445 => x"ff",
          4446 => x"81",
          4447 => x"79",
          4448 => x"58",
          4449 => x"d3",
          4450 => x"c0",
          4451 => x"33",
          4452 => x"2e",
          4453 => x"99",
          4454 => x"75",
          4455 => x"c6",
          4456 => x"54",
          4457 => x"15",
          4458 => x"81",
          4459 => x"9c",
          4460 => x"c8",
          4461 => x"d3",
          4462 => x"81",
          4463 => x"8c",
          4464 => x"ff",
          4465 => x"81",
          4466 => x"55",
          4467 => x"84",
          4468 => x"0d",
          4469 => x"0d",
          4470 => x"05",
          4471 => x"05",
          4472 => x"33",
          4473 => x"53",
          4474 => x"05",
          4475 => x"51",
          4476 => x"81",
          4477 => x"55",
          4478 => x"08",
          4479 => x"78",
          4480 => x"95",
          4481 => x"51",
          4482 => x"81",
          4483 => x"55",
          4484 => x"08",
          4485 => x"80",
          4486 => x"81",
          4487 => x"86",
          4488 => x"38",
          4489 => x"61",
          4490 => x"12",
          4491 => x"7a",
          4492 => x"51",
          4493 => x"74",
          4494 => x"78",
          4495 => x"83",
          4496 => x"51",
          4497 => x"3f",
          4498 => x"08",
          4499 => x"d3",
          4500 => x"3d",
          4501 => x"3d",
          4502 => x"82",
          4503 => x"d0",
          4504 => x"3d",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"84",
          4508 => x"38",
          4509 => x"52",
          4510 => x"05",
          4511 => x"3f",
          4512 => x"08",
          4513 => x"84",
          4514 => x"02",
          4515 => x"33",
          4516 => x"54",
          4517 => x"a6",
          4518 => x"22",
          4519 => x"71",
          4520 => x"53",
          4521 => x"51",
          4522 => x"3f",
          4523 => x"0b",
          4524 => x"76",
          4525 => x"b8",
          4526 => x"84",
          4527 => x"81",
          4528 => x"93",
          4529 => x"ea",
          4530 => x"6b",
          4531 => x"53",
          4532 => x"05",
          4533 => x"51",
          4534 => x"81",
          4535 => x"81",
          4536 => x"30",
          4537 => x"84",
          4538 => x"25",
          4539 => x"79",
          4540 => x"85",
          4541 => x"75",
          4542 => x"73",
          4543 => x"f9",
          4544 => x"80",
          4545 => x"8d",
          4546 => x"54",
          4547 => x"3f",
          4548 => x"08",
          4549 => x"84",
          4550 => x"38",
          4551 => x"51",
          4552 => x"81",
          4553 => x"57",
          4554 => x"08",
          4555 => x"d3",
          4556 => x"d3",
          4557 => x"5b",
          4558 => x"18",
          4559 => x"18",
          4560 => x"74",
          4561 => x"81",
          4562 => x"78",
          4563 => x"8b",
          4564 => x"54",
          4565 => x"75",
          4566 => x"38",
          4567 => x"1b",
          4568 => x"55",
          4569 => x"2e",
          4570 => x"39",
          4571 => x"09",
          4572 => x"38",
          4573 => x"80",
          4574 => x"70",
          4575 => x"25",
          4576 => x"80",
          4577 => x"38",
          4578 => x"bc",
          4579 => x"11",
          4580 => x"ff",
          4581 => x"81",
          4582 => x"57",
          4583 => x"08",
          4584 => x"70",
          4585 => x"80",
          4586 => x"83",
          4587 => x"80",
          4588 => x"84",
          4589 => x"a7",
          4590 => x"b4",
          4591 => x"ad",
          4592 => x"d3",
          4593 => x"0c",
          4594 => x"84",
          4595 => x"0d",
          4596 => x"0d",
          4597 => x"3d",
          4598 => x"52",
          4599 => x"ce",
          4600 => x"d3",
          4601 => x"d3",
          4602 => x"54",
          4603 => x"08",
          4604 => x"8b",
          4605 => x"8b",
          4606 => x"59",
          4607 => x"3f",
          4608 => x"33",
          4609 => x"06",
          4610 => x"57",
          4611 => x"81",
          4612 => x"58",
          4613 => x"06",
          4614 => x"4e",
          4615 => x"ff",
          4616 => x"81",
          4617 => x"80",
          4618 => x"6c",
          4619 => x"53",
          4620 => x"ae",
          4621 => x"d3",
          4622 => x"2e",
          4623 => x"88",
          4624 => x"6d",
          4625 => x"55",
          4626 => x"d3",
          4627 => x"ff",
          4628 => x"83",
          4629 => x"51",
          4630 => x"26",
          4631 => x"15",
          4632 => x"ff",
          4633 => x"80",
          4634 => x"87",
          4635 => x"f8",
          4636 => x"74",
          4637 => x"38",
          4638 => x"c3",
          4639 => x"ae",
          4640 => x"d3",
          4641 => x"38",
          4642 => x"27",
          4643 => x"89",
          4644 => x"8b",
          4645 => x"27",
          4646 => x"55",
          4647 => x"81",
          4648 => x"8f",
          4649 => x"2a",
          4650 => x"70",
          4651 => x"34",
          4652 => x"74",
          4653 => x"05",
          4654 => x"17",
          4655 => x"70",
          4656 => x"52",
          4657 => x"73",
          4658 => x"c8",
          4659 => x"33",
          4660 => x"73",
          4661 => x"81",
          4662 => x"80",
          4663 => x"02",
          4664 => x"76",
          4665 => x"51",
          4666 => x"2e",
          4667 => x"87",
          4668 => x"57",
          4669 => x"79",
          4670 => x"80",
          4671 => x"70",
          4672 => x"ba",
          4673 => x"d3",
          4674 => x"81",
          4675 => x"80",
          4676 => x"52",
          4677 => x"bf",
          4678 => x"d3",
          4679 => x"81",
          4680 => x"8d",
          4681 => x"c4",
          4682 => x"e5",
          4683 => x"c6",
          4684 => x"84",
          4685 => x"09",
          4686 => x"cc",
          4687 => x"76",
          4688 => x"c4",
          4689 => x"74",
          4690 => x"b0",
          4691 => x"84",
          4692 => x"d3",
          4693 => x"38",
          4694 => x"d3",
          4695 => x"67",
          4696 => x"db",
          4697 => x"88",
          4698 => x"34",
          4699 => x"52",
          4700 => x"ab",
          4701 => x"54",
          4702 => x"15",
          4703 => x"ff",
          4704 => x"81",
          4705 => x"54",
          4706 => x"81",
          4707 => x"9c",
          4708 => x"f2",
          4709 => x"62",
          4710 => x"80",
          4711 => x"93",
          4712 => x"55",
          4713 => x"5e",
          4714 => x"3f",
          4715 => x"08",
          4716 => x"84",
          4717 => x"38",
          4718 => x"58",
          4719 => x"38",
          4720 => x"97",
          4721 => x"08",
          4722 => x"38",
          4723 => x"70",
          4724 => x"81",
          4725 => x"55",
          4726 => x"87",
          4727 => x"39",
          4728 => x"90",
          4729 => x"82",
          4730 => x"8a",
          4731 => x"89",
          4732 => x"7f",
          4733 => x"56",
          4734 => x"3f",
          4735 => x"06",
          4736 => x"72",
          4737 => x"81",
          4738 => x"05",
          4739 => x"7c",
          4740 => x"55",
          4741 => x"27",
          4742 => x"16",
          4743 => x"83",
          4744 => x"76",
          4745 => x"80",
          4746 => x"79",
          4747 => x"99",
          4748 => x"7f",
          4749 => x"14",
          4750 => x"83",
          4751 => x"81",
          4752 => x"81",
          4753 => x"38",
          4754 => x"08",
          4755 => x"95",
          4756 => x"84",
          4757 => x"81",
          4758 => x"7b",
          4759 => x"06",
          4760 => x"39",
          4761 => x"56",
          4762 => x"09",
          4763 => x"b9",
          4764 => x"80",
          4765 => x"80",
          4766 => x"78",
          4767 => x"7a",
          4768 => x"38",
          4769 => x"73",
          4770 => x"81",
          4771 => x"ff",
          4772 => x"74",
          4773 => x"ff",
          4774 => x"81",
          4775 => x"58",
          4776 => x"08",
          4777 => x"74",
          4778 => x"16",
          4779 => x"73",
          4780 => x"39",
          4781 => x"7e",
          4782 => x"0c",
          4783 => x"2e",
          4784 => x"88",
          4785 => x"8c",
          4786 => x"1a",
          4787 => x"07",
          4788 => x"1b",
          4789 => x"08",
          4790 => x"16",
          4791 => x"75",
          4792 => x"38",
          4793 => x"90",
          4794 => x"15",
          4795 => x"54",
          4796 => x"34",
          4797 => x"81",
          4798 => x"90",
          4799 => x"e9",
          4800 => x"6d",
          4801 => x"80",
          4802 => x"9d",
          4803 => x"5c",
          4804 => x"3f",
          4805 => x"0b",
          4806 => x"08",
          4807 => x"38",
          4808 => x"08",
          4809 => x"d3",
          4810 => x"08",
          4811 => x"80",
          4812 => x"80",
          4813 => x"d3",
          4814 => x"ff",
          4815 => x"52",
          4816 => x"a0",
          4817 => x"d3",
          4818 => x"ff",
          4819 => x"06",
          4820 => x"56",
          4821 => x"38",
          4822 => x"70",
          4823 => x"55",
          4824 => x"8b",
          4825 => x"3d",
          4826 => x"83",
          4827 => x"ff",
          4828 => x"81",
          4829 => x"99",
          4830 => x"74",
          4831 => x"38",
          4832 => x"80",
          4833 => x"ff",
          4834 => x"55",
          4835 => x"83",
          4836 => x"78",
          4837 => x"38",
          4838 => x"26",
          4839 => x"81",
          4840 => x"8b",
          4841 => x"79",
          4842 => x"80",
          4843 => x"93",
          4844 => x"39",
          4845 => x"6e",
          4846 => x"89",
          4847 => x"48",
          4848 => x"83",
          4849 => x"61",
          4850 => x"25",
          4851 => x"55",
          4852 => x"8a",
          4853 => x"3d",
          4854 => x"81",
          4855 => x"ff",
          4856 => x"81",
          4857 => x"84",
          4858 => x"38",
          4859 => x"70",
          4860 => x"d3",
          4861 => x"56",
          4862 => x"38",
          4863 => x"55",
          4864 => x"75",
          4865 => x"38",
          4866 => x"70",
          4867 => x"ff",
          4868 => x"83",
          4869 => x"78",
          4870 => x"89",
          4871 => x"81",
          4872 => x"06",
          4873 => x"80",
          4874 => x"77",
          4875 => x"74",
          4876 => x"8d",
          4877 => x"06",
          4878 => x"2e",
          4879 => x"77",
          4880 => x"93",
          4881 => x"74",
          4882 => x"cb",
          4883 => x"7d",
          4884 => x"81",
          4885 => x"38",
          4886 => x"66",
          4887 => x"81",
          4888 => x"9c",
          4889 => x"74",
          4890 => x"38",
          4891 => x"98",
          4892 => x"9c",
          4893 => x"82",
          4894 => x"57",
          4895 => x"80",
          4896 => x"76",
          4897 => x"38",
          4898 => x"51",
          4899 => x"3f",
          4900 => x"08",
          4901 => x"87",
          4902 => x"2a",
          4903 => x"5c",
          4904 => x"d3",
          4905 => x"80",
          4906 => x"44",
          4907 => x"0a",
          4908 => x"ec",
          4909 => x"39",
          4910 => x"66",
          4911 => x"81",
          4912 => x"8c",
          4913 => x"74",
          4914 => x"38",
          4915 => x"98",
          4916 => x"8c",
          4917 => x"82",
          4918 => x"57",
          4919 => x"80",
          4920 => x"76",
          4921 => x"38",
          4922 => x"51",
          4923 => x"3f",
          4924 => x"08",
          4925 => x"57",
          4926 => x"08",
          4927 => x"96",
          4928 => x"81",
          4929 => x"10",
          4930 => x"08",
          4931 => x"72",
          4932 => x"59",
          4933 => x"ff",
          4934 => x"5d",
          4935 => x"44",
          4936 => x"11",
          4937 => x"70",
          4938 => x"71",
          4939 => x"06",
          4940 => x"52",
          4941 => x"40",
          4942 => x"09",
          4943 => x"38",
          4944 => x"18",
          4945 => x"39",
          4946 => x"79",
          4947 => x"70",
          4948 => x"58",
          4949 => x"76",
          4950 => x"38",
          4951 => x"7d",
          4952 => x"70",
          4953 => x"55",
          4954 => x"3f",
          4955 => x"08",
          4956 => x"2e",
          4957 => x"9b",
          4958 => x"84",
          4959 => x"f5",
          4960 => x"38",
          4961 => x"38",
          4962 => x"59",
          4963 => x"38",
          4964 => x"7d",
          4965 => x"81",
          4966 => x"38",
          4967 => x"0b",
          4968 => x"08",
          4969 => x"78",
          4970 => x"1a",
          4971 => x"c0",
          4972 => x"74",
          4973 => x"39",
          4974 => x"55",
          4975 => x"8f",
          4976 => x"fd",
          4977 => x"d3",
          4978 => x"f5",
          4979 => x"78",
          4980 => x"79",
          4981 => x"80",
          4982 => x"f1",
          4983 => x"39",
          4984 => x"81",
          4985 => x"06",
          4986 => x"55",
          4987 => x"27",
          4988 => x"81",
          4989 => x"56",
          4990 => x"38",
          4991 => x"80",
          4992 => x"ff",
          4993 => x"8b",
          4994 => x"b4",
          4995 => x"ff",
          4996 => x"84",
          4997 => x"1b",
          4998 => x"b3",
          4999 => x"1c",
          5000 => x"ff",
          5001 => x"8e",
          5002 => x"a1",
          5003 => x"0b",
          5004 => x"7d",
          5005 => x"30",
          5006 => x"84",
          5007 => x"51",
          5008 => x"51",
          5009 => x"3f",
          5010 => x"83",
          5011 => x"90",
          5012 => x"ff",
          5013 => x"93",
          5014 => x"a0",
          5015 => x"39",
          5016 => x"1b",
          5017 => x"85",
          5018 => x"95",
          5019 => x"52",
          5020 => x"ff",
          5021 => x"81",
          5022 => x"1b",
          5023 => x"cf",
          5024 => x"9c",
          5025 => x"a0",
          5026 => x"83",
          5027 => x"06",
          5028 => x"82",
          5029 => x"52",
          5030 => x"51",
          5031 => x"3f",
          5032 => x"1b",
          5033 => x"c5",
          5034 => x"ac",
          5035 => x"a0",
          5036 => x"52",
          5037 => x"ff",
          5038 => x"86",
          5039 => x"51",
          5040 => x"3f",
          5041 => x"80",
          5042 => x"a9",
          5043 => x"1c",
          5044 => x"81",
          5045 => x"80",
          5046 => x"ae",
          5047 => x"b2",
          5048 => x"1b",
          5049 => x"85",
          5050 => x"ff",
          5051 => x"96",
          5052 => x"9f",
          5053 => x"80",
          5054 => x"34",
          5055 => x"1c",
          5056 => x"81",
          5057 => x"ab",
          5058 => x"a0",
          5059 => x"d4",
          5060 => x"fe",
          5061 => x"59",
          5062 => x"3f",
          5063 => x"53",
          5064 => x"51",
          5065 => x"3f",
          5066 => x"d3",
          5067 => x"e7",
          5068 => x"2e",
          5069 => x"80",
          5070 => x"54",
          5071 => x"53",
          5072 => x"51",
          5073 => x"3f",
          5074 => x"80",
          5075 => x"ff",
          5076 => x"84",
          5077 => x"d2",
          5078 => x"ff",
          5079 => x"86",
          5080 => x"f2",
          5081 => x"1b",
          5082 => x"81",
          5083 => x"52",
          5084 => x"51",
          5085 => x"3f",
          5086 => x"ec",
          5087 => x"9e",
          5088 => x"d4",
          5089 => x"51",
          5090 => x"3f",
          5091 => x"87",
          5092 => x"52",
          5093 => x"9a",
          5094 => x"54",
          5095 => x"7a",
          5096 => x"ff",
          5097 => x"65",
          5098 => x"7a",
          5099 => x"8f",
          5100 => x"80",
          5101 => x"2e",
          5102 => x"9a",
          5103 => x"7a",
          5104 => x"a9",
          5105 => x"84",
          5106 => x"9e",
          5107 => x"0a",
          5108 => x"51",
          5109 => x"ff",
          5110 => x"7d",
          5111 => x"38",
          5112 => x"52",
          5113 => x"9e",
          5114 => x"55",
          5115 => x"62",
          5116 => x"74",
          5117 => x"75",
          5118 => x"7e",
          5119 => x"fe",
          5120 => x"84",
          5121 => x"38",
          5122 => x"81",
          5123 => x"52",
          5124 => x"9e",
          5125 => x"16",
          5126 => x"56",
          5127 => x"38",
          5128 => x"77",
          5129 => x"8d",
          5130 => x"7d",
          5131 => x"38",
          5132 => x"57",
          5133 => x"83",
          5134 => x"76",
          5135 => x"7a",
          5136 => x"ff",
          5137 => x"81",
          5138 => x"81",
          5139 => x"16",
          5140 => x"56",
          5141 => x"38",
          5142 => x"83",
          5143 => x"86",
          5144 => x"ff",
          5145 => x"38",
          5146 => x"82",
          5147 => x"81",
          5148 => x"06",
          5149 => x"fe",
          5150 => x"53",
          5151 => x"51",
          5152 => x"3f",
          5153 => x"52",
          5154 => x"9c",
          5155 => x"be",
          5156 => x"75",
          5157 => x"81",
          5158 => x"0b",
          5159 => x"77",
          5160 => x"75",
          5161 => x"60",
          5162 => x"80",
          5163 => x"75",
          5164 => x"c4",
          5165 => x"85",
          5166 => x"d3",
          5167 => x"2a",
          5168 => x"75",
          5169 => x"81",
          5170 => x"87",
          5171 => x"52",
          5172 => x"51",
          5173 => x"3f",
          5174 => x"ca",
          5175 => x"9c",
          5176 => x"54",
          5177 => x"52",
          5178 => x"98",
          5179 => x"56",
          5180 => x"08",
          5181 => x"53",
          5182 => x"51",
          5183 => x"3f",
          5184 => x"d3",
          5185 => x"38",
          5186 => x"56",
          5187 => x"56",
          5188 => x"d3",
          5189 => x"75",
          5190 => x"0c",
          5191 => x"04",
          5192 => x"73",
          5193 => x"26",
          5194 => x"71",
          5195 => x"bd",
          5196 => x"71",
          5197 => x"c5",
          5198 => x"80",
          5199 => x"b8",
          5200 => x"39",
          5201 => x"51",
          5202 => x"81",
          5203 => x"80",
          5204 => x"c5",
          5205 => x"e4",
          5206 => x"80",
          5207 => x"39",
          5208 => x"51",
          5209 => x"81",
          5210 => x"80",
          5211 => x"c6",
          5212 => x"c8",
          5213 => x"d4",
          5214 => x"39",
          5215 => x"51",
          5216 => x"c7",
          5217 => x"39",
          5218 => x"51",
          5219 => x"c7",
          5220 => x"39",
          5221 => x"51",
          5222 => x"c7",
          5223 => x"39",
          5224 => x"51",
          5225 => x"c8",
          5226 => x"39",
          5227 => x"51",
          5228 => x"c8",
          5229 => x"39",
          5230 => x"51",
          5231 => x"3f",
          5232 => x"04",
          5233 => x"77",
          5234 => x"74",
          5235 => x"8a",
          5236 => x"75",
          5237 => x"51",
          5238 => x"e8",
          5239 => x"fe",
          5240 => x"81",
          5241 => x"52",
          5242 => x"ef",
          5243 => x"d3",
          5244 => x"79",
          5245 => x"81",
          5246 => x"ff",
          5247 => x"87",
          5248 => x"f5",
          5249 => x"7f",
          5250 => x"05",
          5251 => x"33",
          5252 => x"66",
          5253 => x"5a",
          5254 => x"78",
          5255 => x"98",
          5256 => x"fa",
          5257 => x"a0",
          5258 => x"8e",
          5259 => x"74",
          5260 => x"fc",
          5261 => x"2e",
          5262 => x"a0",
          5263 => x"80",
          5264 => x"16",
          5265 => x"27",
          5266 => x"22",
          5267 => x"a4",
          5268 => x"ca",
          5269 => x"81",
          5270 => x"ff",
          5271 => x"82",
          5272 => x"c3",
          5273 => x"53",
          5274 => x"8e",
          5275 => x"52",
          5276 => x"51",
          5277 => x"3f",
          5278 => x"c9",
          5279 => x"86",
          5280 => x"15",
          5281 => x"74",
          5282 => x"78",
          5283 => x"72",
          5284 => x"c9",
          5285 => x"8c",
          5286 => x"39",
          5287 => x"51",
          5288 => x"3f",
          5289 => x"a0",
          5290 => x"8f",
          5291 => x"39",
          5292 => x"51",
          5293 => x"3f",
          5294 => x"77",
          5295 => x"74",
          5296 => x"79",
          5297 => x"55",
          5298 => x"27",
          5299 => x"80",
          5300 => x"73",
          5301 => x"85",
          5302 => x"83",
          5303 => x"fe",
          5304 => x"81",
          5305 => x"39",
          5306 => x"51",
          5307 => x"3f",
          5308 => x"1a",
          5309 => x"fd",
          5310 => x"d3",
          5311 => x"2b",
          5312 => x"51",
          5313 => x"2e",
          5314 => x"a5",
          5315 => x"fd",
          5316 => x"84",
          5317 => x"70",
          5318 => x"a0",
          5319 => x"70",
          5320 => x"2a",
          5321 => x"51",
          5322 => x"2e",
          5323 => x"dd",
          5324 => x"2e",
          5325 => x"85",
          5326 => x"8c",
          5327 => x"53",
          5328 => x"fd",
          5329 => x"53",
          5330 => x"84",
          5331 => x"0d",
          5332 => x"0d",
          5333 => x"05",
          5334 => x"33",
          5335 => x"70",
          5336 => x"25",
          5337 => x"74",
          5338 => x"51",
          5339 => x"56",
          5340 => x"80",
          5341 => x"53",
          5342 => x"3d",
          5343 => x"c0",
          5344 => x"d3",
          5345 => x"81",
          5346 => x"b8",
          5347 => x"84",
          5348 => x"98",
          5349 => x"d3",
          5350 => x"96",
          5351 => x"54",
          5352 => x"77",
          5353 => x"c4",
          5354 => x"d3",
          5355 => x"81",
          5356 => x"90",
          5357 => x"74",
          5358 => x"38",
          5359 => x"19",
          5360 => x"39",
          5361 => x"05",
          5362 => x"3f",
          5363 => x"77",
          5364 => x"51",
          5365 => x"2e",
          5366 => x"80",
          5367 => x"81",
          5368 => x"87",
          5369 => x"08",
          5370 => x"fb",
          5371 => x"57",
          5372 => x"84",
          5373 => x"0d",
          5374 => x"0d",
          5375 => x"05",
          5376 => x"57",
          5377 => x"80",
          5378 => x"79",
          5379 => x"3f",
          5380 => x"08",
          5381 => x"80",
          5382 => x"75",
          5383 => x"38",
          5384 => x"55",
          5385 => x"d3",
          5386 => x"52",
          5387 => x"2d",
          5388 => x"08",
          5389 => x"77",
          5390 => x"d3",
          5391 => x"3d",
          5392 => x"3d",
          5393 => x"05",
          5394 => x"d4",
          5395 => x"dc",
          5396 => x"88",
          5397 => x"d0",
          5398 => x"ff",
          5399 => x"81",
          5400 => x"81",
          5401 => x"81",
          5402 => x"52",
          5403 => x"51",
          5404 => x"3f",
          5405 => x"85",
          5406 => x"94",
          5407 => x"0d",
          5408 => x"0d",
          5409 => x"80",
          5410 => x"80",
          5411 => x"51",
          5412 => x"3f",
          5413 => x"51",
          5414 => x"3f",
          5415 => x"f6",
          5416 => x"81",
          5417 => x"06",
          5418 => x"80",
          5419 => x"81",
          5420 => x"ed",
          5421 => x"b4",
          5422 => x"e5",
          5423 => x"fe",
          5424 => x"72",
          5425 => x"81",
          5426 => x"71",
          5427 => x"38",
          5428 => x"f5",
          5429 => x"ca",
          5430 => x"f7",
          5431 => x"51",
          5432 => x"3f",
          5433 => x"70",
          5434 => x"52",
          5435 => x"95",
          5436 => x"fe",
          5437 => x"81",
          5438 => x"fe",
          5439 => x"80",
          5440 => x"9d",
          5441 => x"2a",
          5442 => x"51",
          5443 => x"2e",
          5444 => x"51",
          5445 => x"3f",
          5446 => x"51",
          5447 => x"3f",
          5448 => x"f4",
          5449 => x"85",
          5450 => x"06",
          5451 => x"80",
          5452 => x"81",
          5453 => x"e9",
          5454 => x"80",
          5455 => x"e1",
          5456 => x"fe",
          5457 => x"72",
          5458 => x"81",
          5459 => x"71",
          5460 => x"38",
          5461 => x"f4",
          5462 => x"cb",
          5463 => x"f6",
          5464 => x"51",
          5465 => x"3f",
          5466 => x"70",
          5467 => x"52",
          5468 => x"95",
          5469 => x"fe",
          5470 => x"81",
          5471 => x"fe",
          5472 => x"80",
          5473 => x"99",
          5474 => x"2a",
          5475 => x"51",
          5476 => x"2e",
          5477 => x"51",
          5478 => x"3f",
          5479 => x"51",
          5480 => x"3f",
          5481 => x"f3",
          5482 => x"ff",
          5483 => x"3d",
          5484 => x"3d",
          5485 => x"08",
          5486 => x"57",
          5487 => x"80",
          5488 => x"39",
          5489 => x"85",
          5490 => x"80",
          5491 => x"14",
          5492 => x"33",
          5493 => x"06",
          5494 => x"74",
          5495 => x"38",
          5496 => x"80",
          5497 => x"72",
          5498 => x"81",
          5499 => x"72",
          5500 => x"81",
          5501 => x"80",
          5502 => x"05",
          5503 => x"56",
          5504 => x"81",
          5505 => x"77",
          5506 => x"08",
          5507 => x"ed",
          5508 => x"d3",
          5509 => x"38",
          5510 => x"53",
          5511 => x"ff",
          5512 => x"16",
          5513 => x"06",
          5514 => x"76",
          5515 => x"ff",
          5516 => x"d3",
          5517 => x"3d",
          5518 => x"3d",
          5519 => x"71",
          5520 => x"0c",
          5521 => x"52",
          5522 => x"8a",
          5523 => x"d3",
          5524 => x"ff",
          5525 => x"7c",
          5526 => x"06",
          5527 => x"cb",
          5528 => x"3d",
          5529 => x"ff",
          5530 => x"7b",
          5531 => x"81",
          5532 => x"ff",
          5533 => x"81",
          5534 => x"7c",
          5535 => x"81",
          5536 => x"8e",
          5537 => x"70",
          5538 => x"cc",
          5539 => x"fe",
          5540 => x"3d",
          5541 => x"80",
          5542 => x"52",
          5543 => x"eb",
          5544 => x"f8",
          5545 => x"ff",
          5546 => x"b7",
          5547 => x"05",
          5548 => x"3f",
          5549 => x"08",
          5550 => x"90",
          5551 => x"78",
          5552 => x"8a",
          5553 => x"80",
          5554 => x"dc",
          5555 => x"2e",
          5556 => x"78",
          5557 => x"38",
          5558 => x"81",
          5559 => x"82",
          5560 => x"78",
          5561 => x"a2",
          5562 => x"39",
          5563 => x"82",
          5564 => x"94",
          5565 => x"38",
          5566 => x"78",
          5567 => x"85",
          5568 => x"80",
          5569 => x"38",
          5570 => x"83",
          5571 => x"bc",
          5572 => x"38",
          5573 => x"78",
          5574 => x"86",
          5575 => x"80",
          5576 => x"8c",
          5577 => x"39",
          5578 => x"2e",
          5579 => x"78",
          5580 => x"a9",
          5581 => x"d1",
          5582 => x"38",
          5583 => x"24",
          5584 => x"80",
          5585 => x"c4",
          5586 => x"39",
          5587 => x"2e",
          5588 => x"78",
          5589 => x"8a",
          5590 => x"97",
          5591 => x"83",
          5592 => x"38",
          5593 => x"24",
          5594 => x"80",
          5595 => x"9d",
          5596 => x"82",
          5597 => x"38",
          5598 => x"78",
          5599 => x"8b",
          5600 => x"81",
          5601 => x"82",
          5602 => x"39",
          5603 => x"f4",
          5604 => x"f8",
          5605 => x"83",
          5606 => x"d3",
          5607 => x"38",
          5608 => x"51",
          5609 => x"b7",
          5610 => x"11",
          5611 => x"05",
          5612 => x"df",
          5613 => x"84",
          5614 => x"88",
          5615 => x"25",
          5616 => x"43",
          5617 => x"05",
          5618 => x"80",
          5619 => x"51",
          5620 => x"3f",
          5621 => x"08",
          5622 => x"59",
          5623 => x"81",
          5624 => x"fe",
          5625 => x"81",
          5626 => x"39",
          5627 => x"51",
          5628 => x"b7",
          5629 => x"11",
          5630 => x"05",
          5631 => x"93",
          5632 => x"84",
          5633 => x"fd",
          5634 => x"53",
          5635 => x"80",
          5636 => x"51",
          5637 => x"3f",
          5638 => x"08",
          5639 => x"f4",
          5640 => x"39",
          5641 => x"f4",
          5642 => x"f8",
          5643 => x"82",
          5644 => x"d3",
          5645 => x"2e",
          5646 => x"89",
          5647 => x"38",
          5648 => x"f0",
          5649 => x"f8",
          5650 => x"82",
          5651 => x"d3",
          5652 => x"38",
          5653 => x"08",
          5654 => x"81",
          5655 => x"79",
          5656 => x"d0",
          5657 => x"cb",
          5658 => x"79",
          5659 => x"b4",
          5660 => x"b4",
          5661 => x"b5",
          5662 => x"d3",
          5663 => x"93",
          5664 => x"cc",
          5665 => x"b2",
          5666 => x"fb",
          5667 => x"3d",
          5668 => x"51",
          5669 => x"3f",
          5670 => x"08",
          5671 => x"f8",
          5672 => x"fe",
          5673 => x"81",
          5674 => x"84",
          5675 => x"51",
          5676 => x"80",
          5677 => x"3d",
          5678 => x"51",
          5679 => x"3f",
          5680 => x"08",
          5681 => x"f8",
          5682 => x"fe",
          5683 => x"81",
          5684 => x"b8",
          5685 => x"05",
          5686 => x"ea",
          5687 => x"d3",
          5688 => x"3d",
          5689 => x"52",
          5690 => x"c8",
          5691 => x"80",
          5692 => x"b8",
          5693 => x"80",
          5694 => x"84",
          5695 => x"06",
          5696 => x"79",
          5697 => x"f5",
          5698 => x"d3",
          5699 => x"2e",
          5700 => x"81",
          5701 => x"51",
          5702 => x"fa",
          5703 => x"3d",
          5704 => x"53",
          5705 => x"51",
          5706 => x"3f",
          5707 => x"08",
          5708 => x"d6",
          5709 => x"fe",
          5710 => x"fe",
          5711 => x"ff",
          5712 => x"81",
          5713 => x"80",
          5714 => x"38",
          5715 => x"ec",
          5716 => x"f8",
          5717 => x"80",
          5718 => x"d3",
          5719 => x"38",
          5720 => x"08",
          5721 => x"80",
          5722 => x"ce",
          5723 => x"5c",
          5724 => x"27",
          5725 => x"59",
          5726 => x"84",
          5727 => x"7a",
          5728 => x"38",
          5729 => x"51",
          5730 => x"b7",
          5731 => x"11",
          5732 => x"05",
          5733 => x"fb",
          5734 => x"84",
          5735 => x"38",
          5736 => x"33",
          5737 => x"2e",
          5738 => x"d0",
          5739 => x"b3",
          5740 => x"ae",
          5741 => x"80",
          5742 => x"81",
          5743 => x"44",
          5744 => x"d0",
          5745 => x"78",
          5746 => x"d0",
          5747 => x"78",
          5748 => x"38",
          5749 => x"08",
          5750 => x"81",
          5751 => x"fc",
          5752 => x"b7",
          5753 => x"11",
          5754 => x"05",
          5755 => x"a3",
          5756 => x"84",
          5757 => x"38",
          5758 => x"33",
          5759 => x"2e",
          5760 => x"d0",
          5761 => x"b2",
          5762 => x"ae",
          5763 => x"80",
          5764 => x"81",
          5765 => x"43",
          5766 => x"d0",
          5767 => x"78",
          5768 => x"d0",
          5769 => x"78",
          5770 => x"38",
          5771 => x"08",
          5772 => x"81",
          5773 => x"88",
          5774 => x"3d",
          5775 => x"53",
          5776 => x"51",
          5777 => x"3f",
          5778 => x"08",
          5779 => x"38",
          5780 => x"59",
          5781 => x"83",
          5782 => x"79",
          5783 => x"38",
          5784 => x"88",
          5785 => x"2e",
          5786 => x"42",
          5787 => x"51",
          5788 => x"3f",
          5789 => x"54",
          5790 => x"52",
          5791 => x"83",
          5792 => x"9c",
          5793 => x"39",
          5794 => x"f4",
          5795 => x"f8",
          5796 => x"fd",
          5797 => x"d3",
          5798 => x"2e",
          5799 => x"b7",
          5800 => x"11",
          5801 => x"05",
          5802 => x"e7",
          5803 => x"84",
          5804 => x"a5",
          5805 => x"02",
          5806 => x"33",
          5807 => x"81",
          5808 => x"3d",
          5809 => x"53",
          5810 => x"51",
          5811 => x"3f",
          5812 => x"08",
          5813 => x"b2",
          5814 => x"33",
          5815 => x"cd",
          5816 => x"fb",
          5817 => x"f8",
          5818 => x"fe",
          5819 => x"79",
          5820 => x"59",
          5821 => x"f7",
          5822 => x"79",
          5823 => x"b7",
          5824 => x"11",
          5825 => x"05",
          5826 => x"87",
          5827 => x"84",
          5828 => x"91",
          5829 => x"02",
          5830 => x"33",
          5831 => x"81",
          5832 => x"b5",
          5833 => x"b4",
          5834 => x"8e",
          5835 => x"39",
          5836 => x"e8",
          5837 => x"f8",
          5838 => x"fe",
          5839 => x"d3",
          5840 => x"2e",
          5841 => x"b7",
          5842 => x"11",
          5843 => x"05",
          5844 => x"b1",
          5845 => x"84",
          5846 => x"a6",
          5847 => x"02",
          5848 => x"79",
          5849 => x"5b",
          5850 => x"b7",
          5851 => x"11",
          5852 => x"05",
          5853 => x"8d",
          5854 => x"84",
          5855 => x"f6",
          5856 => x"70",
          5857 => x"81",
          5858 => x"fe",
          5859 => x"80",
          5860 => x"51",
          5861 => x"3f",
          5862 => x"33",
          5863 => x"2e",
          5864 => x"78",
          5865 => x"38",
          5866 => x"41",
          5867 => x"3d",
          5868 => x"53",
          5869 => x"51",
          5870 => x"3f",
          5871 => x"08",
          5872 => x"38",
          5873 => x"be",
          5874 => x"70",
          5875 => x"23",
          5876 => x"ae",
          5877 => x"b4",
          5878 => x"de",
          5879 => x"39",
          5880 => x"e8",
          5881 => x"f8",
          5882 => x"fd",
          5883 => x"d3",
          5884 => x"2e",
          5885 => x"b7",
          5886 => x"11",
          5887 => x"05",
          5888 => x"81",
          5889 => x"84",
          5890 => x"a1",
          5891 => x"71",
          5892 => x"84",
          5893 => x"3d",
          5894 => x"53",
          5895 => x"51",
          5896 => x"3f",
          5897 => x"08",
          5898 => x"de",
          5899 => x"08",
          5900 => x"cd",
          5901 => x"f8",
          5902 => x"f8",
          5903 => x"fe",
          5904 => x"79",
          5905 => x"59",
          5906 => x"f4",
          5907 => x"79",
          5908 => x"b7",
          5909 => x"11",
          5910 => x"05",
          5911 => x"a5",
          5912 => x"84",
          5913 => x"99",
          5914 => x"60",
          5915 => x"c8",
          5916 => x"aa",
          5917 => x"71",
          5918 => x"84",
          5919 => x"ad",
          5920 => x"b4",
          5921 => x"b2",
          5922 => x"39",
          5923 => x"51",
          5924 => x"3f",
          5925 => x"f1",
          5926 => x"ee",
          5927 => x"ec",
          5928 => x"96",
          5929 => x"fe",
          5930 => x"f3",
          5931 => x"80",
          5932 => x"c0",
          5933 => x"84",
          5934 => x"87",
          5935 => x"0c",
          5936 => x"51",
          5937 => x"3f",
          5938 => x"81",
          5939 => x"fe",
          5940 => x"8c",
          5941 => x"87",
          5942 => x"0c",
          5943 => x"0b",
          5944 => x"94",
          5945 => x"39",
          5946 => x"f4",
          5947 => x"f8",
          5948 => x"f9",
          5949 => x"d3",
          5950 => x"2e",
          5951 => x"63",
          5952 => x"ac",
          5953 => x"96",
          5954 => x"78",
          5955 => x"fe",
          5956 => x"fe",
          5957 => x"fe",
          5958 => x"81",
          5959 => x"80",
          5960 => x"38",
          5961 => x"ce",
          5962 => x"f6",
          5963 => x"59",
          5964 => x"d3",
          5965 => x"81",
          5966 => x"80",
          5967 => x"38",
          5968 => x"08",
          5969 => x"e4",
          5970 => x"d2",
          5971 => x"39",
          5972 => x"51",
          5973 => x"3f",
          5974 => x"3f",
          5975 => x"81",
          5976 => x"fe",
          5977 => x"80",
          5978 => x"39",
          5979 => x"3f",
          5980 => x"64",
          5981 => x"59",
          5982 => x"f2",
          5983 => x"80",
          5984 => x"38",
          5985 => x"80",
          5986 => x"3d",
          5987 => x"51",
          5988 => x"3f",
          5989 => x"56",
          5990 => x"08",
          5991 => x"b4",
          5992 => x"81",
          5993 => x"a3",
          5994 => x"5a",
          5995 => x"3f",
          5996 => x"58",
          5997 => x"57",
          5998 => x"81",
          5999 => x"05",
          6000 => x"82",
          6001 => x"82",
          6002 => x"79",
          6003 => x"3f",
          6004 => x"08",
          6005 => x"32",
          6006 => x"07",
          6007 => x"38",
          6008 => x"09",
          6009 => x"a2",
          6010 => x"c8",
          6011 => x"ae",
          6012 => x"39",
          6013 => x"80",
          6014 => x"b8",
          6015 => x"86",
          6016 => x"c0",
          6017 => x"9b",
          6018 => x"0b",
          6019 => x"9c",
          6020 => x"83",
          6021 => x"94",
          6022 => x"80",
          6023 => x"c0",
          6024 => x"9f",
          6025 => x"d3",
          6026 => x"bb",
          6027 => x"98",
          6028 => x"b1",
          6029 => x"d2",
          6030 => x"d8",
          6031 => x"e1",
          6032 => x"e4",
          6033 => x"f2",
          6034 => x"80",
          6035 => x"b5",
          6036 => x"eb",
          6037 => x"e2",
          6038 => x"00",
          6039 => x"ff",
          6040 => x"ff",
          6041 => x"00",
          6042 => x"ff",
          6043 => x"14",
          6044 => x"14",
          6045 => x"14",
          6046 => x"14",
          6047 => x"14",
          6048 => x"51",
          6049 => x"51",
          6050 => x"51",
          6051 => x"51",
          6052 => x"51",
          6053 => x"51",
          6054 => x"51",
          6055 => x"51",
          6056 => x"51",
          6057 => x"51",
          6058 => x"51",
          6059 => x"51",
          6060 => x"51",
          6061 => x"51",
          6062 => x"51",
          6063 => x"51",
          6064 => x"51",
          6065 => x"51",
          6066 => x"51",
          6067 => x"51",
          6068 => x"2f",
          6069 => x"25",
          6070 => x"64",
          6071 => x"3a",
          6072 => x"25",
          6073 => x"0a",
          6074 => x"43",
          6075 => x"6e",
          6076 => x"75",
          6077 => x"69",
          6078 => x"00",
          6079 => x"66",
          6080 => x"20",
          6081 => x"20",
          6082 => x"66",
          6083 => x"00",
          6084 => x"44",
          6085 => x"63",
          6086 => x"69",
          6087 => x"65",
          6088 => x"74",
          6089 => x"0a",
          6090 => x"20",
          6091 => x"53",
          6092 => x"52",
          6093 => x"28",
          6094 => x"72",
          6095 => x"30",
          6096 => x"20",
          6097 => x"65",
          6098 => x"38",
          6099 => x"0a",
          6100 => x"20",
          6101 => x"41",
          6102 => x"53",
          6103 => x"74",
          6104 => x"38",
          6105 => x"53",
          6106 => x"3d",
          6107 => x"58",
          6108 => x"00",
          6109 => x"20",
          6110 => x"4d",
          6111 => x"74",
          6112 => x"3d",
          6113 => x"58",
          6114 => x"69",
          6115 => x"25",
          6116 => x"29",
          6117 => x"00",
          6118 => x"20",
          6119 => x"43",
          6120 => x"00",
          6121 => x"20",
          6122 => x"32",
          6123 => x"00",
          6124 => x"20",
          6125 => x"49",
          6126 => x"00",
          6127 => x"20",
          6128 => x"20",
          6129 => x"64",
          6130 => x"65",
          6131 => x"65",
          6132 => x"30",
          6133 => x"2e",
          6134 => x"00",
          6135 => x"20",
          6136 => x"54",
          6137 => x"55",
          6138 => x"43",
          6139 => x"52",
          6140 => x"45",
          6141 => x"00",
          6142 => x"20",
          6143 => x"4d",
          6144 => x"20",
          6145 => x"6d",
          6146 => x"3d",
          6147 => x"58",
          6148 => x"00",
          6149 => x"64",
          6150 => x"73",
          6151 => x"0a",
          6152 => x"20",
          6153 => x"55",
          6154 => x"73",
          6155 => x"56",
          6156 => x"6f",
          6157 => x"64",
          6158 => x"73",
          6159 => x"20",
          6160 => x"58",
          6161 => x"00",
          6162 => x"20",
          6163 => x"55",
          6164 => x"6d",
          6165 => x"20",
          6166 => x"72",
          6167 => x"64",
          6168 => x"73",
          6169 => x"20",
          6170 => x"58",
          6171 => x"00",
          6172 => x"20",
          6173 => x"61",
          6174 => x"53",
          6175 => x"74",
          6176 => x"64",
          6177 => x"73",
          6178 => x"20",
          6179 => x"20",
          6180 => x"58",
          6181 => x"00",
          6182 => x"20",
          6183 => x"55",
          6184 => x"20",
          6185 => x"20",
          6186 => x"20",
          6187 => x"20",
          6188 => x"20",
          6189 => x"20",
          6190 => x"58",
          6191 => x"00",
          6192 => x"20",
          6193 => x"73",
          6194 => x"20",
          6195 => x"63",
          6196 => x"72",
          6197 => x"20",
          6198 => x"20",
          6199 => x"20",
          6200 => x"58",
          6201 => x"00",
          6202 => x"61",
          6203 => x"00",
          6204 => x"64",
          6205 => x"00",
          6206 => x"65",
          6207 => x"00",
          6208 => x"4f",
          6209 => x"4f",
          6210 => x"00",
          6211 => x"6b",
          6212 => x"6e",
          6213 => x"00",
          6214 => x"2b",
          6215 => x"3c",
          6216 => x"5b",
          6217 => x"00",
          6218 => x"54",
          6219 => x"54",
          6220 => x"00",
          6221 => x"90",
          6222 => x"4f",
          6223 => x"30",
          6224 => x"20",
          6225 => x"45",
          6226 => x"20",
          6227 => x"33",
          6228 => x"20",
          6229 => x"20",
          6230 => x"45",
          6231 => x"20",
          6232 => x"20",
          6233 => x"20",
          6234 => x"61",
          6235 => x"00",
          6236 => x"00",
          6237 => x"00",
          6238 => x"45",
          6239 => x"8f",
          6240 => x"45",
          6241 => x"8e",
          6242 => x"92",
          6243 => x"55",
          6244 => x"9a",
          6245 => x"9e",
          6246 => x"4f",
          6247 => x"a6",
          6248 => x"aa",
          6249 => x"ae",
          6250 => x"b2",
          6251 => x"b6",
          6252 => x"ba",
          6253 => x"be",
          6254 => x"c2",
          6255 => x"c6",
          6256 => x"ca",
          6257 => x"ce",
          6258 => x"d2",
          6259 => x"d6",
          6260 => x"da",
          6261 => x"de",
          6262 => x"e2",
          6263 => x"e6",
          6264 => x"ea",
          6265 => x"ee",
          6266 => x"f2",
          6267 => x"f6",
          6268 => x"fa",
          6269 => x"fe",
          6270 => x"2c",
          6271 => x"5d",
          6272 => x"2a",
          6273 => x"3f",
          6274 => x"00",
          6275 => x"00",
          6276 => x"00",
          6277 => x"02",
          6278 => x"00",
          6279 => x"00",
          6280 => x"00",
          6281 => x"00",
          6282 => x"00",
          6283 => x"6e",
          6284 => x"00",
          6285 => x"6f",
          6286 => x"00",
          6287 => x"6e",
          6288 => x"00",
          6289 => x"6f",
          6290 => x"00",
          6291 => x"78",
          6292 => x"00",
          6293 => x"6c",
          6294 => x"00",
          6295 => x"75",
          6296 => x"00",
          6297 => x"62",
          6298 => x"68",
          6299 => x"77",
          6300 => x"64",
          6301 => x"65",
          6302 => x"64",
          6303 => x"65",
          6304 => x"6c",
          6305 => x"00",
          6306 => x"70",
          6307 => x"73",
          6308 => x"74",
          6309 => x"73",
          6310 => x"00",
          6311 => x"66",
          6312 => x"00",
          6313 => x"73",
          6314 => x"00",
          6315 => x"73",
          6316 => x"72",
          6317 => x"0a",
          6318 => x"74",
          6319 => x"61",
          6320 => x"72",
          6321 => x"2e",
          6322 => x"00",
          6323 => x"73",
          6324 => x"6f",
          6325 => x"65",
          6326 => x"2e",
          6327 => x"00",
          6328 => x"20",
          6329 => x"65",
          6330 => x"75",
          6331 => x"0a",
          6332 => x"20",
          6333 => x"68",
          6334 => x"75",
          6335 => x"0a",
          6336 => x"76",
          6337 => x"64",
          6338 => x"6c",
          6339 => x"6d",
          6340 => x"00",
          6341 => x"63",
          6342 => x"20",
          6343 => x"69",
          6344 => x"0a",
          6345 => x"6c",
          6346 => x"6c",
          6347 => x"64",
          6348 => x"78",
          6349 => x"73",
          6350 => x"00",
          6351 => x"6c",
          6352 => x"61",
          6353 => x"65",
          6354 => x"76",
          6355 => x"64",
          6356 => x"00",
          6357 => x"20",
          6358 => x"77",
          6359 => x"65",
          6360 => x"6f",
          6361 => x"74",
          6362 => x"0a",
          6363 => x"69",
          6364 => x"6e",
          6365 => x"65",
          6366 => x"73",
          6367 => x"76",
          6368 => x"64",
          6369 => x"00",
          6370 => x"73",
          6371 => x"6f",
          6372 => x"6e",
          6373 => x"65",
          6374 => x"00",
          6375 => x"20",
          6376 => x"70",
          6377 => x"62",
          6378 => x"66",
          6379 => x"73",
          6380 => x"65",
          6381 => x"6f",
          6382 => x"20",
          6383 => x"64",
          6384 => x"2e",
          6385 => x"00",
          6386 => x"72",
          6387 => x"20",
          6388 => x"72",
          6389 => x"2e",
          6390 => x"00",
          6391 => x"6d",
          6392 => x"74",
          6393 => x"70",
          6394 => x"74",
          6395 => x"20",
          6396 => x"63",
          6397 => x"65",
          6398 => x"00",
          6399 => x"6c",
          6400 => x"73",
          6401 => x"63",
          6402 => x"2e",
          6403 => x"00",
          6404 => x"73",
          6405 => x"69",
          6406 => x"6e",
          6407 => x"65",
          6408 => x"79",
          6409 => x"00",
          6410 => x"6f",
          6411 => x"6e",
          6412 => x"70",
          6413 => x"66",
          6414 => x"73",
          6415 => x"00",
          6416 => x"72",
          6417 => x"74",
          6418 => x"20",
          6419 => x"6f",
          6420 => x"63",
          6421 => x"00",
          6422 => x"63",
          6423 => x"73",
          6424 => x"00",
          6425 => x"6b",
          6426 => x"6e",
          6427 => x"72",
          6428 => x"0a",
          6429 => x"6c",
          6430 => x"79",
          6431 => x"20",
          6432 => x"61",
          6433 => x"6c",
          6434 => x"79",
          6435 => x"2f",
          6436 => x"2e",
          6437 => x"00",
          6438 => x"38",
          6439 => x"00",
          6440 => x"20",
          6441 => x"34",
          6442 => x"00",
          6443 => x"20",
          6444 => x"20",
          6445 => x"00",
          6446 => x"32",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"0a",
          6451 => x"61",
          6452 => x"00",
          6453 => x"55",
          6454 => x"00",
          6455 => x"2a",
          6456 => x"20",
          6457 => x"00",
          6458 => x"2f",
          6459 => x"32",
          6460 => x"00",
          6461 => x"2e",
          6462 => x"00",
          6463 => x"50",
          6464 => x"72",
          6465 => x"25",
          6466 => x"29",
          6467 => x"20",
          6468 => x"2a",
          6469 => x"00",
          6470 => x"55",
          6471 => x"49",
          6472 => x"72",
          6473 => x"74",
          6474 => x"6e",
          6475 => x"72",
          6476 => x"00",
          6477 => x"6d",
          6478 => x"69",
          6479 => x"72",
          6480 => x"74",
          6481 => x"00",
          6482 => x"32",
          6483 => x"74",
          6484 => x"75",
          6485 => x"00",
          6486 => x"43",
          6487 => x"52",
          6488 => x"6e",
          6489 => x"72",
          6490 => x"0a",
          6491 => x"43",
          6492 => x"57",
          6493 => x"6e",
          6494 => x"72",
          6495 => x"0a",
          6496 => x"52",
          6497 => x"52",
          6498 => x"6e",
          6499 => x"72",
          6500 => x"0a",
          6501 => x"52",
          6502 => x"54",
          6503 => x"6e",
          6504 => x"72",
          6505 => x"0a",
          6506 => x"52",
          6507 => x"52",
          6508 => x"6e",
          6509 => x"72",
          6510 => x"0a",
          6511 => x"52",
          6512 => x"54",
          6513 => x"6e",
          6514 => x"72",
          6515 => x"0a",
          6516 => x"74",
          6517 => x"67",
          6518 => x"20",
          6519 => x"65",
          6520 => x"2e",
          6521 => x"00",
          6522 => x"61",
          6523 => x"6e",
          6524 => x"69",
          6525 => x"2e",
          6526 => x"00",
          6527 => x"00",
          6528 => x"69",
          6529 => x"20",
          6530 => x"69",
          6531 => x"69",
          6532 => x"73",
          6533 => x"64",
          6534 => x"72",
          6535 => x"2c",
          6536 => x"65",
          6537 => x"20",
          6538 => x"74",
          6539 => x"6e",
          6540 => x"6c",
          6541 => x"00",
          6542 => x"00",
          6543 => x"64",
          6544 => x"73",
          6545 => x"64",
          6546 => x"00",
          6547 => x"69",
          6548 => x"6c",
          6549 => x"64",
          6550 => x"00",
          6551 => x"69",
          6552 => x"20",
          6553 => x"69",
          6554 => x"69",
          6555 => x"73",
          6556 => x"00",
          6557 => x"3d",
          6558 => x"00",
          6559 => x"3a",
          6560 => x"65",
          6561 => x"6e",
          6562 => x"2e",
          6563 => x"6d",
          6564 => x"65",
          6565 => x"79",
          6566 => x"00",
          6567 => x"6f",
          6568 => x"65",
          6569 => x"0a",
          6570 => x"38",
          6571 => x"30",
          6572 => x"00",
          6573 => x"3f",
          6574 => x"00",
          6575 => x"38",
          6576 => x"30",
          6577 => x"00",
          6578 => x"38",
          6579 => x"30",
          6580 => x"00",
          6581 => x"73",
          6582 => x"69",
          6583 => x"69",
          6584 => x"72",
          6585 => x"74",
          6586 => x"00",
          6587 => x"61",
          6588 => x"6e",
          6589 => x"6e",
          6590 => x"72",
          6591 => x"73",
          6592 => x"00",
          6593 => x"73",
          6594 => x"65",
          6595 => x"61",
          6596 => x"66",
          6597 => x"0a",
          6598 => x"61",
          6599 => x"6e",
          6600 => x"61",
          6601 => x"66",
          6602 => x"0a",
          6603 => x"65",
          6604 => x"69",
          6605 => x"63",
          6606 => x"20",
          6607 => x"30",
          6608 => x"2e",
          6609 => x"00",
          6610 => x"6c",
          6611 => x"67",
          6612 => x"64",
          6613 => x"20",
          6614 => x"78",
          6615 => x"2e",
          6616 => x"00",
          6617 => x"6c",
          6618 => x"65",
          6619 => x"6e",
          6620 => x"63",
          6621 => x"20",
          6622 => x"29",
          6623 => x"00",
          6624 => x"73",
          6625 => x"74",
          6626 => x"20",
          6627 => x"6c",
          6628 => x"74",
          6629 => x"2e",
          6630 => x"00",
          6631 => x"6c",
          6632 => x"65",
          6633 => x"74",
          6634 => x"2e",
          6635 => x"00",
          6636 => x"55",
          6637 => x"6e",
          6638 => x"3a",
          6639 => x"5c",
          6640 => x"25",
          6641 => x"00",
          6642 => x"64",
          6643 => x"6d",
          6644 => x"64",
          6645 => x"00",
          6646 => x"6e",
          6647 => x"67",
          6648 => x"0a",
          6649 => x"61",
          6650 => x"6e",
          6651 => x"6e",
          6652 => x"72",
          6653 => x"73",
          6654 => x"0a",
          6655 => x"00",
          6656 => x"00",
          6657 => x"7f",
          6658 => x"00",
          6659 => x"7f",
          6660 => x"00",
          6661 => x"7f",
          6662 => x"00",
          6663 => x"00",
          6664 => x"78",
          6665 => x"00",
          6666 => x"e1",
          6667 => x"01",
          6668 => x"01",
          6669 => x"01",
          6670 => x"00",
          6671 => x"00",
          6672 => x"00",
          6673 => x"62",
          6674 => x"01",
          6675 => x"00",
          6676 => x"00",
          6677 => x"62",
          6678 => x"01",
          6679 => x"00",
          6680 => x"00",
          6681 => x"62",
          6682 => x"03",
          6683 => x"00",
          6684 => x"00",
          6685 => x"62",
          6686 => x"03",
          6687 => x"00",
          6688 => x"00",
          6689 => x"62",
          6690 => x"03",
          6691 => x"00",
          6692 => x"00",
          6693 => x"62",
          6694 => x"04",
          6695 => x"00",
          6696 => x"00",
          6697 => x"62",
          6698 => x"04",
          6699 => x"00",
          6700 => x"00",
          6701 => x"62",
          6702 => x"04",
          6703 => x"00",
          6704 => x"00",
          6705 => x"62",
          6706 => x"04",
          6707 => x"00",
          6708 => x"00",
          6709 => x"62",
          6710 => x"04",
          6711 => x"00",
          6712 => x"00",
          6713 => x"62",
          6714 => x"05",
          6715 => x"00",
          6716 => x"00",
          6717 => x"62",
          6718 => x"05",
          6719 => x"00",
          6720 => x"00",
          6721 => x"62",
          6722 => x"05",
          6723 => x"00",
          6724 => x"00",
          6725 => x"62",
          6726 => x"05",
          6727 => x"00",
          6728 => x"00",
          6729 => x"62",
          6730 => x"07",
          6731 => x"00",
          6732 => x"00",
          6733 => x"62",
          6734 => x"07",
          6735 => x"00",
          6736 => x"00",
          6737 => x"62",
          6738 => x"08",
          6739 => x"00",
          6740 => x"00",
          6741 => x"62",
          6742 => x"08",
          6743 => x"00",
          6744 => x"00",
          6745 => x"62",
          6746 => x"08",
          6747 => x"00",
          6748 => x"00",
          6749 => x"62",
          6750 => x"08",
          6751 => x"00",
          6752 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"a4",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8c",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"81",
           386 => x"a0",
           387 => x"d3",
           388 => x"a0",
           389 => x"d3",
           390 => x"dc",
           391 => x"90",
           392 => x"90",
           393 => x"90",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"81",
           399 => x"82",
           400 => x"81",
           401 => x"b1",
           402 => x"d3",
           403 => x"a0",
           404 => x"d3",
           405 => x"f5",
           406 => x"90",
           407 => x"90",
           408 => x"90",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"81",
           414 => x"82",
           415 => x"81",
           416 => x"b5",
           417 => x"d3",
           418 => x"a0",
           419 => x"d3",
           420 => x"9d",
           421 => x"90",
           422 => x"90",
           423 => x"90",
           424 => x"2d",
           425 => x"08",
           426 => x"04",
           427 => x"0c",
           428 => x"81",
           429 => x"82",
           430 => x"81",
           431 => x"a2",
           432 => x"d3",
           433 => x"a0",
           434 => x"d3",
           435 => x"8c",
           436 => x"90",
           437 => x"90",
           438 => x"90",
           439 => x"2d",
           440 => x"08",
           441 => x"04",
           442 => x"0c",
           443 => x"81",
           444 => x"82",
           445 => x"81",
           446 => x"9e",
           447 => x"d3",
           448 => x"a0",
           449 => x"d3",
           450 => x"e7",
           451 => x"d3",
           452 => x"a0",
           453 => x"d3",
           454 => x"f4",
           455 => x"d3",
           456 => x"a0",
           457 => x"d3",
           458 => x"ec",
           459 => x"d3",
           460 => x"a0",
           461 => x"d3",
           462 => x"ef",
           463 => x"d3",
           464 => x"a0",
           465 => x"d3",
           466 => x"f9",
           467 => x"d3",
           468 => x"a0",
           469 => x"d3",
           470 => x"82",
           471 => x"d3",
           472 => x"a0",
           473 => x"d3",
           474 => x"f3",
           475 => x"d3",
           476 => x"a0",
           477 => x"d3",
           478 => x"fc",
           479 => x"d3",
           480 => x"a0",
           481 => x"d3",
           482 => x"fd",
           483 => x"d3",
           484 => x"a0",
           485 => x"d3",
           486 => x"fe",
           487 => x"d3",
           488 => x"a0",
           489 => x"d3",
           490 => x"86",
           491 => x"d3",
           492 => x"a0",
           493 => x"d3",
           494 => x"83",
           495 => x"d3",
           496 => x"a0",
           497 => x"d3",
           498 => x"88",
           499 => x"d3",
           500 => x"a0",
           501 => x"d3",
           502 => x"ff",
           503 => x"d3",
           504 => x"a0",
           505 => x"d3",
           506 => x"8b",
           507 => x"d3",
           508 => x"a0",
           509 => x"d3",
           510 => x"8c",
           511 => x"d3",
           512 => x"a0",
           513 => x"d3",
           514 => x"f5",
           515 => x"d3",
           516 => x"a0",
           517 => x"d3",
           518 => x"f4",
           519 => x"d3",
           520 => x"a0",
           521 => x"d3",
           522 => x"f6",
           523 => x"d3",
           524 => x"a0",
           525 => x"d3",
           526 => x"ff",
           527 => x"d3",
           528 => x"a0",
           529 => x"d3",
           530 => x"8d",
           531 => x"d3",
           532 => x"a0",
           533 => x"d3",
           534 => x"8f",
           535 => x"d3",
           536 => x"a0",
           537 => x"d3",
           538 => x"93",
           539 => x"d3",
           540 => x"a0",
           541 => x"d3",
           542 => x"e6",
           543 => x"d3",
           544 => x"a0",
           545 => x"d3",
           546 => x"95",
           547 => x"d3",
           548 => x"a0",
           549 => x"d3",
           550 => x"93",
           551 => x"90",
           552 => x"90",
           553 => x"90",
           554 => x"2d",
           555 => x"08",
           556 => x"04",
           557 => x"0c",
           558 => x"81",
           559 => x"82",
           560 => x"81",
           561 => x"9b",
           562 => x"d3",
           563 => x"a0",
           564 => x"d3",
           565 => x"b3",
           566 => x"90",
           567 => x"90",
           568 => x"90",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"04",
           585 => x"81",
           586 => x"83",
           587 => x"05",
           588 => x"10",
           589 => x"72",
           590 => x"51",
           591 => x"72",
           592 => x"06",
           593 => x"72",
           594 => x"10",
           595 => x"10",
           596 => x"ed",
           597 => x"53",
           598 => x"d3",
           599 => x"ea",
           600 => x"38",
           601 => x"84",
           602 => x"0b",
           603 => x"db",
           604 => x"51",
           605 => x"04",
           606 => x"90",
           607 => x"d3",
           608 => x"3d",
           609 => x"81",
           610 => x"8c",
           611 => x"81",
           612 => x"88",
           613 => x"83",
           614 => x"d3",
           615 => x"81",
           616 => x"54",
           617 => x"81",
           618 => x"04",
           619 => x"08",
           620 => x"90",
           621 => x"0d",
           622 => x"d3",
           623 => x"05",
           624 => x"d3",
           625 => x"05",
           626 => x"a1",
           627 => x"84",
           628 => x"d3",
           629 => x"85",
           630 => x"d3",
           631 => x"81",
           632 => x"02",
           633 => x"0c",
           634 => x"80",
           635 => x"90",
           636 => x"0c",
           637 => x"08",
           638 => x"80",
           639 => x"81",
           640 => x"88",
           641 => x"81",
           642 => x"88",
           643 => x"0b",
           644 => x"08",
           645 => x"81",
           646 => x"fc",
           647 => x"38",
           648 => x"d3",
           649 => x"05",
           650 => x"90",
           651 => x"08",
           652 => x"08",
           653 => x"81",
           654 => x"8c",
           655 => x"25",
           656 => x"d3",
           657 => x"05",
           658 => x"d3",
           659 => x"05",
           660 => x"81",
           661 => x"f0",
           662 => x"d3",
           663 => x"05",
           664 => x"81",
           665 => x"90",
           666 => x"0c",
           667 => x"08",
           668 => x"81",
           669 => x"fc",
           670 => x"53",
           671 => x"08",
           672 => x"52",
           673 => x"08",
           674 => x"51",
           675 => x"81",
           676 => x"70",
           677 => x"08",
           678 => x"54",
           679 => x"08",
           680 => x"80",
           681 => x"81",
           682 => x"f8",
           683 => x"81",
           684 => x"f8",
           685 => x"d3",
           686 => x"05",
           687 => x"d3",
           688 => x"89",
           689 => x"d3",
           690 => x"81",
           691 => x"02",
           692 => x"0c",
           693 => x"80",
           694 => x"90",
           695 => x"0c",
           696 => x"08",
           697 => x"80",
           698 => x"81",
           699 => x"88",
           700 => x"81",
           701 => x"88",
           702 => x"0b",
           703 => x"08",
           704 => x"81",
           705 => x"8c",
           706 => x"25",
           707 => x"d3",
           708 => x"05",
           709 => x"d3",
           710 => x"05",
           711 => x"81",
           712 => x"8c",
           713 => x"81",
           714 => x"88",
           715 => x"bd",
           716 => x"84",
           717 => x"d3",
           718 => x"05",
           719 => x"d3",
           720 => x"05",
           721 => x"90",
           722 => x"90",
           723 => x"08",
           724 => x"90",
           725 => x"0c",
           726 => x"08",
           727 => x"70",
           728 => x"0c",
           729 => x"0d",
           730 => x"0c",
           731 => x"90",
           732 => x"d3",
           733 => x"3d",
           734 => x"81",
           735 => x"fc",
           736 => x"0b",
           737 => x"08",
           738 => x"81",
           739 => x"8c",
           740 => x"d3",
           741 => x"05",
           742 => x"38",
           743 => x"08",
           744 => x"80",
           745 => x"80",
           746 => x"90",
           747 => x"08",
           748 => x"81",
           749 => x"8c",
           750 => x"81",
           751 => x"8c",
           752 => x"d3",
           753 => x"05",
           754 => x"d3",
           755 => x"05",
           756 => x"39",
           757 => x"08",
           758 => x"80",
           759 => x"38",
           760 => x"08",
           761 => x"81",
           762 => x"88",
           763 => x"ad",
           764 => x"90",
           765 => x"08",
           766 => x"08",
           767 => x"31",
           768 => x"08",
           769 => x"81",
           770 => x"f8",
           771 => x"d3",
           772 => x"05",
           773 => x"d3",
           774 => x"05",
           775 => x"90",
           776 => x"08",
           777 => x"d3",
           778 => x"05",
           779 => x"90",
           780 => x"08",
           781 => x"d3",
           782 => x"05",
           783 => x"39",
           784 => x"08",
           785 => x"80",
           786 => x"81",
           787 => x"88",
           788 => x"81",
           789 => x"f4",
           790 => x"91",
           791 => x"90",
           792 => x"08",
           793 => x"90",
           794 => x"0c",
           795 => x"90",
           796 => x"08",
           797 => x"0c",
           798 => x"81",
           799 => x"04",
           800 => x"76",
           801 => x"8c",
           802 => x"33",
           803 => x"55",
           804 => x"8a",
           805 => x"06",
           806 => x"2e",
           807 => x"12",
           808 => x"2e",
           809 => x"73",
           810 => x"55",
           811 => x"52",
           812 => x"09",
           813 => x"38",
           814 => x"84",
           815 => x"0d",
           816 => x"88",
           817 => x"70",
           818 => x"07",
           819 => x"8f",
           820 => x"38",
           821 => x"84",
           822 => x"72",
           823 => x"05",
           824 => x"71",
           825 => x"53",
           826 => x"70",
           827 => x"0c",
           828 => x"71",
           829 => x"38",
           830 => x"90",
           831 => x"70",
           832 => x"0c",
           833 => x"71",
           834 => x"38",
           835 => x"8e",
           836 => x"0d",
           837 => x"72",
           838 => x"53",
           839 => x"93",
           840 => x"73",
           841 => x"54",
           842 => x"2e",
           843 => x"73",
           844 => x"71",
           845 => x"ff",
           846 => x"70",
           847 => x"38",
           848 => x"70",
           849 => x"81",
           850 => x"81",
           851 => x"71",
           852 => x"ff",
           853 => x"54",
           854 => x"38",
           855 => x"73",
           856 => x"75",
           857 => x"71",
           858 => x"d3",
           859 => x"52",
           860 => x"04",
           861 => x"f7",
           862 => x"14",
           863 => x"84",
           864 => x"06",
           865 => x"70",
           866 => x"14",
           867 => x"08",
           868 => x"71",
           869 => x"dc",
           870 => x"54",
           871 => x"39",
           872 => x"d3",
           873 => x"3d",
           874 => x"3d",
           875 => x"83",
           876 => x"2b",
           877 => x"3f",
           878 => x"08",
           879 => x"72",
           880 => x"54",
           881 => x"25",
           882 => x"81",
           883 => x"84",
           884 => x"fb",
           885 => x"70",
           886 => x"53",
           887 => x"2e",
           888 => x"71",
           889 => x"a0",
           890 => x"06",
           891 => x"12",
           892 => x"71",
           893 => x"81",
           894 => x"73",
           895 => x"ff",
           896 => x"55",
           897 => x"83",
           898 => x"70",
           899 => x"38",
           900 => x"73",
           901 => x"51",
           902 => x"09",
           903 => x"38",
           904 => x"81",
           905 => x"72",
           906 => x"51",
           907 => x"84",
           908 => x"0d",
           909 => x"0d",
           910 => x"08",
           911 => x"38",
           912 => x"05",
           913 => x"98",
           914 => x"d3",
           915 => x"38",
           916 => x"39",
           917 => x"81",
           918 => x"86",
           919 => x"fc",
           920 => x"82",
           921 => x"05",
           922 => x"52",
           923 => x"81",
           924 => x"13",
           925 => x"51",
           926 => x"9e",
           927 => x"38",
           928 => x"51",
           929 => x"97",
           930 => x"38",
           931 => x"51",
           932 => x"bb",
           933 => x"38",
           934 => x"51",
           935 => x"bb",
           936 => x"38",
           937 => x"55",
           938 => x"87",
           939 => x"d9",
           940 => x"22",
           941 => x"73",
           942 => x"80",
           943 => x"0b",
           944 => x"9c",
           945 => x"87",
           946 => x"0c",
           947 => x"87",
           948 => x"0c",
           949 => x"87",
           950 => x"0c",
           951 => x"87",
           952 => x"0c",
           953 => x"87",
           954 => x"0c",
           955 => x"87",
           956 => x"0c",
           957 => x"98",
           958 => x"87",
           959 => x"0c",
           960 => x"c0",
           961 => x"80",
           962 => x"d3",
           963 => x"3d",
           964 => x"3d",
           965 => x"87",
           966 => x"5d",
           967 => x"87",
           968 => x"08",
           969 => x"23",
           970 => x"b8",
           971 => x"82",
           972 => x"c0",
           973 => x"5a",
           974 => x"34",
           975 => x"b0",
           976 => x"84",
           977 => x"c0",
           978 => x"5a",
           979 => x"34",
           980 => x"a8",
           981 => x"86",
           982 => x"c0",
           983 => x"5c",
           984 => x"23",
           985 => x"a0",
           986 => x"8a",
           987 => x"7d",
           988 => x"ff",
           989 => x"7b",
           990 => x"06",
           991 => x"33",
           992 => x"33",
           993 => x"33",
           994 => x"33",
           995 => x"33",
           996 => x"ff",
           997 => x"81",
           998 => x"92",
           999 => x"3d",
          1000 => x"3d",
          1001 => x"05",
          1002 => x"70",
          1003 => x"52",
          1004 => x"0b",
          1005 => x"34",
          1006 => x"04",
          1007 => x"77",
          1008 => x"cf",
          1009 => x"81",
          1010 => x"55",
          1011 => x"94",
          1012 => x"80",
          1013 => x"87",
          1014 => x"51",
          1015 => x"96",
          1016 => x"06",
          1017 => x"70",
          1018 => x"38",
          1019 => x"70",
          1020 => x"51",
          1021 => x"72",
          1022 => x"81",
          1023 => x"70",
          1024 => x"38",
          1025 => x"70",
          1026 => x"51",
          1027 => x"38",
          1028 => x"06",
          1029 => x"94",
          1030 => x"80",
          1031 => x"87",
          1032 => x"52",
          1033 => x"75",
          1034 => x"0c",
          1035 => x"04",
          1036 => x"02",
          1037 => x"0b",
          1038 => x"fc",
          1039 => x"ff",
          1040 => x"56",
          1041 => x"84",
          1042 => x"2e",
          1043 => x"c0",
          1044 => x"70",
          1045 => x"2a",
          1046 => x"53",
          1047 => x"80",
          1048 => x"71",
          1049 => x"81",
          1050 => x"70",
          1051 => x"81",
          1052 => x"06",
          1053 => x"80",
          1054 => x"71",
          1055 => x"81",
          1056 => x"70",
          1057 => x"73",
          1058 => x"51",
          1059 => x"80",
          1060 => x"2e",
          1061 => x"c0",
          1062 => x"75",
          1063 => x"3d",
          1064 => x"3d",
          1065 => x"80",
          1066 => x"81",
          1067 => x"53",
          1068 => x"2e",
          1069 => x"71",
          1070 => x"81",
          1071 => x"81",
          1072 => x"70",
          1073 => x"59",
          1074 => x"87",
          1075 => x"51",
          1076 => x"86",
          1077 => x"94",
          1078 => x"08",
          1079 => x"70",
          1080 => x"54",
          1081 => x"2e",
          1082 => x"91",
          1083 => x"06",
          1084 => x"d7",
          1085 => x"32",
          1086 => x"51",
          1087 => x"2e",
          1088 => x"93",
          1089 => x"06",
          1090 => x"ff",
          1091 => x"81",
          1092 => x"87",
          1093 => x"52",
          1094 => x"86",
          1095 => x"94",
          1096 => x"72",
          1097 => x"74",
          1098 => x"ff",
          1099 => x"57",
          1100 => x"38",
          1101 => x"84",
          1102 => x"0d",
          1103 => x"0d",
          1104 => x"cf",
          1105 => x"81",
          1106 => x"52",
          1107 => x"84",
          1108 => x"2e",
          1109 => x"c0",
          1110 => x"70",
          1111 => x"2a",
          1112 => x"51",
          1113 => x"80",
          1114 => x"71",
          1115 => x"51",
          1116 => x"80",
          1117 => x"2e",
          1118 => x"c0",
          1119 => x"71",
          1120 => x"ff",
          1121 => x"84",
          1122 => x"3d",
          1123 => x"3d",
          1124 => x"81",
          1125 => x"70",
          1126 => x"52",
          1127 => x"94",
          1128 => x"80",
          1129 => x"87",
          1130 => x"52",
          1131 => x"82",
          1132 => x"06",
          1133 => x"ff",
          1134 => x"2e",
          1135 => x"81",
          1136 => x"87",
          1137 => x"52",
          1138 => x"86",
          1139 => x"94",
          1140 => x"08",
          1141 => x"70",
          1142 => x"53",
          1143 => x"d3",
          1144 => x"3d",
          1145 => x"3d",
          1146 => x"9e",
          1147 => x"9c",
          1148 => x"51",
          1149 => x"2e",
          1150 => x"87",
          1151 => x"08",
          1152 => x"0c",
          1153 => x"a0",
          1154 => x"84",
          1155 => x"9e",
          1156 => x"d0",
          1157 => x"c0",
          1158 => x"81",
          1159 => x"87",
          1160 => x"08",
          1161 => x"0c",
          1162 => x"98",
          1163 => x"94",
          1164 => x"9e",
          1165 => x"d0",
          1166 => x"c0",
          1167 => x"81",
          1168 => x"87",
          1169 => x"08",
          1170 => x"0c",
          1171 => x"80",
          1172 => x"81",
          1173 => x"87",
          1174 => x"08",
          1175 => x"0c",
          1176 => x"d0",
          1177 => x"0b",
          1178 => x"88",
          1179 => x"80",
          1180 => x"52",
          1181 => x"83",
          1182 => x"71",
          1183 => x"34",
          1184 => x"c0",
          1185 => x"70",
          1186 => x"06",
          1187 => x"70",
          1188 => x"38",
          1189 => x"81",
          1190 => x"80",
          1191 => x"9e",
          1192 => x"80",
          1193 => x"51",
          1194 => x"80",
          1195 => x"81",
          1196 => x"d0",
          1197 => x"0b",
          1198 => x"88",
          1199 => x"80",
          1200 => x"52",
          1201 => x"83",
          1202 => x"71",
          1203 => x"34",
          1204 => x"c0",
          1205 => x"70",
          1206 => x"51",
          1207 => x"80",
          1208 => x"81",
          1209 => x"d0",
          1210 => x"0b",
          1211 => x"88",
          1212 => x"80",
          1213 => x"52",
          1214 => x"83",
          1215 => x"71",
          1216 => x"34",
          1217 => x"c0",
          1218 => x"70",
          1219 => x"51",
          1220 => x"80",
          1221 => x"81",
          1222 => x"d0",
          1223 => x"0b",
          1224 => x"88",
          1225 => x"80",
          1226 => x"52",
          1227 => x"83",
          1228 => x"71",
          1229 => x"34",
          1230 => x"88",
          1231 => x"e0",
          1232 => x"2c",
          1233 => x"70",
          1234 => x"34",
          1235 => x"c0",
          1236 => x"70",
          1237 => x"52",
          1238 => x"2e",
          1239 => x"52",
          1240 => x"b6",
          1241 => x"87",
          1242 => x"08",
          1243 => x"51",
          1244 => x"80",
          1245 => x"81",
          1246 => x"d0",
          1247 => x"c0",
          1248 => x"70",
          1249 => x"51",
          1250 => x"b8",
          1251 => x"0d",
          1252 => x"0d",
          1253 => x"51",
          1254 => x"81",
          1255 => x"54",
          1256 => x"88",
          1257 => x"fc",
          1258 => x"3f",
          1259 => x"51",
          1260 => x"81",
          1261 => x"54",
          1262 => x"92",
          1263 => x"84",
          1264 => x"d0",
          1265 => x"81",
          1266 => x"89",
          1267 => x"d0",
          1268 => x"73",
          1269 => x"38",
          1270 => x"08",
          1271 => x"88",
          1272 => x"be",
          1273 => x"b7",
          1274 => x"af",
          1275 => x"8b",
          1276 => x"b0",
          1277 => x"80",
          1278 => x"81",
          1279 => x"53",
          1280 => x"08",
          1281 => x"f4",
          1282 => x"3f",
          1283 => x"33",
          1284 => x"2e",
          1285 => x"bf",
          1286 => x"9f",
          1287 => x"b2",
          1288 => x"80",
          1289 => x"81",
          1290 => x"83",
          1291 => x"d0",
          1292 => x"73",
          1293 => x"38",
          1294 => x"51",
          1295 => x"81",
          1296 => x"54",
          1297 => x"8d",
          1298 => x"b5",
          1299 => x"bf",
          1300 => x"cb",
          1301 => x"b6",
          1302 => x"80",
          1303 => x"81",
          1304 => x"82",
          1305 => x"d0",
          1306 => x"73",
          1307 => x"38",
          1308 => x"33",
          1309 => x"f8",
          1310 => x"3f",
          1311 => x"51",
          1312 => x"81",
          1313 => x"52",
          1314 => x"51",
          1315 => x"81",
          1316 => x"52",
          1317 => x"51",
          1318 => x"81",
          1319 => x"52",
          1320 => x"51",
          1321 => x"81",
          1322 => x"52",
          1323 => x"51",
          1324 => x"81",
          1325 => x"52",
          1326 => x"51",
          1327 => x"85",
          1328 => x"fe",
          1329 => x"92",
          1330 => x"05",
          1331 => x"26",
          1332 => x"84",
          1333 => x"ec",
          1334 => x"08",
          1335 => x"e8",
          1336 => x"81",
          1337 => x"97",
          1338 => x"f8",
          1339 => x"81",
          1340 => x"8b",
          1341 => x"84",
          1342 => x"81",
          1343 => x"f7",
          1344 => x"3d",
          1345 => x"88",
          1346 => x"80",
          1347 => x"96",
          1348 => x"ff",
          1349 => x"c0",
          1350 => x"08",
          1351 => x"72",
          1352 => x"07",
          1353 => x"bc",
          1354 => x"83",
          1355 => x"ff",
          1356 => x"c0",
          1357 => x"08",
          1358 => x"0c",
          1359 => x"0c",
          1360 => x"81",
          1361 => x"06",
          1362 => x"bc",
          1363 => x"51",
          1364 => x"04",
          1365 => x"08",
          1366 => x"84",
          1367 => x"3d",
          1368 => x"05",
          1369 => x"8a",
          1370 => x"06",
          1371 => x"51",
          1372 => x"d3",
          1373 => x"71",
          1374 => x"38",
          1375 => x"81",
          1376 => x"81",
          1377 => x"9c",
          1378 => x"81",
          1379 => x"52",
          1380 => x"85",
          1381 => x"71",
          1382 => x"0d",
          1383 => x"0d",
          1384 => x"33",
          1385 => x"08",
          1386 => x"94",
          1387 => x"ff",
          1388 => x"81",
          1389 => x"84",
          1390 => x"fd",
          1391 => x"54",
          1392 => x"81",
          1393 => x"53",
          1394 => x"8e",
          1395 => x"ff",
          1396 => x"14",
          1397 => x"3f",
          1398 => x"3d",
          1399 => x"3d",
          1400 => x"d3",
          1401 => x"81",
          1402 => x"56",
          1403 => x"70",
          1404 => x"53",
          1405 => x"2e",
          1406 => x"81",
          1407 => x"81",
          1408 => x"da",
          1409 => x"74",
          1410 => x"0c",
          1411 => x"04",
          1412 => x"66",
          1413 => x"78",
          1414 => x"5a",
          1415 => x"80",
          1416 => x"38",
          1417 => x"09",
          1418 => x"de",
          1419 => x"7a",
          1420 => x"5c",
          1421 => x"5b",
          1422 => x"09",
          1423 => x"38",
          1424 => x"39",
          1425 => x"09",
          1426 => x"38",
          1427 => x"70",
          1428 => x"33",
          1429 => x"2e",
          1430 => x"92",
          1431 => x"19",
          1432 => x"70",
          1433 => x"33",
          1434 => x"53",
          1435 => x"16",
          1436 => x"26",
          1437 => x"88",
          1438 => x"05",
          1439 => x"05",
          1440 => x"05",
          1441 => x"5b",
          1442 => x"80",
          1443 => x"30",
          1444 => x"80",
          1445 => x"cc",
          1446 => x"70",
          1447 => x"25",
          1448 => x"54",
          1449 => x"53",
          1450 => x"8c",
          1451 => x"07",
          1452 => x"05",
          1453 => x"5a",
          1454 => x"83",
          1455 => x"54",
          1456 => x"27",
          1457 => x"16",
          1458 => x"06",
          1459 => x"80",
          1460 => x"aa",
          1461 => x"cf",
          1462 => x"73",
          1463 => x"81",
          1464 => x"80",
          1465 => x"38",
          1466 => x"2e",
          1467 => x"81",
          1468 => x"80",
          1469 => x"8a",
          1470 => x"39",
          1471 => x"2e",
          1472 => x"73",
          1473 => x"8a",
          1474 => x"d3",
          1475 => x"80",
          1476 => x"80",
          1477 => x"ee",
          1478 => x"39",
          1479 => x"71",
          1480 => x"53",
          1481 => x"54",
          1482 => x"2e",
          1483 => x"15",
          1484 => x"33",
          1485 => x"72",
          1486 => x"81",
          1487 => x"39",
          1488 => x"56",
          1489 => x"27",
          1490 => x"51",
          1491 => x"75",
          1492 => x"72",
          1493 => x"38",
          1494 => x"df",
          1495 => x"16",
          1496 => x"7b",
          1497 => x"38",
          1498 => x"f2",
          1499 => x"77",
          1500 => x"12",
          1501 => x"53",
          1502 => x"5c",
          1503 => x"5c",
          1504 => x"5c",
          1505 => x"5c",
          1506 => x"51",
          1507 => x"fd",
          1508 => x"82",
          1509 => x"06",
          1510 => x"80",
          1511 => x"77",
          1512 => x"53",
          1513 => x"18",
          1514 => x"72",
          1515 => x"c4",
          1516 => x"70",
          1517 => x"25",
          1518 => x"55",
          1519 => x"8d",
          1520 => x"2e",
          1521 => x"30",
          1522 => x"5b",
          1523 => x"8f",
          1524 => x"7b",
          1525 => x"e3",
          1526 => x"d3",
          1527 => x"ff",
          1528 => x"75",
          1529 => x"91",
          1530 => x"84",
          1531 => x"74",
          1532 => x"a7",
          1533 => x"80",
          1534 => x"38",
          1535 => x"72",
          1536 => x"54",
          1537 => x"72",
          1538 => x"05",
          1539 => x"17",
          1540 => x"77",
          1541 => x"51",
          1542 => x"9f",
          1543 => x"72",
          1544 => x"79",
          1545 => x"81",
          1546 => x"72",
          1547 => x"38",
          1548 => x"05",
          1549 => x"ad",
          1550 => x"17",
          1551 => x"81",
          1552 => x"b0",
          1553 => x"38",
          1554 => x"81",
          1555 => x"06",
          1556 => x"9f",
          1557 => x"55",
          1558 => x"97",
          1559 => x"f9",
          1560 => x"81",
          1561 => x"8b",
          1562 => x"16",
          1563 => x"73",
          1564 => x"96",
          1565 => x"e0",
          1566 => x"17",
          1567 => x"33",
          1568 => x"f9",
          1569 => x"f2",
          1570 => x"16",
          1571 => x"7b",
          1572 => x"38",
          1573 => x"c6",
          1574 => x"96",
          1575 => x"fd",
          1576 => x"3d",
          1577 => x"05",
          1578 => x"52",
          1579 => x"e0",
          1580 => x"0d",
          1581 => x"0d",
          1582 => x"9c",
          1583 => x"88",
          1584 => x"51",
          1585 => x"81",
          1586 => x"53",
          1587 => x"80",
          1588 => x"9c",
          1589 => x"0d",
          1590 => x"0d",
          1591 => x"08",
          1592 => x"94",
          1593 => x"88",
          1594 => x"52",
          1595 => x"3f",
          1596 => x"94",
          1597 => x"0d",
          1598 => x"0d",
          1599 => x"d3",
          1600 => x"56",
          1601 => x"80",
          1602 => x"2e",
          1603 => x"81",
          1604 => x"52",
          1605 => x"d3",
          1606 => x"ff",
          1607 => x"80",
          1608 => x"38",
          1609 => x"b9",
          1610 => x"32",
          1611 => x"80",
          1612 => x"52",
          1613 => x"8b",
          1614 => x"2e",
          1615 => x"14",
          1616 => x"9f",
          1617 => x"38",
          1618 => x"73",
          1619 => x"38",
          1620 => x"72",
          1621 => x"14",
          1622 => x"f8",
          1623 => x"af",
          1624 => x"52",
          1625 => x"8a",
          1626 => x"3f",
          1627 => x"81",
          1628 => x"87",
          1629 => x"fe",
          1630 => x"d3",
          1631 => x"81",
          1632 => x"77",
          1633 => x"53",
          1634 => x"72",
          1635 => x"0c",
          1636 => x"04",
          1637 => x"7a",
          1638 => x"80",
          1639 => x"58",
          1640 => x"33",
          1641 => x"a0",
          1642 => x"06",
          1643 => x"13",
          1644 => x"39",
          1645 => x"09",
          1646 => x"38",
          1647 => x"11",
          1648 => x"08",
          1649 => x"54",
          1650 => x"2e",
          1651 => x"80",
          1652 => x"08",
          1653 => x"0c",
          1654 => x"33",
          1655 => x"80",
          1656 => x"38",
          1657 => x"80",
          1658 => x"38",
          1659 => x"57",
          1660 => x"0c",
          1661 => x"33",
          1662 => x"39",
          1663 => x"74",
          1664 => x"38",
          1665 => x"80",
          1666 => x"89",
          1667 => x"38",
          1668 => x"d0",
          1669 => x"55",
          1670 => x"80",
          1671 => x"39",
          1672 => x"d9",
          1673 => x"80",
          1674 => x"27",
          1675 => x"80",
          1676 => x"89",
          1677 => x"70",
          1678 => x"55",
          1679 => x"70",
          1680 => x"55",
          1681 => x"27",
          1682 => x"14",
          1683 => x"06",
          1684 => x"74",
          1685 => x"73",
          1686 => x"38",
          1687 => x"14",
          1688 => x"05",
          1689 => x"08",
          1690 => x"54",
          1691 => x"39",
          1692 => x"84",
          1693 => x"55",
          1694 => x"81",
          1695 => x"d3",
          1696 => x"3d",
          1697 => x"3d",
          1698 => x"5a",
          1699 => x"7a",
          1700 => x"08",
          1701 => x"53",
          1702 => x"09",
          1703 => x"38",
          1704 => x"0c",
          1705 => x"ad",
          1706 => x"06",
          1707 => x"76",
          1708 => x"0c",
          1709 => x"33",
          1710 => x"73",
          1711 => x"81",
          1712 => x"38",
          1713 => x"05",
          1714 => x"08",
          1715 => x"53",
          1716 => x"2e",
          1717 => x"57",
          1718 => x"2e",
          1719 => x"39",
          1720 => x"13",
          1721 => x"08",
          1722 => x"53",
          1723 => x"55",
          1724 => x"80",
          1725 => x"14",
          1726 => x"88",
          1727 => x"27",
          1728 => x"eb",
          1729 => x"53",
          1730 => x"89",
          1731 => x"38",
          1732 => x"55",
          1733 => x"8a",
          1734 => x"a0",
          1735 => x"c2",
          1736 => x"74",
          1737 => x"e0",
          1738 => x"ff",
          1739 => x"d0",
          1740 => x"ff",
          1741 => x"90",
          1742 => x"38",
          1743 => x"81",
          1744 => x"53",
          1745 => x"ca",
          1746 => x"27",
          1747 => x"77",
          1748 => x"08",
          1749 => x"0c",
          1750 => x"33",
          1751 => x"ff",
          1752 => x"80",
          1753 => x"74",
          1754 => x"79",
          1755 => x"74",
          1756 => x"0c",
          1757 => x"04",
          1758 => x"02",
          1759 => x"51",
          1760 => x"72",
          1761 => x"81",
          1762 => x"33",
          1763 => x"d3",
          1764 => x"3d",
          1765 => x"3d",
          1766 => x"05",
          1767 => x"05",
          1768 => x"56",
          1769 => x"72",
          1770 => x"e0",
          1771 => x"2b",
          1772 => x"8c",
          1773 => x"88",
          1774 => x"2e",
          1775 => x"88",
          1776 => x"0c",
          1777 => x"8c",
          1778 => x"71",
          1779 => x"87",
          1780 => x"0c",
          1781 => x"08",
          1782 => x"51",
          1783 => x"2e",
          1784 => x"c0",
          1785 => x"51",
          1786 => x"71",
          1787 => x"80",
          1788 => x"92",
          1789 => x"98",
          1790 => x"70",
          1791 => x"38",
          1792 => x"c0",
          1793 => x"d0",
          1794 => x"51",
          1795 => x"84",
          1796 => x"0d",
          1797 => x"0d",
          1798 => x"02",
          1799 => x"05",
          1800 => x"58",
          1801 => x"52",
          1802 => x"3f",
          1803 => x"08",
          1804 => x"54",
          1805 => x"be",
          1806 => x"75",
          1807 => x"c0",
          1808 => x"87",
          1809 => x"12",
          1810 => x"84",
          1811 => x"40",
          1812 => x"85",
          1813 => x"98",
          1814 => x"7d",
          1815 => x"0c",
          1816 => x"85",
          1817 => x"06",
          1818 => x"71",
          1819 => x"38",
          1820 => x"71",
          1821 => x"05",
          1822 => x"19",
          1823 => x"a2",
          1824 => x"71",
          1825 => x"38",
          1826 => x"83",
          1827 => x"38",
          1828 => x"8a",
          1829 => x"98",
          1830 => x"71",
          1831 => x"c0",
          1832 => x"52",
          1833 => x"87",
          1834 => x"80",
          1835 => x"81",
          1836 => x"c0",
          1837 => x"53",
          1838 => x"82",
          1839 => x"71",
          1840 => x"1a",
          1841 => x"84",
          1842 => x"19",
          1843 => x"06",
          1844 => x"79",
          1845 => x"38",
          1846 => x"80",
          1847 => x"87",
          1848 => x"26",
          1849 => x"73",
          1850 => x"06",
          1851 => x"2e",
          1852 => x"52",
          1853 => x"81",
          1854 => x"8f",
          1855 => x"f3",
          1856 => x"62",
          1857 => x"05",
          1858 => x"57",
          1859 => x"83",
          1860 => x"52",
          1861 => x"3f",
          1862 => x"08",
          1863 => x"54",
          1864 => x"2e",
          1865 => x"81",
          1866 => x"74",
          1867 => x"c0",
          1868 => x"87",
          1869 => x"12",
          1870 => x"84",
          1871 => x"5f",
          1872 => x"0b",
          1873 => x"8c",
          1874 => x"0c",
          1875 => x"80",
          1876 => x"70",
          1877 => x"81",
          1878 => x"54",
          1879 => x"8c",
          1880 => x"81",
          1881 => x"7c",
          1882 => x"58",
          1883 => x"70",
          1884 => x"52",
          1885 => x"8a",
          1886 => x"98",
          1887 => x"71",
          1888 => x"c0",
          1889 => x"52",
          1890 => x"87",
          1891 => x"80",
          1892 => x"81",
          1893 => x"c0",
          1894 => x"53",
          1895 => x"82",
          1896 => x"71",
          1897 => x"19",
          1898 => x"81",
          1899 => x"ff",
          1900 => x"19",
          1901 => x"78",
          1902 => x"38",
          1903 => x"80",
          1904 => x"87",
          1905 => x"26",
          1906 => x"73",
          1907 => x"06",
          1908 => x"2e",
          1909 => x"52",
          1910 => x"81",
          1911 => x"8f",
          1912 => x"f6",
          1913 => x"02",
          1914 => x"05",
          1915 => x"05",
          1916 => x"71",
          1917 => x"57",
          1918 => x"81",
          1919 => x"81",
          1920 => x"54",
          1921 => x"38",
          1922 => x"c0",
          1923 => x"81",
          1924 => x"2e",
          1925 => x"71",
          1926 => x"38",
          1927 => x"87",
          1928 => x"11",
          1929 => x"80",
          1930 => x"80",
          1931 => x"83",
          1932 => x"38",
          1933 => x"72",
          1934 => x"2a",
          1935 => x"51",
          1936 => x"80",
          1937 => x"87",
          1938 => x"08",
          1939 => x"38",
          1940 => x"8c",
          1941 => x"96",
          1942 => x"0c",
          1943 => x"8c",
          1944 => x"08",
          1945 => x"51",
          1946 => x"38",
          1947 => x"56",
          1948 => x"80",
          1949 => x"85",
          1950 => x"77",
          1951 => x"83",
          1952 => x"75",
          1953 => x"d3",
          1954 => x"3d",
          1955 => x"3d",
          1956 => x"11",
          1957 => x"71",
          1958 => x"81",
          1959 => x"53",
          1960 => x"0d",
          1961 => x"0d",
          1962 => x"33",
          1963 => x"71",
          1964 => x"88",
          1965 => x"14",
          1966 => x"07",
          1967 => x"33",
          1968 => x"d3",
          1969 => x"53",
          1970 => x"52",
          1971 => x"04",
          1972 => x"73",
          1973 => x"92",
          1974 => x"52",
          1975 => x"81",
          1976 => x"70",
          1977 => x"70",
          1978 => x"3d",
          1979 => x"3d",
          1980 => x"52",
          1981 => x"70",
          1982 => x"34",
          1983 => x"51",
          1984 => x"81",
          1985 => x"70",
          1986 => x"70",
          1987 => x"05",
          1988 => x"88",
          1989 => x"72",
          1990 => x"0d",
          1991 => x"0d",
          1992 => x"54",
          1993 => x"80",
          1994 => x"71",
          1995 => x"53",
          1996 => x"81",
          1997 => x"ff",
          1998 => x"39",
          1999 => x"04",
          2000 => x"75",
          2001 => x"52",
          2002 => x"70",
          2003 => x"34",
          2004 => x"70",
          2005 => x"3d",
          2006 => x"3d",
          2007 => x"79",
          2008 => x"74",
          2009 => x"56",
          2010 => x"81",
          2011 => x"71",
          2012 => x"16",
          2013 => x"52",
          2014 => x"86",
          2015 => x"2e",
          2016 => x"81",
          2017 => x"86",
          2018 => x"fe",
          2019 => x"76",
          2020 => x"39",
          2021 => x"8a",
          2022 => x"51",
          2023 => x"71",
          2024 => x"33",
          2025 => x"0c",
          2026 => x"04",
          2027 => x"d3",
          2028 => x"80",
          2029 => x"84",
          2030 => x"3d",
          2031 => x"80",
          2032 => x"33",
          2033 => x"7a",
          2034 => x"38",
          2035 => x"16",
          2036 => x"16",
          2037 => x"17",
          2038 => x"fa",
          2039 => x"d3",
          2040 => x"2e",
          2041 => x"b7",
          2042 => x"84",
          2043 => x"34",
          2044 => x"70",
          2045 => x"31",
          2046 => x"59",
          2047 => x"77",
          2048 => x"82",
          2049 => x"74",
          2050 => x"81",
          2051 => x"81",
          2052 => x"53",
          2053 => x"16",
          2054 => x"e3",
          2055 => x"81",
          2056 => x"d3",
          2057 => x"3d",
          2058 => x"3d",
          2059 => x"56",
          2060 => x"74",
          2061 => x"2e",
          2062 => x"51",
          2063 => x"81",
          2064 => x"57",
          2065 => x"08",
          2066 => x"54",
          2067 => x"16",
          2068 => x"33",
          2069 => x"3f",
          2070 => x"08",
          2071 => x"38",
          2072 => x"57",
          2073 => x"0c",
          2074 => x"84",
          2075 => x"0d",
          2076 => x"0d",
          2077 => x"57",
          2078 => x"81",
          2079 => x"58",
          2080 => x"08",
          2081 => x"76",
          2082 => x"83",
          2083 => x"06",
          2084 => x"84",
          2085 => x"78",
          2086 => x"81",
          2087 => x"38",
          2088 => x"81",
          2089 => x"52",
          2090 => x"52",
          2091 => x"3f",
          2092 => x"52",
          2093 => x"51",
          2094 => x"84",
          2095 => x"d2",
          2096 => x"fc",
          2097 => x"8a",
          2098 => x"52",
          2099 => x"51",
          2100 => x"90",
          2101 => x"84",
          2102 => x"fc",
          2103 => x"17",
          2104 => x"a0",
          2105 => x"86",
          2106 => x"08",
          2107 => x"b0",
          2108 => x"55",
          2109 => x"81",
          2110 => x"f8",
          2111 => x"84",
          2112 => x"53",
          2113 => x"17",
          2114 => x"d7",
          2115 => x"84",
          2116 => x"83",
          2117 => x"77",
          2118 => x"0c",
          2119 => x"04",
          2120 => x"77",
          2121 => x"12",
          2122 => x"55",
          2123 => x"56",
          2124 => x"8d",
          2125 => x"22",
          2126 => x"ac",
          2127 => x"57",
          2128 => x"d3",
          2129 => x"3d",
          2130 => x"3d",
          2131 => x"70",
          2132 => x"57",
          2133 => x"81",
          2134 => x"98",
          2135 => x"81",
          2136 => x"74",
          2137 => x"72",
          2138 => x"f5",
          2139 => x"24",
          2140 => x"81",
          2141 => x"81",
          2142 => x"83",
          2143 => x"38",
          2144 => x"76",
          2145 => x"70",
          2146 => x"16",
          2147 => x"74",
          2148 => x"96",
          2149 => x"84",
          2150 => x"38",
          2151 => x"06",
          2152 => x"33",
          2153 => x"89",
          2154 => x"08",
          2155 => x"54",
          2156 => x"fc",
          2157 => x"d3",
          2158 => x"fe",
          2159 => x"ff",
          2160 => x"11",
          2161 => x"2b",
          2162 => x"81",
          2163 => x"2a",
          2164 => x"51",
          2165 => x"e2",
          2166 => x"ff",
          2167 => x"da",
          2168 => x"2a",
          2169 => x"05",
          2170 => x"fc",
          2171 => x"d3",
          2172 => x"c6",
          2173 => x"83",
          2174 => x"05",
          2175 => x"f9",
          2176 => x"d3",
          2177 => x"ff",
          2178 => x"ae",
          2179 => x"2a",
          2180 => x"05",
          2181 => x"fc",
          2182 => x"d3",
          2183 => x"38",
          2184 => x"83",
          2185 => x"05",
          2186 => x"f8",
          2187 => x"d3",
          2188 => x"0a",
          2189 => x"39",
          2190 => x"81",
          2191 => x"89",
          2192 => x"f8",
          2193 => x"7c",
          2194 => x"56",
          2195 => x"77",
          2196 => x"38",
          2197 => x"08",
          2198 => x"38",
          2199 => x"72",
          2200 => x"9d",
          2201 => x"24",
          2202 => x"81",
          2203 => x"82",
          2204 => x"83",
          2205 => x"38",
          2206 => x"76",
          2207 => x"70",
          2208 => x"18",
          2209 => x"76",
          2210 => x"9e",
          2211 => x"84",
          2212 => x"d3",
          2213 => x"d9",
          2214 => x"ff",
          2215 => x"05",
          2216 => x"81",
          2217 => x"54",
          2218 => x"80",
          2219 => x"77",
          2220 => x"f0",
          2221 => x"8f",
          2222 => x"51",
          2223 => x"34",
          2224 => x"17",
          2225 => x"2a",
          2226 => x"05",
          2227 => x"fa",
          2228 => x"d3",
          2229 => x"81",
          2230 => x"81",
          2231 => x"83",
          2232 => x"b4",
          2233 => x"2a",
          2234 => x"8f",
          2235 => x"2a",
          2236 => x"f0",
          2237 => x"06",
          2238 => x"72",
          2239 => x"ec",
          2240 => x"2a",
          2241 => x"05",
          2242 => x"fa",
          2243 => x"d3",
          2244 => x"81",
          2245 => x"80",
          2246 => x"83",
          2247 => x"52",
          2248 => x"fe",
          2249 => x"b4",
          2250 => x"a4",
          2251 => x"76",
          2252 => x"17",
          2253 => x"75",
          2254 => x"3f",
          2255 => x"08",
          2256 => x"84",
          2257 => x"77",
          2258 => x"77",
          2259 => x"fc",
          2260 => x"b4",
          2261 => x"51",
          2262 => x"c9",
          2263 => x"84",
          2264 => x"06",
          2265 => x"72",
          2266 => x"3f",
          2267 => x"17",
          2268 => x"d3",
          2269 => x"3d",
          2270 => x"3d",
          2271 => x"7e",
          2272 => x"56",
          2273 => x"75",
          2274 => x"74",
          2275 => x"27",
          2276 => x"80",
          2277 => x"ff",
          2278 => x"75",
          2279 => x"3f",
          2280 => x"08",
          2281 => x"84",
          2282 => x"38",
          2283 => x"54",
          2284 => x"81",
          2285 => x"39",
          2286 => x"08",
          2287 => x"39",
          2288 => x"51",
          2289 => x"81",
          2290 => x"58",
          2291 => x"08",
          2292 => x"c7",
          2293 => x"84",
          2294 => x"d2",
          2295 => x"84",
          2296 => x"cf",
          2297 => x"74",
          2298 => x"fc",
          2299 => x"d3",
          2300 => x"38",
          2301 => x"fe",
          2302 => x"08",
          2303 => x"74",
          2304 => x"38",
          2305 => x"17",
          2306 => x"33",
          2307 => x"73",
          2308 => x"77",
          2309 => x"26",
          2310 => x"80",
          2311 => x"d3",
          2312 => x"3d",
          2313 => x"3d",
          2314 => x"71",
          2315 => x"5b",
          2316 => x"8c",
          2317 => x"77",
          2318 => x"38",
          2319 => x"78",
          2320 => x"81",
          2321 => x"79",
          2322 => x"f9",
          2323 => x"55",
          2324 => x"84",
          2325 => x"e0",
          2326 => x"84",
          2327 => x"d3",
          2328 => x"2e",
          2329 => x"98",
          2330 => x"d3",
          2331 => x"82",
          2332 => x"58",
          2333 => x"70",
          2334 => x"80",
          2335 => x"38",
          2336 => x"09",
          2337 => x"e2",
          2338 => x"56",
          2339 => x"76",
          2340 => x"82",
          2341 => x"7a",
          2342 => x"3f",
          2343 => x"d3",
          2344 => x"2e",
          2345 => x"86",
          2346 => x"84",
          2347 => x"d3",
          2348 => x"70",
          2349 => x"07",
          2350 => x"7c",
          2351 => x"84",
          2352 => x"51",
          2353 => x"81",
          2354 => x"d3",
          2355 => x"2e",
          2356 => x"17",
          2357 => x"74",
          2358 => x"73",
          2359 => x"27",
          2360 => x"58",
          2361 => x"80",
          2362 => x"56",
          2363 => x"98",
          2364 => x"26",
          2365 => x"56",
          2366 => x"81",
          2367 => x"52",
          2368 => x"c6",
          2369 => x"84",
          2370 => x"b8",
          2371 => x"81",
          2372 => x"81",
          2373 => x"06",
          2374 => x"d3",
          2375 => x"81",
          2376 => x"09",
          2377 => x"72",
          2378 => x"70",
          2379 => x"51",
          2380 => x"80",
          2381 => x"78",
          2382 => x"06",
          2383 => x"73",
          2384 => x"39",
          2385 => x"52",
          2386 => x"f7",
          2387 => x"84",
          2388 => x"84",
          2389 => x"81",
          2390 => x"07",
          2391 => x"55",
          2392 => x"2e",
          2393 => x"80",
          2394 => x"75",
          2395 => x"76",
          2396 => x"3f",
          2397 => x"08",
          2398 => x"38",
          2399 => x"0c",
          2400 => x"fe",
          2401 => x"08",
          2402 => x"74",
          2403 => x"ff",
          2404 => x"0c",
          2405 => x"81",
          2406 => x"84",
          2407 => x"39",
          2408 => x"81",
          2409 => x"8c",
          2410 => x"8c",
          2411 => x"84",
          2412 => x"39",
          2413 => x"55",
          2414 => x"84",
          2415 => x"0d",
          2416 => x"0d",
          2417 => x"55",
          2418 => x"81",
          2419 => x"58",
          2420 => x"d3",
          2421 => x"d8",
          2422 => x"74",
          2423 => x"3f",
          2424 => x"08",
          2425 => x"08",
          2426 => x"59",
          2427 => x"77",
          2428 => x"70",
          2429 => x"c8",
          2430 => x"84",
          2431 => x"56",
          2432 => x"58",
          2433 => x"97",
          2434 => x"75",
          2435 => x"52",
          2436 => x"51",
          2437 => x"81",
          2438 => x"80",
          2439 => x"8a",
          2440 => x"32",
          2441 => x"72",
          2442 => x"2a",
          2443 => x"56",
          2444 => x"84",
          2445 => x"0d",
          2446 => x"0d",
          2447 => x"08",
          2448 => x"74",
          2449 => x"26",
          2450 => x"74",
          2451 => x"72",
          2452 => x"74",
          2453 => x"88",
          2454 => x"73",
          2455 => x"33",
          2456 => x"27",
          2457 => x"16",
          2458 => x"9b",
          2459 => x"2a",
          2460 => x"88",
          2461 => x"58",
          2462 => x"80",
          2463 => x"16",
          2464 => x"0c",
          2465 => x"8a",
          2466 => x"89",
          2467 => x"72",
          2468 => x"38",
          2469 => x"51",
          2470 => x"81",
          2471 => x"54",
          2472 => x"08",
          2473 => x"38",
          2474 => x"d3",
          2475 => x"8b",
          2476 => x"08",
          2477 => x"08",
          2478 => x"82",
          2479 => x"74",
          2480 => x"cb",
          2481 => x"75",
          2482 => x"3f",
          2483 => x"08",
          2484 => x"73",
          2485 => x"98",
          2486 => x"82",
          2487 => x"2e",
          2488 => x"39",
          2489 => x"39",
          2490 => x"13",
          2491 => x"74",
          2492 => x"16",
          2493 => x"18",
          2494 => x"77",
          2495 => x"0c",
          2496 => x"04",
          2497 => x"7a",
          2498 => x"12",
          2499 => x"59",
          2500 => x"80",
          2501 => x"86",
          2502 => x"98",
          2503 => x"14",
          2504 => x"55",
          2505 => x"81",
          2506 => x"83",
          2507 => x"77",
          2508 => x"81",
          2509 => x"0c",
          2510 => x"55",
          2511 => x"76",
          2512 => x"17",
          2513 => x"74",
          2514 => x"9b",
          2515 => x"39",
          2516 => x"ff",
          2517 => x"2a",
          2518 => x"81",
          2519 => x"52",
          2520 => x"e6",
          2521 => x"84",
          2522 => x"55",
          2523 => x"d3",
          2524 => x"80",
          2525 => x"55",
          2526 => x"08",
          2527 => x"f4",
          2528 => x"08",
          2529 => x"08",
          2530 => x"38",
          2531 => x"77",
          2532 => x"84",
          2533 => x"39",
          2534 => x"52",
          2535 => x"86",
          2536 => x"84",
          2537 => x"55",
          2538 => x"08",
          2539 => x"c4",
          2540 => x"81",
          2541 => x"81",
          2542 => x"81",
          2543 => x"84",
          2544 => x"b0",
          2545 => x"84",
          2546 => x"51",
          2547 => x"81",
          2548 => x"a0",
          2549 => x"15",
          2550 => x"75",
          2551 => x"3f",
          2552 => x"08",
          2553 => x"76",
          2554 => x"77",
          2555 => x"9c",
          2556 => x"55",
          2557 => x"84",
          2558 => x"0d",
          2559 => x"0d",
          2560 => x"08",
          2561 => x"80",
          2562 => x"fc",
          2563 => x"d3",
          2564 => x"81",
          2565 => x"80",
          2566 => x"d3",
          2567 => x"98",
          2568 => x"78",
          2569 => x"3f",
          2570 => x"08",
          2571 => x"84",
          2572 => x"38",
          2573 => x"08",
          2574 => x"70",
          2575 => x"58",
          2576 => x"2e",
          2577 => x"83",
          2578 => x"81",
          2579 => x"55",
          2580 => x"81",
          2581 => x"07",
          2582 => x"2e",
          2583 => x"16",
          2584 => x"2e",
          2585 => x"88",
          2586 => x"81",
          2587 => x"56",
          2588 => x"51",
          2589 => x"81",
          2590 => x"54",
          2591 => x"08",
          2592 => x"9b",
          2593 => x"2e",
          2594 => x"83",
          2595 => x"73",
          2596 => x"0c",
          2597 => x"04",
          2598 => x"76",
          2599 => x"54",
          2600 => x"81",
          2601 => x"83",
          2602 => x"76",
          2603 => x"53",
          2604 => x"2e",
          2605 => x"90",
          2606 => x"51",
          2607 => x"81",
          2608 => x"90",
          2609 => x"53",
          2610 => x"84",
          2611 => x"0d",
          2612 => x"0d",
          2613 => x"83",
          2614 => x"54",
          2615 => x"55",
          2616 => x"3f",
          2617 => x"51",
          2618 => x"2e",
          2619 => x"8b",
          2620 => x"2a",
          2621 => x"51",
          2622 => x"86",
          2623 => x"f7",
          2624 => x"7d",
          2625 => x"75",
          2626 => x"98",
          2627 => x"2e",
          2628 => x"98",
          2629 => x"78",
          2630 => x"3f",
          2631 => x"08",
          2632 => x"84",
          2633 => x"38",
          2634 => x"70",
          2635 => x"73",
          2636 => x"58",
          2637 => x"8b",
          2638 => x"bf",
          2639 => x"ff",
          2640 => x"53",
          2641 => x"34",
          2642 => x"08",
          2643 => x"e5",
          2644 => x"81",
          2645 => x"2e",
          2646 => x"70",
          2647 => x"57",
          2648 => x"9e",
          2649 => x"2e",
          2650 => x"d3",
          2651 => x"df",
          2652 => x"72",
          2653 => x"81",
          2654 => x"76",
          2655 => x"2e",
          2656 => x"52",
          2657 => x"fc",
          2658 => x"84",
          2659 => x"d3",
          2660 => x"38",
          2661 => x"fe",
          2662 => x"39",
          2663 => x"16",
          2664 => x"d3",
          2665 => x"3d",
          2666 => x"3d",
          2667 => x"08",
          2668 => x"52",
          2669 => x"c5",
          2670 => x"84",
          2671 => x"d3",
          2672 => x"38",
          2673 => x"52",
          2674 => x"de",
          2675 => x"84",
          2676 => x"d3",
          2677 => x"38",
          2678 => x"d3",
          2679 => x"9c",
          2680 => x"ea",
          2681 => x"53",
          2682 => x"9c",
          2683 => x"ea",
          2684 => x"0b",
          2685 => x"74",
          2686 => x"0c",
          2687 => x"04",
          2688 => x"75",
          2689 => x"12",
          2690 => x"53",
          2691 => x"9a",
          2692 => x"84",
          2693 => x"9c",
          2694 => x"e5",
          2695 => x"0b",
          2696 => x"85",
          2697 => x"fa",
          2698 => x"7a",
          2699 => x"0b",
          2700 => x"98",
          2701 => x"2e",
          2702 => x"80",
          2703 => x"55",
          2704 => x"17",
          2705 => x"33",
          2706 => x"51",
          2707 => x"2e",
          2708 => x"85",
          2709 => x"06",
          2710 => x"e5",
          2711 => x"2e",
          2712 => x"8b",
          2713 => x"70",
          2714 => x"34",
          2715 => x"71",
          2716 => x"05",
          2717 => x"15",
          2718 => x"27",
          2719 => x"15",
          2720 => x"80",
          2721 => x"34",
          2722 => x"52",
          2723 => x"88",
          2724 => x"17",
          2725 => x"52",
          2726 => x"3f",
          2727 => x"08",
          2728 => x"12",
          2729 => x"3f",
          2730 => x"08",
          2731 => x"98",
          2732 => x"da",
          2733 => x"84",
          2734 => x"23",
          2735 => x"04",
          2736 => x"7f",
          2737 => x"5b",
          2738 => x"33",
          2739 => x"73",
          2740 => x"38",
          2741 => x"80",
          2742 => x"38",
          2743 => x"8c",
          2744 => x"08",
          2745 => x"aa",
          2746 => x"41",
          2747 => x"33",
          2748 => x"73",
          2749 => x"81",
          2750 => x"81",
          2751 => x"dc",
          2752 => x"70",
          2753 => x"07",
          2754 => x"73",
          2755 => x"88",
          2756 => x"70",
          2757 => x"73",
          2758 => x"38",
          2759 => x"ab",
          2760 => x"52",
          2761 => x"91",
          2762 => x"84",
          2763 => x"98",
          2764 => x"61",
          2765 => x"5a",
          2766 => x"a0",
          2767 => x"e7",
          2768 => x"70",
          2769 => x"79",
          2770 => x"73",
          2771 => x"81",
          2772 => x"38",
          2773 => x"33",
          2774 => x"ae",
          2775 => x"70",
          2776 => x"82",
          2777 => x"51",
          2778 => x"54",
          2779 => x"79",
          2780 => x"74",
          2781 => x"57",
          2782 => x"af",
          2783 => x"70",
          2784 => x"51",
          2785 => x"dc",
          2786 => x"73",
          2787 => x"38",
          2788 => x"82",
          2789 => x"19",
          2790 => x"54",
          2791 => x"82",
          2792 => x"54",
          2793 => x"78",
          2794 => x"81",
          2795 => x"54",
          2796 => x"81",
          2797 => x"af",
          2798 => x"77",
          2799 => x"70",
          2800 => x"25",
          2801 => x"07",
          2802 => x"51",
          2803 => x"2e",
          2804 => x"39",
          2805 => x"80",
          2806 => x"33",
          2807 => x"73",
          2808 => x"81",
          2809 => x"81",
          2810 => x"dc",
          2811 => x"70",
          2812 => x"07",
          2813 => x"73",
          2814 => x"b5",
          2815 => x"2e",
          2816 => x"83",
          2817 => x"76",
          2818 => x"07",
          2819 => x"2e",
          2820 => x"8b",
          2821 => x"77",
          2822 => x"30",
          2823 => x"71",
          2824 => x"53",
          2825 => x"55",
          2826 => x"38",
          2827 => x"5c",
          2828 => x"75",
          2829 => x"73",
          2830 => x"38",
          2831 => x"06",
          2832 => x"11",
          2833 => x"75",
          2834 => x"3f",
          2835 => x"08",
          2836 => x"38",
          2837 => x"33",
          2838 => x"54",
          2839 => x"e6",
          2840 => x"d3",
          2841 => x"2e",
          2842 => x"ff",
          2843 => x"74",
          2844 => x"38",
          2845 => x"75",
          2846 => x"17",
          2847 => x"57",
          2848 => x"a7",
          2849 => x"81",
          2850 => x"e5",
          2851 => x"d3",
          2852 => x"38",
          2853 => x"54",
          2854 => x"89",
          2855 => x"70",
          2856 => x"57",
          2857 => x"54",
          2858 => x"81",
          2859 => x"f7",
          2860 => x"7e",
          2861 => x"2e",
          2862 => x"33",
          2863 => x"e5",
          2864 => x"06",
          2865 => x"7a",
          2866 => x"a0",
          2867 => x"38",
          2868 => x"55",
          2869 => x"84",
          2870 => x"39",
          2871 => x"8b",
          2872 => x"7b",
          2873 => x"7a",
          2874 => x"3f",
          2875 => x"08",
          2876 => x"84",
          2877 => x"38",
          2878 => x"52",
          2879 => x"aa",
          2880 => x"84",
          2881 => x"d3",
          2882 => x"c2",
          2883 => x"08",
          2884 => x"55",
          2885 => x"ff",
          2886 => x"15",
          2887 => x"54",
          2888 => x"34",
          2889 => x"70",
          2890 => x"81",
          2891 => x"58",
          2892 => x"8b",
          2893 => x"74",
          2894 => x"3f",
          2895 => x"08",
          2896 => x"38",
          2897 => x"51",
          2898 => x"ff",
          2899 => x"ab",
          2900 => x"55",
          2901 => x"bb",
          2902 => x"2e",
          2903 => x"80",
          2904 => x"85",
          2905 => x"06",
          2906 => x"58",
          2907 => x"80",
          2908 => x"75",
          2909 => x"73",
          2910 => x"b5",
          2911 => x"0b",
          2912 => x"80",
          2913 => x"39",
          2914 => x"54",
          2915 => x"85",
          2916 => x"75",
          2917 => x"81",
          2918 => x"73",
          2919 => x"1b",
          2920 => x"2a",
          2921 => x"51",
          2922 => x"80",
          2923 => x"90",
          2924 => x"ff",
          2925 => x"05",
          2926 => x"f5",
          2927 => x"d3",
          2928 => x"1c",
          2929 => x"39",
          2930 => x"84",
          2931 => x"0d",
          2932 => x"0d",
          2933 => x"7b",
          2934 => x"73",
          2935 => x"55",
          2936 => x"2e",
          2937 => x"75",
          2938 => x"57",
          2939 => x"26",
          2940 => x"ba",
          2941 => x"70",
          2942 => x"ba",
          2943 => x"06",
          2944 => x"73",
          2945 => x"70",
          2946 => x"51",
          2947 => x"89",
          2948 => x"82",
          2949 => x"ff",
          2950 => x"56",
          2951 => x"2e",
          2952 => x"80",
          2953 => x"e8",
          2954 => x"08",
          2955 => x"76",
          2956 => x"58",
          2957 => x"81",
          2958 => x"ff",
          2959 => x"53",
          2960 => x"26",
          2961 => x"13",
          2962 => x"06",
          2963 => x"9f",
          2964 => x"99",
          2965 => x"e0",
          2966 => x"ff",
          2967 => x"72",
          2968 => x"2a",
          2969 => x"72",
          2970 => x"06",
          2971 => x"ff",
          2972 => x"30",
          2973 => x"70",
          2974 => x"07",
          2975 => x"9f",
          2976 => x"54",
          2977 => x"80",
          2978 => x"81",
          2979 => x"59",
          2980 => x"25",
          2981 => x"8b",
          2982 => x"24",
          2983 => x"76",
          2984 => x"78",
          2985 => x"81",
          2986 => x"51",
          2987 => x"84",
          2988 => x"0d",
          2989 => x"0d",
          2990 => x"0b",
          2991 => x"ff",
          2992 => x"0c",
          2993 => x"51",
          2994 => x"84",
          2995 => x"84",
          2996 => x"38",
          2997 => x"51",
          2998 => x"81",
          2999 => x"83",
          3000 => x"54",
          3001 => x"82",
          3002 => x"09",
          3003 => x"e3",
          3004 => x"b4",
          3005 => x"57",
          3006 => x"2e",
          3007 => x"83",
          3008 => x"74",
          3009 => x"70",
          3010 => x"25",
          3011 => x"51",
          3012 => x"38",
          3013 => x"2e",
          3014 => x"b5",
          3015 => x"81",
          3016 => x"80",
          3017 => x"e0",
          3018 => x"d3",
          3019 => x"81",
          3020 => x"80",
          3021 => x"85",
          3022 => x"ac",
          3023 => x"16",
          3024 => x"3f",
          3025 => x"08",
          3026 => x"84",
          3027 => x"83",
          3028 => x"74",
          3029 => x"0c",
          3030 => x"04",
          3031 => x"61",
          3032 => x"80",
          3033 => x"58",
          3034 => x"0c",
          3035 => x"e1",
          3036 => x"84",
          3037 => x"56",
          3038 => x"d3",
          3039 => x"86",
          3040 => x"d3",
          3041 => x"29",
          3042 => x"05",
          3043 => x"53",
          3044 => x"80",
          3045 => x"38",
          3046 => x"76",
          3047 => x"74",
          3048 => x"72",
          3049 => x"38",
          3050 => x"51",
          3051 => x"81",
          3052 => x"81",
          3053 => x"81",
          3054 => x"72",
          3055 => x"80",
          3056 => x"38",
          3057 => x"70",
          3058 => x"53",
          3059 => x"86",
          3060 => x"a7",
          3061 => x"34",
          3062 => x"34",
          3063 => x"14",
          3064 => x"b2",
          3065 => x"84",
          3066 => x"06",
          3067 => x"54",
          3068 => x"72",
          3069 => x"76",
          3070 => x"38",
          3071 => x"70",
          3072 => x"53",
          3073 => x"85",
          3074 => x"70",
          3075 => x"5b",
          3076 => x"81",
          3077 => x"81",
          3078 => x"76",
          3079 => x"81",
          3080 => x"38",
          3081 => x"56",
          3082 => x"83",
          3083 => x"70",
          3084 => x"80",
          3085 => x"83",
          3086 => x"dc",
          3087 => x"d3",
          3088 => x"76",
          3089 => x"05",
          3090 => x"16",
          3091 => x"56",
          3092 => x"d7",
          3093 => x"8d",
          3094 => x"72",
          3095 => x"54",
          3096 => x"57",
          3097 => x"95",
          3098 => x"73",
          3099 => x"3f",
          3100 => x"08",
          3101 => x"57",
          3102 => x"89",
          3103 => x"56",
          3104 => x"d7",
          3105 => x"76",
          3106 => x"f1",
          3107 => x"76",
          3108 => x"e9",
          3109 => x"51",
          3110 => x"81",
          3111 => x"83",
          3112 => x"53",
          3113 => x"2e",
          3114 => x"84",
          3115 => x"ca",
          3116 => x"da",
          3117 => x"84",
          3118 => x"ff",
          3119 => x"8d",
          3120 => x"14",
          3121 => x"3f",
          3122 => x"08",
          3123 => x"15",
          3124 => x"14",
          3125 => x"34",
          3126 => x"33",
          3127 => x"81",
          3128 => x"54",
          3129 => x"72",
          3130 => x"91",
          3131 => x"ff",
          3132 => x"29",
          3133 => x"33",
          3134 => x"72",
          3135 => x"72",
          3136 => x"38",
          3137 => x"06",
          3138 => x"2e",
          3139 => x"56",
          3140 => x"80",
          3141 => x"da",
          3142 => x"d3",
          3143 => x"81",
          3144 => x"88",
          3145 => x"8f",
          3146 => x"56",
          3147 => x"38",
          3148 => x"51",
          3149 => x"81",
          3150 => x"83",
          3151 => x"55",
          3152 => x"80",
          3153 => x"da",
          3154 => x"d3",
          3155 => x"80",
          3156 => x"da",
          3157 => x"d3",
          3158 => x"ff",
          3159 => x"8d",
          3160 => x"2e",
          3161 => x"88",
          3162 => x"14",
          3163 => x"05",
          3164 => x"75",
          3165 => x"38",
          3166 => x"52",
          3167 => x"51",
          3168 => x"3f",
          3169 => x"08",
          3170 => x"84",
          3171 => x"82",
          3172 => x"d3",
          3173 => x"ff",
          3174 => x"26",
          3175 => x"57",
          3176 => x"f5",
          3177 => x"82",
          3178 => x"f5",
          3179 => x"81",
          3180 => x"8d",
          3181 => x"2e",
          3182 => x"82",
          3183 => x"16",
          3184 => x"16",
          3185 => x"70",
          3186 => x"7a",
          3187 => x"0c",
          3188 => x"83",
          3189 => x"06",
          3190 => x"de",
          3191 => x"ae",
          3192 => x"84",
          3193 => x"ff",
          3194 => x"56",
          3195 => x"38",
          3196 => x"38",
          3197 => x"51",
          3198 => x"81",
          3199 => x"a8",
          3200 => x"82",
          3201 => x"39",
          3202 => x"80",
          3203 => x"38",
          3204 => x"15",
          3205 => x"53",
          3206 => x"8d",
          3207 => x"15",
          3208 => x"76",
          3209 => x"51",
          3210 => x"13",
          3211 => x"8d",
          3212 => x"15",
          3213 => x"c5",
          3214 => x"90",
          3215 => x"0b",
          3216 => x"ff",
          3217 => x"15",
          3218 => x"2e",
          3219 => x"81",
          3220 => x"e4",
          3221 => x"b6",
          3222 => x"84",
          3223 => x"ff",
          3224 => x"81",
          3225 => x"06",
          3226 => x"81",
          3227 => x"51",
          3228 => x"81",
          3229 => x"80",
          3230 => x"d3",
          3231 => x"15",
          3232 => x"14",
          3233 => x"3f",
          3234 => x"08",
          3235 => x"06",
          3236 => x"d4",
          3237 => x"81",
          3238 => x"38",
          3239 => x"d8",
          3240 => x"d3",
          3241 => x"8b",
          3242 => x"2e",
          3243 => x"b3",
          3244 => x"14",
          3245 => x"3f",
          3246 => x"08",
          3247 => x"e4",
          3248 => x"81",
          3249 => x"84",
          3250 => x"d7",
          3251 => x"d3",
          3252 => x"15",
          3253 => x"14",
          3254 => x"3f",
          3255 => x"08",
          3256 => x"76",
          3257 => x"d3",
          3258 => x"05",
          3259 => x"d3",
          3260 => x"86",
          3261 => x"0b",
          3262 => x"80",
          3263 => x"d3",
          3264 => x"3d",
          3265 => x"3d",
          3266 => x"89",
          3267 => x"2e",
          3268 => x"08",
          3269 => x"2e",
          3270 => x"33",
          3271 => x"2e",
          3272 => x"13",
          3273 => x"22",
          3274 => x"76",
          3275 => x"06",
          3276 => x"13",
          3277 => x"c0",
          3278 => x"84",
          3279 => x"52",
          3280 => x"71",
          3281 => x"55",
          3282 => x"53",
          3283 => x"0c",
          3284 => x"d3",
          3285 => x"3d",
          3286 => x"3d",
          3287 => x"05",
          3288 => x"89",
          3289 => x"52",
          3290 => x"3f",
          3291 => x"0b",
          3292 => x"08",
          3293 => x"81",
          3294 => x"84",
          3295 => x"a0",
          3296 => x"55",
          3297 => x"2e",
          3298 => x"74",
          3299 => x"73",
          3300 => x"38",
          3301 => x"78",
          3302 => x"54",
          3303 => x"92",
          3304 => x"89",
          3305 => x"84",
          3306 => x"b0",
          3307 => x"84",
          3308 => x"81",
          3309 => x"88",
          3310 => x"eb",
          3311 => x"02",
          3312 => x"e7",
          3313 => x"59",
          3314 => x"80",
          3315 => x"38",
          3316 => x"70",
          3317 => x"d0",
          3318 => x"3d",
          3319 => x"58",
          3320 => x"81",
          3321 => x"55",
          3322 => x"08",
          3323 => x"7a",
          3324 => x"8c",
          3325 => x"56",
          3326 => x"81",
          3327 => x"55",
          3328 => x"08",
          3329 => x"80",
          3330 => x"70",
          3331 => x"57",
          3332 => x"83",
          3333 => x"77",
          3334 => x"73",
          3335 => x"ab",
          3336 => x"2e",
          3337 => x"84",
          3338 => x"06",
          3339 => x"51",
          3340 => x"81",
          3341 => x"55",
          3342 => x"b2",
          3343 => x"06",
          3344 => x"b8",
          3345 => x"2a",
          3346 => x"51",
          3347 => x"2e",
          3348 => x"55",
          3349 => x"77",
          3350 => x"74",
          3351 => x"77",
          3352 => x"81",
          3353 => x"73",
          3354 => x"af",
          3355 => x"7a",
          3356 => x"3f",
          3357 => x"08",
          3358 => x"b2",
          3359 => x"8e",
          3360 => x"ea",
          3361 => x"a0",
          3362 => x"34",
          3363 => x"52",
          3364 => x"bd",
          3365 => x"62",
          3366 => x"d4",
          3367 => x"54",
          3368 => x"15",
          3369 => x"2e",
          3370 => x"7a",
          3371 => x"51",
          3372 => x"75",
          3373 => x"d4",
          3374 => x"be",
          3375 => x"84",
          3376 => x"d3",
          3377 => x"ca",
          3378 => x"74",
          3379 => x"02",
          3380 => x"70",
          3381 => x"81",
          3382 => x"56",
          3383 => x"86",
          3384 => x"82",
          3385 => x"81",
          3386 => x"06",
          3387 => x"80",
          3388 => x"75",
          3389 => x"73",
          3390 => x"38",
          3391 => x"92",
          3392 => x"7a",
          3393 => x"3f",
          3394 => x"08",
          3395 => x"8c",
          3396 => x"55",
          3397 => x"08",
          3398 => x"77",
          3399 => x"81",
          3400 => x"73",
          3401 => x"38",
          3402 => x"07",
          3403 => x"11",
          3404 => x"0c",
          3405 => x"0c",
          3406 => x"52",
          3407 => x"3f",
          3408 => x"08",
          3409 => x"08",
          3410 => x"63",
          3411 => x"5a",
          3412 => x"81",
          3413 => x"81",
          3414 => x"8c",
          3415 => x"7a",
          3416 => x"17",
          3417 => x"23",
          3418 => x"34",
          3419 => x"1a",
          3420 => x"9c",
          3421 => x"0b",
          3422 => x"77",
          3423 => x"81",
          3424 => x"73",
          3425 => x"8d",
          3426 => x"84",
          3427 => x"81",
          3428 => x"d3",
          3429 => x"1a",
          3430 => x"22",
          3431 => x"7b",
          3432 => x"a8",
          3433 => x"78",
          3434 => x"3f",
          3435 => x"08",
          3436 => x"84",
          3437 => x"83",
          3438 => x"81",
          3439 => x"ff",
          3440 => x"06",
          3441 => x"55",
          3442 => x"56",
          3443 => x"76",
          3444 => x"51",
          3445 => x"27",
          3446 => x"70",
          3447 => x"5a",
          3448 => x"76",
          3449 => x"74",
          3450 => x"83",
          3451 => x"73",
          3452 => x"38",
          3453 => x"51",
          3454 => x"81",
          3455 => x"85",
          3456 => x"8e",
          3457 => x"2a",
          3458 => x"08",
          3459 => x"0c",
          3460 => x"79",
          3461 => x"73",
          3462 => x"0c",
          3463 => x"04",
          3464 => x"60",
          3465 => x"40",
          3466 => x"80",
          3467 => x"3d",
          3468 => x"78",
          3469 => x"3f",
          3470 => x"08",
          3471 => x"84",
          3472 => x"91",
          3473 => x"74",
          3474 => x"38",
          3475 => x"c4",
          3476 => x"33",
          3477 => x"87",
          3478 => x"2e",
          3479 => x"95",
          3480 => x"91",
          3481 => x"56",
          3482 => x"81",
          3483 => x"34",
          3484 => x"a0",
          3485 => x"08",
          3486 => x"31",
          3487 => x"27",
          3488 => x"5c",
          3489 => x"82",
          3490 => x"19",
          3491 => x"ff",
          3492 => x"74",
          3493 => x"7e",
          3494 => x"ff",
          3495 => x"2a",
          3496 => x"79",
          3497 => x"87",
          3498 => x"08",
          3499 => x"98",
          3500 => x"78",
          3501 => x"3f",
          3502 => x"08",
          3503 => x"27",
          3504 => x"74",
          3505 => x"a3",
          3506 => x"1a",
          3507 => x"08",
          3508 => x"d4",
          3509 => x"d3",
          3510 => x"2e",
          3511 => x"81",
          3512 => x"1a",
          3513 => x"59",
          3514 => x"2e",
          3515 => x"77",
          3516 => x"11",
          3517 => x"55",
          3518 => x"85",
          3519 => x"31",
          3520 => x"76",
          3521 => x"81",
          3522 => x"ca",
          3523 => x"d3",
          3524 => x"d7",
          3525 => x"11",
          3526 => x"74",
          3527 => x"38",
          3528 => x"77",
          3529 => x"78",
          3530 => x"84",
          3531 => x"16",
          3532 => x"08",
          3533 => x"2b",
          3534 => x"cf",
          3535 => x"89",
          3536 => x"39",
          3537 => x"0c",
          3538 => x"83",
          3539 => x"80",
          3540 => x"55",
          3541 => x"83",
          3542 => x"9c",
          3543 => x"7e",
          3544 => x"3f",
          3545 => x"08",
          3546 => x"75",
          3547 => x"08",
          3548 => x"1f",
          3549 => x"7c",
          3550 => x"3f",
          3551 => x"7e",
          3552 => x"0c",
          3553 => x"1b",
          3554 => x"1c",
          3555 => x"fd",
          3556 => x"56",
          3557 => x"84",
          3558 => x"0d",
          3559 => x"0d",
          3560 => x"64",
          3561 => x"58",
          3562 => x"90",
          3563 => x"52",
          3564 => x"d2",
          3565 => x"84",
          3566 => x"d3",
          3567 => x"38",
          3568 => x"55",
          3569 => x"86",
          3570 => x"83",
          3571 => x"18",
          3572 => x"2a",
          3573 => x"51",
          3574 => x"56",
          3575 => x"83",
          3576 => x"39",
          3577 => x"19",
          3578 => x"83",
          3579 => x"0b",
          3580 => x"81",
          3581 => x"39",
          3582 => x"7c",
          3583 => x"74",
          3584 => x"38",
          3585 => x"7b",
          3586 => x"ec",
          3587 => x"08",
          3588 => x"06",
          3589 => x"81",
          3590 => x"8a",
          3591 => x"05",
          3592 => x"06",
          3593 => x"bf",
          3594 => x"38",
          3595 => x"55",
          3596 => x"7a",
          3597 => x"98",
          3598 => x"77",
          3599 => x"3f",
          3600 => x"08",
          3601 => x"84",
          3602 => x"82",
          3603 => x"81",
          3604 => x"38",
          3605 => x"ff",
          3606 => x"98",
          3607 => x"18",
          3608 => x"74",
          3609 => x"7e",
          3610 => x"08",
          3611 => x"2e",
          3612 => x"8d",
          3613 => x"ce",
          3614 => x"d3",
          3615 => x"ee",
          3616 => x"08",
          3617 => x"d1",
          3618 => x"d3",
          3619 => x"2e",
          3620 => x"81",
          3621 => x"1b",
          3622 => x"5a",
          3623 => x"2e",
          3624 => x"78",
          3625 => x"11",
          3626 => x"55",
          3627 => x"85",
          3628 => x"31",
          3629 => x"76",
          3630 => x"81",
          3631 => x"c8",
          3632 => x"d3",
          3633 => x"a6",
          3634 => x"11",
          3635 => x"56",
          3636 => x"27",
          3637 => x"80",
          3638 => x"08",
          3639 => x"2b",
          3640 => x"b4",
          3641 => x"b5",
          3642 => x"80",
          3643 => x"34",
          3644 => x"56",
          3645 => x"8c",
          3646 => x"19",
          3647 => x"38",
          3648 => x"b6",
          3649 => x"84",
          3650 => x"38",
          3651 => x"12",
          3652 => x"9c",
          3653 => x"18",
          3654 => x"06",
          3655 => x"31",
          3656 => x"76",
          3657 => x"7b",
          3658 => x"08",
          3659 => x"cd",
          3660 => x"d3",
          3661 => x"b6",
          3662 => x"7c",
          3663 => x"08",
          3664 => x"1f",
          3665 => x"cb",
          3666 => x"55",
          3667 => x"16",
          3668 => x"31",
          3669 => x"7f",
          3670 => x"94",
          3671 => x"70",
          3672 => x"8c",
          3673 => x"58",
          3674 => x"76",
          3675 => x"75",
          3676 => x"19",
          3677 => x"39",
          3678 => x"80",
          3679 => x"74",
          3680 => x"80",
          3681 => x"d3",
          3682 => x"3d",
          3683 => x"3d",
          3684 => x"3d",
          3685 => x"70",
          3686 => x"ea",
          3687 => x"84",
          3688 => x"d3",
          3689 => x"fb",
          3690 => x"33",
          3691 => x"70",
          3692 => x"55",
          3693 => x"2e",
          3694 => x"a0",
          3695 => x"78",
          3696 => x"3f",
          3697 => x"08",
          3698 => x"84",
          3699 => x"38",
          3700 => x"8b",
          3701 => x"07",
          3702 => x"8b",
          3703 => x"16",
          3704 => x"52",
          3705 => x"dd",
          3706 => x"16",
          3707 => x"15",
          3708 => x"3f",
          3709 => x"0a",
          3710 => x"51",
          3711 => x"76",
          3712 => x"51",
          3713 => x"78",
          3714 => x"83",
          3715 => x"51",
          3716 => x"81",
          3717 => x"90",
          3718 => x"bf",
          3719 => x"73",
          3720 => x"76",
          3721 => x"0c",
          3722 => x"04",
          3723 => x"76",
          3724 => x"fe",
          3725 => x"d3",
          3726 => x"81",
          3727 => x"9c",
          3728 => x"fc",
          3729 => x"51",
          3730 => x"81",
          3731 => x"53",
          3732 => x"08",
          3733 => x"d3",
          3734 => x"0c",
          3735 => x"84",
          3736 => x"0d",
          3737 => x"0d",
          3738 => x"e6",
          3739 => x"52",
          3740 => x"d3",
          3741 => x"8b",
          3742 => x"84",
          3743 => x"b4",
          3744 => x"71",
          3745 => x"0c",
          3746 => x"04",
          3747 => x"80",
          3748 => x"d0",
          3749 => x"3d",
          3750 => x"3f",
          3751 => x"08",
          3752 => x"84",
          3753 => x"38",
          3754 => x"52",
          3755 => x"05",
          3756 => x"3f",
          3757 => x"08",
          3758 => x"84",
          3759 => x"02",
          3760 => x"33",
          3761 => x"55",
          3762 => x"25",
          3763 => x"7a",
          3764 => x"54",
          3765 => x"a2",
          3766 => x"84",
          3767 => x"06",
          3768 => x"73",
          3769 => x"38",
          3770 => x"70",
          3771 => x"a8",
          3772 => x"84",
          3773 => x"0c",
          3774 => x"d3",
          3775 => x"2e",
          3776 => x"83",
          3777 => x"74",
          3778 => x"0c",
          3779 => x"04",
          3780 => x"6f",
          3781 => x"80",
          3782 => x"53",
          3783 => x"b8",
          3784 => x"3d",
          3785 => x"3f",
          3786 => x"08",
          3787 => x"84",
          3788 => x"38",
          3789 => x"7c",
          3790 => x"47",
          3791 => x"54",
          3792 => x"81",
          3793 => x"52",
          3794 => x"52",
          3795 => x"3f",
          3796 => x"08",
          3797 => x"84",
          3798 => x"38",
          3799 => x"51",
          3800 => x"81",
          3801 => x"57",
          3802 => x"08",
          3803 => x"69",
          3804 => x"da",
          3805 => x"d3",
          3806 => x"76",
          3807 => x"d5",
          3808 => x"d3",
          3809 => x"81",
          3810 => x"82",
          3811 => x"52",
          3812 => x"eb",
          3813 => x"84",
          3814 => x"d3",
          3815 => x"38",
          3816 => x"51",
          3817 => x"73",
          3818 => x"08",
          3819 => x"76",
          3820 => x"d6",
          3821 => x"d3",
          3822 => x"81",
          3823 => x"80",
          3824 => x"76",
          3825 => x"81",
          3826 => x"82",
          3827 => x"39",
          3828 => x"38",
          3829 => x"bc",
          3830 => x"51",
          3831 => x"76",
          3832 => x"11",
          3833 => x"51",
          3834 => x"73",
          3835 => x"38",
          3836 => x"55",
          3837 => x"16",
          3838 => x"56",
          3839 => x"38",
          3840 => x"73",
          3841 => x"90",
          3842 => x"2e",
          3843 => x"16",
          3844 => x"ff",
          3845 => x"ff",
          3846 => x"58",
          3847 => x"74",
          3848 => x"75",
          3849 => x"18",
          3850 => x"58",
          3851 => x"fe",
          3852 => x"7b",
          3853 => x"06",
          3854 => x"18",
          3855 => x"58",
          3856 => x"80",
          3857 => x"b4",
          3858 => x"29",
          3859 => x"05",
          3860 => x"33",
          3861 => x"56",
          3862 => x"2e",
          3863 => x"16",
          3864 => x"33",
          3865 => x"73",
          3866 => x"16",
          3867 => x"26",
          3868 => x"55",
          3869 => x"91",
          3870 => x"54",
          3871 => x"70",
          3872 => x"34",
          3873 => x"ec",
          3874 => x"70",
          3875 => x"34",
          3876 => x"09",
          3877 => x"38",
          3878 => x"39",
          3879 => x"19",
          3880 => x"33",
          3881 => x"05",
          3882 => x"78",
          3883 => x"80",
          3884 => x"81",
          3885 => x"9e",
          3886 => x"f7",
          3887 => x"7d",
          3888 => x"05",
          3889 => x"57",
          3890 => x"3f",
          3891 => x"08",
          3892 => x"84",
          3893 => x"38",
          3894 => x"53",
          3895 => x"38",
          3896 => x"54",
          3897 => x"92",
          3898 => x"33",
          3899 => x"70",
          3900 => x"54",
          3901 => x"38",
          3902 => x"15",
          3903 => x"70",
          3904 => x"58",
          3905 => x"82",
          3906 => x"8a",
          3907 => x"89",
          3908 => x"53",
          3909 => x"b7",
          3910 => x"ff",
          3911 => x"98",
          3912 => x"d3",
          3913 => x"15",
          3914 => x"53",
          3915 => x"98",
          3916 => x"d3",
          3917 => x"26",
          3918 => x"30",
          3919 => x"70",
          3920 => x"77",
          3921 => x"18",
          3922 => x"51",
          3923 => x"88",
          3924 => x"73",
          3925 => x"52",
          3926 => x"ca",
          3927 => x"84",
          3928 => x"d3",
          3929 => x"2e",
          3930 => x"81",
          3931 => x"ff",
          3932 => x"38",
          3933 => x"08",
          3934 => x"73",
          3935 => x"73",
          3936 => x"9c",
          3937 => x"27",
          3938 => x"75",
          3939 => x"16",
          3940 => x"17",
          3941 => x"33",
          3942 => x"70",
          3943 => x"55",
          3944 => x"80",
          3945 => x"73",
          3946 => x"cc",
          3947 => x"d3",
          3948 => x"81",
          3949 => x"94",
          3950 => x"84",
          3951 => x"39",
          3952 => x"51",
          3953 => x"81",
          3954 => x"54",
          3955 => x"be",
          3956 => x"27",
          3957 => x"53",
          3958 => x"08",
          3959 => x"73",
          3960 => x"ff",
          3961 => x"15",
          3962 => x"16",
          3963 => x"ff",
          3964 => x"80",
          3965 => x"73",
          3966 => x"c6",
          3967 => x"d3",
          3968 => x"38",
          3969 => x"16",
          3970 => x"80",
          3971 => x"0b",
          3972 => x"81",
          3973 => x"75",
          3974 => x"d3",
          3975 => x"58",
          3976 => x"54",
          3977 => x"74",
          3978 => x"73",
          3979 => x"90",
          3980 => x"c0",
          3981 => x"90",
          3982 => x"83",
          3983 => x"72",
          3984 => x"38",
          3985 => x"08",
          3986 => x"77",
          3987 => x"80",
          3988 => x"d3",
          3989 => x"3d",
          3990 => x"3d",
          3991 => x"89",
          3992 => x"2e",
          3993 => x"80",
          3994 => x"fc",
          3995 => x"3d",
          3996 => x"e1",
          3997 => x"d3",
          3998 => x"81",
          3999 => x"80",
          4000 => x"76",
          4001 => x"75",
          4002 => x"3f",
          4003 => x"08",
          4004 => x"84",
          4005 => x"38",
          4006 => x"70",
          4007 => x"57",
          4008 => x"a2",
          4009 => x"33",
          4010 => x"70",
          4011 => x"55",
          4012 => x"2e",
          4013 => x"16",
          4014 => x"51",
          4015 => x"81",
          4016 => x"88",
          4017 => x"54",
          4018 => x"84",
          4019 => x"52",
          4020 => x"e5",
          4021 => x"84",
          4022 => x"84",
          4023 => x"06",
          4024 => x"55",
          4025 => x"80",
          4026 => x"80",
          4027 => x"54",
          4028 => x"84",
          4029 => x"0d",
          4030 => x"0d",
          4031 => x"fc",
          4032 => x"52",
          4033 => x"3f",
          4034 => x"08",
          4035 => x"d3",
          4036 => x"0c",
          4037 => x"04",
          4038 => x"77",
          4039 => x"fc",
          4040 => x"53",
          4041 => x"de",
          4042 => x"84",
          4043 => x"d3",
          4044 => x"df",
          4045 => x"38",
          4046 => x"08",
          4047 => x"cd",
          4048 => x"d3",
          4049 => x"80",
          4050 => x"d3",
          4051 => x"73",
          4052 => x"3f",
          4053 => x"08",
          4054 => x"84",
          4055 => x"09",
          4056 => x"38",
          4057 => x"39",
          4058 => x"08",
          4059 => x"52",
          4060 => x"b3",
          4061 => x"73",
          4062 => x"3f",
          4063 => x"08",
          4064 => x"30",
          4065 => x"9f",
          4066 => x"d3",
          4067 => x"51",
          4068 => x"72",
          4069 => x"0c",
          4070 => x"04",
          4071 => x"65",
          4072 => x"89",
          4073 => x"96",
          4074 => x"df",
          4075 => x"d3",
          4076 => x"81",
          4077 => x"b2",
          4078 => x"75",
          4079 => x"3f",
          4080 => x"08",
          4081 => x"84",
          4082 => x"02",
          4083 => x"33",
          4084 => x"55",
          4085 => x"25",
          4086 => x"55",
          4087 => x"80",
          4088 => x"76",
          4089 => x"d4",
          4090 => x"81",
          4091 => x"94",
          4092 => x"f0",
          4093 => x"65",
          4094 => x"53",
          4095 => x"05",
          4096 => x"51",
          4097 => x"81",
          4098 => x"5b",
          4099 => x"08",
          4100 => x"7c",
          4101 => x"08",
          4102 => x"fe",
          4103 => x"08",
          4104 => x"55",
          4105 => x"91",
          4106 => x"0c",
          4107 => x"81",
          4108 => x"39",
          4109 => x"c7",
          4110 => x"84",
          4111 => x"55",
          4112 => x"2e",
          4113 => x"bf",
          4114 => x"5f",
          4115 => x"92",
          4116 => x"51",
          4117 => x"81",
          4118 => x"ff",
          4119 => x"81",
          4120 => x"81",
          4121 => x"81",
          4122 => x"30",
          4123 => x"84",
          4124 => x"25",
          4125 => x"19",
          4126 => x"5a",
          4127 => x"08",
          4128 => x"38",
          4129 => x"a4",
          4130 => x"d3",
          4131 => x"58",
          4132 => x"77",
          4133 => x"7d",
          4134 => x"bf",
          4135 => x"d3",
          4136 => x"81",
          4137 => x"80",
          4138 => x"70",
          4139 => x"ff",
          4140 => x"56",
          4141 => x"2e",
          4142 => x"9e",
          4143 => x"51",
          4144 => x"3f",
          4145 => x"08",
          4146 => x"06",
          4147 => x"80",
          4148 => x"19",
          4149 => x"54",
          4150 => x"14",
          4151 => x"c5",
          4152 => x"84",
          4153 => x"06",
          4154 => x"80",
          4155 => x"19",
          4156 => x"54",
          4157 => x"06",
          4158 => x"79",
          4159 => x"78",
          4160 => x"79",
          4161 => x"84",
          4162 => x"07",
          4163 => x"84",
          4164 => x"81",
          4165 => x"92",
          4166 => x"f9",
          4167 => x"8a",
          4168 => x"53",
          4169 => x"e3",
          4170 => x"d3",
          4171 => x"81",
          4172 => x"81",
          4173 => x"17",
          4174 => x"81",
          4175 => x"17",
          4176 => x"2a",
          4177 => x"51",
          4178 => x"55",
          4179 => x"81",
          4180 => x"17",
          4181 => x"8c",
          4182 => x"81",
          4183 => x"9b",
          4184 => x"84",
          4185 => x"17",
          4186 => x"51",
          4187 => x"81",
          4188 => x"74",
          4189 => x"56",
          4190 => x"98",
          4191 => x"76",
          4192 => x"c6",
          4193 => x"84",
          4194 => x"09",
          4195 => x"38",
          4196 => x"d3",
          4197 => x"2e",
          4198 => x"85",
          4199 => x"a3",
          4200 => x"38",
          4201 => x"d3",
          4202 => x"15",
          4203 => x"38",
          4204 => x"53",
          4205 => x"08",
          4206 => x"c3",
          4207 => x"d3",
          4208 => x"94",
          4209 => x"18",
          4210 => x"33",
          4211 => x"54",
          4212 => x"34",
          4213 => x"85",
          4214 => x"18",
          4215 => x"74",
          4216 => x"0c",
          4217 => x"04",
          4218 => x"82",
          4219 => x"ff",
          4220 => x"a1",
          4221 => x"e4",
          4222 => x"84",
          4223 => x"d3",
          4224 => x"f5",
          4225 => x"a1",
          4226 => x"95",
          4227 => x"58",
          4228 => x"81",
          4229 => x"55",
          4230 => x"08",
          4231 => x"02",
          4232 => x"33",
          4233 => x"70",
          4234 => x"55",
          4235 => x"73",
          4236 => x"75",
          4237 => x"80",
          4238 => x"bd",
          4239 => x"d6",
          4240 => x"81",
          4241 => x"87",
          4242 => x"ad",
          4243 => x"78",
          4244 => x"3f",
          4245 => x"08",
          4246 => x"70",
          4247 => x"55",
          4248 => x"2e",
          4249 => x"78",
          4250 => x"84",
          4251 => x"08",
          4252 => x"38",
          4253 => x"d3",
          4254 => x"76",
          4255 => x"70",
          4256 => x"b5",
          4257 => x"84",
          4258 => x"d3",
          4259 => x"e9",
          4260 => x"84",
          4261 => x"51",
          4262 => x"81",
          4263 => x"55",
          4264 => x"08",
          4265 => x"55",
          4266 => x"81",
          4267 => x"84",
          4268 => x"81",
          4269 => x"80",
          4270 => x"51",
          4271 => x"81",
          4272 => x"81",
          4273 => x"30",
          4274 => x"84",
          4275 => x"25",
          4276 => x"75",
          4277 => x"38",
          4278 => x"8f",
          4279 => x"75",
          4280 => x"c1",
          4281 => x"d3",
          4282 => x"74",
          4283 => x"51",
          4284 => x"3f",
          4285 => x"08",
          4286 => x"d3",
          4287 => x"3d",
          4288 => x"3d",
          4289 => x"99",
          4290 => x"52",
          4291 => x"d8",
          4292 => x"d3",
          4293 => x"81",
          4294 => x"82",
          4295 => x"5e",
          4296 => x"3d",
          4297 => x"cf",
          4298 => x"d3",
          4299 => x"81",
          4300 => x"86",
          4301 => x"82",
          4302 => x"d3",
          4303 => x"2e",
          4304 => x"82",
          4305 => x"80",
          4306 => x"70",
          4307 => x"06",
          4308 => x"54",
          4309 => x"38",
          4310 => x"52",
          4311 => x"52",
          4312 => x"3f",
          4313 => x"08",
          4314 => x"81",
          4315 => x"83",
          4316 => x"81",
          4317 => x"81",
          4318 => x"06",
          4319 => x"54",
          4320 => x"08",
          4321 => x"81",
          4322 => x"81",
          4323 => x"39",
          4324 => x"38",
          4325 => x"08",
          4326 => x"c4",
          4327 => x"d3",
          4328 => x"81",
          4329 => x"81",
          4330 => x"53",
          4331 => x"19",
          4332 => x"8c",
          4333 => x"ae",
          4334 => x"34",
          4335 => x"0b",
          4336 => x"82",
          4337 => x"52",
          4338 => x"51",
          4339 => x"3f",
          4340 => x"b4",
          4341 => x"c9",
          4342 => x"53",
          4343 => x"53",
          4344 => x"51",
          4345 => x"3f",
          4346 => x"0b",
          4347 => x"34",
          4348 => x"80",
          4349 => x"51",
          4350 => x"78",
          4351 => x"83",
          4352 => x"51",
          4353 => x"81",
          4354 => x"54",
          4355 => x"08",
          4356 => x"88",
          4357 => x"64",
          4358 => x"ff",
          4359 => x"75",
          4360 => x"78",
          4361 => x"3f",
          4362 => x"0b",
          4363 => x"78",
          4364 => x"83",
          4365 => x"51",
          4366 => x"3f",
          4367 => x"08",
          4368 => x"80",
          4369 => x"76",
          4370 => x"ae",
          4371 => x"d3",
          4372 => x"3d",
          4373 => x"3d",
          4374 => x"84",
          4375 => x"f1",
          4376 => x"a8",
          4377 => x"05",
          4378 => x"51",
          4379 => x"81",
          4380 => x"55",
          4381 => x"08",
          4382 => x"78",
          4383 => x"08",
          4384 => x"70",
          4385 => x"b8",
          4386 => x"84",
          4387 => x"d3",
          4388 => x"b9",
          4389 => x"9b",
          4390 => x"a0",
          4391 => x"55",
          4392 => x"38",
          4393 => x"3d",
          4394 => x"3d",
          4395 => x"51",
          4396 => x"3f",
          4397 => x"52",
          4398 => x"52",
          4399 => x"dd",
          4400 => x"08",
          4401 => x"cb",
          4402 => x"d3",
          4403 => x"81",
          4404 => x"95",
          4405 => x"2e",
          4406 => x"88",
          4407 => x"3d",
          4408 => x"38",
          4409 => x"e5",
          4410 => x"84",
          4411 => x"09",
          4412 => x"b8",
          4413 => x"c9",
          4414 => x"d3",
          4415 => x"81",
          4416 => x"81",
          4417 => x"56",
          4418 => x"3d",
          4419 => x"52",
          4420 => x"ff",
          4421 => x"02",
          4422 => x"8b",
          4423 => x"16",
          4424 => x"2a",
          4425 => x"51",
          4426 => x"89",
          4427 => x"07",
          4428 => x"17",
          4429 => x"81",
          4430 => x"34",
          4431 => x"70",
          4432 => x"81",
          4433 => x"55",
          4434 => x"80",
          4435 => x"64",
          4436 => x"38",
          4437 => x"51",
          4438 => x"81",
          4439 => x"52",
          4440 => x"b7",
          4441 => x"55",
          4442 => x"08",
          4443 => x"dd",
          4444 => x"84",
          4445 => x"51",
          4446 => x"3f",
          4447 => x"08",
          4448 => x"11",
          4449 => x"81",
          4450 => x"80",
          4451 => x"16",
          4452 => x"ae",
          4453 => x"06",
          4454 => x"53",
          4455 => x"51",
          4456 => x"78",
          4457 => x"83",
          4458 => x"39",
          4459 => x"08",
          4460 => x"51",
          4461 => x"81",
          4462 => x"55",
          4463 => x"08",
          4464 => x"51",
          4465 => x"3f",
          4466 => x"08",
          4467 => x"d3",
          4468 => x"3d",
          4469 => x"3d",
          4470 => x"db",
          4471 => x"84",
          4472 => x"05",
          4473 => x"82",
          4474 => x"d0",
          4475 => x"3d",
          4476 => x"3f",
          4477 => x"08",
          4478 => x"84",
          4479 => x"38",
          4480 => x"52",
          4481 => x"05",
          4482 => x"3f",
          4483 => x"08",
          4484 => x"84",
          4485 => x"02",
          4486 => x"33",
          4487 => x"54",
          4488 => x"aa",
          4489 => x"06",
          4490 => x"8b",
          4491 => x"06",
          4492 => x"07",
          4493 => x"56",
          4494 => x"34",
          4495 => x"0b",
          4496 => x"78",
          4497 => x"a9",
          4498 => x"84",
          4499 => x"81",
          4500 => x"95",
          4501 => x"ef",
          4502 => x"56",
          4503 => x"3d",
          4504 => x"94",
          4505 => x"f4",
          4506 => x"84",
          4507 => x"d3",
          4508 => x"cb",
          4509 => x"63",
          4510 => x"d4",
          4511 => x"c0",
          4512 => x"84",
          4513 => x"d3",
          4514 => x"38",
          4515 => x"05",
          4516 => x"06",
          4517 => x"73",
          4518 => x"16",
          4519 => x"22",
          4520 => x"07",
          4521 => x"1f",
          4522 => x"c2",
          4523 => x"81",
          4524 => x"34",
          4525 => x"b3",
          4526 => x"d3",
          4527 => x"74",
          4528 => x"0c",
          4529 => x"04",
          4530 => x"69",
          4531 => x"80",
          4532 => x"d0",
          4533 => x"3d",
          4534 => x"3f",
          4535 => x"08",
          4536 => x"08",
          4537 => x"d3",
          4538 => x"80",
          4539 => x"57",
          4540 => x"81",
          4541 => x"70",
          4542 => x"55",
          4543 => x"80",
          4544 => x"5d",
          4545 => x"52",
          4546 => x"52",
          4547 => x"a9",
          4548 => x"84",
          4549 => x"d3",
          4550 => x"d1",
          4551 => x"73",
          4552 => x"3f",
          4553 => x"08",
          4554 => x"84",
          4555 => x"81",
          4556 => x"81",
          4557 => x"65",
          4558 => x"78",
          4559 => x"7b",
          4560 => x"55",
          4561 => x"34",
          4562 => x"8a",
          4563 => x"38",
          4564 => x"1a",
          4565 => x"34",
          4566 => x"9e",
          4567 => x"70",
          4568 => x"51",
          4569 => x"a0",
          4570 => x"8e",
          4571 => x"2e",
          4572 => x"86",
          4573 => x"34",
          4574 => x"30",
          4575 => x"80",
          4576 => x"7a",
          4577 => x"c1",
          4578 => x"2e",
          4579 => x"a0",
          4580 => x"51",
          4581 => x"3f",
          4582 => x"08",
          4583 => x"84",
          4584 => x"7b",
          4585 => x"55",
          4586 => x"73",
          4587 => x"38",
          4588 => x"73",
          4589 => x"38",
          4590 => x"15",
          4591 => x"ff",
          4592 => x"81",
          4593 => x"7b",
          4594 => x"d3",
          4595 => x"3d",
          4596 => x"3d",
          4597 => x"9c",
          4598 => x"05",
          4599 => x"51",
          4600 => x"81",
          4601 => x"81",
          4602 => x"56",
          4603 => x"84",
          4604 => x"38",
          4605 => x"52",
          4606 => x"52",
          4607 => x"c0",
          4608 => x"70",
          4609 => x"ff",
          4610 => x"55",
          4611 => x"27",
          4612 => x"78",
          4613 => x"ff",
          4614 => x"05",
          4615 => x"55",
          4616 => x"3f",
          4617 => x"08",
          4618 => x"38",
          4619 => x"70",
          4620 => x"ff",
          4621 => x"81",
          4622 => x"80",
          4623 => x"74",
          4624 => x"07",
          4625 => x"4e",
          4626 => x"81",
          4627 => x"55",
          4628 => x"70",
          4629 => x"06",
          4630 => x"99",
          4631 => x"e0",
          4632 => x"ff",
          4633 => x"54",
          4634 => x"27",
          4635 => x"c1",
          4636 => x"55",
          4637 => x"a3",
          4638 => x"81",
          4639 => x"ff",
          4640 => x"81",
          4641 => x"93",
          4642 => x"75",
          4643 => x"76",
          4644 => x"38",
          4645 => x"77",
          4646 => x"86",
          4647 => x"39",
          4648 => x"27",
          4649 => x"88",
          4650 => x"78",
          4651 => x"5a",
          4652 => x"57",
          4653 => x"81",
          4654 => x"81",
          4655 => x"33",
          4656 => x"06",
          4657 => x"57",
          4658 => x"fe",
          4659 => x"3d",
          4660 => x"55",
          4661 => x"2e",
          4662 => x"76",
          4663 => x"38",
          4664 => x"55",
          4665 => x"33",
          4666 => x"a0",
          4667 => x"06",
          4668 => x"17",
          4669 => x"38",
          4670 => x"43",
          4671 => x"3d",
          4672 => x"ff",
          4673 => x"81",
          4674 => x"54",
          4675 => x"08",
          4676 => x"81",
          4677 => x"ff",
          4678 => x"81",
          4679 => x"54",
          4680 => x"08",
          4681 => x"80",
          4682 => x"54",
          4683 => x"80",
          4684 => x"d3",
          4685 => x"2e",
          4686 => x"80",
          4687 => x"54",
          4688 => x"80",
          4689 => x"52",
          4690 => x"bd",
          4691 => x"d3",
          4692 => x"81",
          4693 => x"b1",
          4694 => x"81",
          4695 => x"52",
          4696 => x"ab",
          4697 => x"54",
          4698 => x"15",
          4699 => x"78",
          4700 => x"ff",
          4701 => x"79",
          4702 => x"83",
          4703 => x"51",
          4704 => x"3f",
          4705 => x"08",
          4706 => x"74",
          4707 => x"0c",
          4708 => x"04",
          4709 => x"60",
          4710 => x"05",
          4711 => x"33",
          4712 => x"05",
          4713 => x"40",
          4714 => x"da",
          4715 => x"84",
          4716 => x"d3",
          4717 => x"bd",
          4718 => x"33",
          4719 => x"b5",
          4720 => x"2e",
          4721 => x"1a",
          4722 => x"90",
          4723 => x"33",
          4724 => x"70",
          4725 => x"55",
          4726 => x"38",
          4727 => x"97",
          4728 => x"82",
          4729 => x"58",
          4730 => x"7e",
          4731 => x"70",
          4732 => x"55",
          4733 => x"56",
          4734 => x"fd",
          4735 => x"7d",
          4736 => x"70",
          4737 => x"2a",
          4738 => x"08",
          4739 => x"08",
          4740 => x"5d",
          4741 => x"77",
          4742 => x"98",
          4743 => x"26",
          4744 => x"57",
          4745 => x"59",
          4746 => x"52",
          4747 => x"ae",
          4748 => x"15",
          4749 => x"98",
          4750 => x"26",
          4751 => x"55",
          4752 => x"08",
          4753 => x"99",
          4754 => x"84",
          4755 => x"ff",
          4756 => x"d3",
          4757 => x"38",
          4758 => x"75",
          4759 => x"81",
          4760 => x"93",
          4761 => x"80",
          4762 => x"2e",
          4763 => x"ff",
          4764 => x"58",
          4765 => x"7d",
          4766 => x"38",
          4767 => x"55",
          4768 => x"b4",
          4769 => x"56",
          4770 => x"09",
          4771 => x"38",
          4772 => x"53",
          4773 => x"51",
          4774 => x"3f",
          4775 => x"08",
          4776 => x"84",
          4777 => x"38",
          4778 => x"ff",
          4779 => x"5c",
          4780 => x"84",
          4781 => x"5c",
          4782 => x"12",
          4783 => x"80",
          4784 => x"78",
          4785 => x"7c",
          4786 => x"90",
          4787 => x"c0",
          4788 => x"90",
          4789 => x"15",
          4790 => x"90",
          4791 => x"54",
          4792 => x"91",
          4793 => x"31",
          4794 => x"84",
          4795 => x"07",
          4796 => x"16",
          4797 => x"73",
          4798 => x"0c",
          4799 => x"04",
          4800 => x"6b",
          4801 => x"05",
          4802 => x"33",
          4803 => x"5a",
          4804 => x"bd",
          4805 => x"80",
          4806 => x"84",
          4807 => x"f8",
          4808 => x"84",
          4809 => x"81",
          4810 => x"70",
          4811 => x"74",
          4812 => x"38",
          4813 => x"81",
          4814 => x"81",
          4815 => x"81",
          4816 => x"ff",
          4817 => x"81",
          4818 => x"81",
          4819 => x"81",
          4820 => x"83",
          4821 => x"c0",
          4822 => x"2a",
          4823 => x"51",
          4824 => x"74",
          4825 => x"99",
          4826 => x"53",
          4827 => x"51",
          4828 => x"3f",
          4829 => x"08",
          4830 => x"55",
          4831 => x"92",
          4832 => x"80",
          4833 => x"38",
          4834 => x"06",
          4835 => x"2e",
          4836 => x"48",
          4837 => x"87",
          4838 => x"79",
          4839 => x"78",
          4840 => x"26",
          4841 => x"19",
          4842 => x"74",
          4843 => x"38",
          4844 => x"e4",
          4845 => x"2a",
          4846 => x"70",
          4847 => x"59",
          4848 => x"7a",
          4849 => x"56",
          4850 => x"80",
          4851 => x"51",
          4852 => x"74",
          4853 => x"99",
          4854 => x"53",
          4855 => x"51",
          4856 => x"3f",
          4857 => x"d3",
          4858 => x"ac",
          4859 => x"2a",
          4860 => x"81",
          4861 => x"43",
          4862 => x"83",
          4863 => x"66",
          4864 => x"60",
          4865 => x"90",
          4866 => x"31",
          4867 => x"80",
          4868 => x"8a",
          4869 => x"56",
          4870 => x"26",
          4871 => x"77",
          4872 => x"81",
          4873 => x"74",
          4874 => x"38",
          4875 => x"55",
          4876 => x"83",
          4877 => x"81",
          4878 => x"80",
          4879 => x"38",
          4880 => x"55",
          4881 => x"5e",
          4882 => x"89",
          4883 => x"5a",
          4884 => x"09",
          4885 => x"e1",
          4886 => x"38",
          4887 => x"57",
          4888 => x"c4",
          4889 => x"5a",
          4890 => x"9d",
          4891 => x"26",
          4892 => x"c4",
          4893 => x"10",
          4894 => x"22",
          4895 => x"74",
          4896 => x"38",
          4897 => x"ee",
          4898 => x"66",
          4899 => x"e9",
          4900 => x"84",
          4901 => x"84",
          4902 => x"89",
          4903 => x"a0",
          4904 => x"81",
          4905 => x"fc",
          4906 => x"56",
          4907 => x"f0",
          4908 => x"80",
          4909 => x"d3",
          4910 => x"38",
          4911 => x"57",
          4912 => x"c4",
          4913 => x"5a",
          4914 => x"9d",
          4915 => x"26",
          4916 => x"c4",
          4917 => x"10",
          4918 => x"22",
          4919 => x"74",
          4920 => x"38",
          4921 => x"ee",
          4922 => x"66",
          4923 => x"89",
          4924 => x"84",
          4925 => x"05",
          4926 => x"84",
          4927 => x"26",
          4928 => x"0b",
          4929 => x"08",
          4930 => x"84",
          4931 => x"11",
          4932 => x"05",
          4933 => x"83",
          4934 => x"2a",
          4935 => x"a0",
          4936 => x"7d",
          4937 => x"69",
          4938 => x"05",
          4939 => x"72",
          4940 => x"5c",
          4941 => x"59",
          4942 => x"2e",
          4943 => x"89",
          4944 => x"60",
          4945 => x"84",
          4946 => x"5d",
          4947 => x"18",
          4948 => x"68",
          4949 => x"74",
          4950 => x"af",
          4951 => x"31",
          4952 => x"53",
          4953 => x"52",
          4954 => x"8d",
          4955 => x"84",
          4956 => x"83",
          4957 => x"06",
          4958 => x"d3",
          4959 => x"ff",
          4960 => x"dd",
          4961 => x"83",
          4962 => x"2a",
          4963 => x"be",
          4964 => x"39",
          4965 => x"09",
          4966 => x"c5",
          4967 => x"f5",
          4968 => x"84",
          4969 => x"38",
          4970 => x"79",
          4971 => x"80",
          4972 => x"38",
          4973 => x"96",
          4974 => x"06",
          4975 => x"2e",
          4976 => x"5e",
          4977 => x"81",
          4978 => x"9f",
          4979 => x"38",
          4980 => x"38",
          4981 => x"81",
          4982 => x"fc",
          4983 => x"ab",
          4984 => x"7d",
          4985 => x"81",
          4986 => x"7d",
          4987 => x"78",
          4988 => x"74",
          4989 => x"8e",
          4990 => x"9c",
          4991 => x"53",
          4992 => x"51",
          4993 => x"3f",
          4994 => x"c2",
          4995 => x"51",
          4996 => x"3f",
          4997 => x"8b",
          4998 => x"a1",
          4999 => x"8d",
          5000 => x"83",
          5001 => x"52",
          5002 => x"ff",
          5003 => x"81",
          5004 => x"34",
          5005 => x"70",
          5006 => x"2a",
          5007 => x"54",
          5008 => x"1b",
          5009 => x"88",
          5010 => x"74",
          5011 => x"26",
          5012 => x"83",
          5013 => x"52",
          5014 => x"ff",
          5015 => x"8a",
          5016 => x"a0",
          5017 => x"a1",
          5018 => x"0b",
          5019 => x"bf",
          5020 => x"51",
          5021 => x"3f",
          5022 => x"9a",
          5023 => x"a0",
          5024 => x"52",
          5025 => x"ff",
          5026 => x"7d",
          5027 => x"81",
          5028 => x"38",
          5029 => x"0a",
          5030 => x"1b",
          5031 => x"ce",
          5032 => x"a4",
          5033 => x"a0",
          5034 => x"52",
          5035 => x"ff",
          5036 => x"81",
          5037 => x"51",
          5038 => x"3f",
          5039 => x"1b",
          5040 => x"8c",
          5041 => x"0b",
          5042 => x"34",
          5043 => x"c2",
          5044 => x"53",
          5045 => x"52",
          5046 => x"51",
          5047 => x"88",
          5048 => x"a7",
          5049 => x"a0",
          5050 => x"83",
          5051 => x"52",
          5052 => x"ff",
          5053 => x"ff",
          5054 => x"1c",
          5055 => x"a6",
          5056 => x"53",
          5057 => x"52",
          5058 => x"ff",
          5059 => x"82",
          5060 => x"83",
          5061 => x"52",
          5062 => x"b4",
          5063 => x"60",
          5064 => x"7e",
          5065 => x"d7",
          5066 => x"81",
          5067 => x"83",
          5068 => x"83",
          5069 => x"06",
          5070 => x"75",
          5071 => x"05",
          5072 => x"7e",
          5073 => x"b7",
          5074 => x"53",
          5075 => x"51",
          5076 => x"3f",
          5077 => x"a4",
          5078 => x"51",
          5079 => x"3f",
          5080 => x"e4",
          5081 => x"e4",
          5082 => x"9f",
          5083 => x"18",
          5084 => x"1b",
          5085 => x"f6",
          5086 => x"83",
          5087 => x"ff",
          5088 => x"82",
          5089 => x"78",
          5090 => x"c4",
          5091 => x"60",
          5092 => x"7a",
          5093 => x"ff",
          5094 => x"75",
          5095 => x"53",
          5096 => x"51",
          5097 => x"3f",
          5098 => x"52",
          5099 => x"9f",
          5100 => x"56",
          5101 => x"83",
          5102 => x"06",
          5103 => x"52",
          5104 => x"9e",
          5105 => x"52",
          5106 => x"ff",
          5107 => x"f0",
          5108 => x"1b",
          5109 => x"87",
          5110 => x"55",
          5111 => x"83",
          5112 => x"74",
          5113 => x"ff",
          5114 => x"7c",
          5115 => x"74",
          5116 => x"38",
          5117 => x"54",
          5118 => x"52",
          5119 => x"99",
          5120 => x"d3",
          5121 => x"87",
          5122 => x"53",
          5123 => x"08",
          5124 => x"ff",
          5125 => x"76",
          5126 => x"31",
          5127 => x"cd",
          5128 => x"58",
          5129 => x"ff",
          5130 => x"55",
          5131 => x"83",
          5132 => x"61",
          5133 => x"26",
          5134 => x"57",
          5135 => x"53",
          5136 => x"51",
          5137 => x"3f",
          5138 => x"08",
          5139 => x"76",
          5140 => x"31",
          5141 => x"db",
          5142 => x"7d",
          5143 => x"38",
          5144 => x"83",
          5145 => x"8a",
          5146 => x"7d",
          5147 => x"38",
          5148 => x"81",
          5149 => x"80",
          5150 => x"80",
          5151 => x"7a",
          5152 => x"bc",
          5153 => x"d5",
          5154 => x"ff",
          5155 => x"83",
          5156 => x"77",
          5157 => x"0b",
          5158 => x"81",
          5159 => x"34",
          5160 => x"34",
          5161 => x"34",
          5162 => x"56",
          5163 => x"52",
          5164 => x"f1",
          5165 => x"0b",
          5166 => x"81",
          5167 => x"82",
          5168 => x"56",
          5169 => x"34",
          5170 => x"08",
          5171 => x"60",
          5172 => x"1b",
          5173 => x"96",
          5174 => x"83",
          5175 => x"ff",
          5176 => x"81",
          5177 => x"7a",
          5178 => x"ff",
          5179 => x"81",
          5180 => x"84",
          5181 => x"80",
          5182 => x"7e",
          5183 => x"e3",
          5184 => x"81",
          5185 => x"90",
          5186 => x"8e",
          5187 => x"81",
          5188 => x"81",
          5189 => x"56",
          5190 => x"84",
          5191 => x"0d",
          5192 => x"0d",
          5193 => x"93",
          5194 => x"38",
          5195 => x"81",
          5196 => x"52",
          5197 => x"81",
          5198 => x"81",
          5199 => x"c5",
          5200 => x"f9",
          5201 => x"cc",
          5202 => x"39",
          5203 => x"51",
          5204 => x"81",
          5205 => x"80",
          5206 => x"c6",
          5207 => x"dd",
          5208 => x"94",
          5209 => x"39",
          5210 => x"51",
          5211 => x"81",
          5212 => x"80",
          5213 => x"c6",
          5214 => x"c1",
          5215 => x"ec",
          5216 => x"81",
          5217 => x"b5",
          5218 => x"9c",
          5219 => x"81",
          5220 => x"a9",
          5221 => x"dc",
          5222 => x"81",
          5223 => x"9d",
          5224 => x"90",
          5225 => x"81",
          5226 => x"91",
          5227 => x"c0",
          5228 => x"81",
          5229 => x"85",
          5230 => x"e4",
          5231 => x"fb",
          5232 => x"0d",
          5233 => x"0d",
          5234 => x"56",
          5235 => x"26",
          5236 => x"52",
          5237 => x"29",
          5238 => x"87",
          5239 => x"51",
          5240 => x"3f",
          5241 => x"08",
          5242 => x"fe",
          5243 => x"81",
          5244 => x"54",
          5245 => x"52",
          5246 => x"51",
          5247 => x"3f",
          5248 => x"04",
          5249 => x"7d",
          5250 => x"8c",
          5251 => x"05",
          5252 => x"15",
          5253 => x"5a",
          5254 => x"5c",
          5255 => x"c9",
          5256 => x"8c",
          5257 => x"c9",
          5258 => x"87",
          5259 => x"55",
          5260 => x"80",
          5261 => x"90",
          5262 => x"79",
          5263 => x"38",
          5264 => x"74",
          5265 => x"78",
          5266 => x"72",
          5267 => x"c9",
          5268 => x"8c",
          5269 => x"39",
          5270 => x"51",
          5271 => x"3f",
          5272 => x"80",
          5273 => x"16",
          5274 => x"27",
          5275 => x"08",
          5276 => x"98",
          5277 => x"a7",
          5278 => x"81",
          5279 => x"ff",
          5280 => x"84",
          5281 => x"39",
          5282 => x"72",
          5283 => x"38",
          5284 => x"81",
          5285 => x"ff",
          5286 => x"89",
          5287 => x"c0",
          5288 => x"97",
          5289 => x"55",
          5290 => x"fa",
          5291 => x"80",
          5292 => x"c4",
          5293 => x"83",
          5294 => x"74",
          5295 => x"38",
          5296 => x"33",
          5297 => x"52",
          5298 => x"74",
          5299 => x"72",
          5300 => x"38",
          5301 => x"26",
          5302 => x"51",
          5303 => x"51",
          5304 => x"3f",
          5305 => x"d3",
          5306 => x"c8",
          5307 => x"cb",
          5308 => x"77",
          5309 => x"fe",
          5310 => x"81",
          5311 => x"98",
          5312 => x"2c",
          5313 => x"a0",
          5314 => x"06",
          5315 => x"fc",
          5316 => x"d3",
          5317 => x"2b",
          5318 => x"70",
          5319 => x"30",
          5320 => x"9f",
          5321 => x"56",
          5322 => x"9b",
          5323 => x"72",
          5324 => x"9b",
          5325 => x"06",
          5326 => x"53",
          5327 => x"1c",
          5328 => x"26",
          5329 => x"ff",
          5330 => x"d3",
          5331 => x"3d",
          5332 => x"3d",
          5333 => x"84",
          5334 => x"05",
          5335 => x"30",
          5336 => x"80",
          5337 => x"ff",
          5338 => x"51",
          5339 => x"5b",
          5340 => x"74",
          5341 => x"81",
          5342 => x"8c",
          5343 => x"57",
          5344 => x"81",
          5345 => x"56",
          5346 => x"08",
          5347 => x"d3",
          5348 => x"c0",
          5349 => x"81",
          5350 => x"59",
          5351 => x"05",
          5352 => x"53",
          5353 => x"51",
          5354 => x"81",
          5355 => x"56",
          5356 => x"08",
          5357 => x"55",
          5358 => x"89",
          5359 => x"75",
          5360 => x"d8",
          5361 => x"d8",
          5362 => x"e0",
          5363 => x"70",
          5364 => x"25",
          5365 => x"80",
          5366 => x"74",
          5367 => x"38",
          5368 => x"53",
          5369 => x"88",
          5370 => x"51",
          5371 => x"75",
          5372 => x"d3",
          5373 => x"3d",
          5374 => x"3d",
          5375 => x"84",
          5376 => x"33",
          5377 => x"57",
          5378 => x"52",
          5379 => x"c2",
          5380 => x"84",
          5381 => x"75",
          5382 => x"38",
          5383 => x"98",
          5384 => x"60",
          5385 => x"81",
          5386 => x"7e",
          5387 => x"77",
          5388 => x"84",
          5389 => x"39",
          5390 => x"81",
          5391 => x"89",
          5392 => x"fc",
          5393 => x"9b",
          5394 => x"c9",
          5395 => x"c9",
          5396 => x"ff",
          5397 => x"81",
          5398 => x"51",
          5399 => x"3f",
          5400 => x"54",
          5401 => x"53",
          5402 => x"33",
          5403 => x"fc",
          5404 => x"ab",
          5405 => x"2e",
          5406 => x"fe",
          5407 => x"3d",
          5408 => x"3d",
          5409 => x"96",
          5410 => x"ff",
          5411 => x"81",
          5412 => x"8e",
          5413 => x"98",
          5414 => x"86",
          5415 => x"fe",
          5416 => x"72",
          5417 => x"81",
          5418 => x"71",
          5419 => x"38",
          5420 => x"f5",
          5421 => x"ca",
          5422 => x"f7",
          5423 => x"51",
          5424 => x"3f",
          5425 => x"70",
          5426 => x"52",
          5427 => x"95",
          5428 => x"fe",
          5429 => x"81",
          5430 => x"fe",
          5431 => x"80",
          5432 => x"be",
          5433 => x"2a",
          5434 => x"51",
          5435 => x"2e",
          5436 => x"51",
          5437 => x"3f",
          5438 => x"51",
          5439 => x"3f",
          5440 => x"f5",
          5441 => x"84",
          5442 => x"06",
          5443 => x"80",
          5444 => x"81",
          5445 => x"8a",
          5446 => x"ec",
          5447 => x"82",
          5448 => x"fe",
          5449 => x"72",
          5450 => x"81",
          5451 => x"71",
          5452 => x"38",
          5453 => x"f4",
          5454 => x"cb",
          5455 => x"f6",
          5456 => x"51",
          5457 => x"3f",
          5458 => x"70",
          5459 => x"52",
          5460 => x"95",
          5461 => x"fe",
          5462 => x"81",
          5463 => x"fe",
          5464 => x"80",
          5465 => x"ba",
          5466 => x"2a",
          5467 => x"51",
          5468 => x"2e",
          5469 => x"51",
          5470 => x"3f",
          5471 => x"51",
          5472 => x"3f",
          5473 => x"f4",
          5474 => x"88",
          5475 => x"06",
          5476 => x"80",
          5477 => x"81",
          5478 => x"86",
          5479 => x"bc",
          5480 => x"fe",
          5481 => x"fe",
          5482 => x"fe",
          5483 => x"84",
          5484 => x"fa",
          5485 => x"70",
          5486 => x"55",
          5487 => x"2e",
          5488 => x"8e",
          5489 => x"0c",
          5490 => x"53",
          5491 => x"81",
          5492 => x"74",
          5493 => x"ff",
          5494 => x"53",
          5495 => x"83",
          5496 => x"74",
          5497 => x"38",
          5498 => x"75",
          5499 => x"53",
          5500 => x"09",
          5501 => x"38",
          5502 => x"81",
          5503 => x"80",
          5504 => x"29",
          5505 => x"05",
          5506 => x"70",
          5507 => x"fe",
          5508 => x"81",
          5509 => x"8b",
          5510 => x"33",
          5511 => x"2e",
          5512 => x"81",
          5513 => x"ff",
          5514 => x"93",
          5515 => x"38",
          5516 => x"81",
          5517 => x"88",
          5518 => x"cb",
          5519 => x"70",
          5520 => x"84",
          5521 => x"81",
          5522 => x"ff",
          5523 => x"81",
          5524 => x"81",
          5525 => x"78",
          5526 => x"81",
          5527 => x"81",
          5528 => x"99",
          5529 => x"59",
          5530 => x"3f",
          5531 => x"52",
          5532 => x"51",
          5533 => x"3f",
          5534 => x"08",
          5535 => x"38",
          5536 => x"51",
          5537 => x"81",
          5538 => x"81",
          5539 => x"fe",
          5540 => x"99",
          5541 => x"5a",
          5542 => x"80",
          5543 => x"fe",
          5544 => x"80",
          5545 => x"51",
          5546 => x"3f",
          5547 => x"f8",
          5548 => x"ff",
          5549 => x"84",
          5550 => x"70",
          5551 => x"59",
          5552 => x"2e",
          5553 => x"78",
          5554 => x"80",
          5555 => x"ab",
          5556 => x"38",
          5557 => x"a4",
          5558 => x"2e",
          5559 => x"78",
          5560 => x"38",
          5561 => x"ff",
          5562 => x"88",
          5563 => x"2e",
          5564 => x"78",
          5565 => x"ad",
          5566 => x"39",
          5567 => x"2e",
          5568 => x"78",
          5569 => x"90",
          5570 => x"2e",
          5571 => x"78",
          5572 => x"8b",
          5573 => x"39",
          5574 => x"2e",
          5575 => x"78",
          5576 => x"88",
          5577 => x"cc",
          5578 => x"f8",
          5579 => x"38",
          5580 => x"24",
          5581 => x"80",
          5582 => x"e2",
          5583 => x"d1",
          5584 => x"78",
          5585 => x"8a",
          5586 => x"a8",
          5587 => x"d4",
          5588 => x"38",
          5589 => x"2e",
          5590 => x"8c",
          5591 => x"81",
          5592 => x"fc",
          5593 => x"83",
          5594 => x"78",
          5595 => x"8b",
          5596 => x"81",
          5597 => x"d9",
          5598 => x"39",
          5599 => x"2e",
          5600 => x"78",
          5601 => x"fe",
          5602 => x"e8",
          5603 => x"fe",
          5604 => x"fe",
          5605 => x"ff",
          5606 => x"81",
          5607 => x"88",
          5608 => x"bc",
          5609 => x"39",
          5610 => x"f0",
          5611 => x"f8",
          5612 => x"83",
          5613 => x"d3",
          5614 => x"2e",
          5615 => x"63",
          5616 => x"80",
          5617 => x"cb",
          5618 => x"02",
          5619 => x"33",
          5620 => x"c2",
          5621 => x"84",
          5622 => x"06",
          5623 => x"38",
          5624 => x"51",
          5625 => x"3f",
          5626 => x"9f",
          5627 => x"dc",
          5628 => x"39",
          5629 => x"f4",
          5630 => x"f8",
          5631 => x"83",
          5632 => x"d3",
          5633 => x"2e",
          5634 => x"80",
          5635 => x"02",
          5636 => x"33",
          5637 => x"cb",
          5638 => x"84",
          5639 => x"cc",
          5640 => x"a6",
          5641 => x"fe",
          5642 => x"fe",
          5643 => x"ff",
          5644 => x"81",
          5645 => x"80",
          5646 => x"63",
          5647 => x"cb",
          5648 => x"fe",
          5649 => x"fe",
          5650 => x"ff",
          5651 => x"81",
          5652 => x"86",
          5653 => x"84",
          5654 => x"53",
          5655 => x"52",
          5656 => x"80",
          5657 => x"80",
          5658 => x"53",
          5659 => x"84",
          5660 => x"d4",
          5661 => x"ff",
          5662 => x"81",
          5663 => x"81",
          5664 => x"cc",
          5665 => x"fa",
          5666 => x"5c",
          5667 => x"b7",
          5668 => x"05",
          5669 => x"bb",
          5670 => x"84",
          5671 => x"fe",
          5672 => x"5b",
          5673 => x"3f",
          5674 => x"d3",
          5675 => x"7a",
          5676 => x"3f",
          5677 => x"b7",
          5678 => x"05",
          5679 => x"93",
          5680 => x"84",
          5681 => x"fe",
          5682 => x"5b",
          5683 => x"3f",
          5684 => x"08",
          5685 => x"f8",
          5686 => x"fe",
          5687 => x"81",
          5688 => x"b8",
          5689 => x"05",
          5690 => x"ea",
          5691 => x"d0",
          5692 => x"d3",
          5693 => x"56",
          5694 => x"d3",
          5695 => x"ff",
          5696 => x"53",
          5697 => x"51",
          5698 => x"81",
          5699 => x"80",
          5700 => x"38",
          5701 => x"08",
          5702 => x"3f",
          5703 => x"b7",
          5704 => x"11",
          5705 => x"05",
          5706 => x"e8",
          5707 => x"84",
          5708 => x"fa",
          5709 => x"3d",
          5710 => x"53",
          5711 => x"51",
          5712 => x"3f",
          5713 => x"08",
          5714 => x"bf",
          5715 => x"fe",
          5716 => x"fe",
          5717 => x"ff",
          5718 => x"81",
          5719 => x"86",
          5720 => x"84",
          5721 => x"cd",
          5722 => x"f8",
          5723 => x"63",
          5724 => x"7b",
          5725 => x"61",
          5726 => x"70",
          5727 => x"0c",
          5728 => x"f5",
          5729 => x"c8",
          5730 => x"39",
          5731 => x"f4",
          5732 => x"f8",
          5733 => x"ff",
          5734 => x"d3",
          5735 => x"c4",
          5736 => x"ad",
          5737 => x"80",
          5738 => x"81",
          5739 => x"44",
          5740 => x"d0",
          5741 => x"78",
          5742 => x"38",
          5743 => x"08",
          5744 => x"81",
          5745 => x"59",
          5746 => x"81",
          5747 => x"59",
          5748 => x"88",
          5749 => x"90",
          5750 => x"39",
          5751 => x"08",
          5752 => x"44",
          5753 => x"f0",
          5754 => x"f8",
          5755 => x"ff",
          5756 => x"d3",
          5757 => x"c3",
          5758 => x"ad",
          5759 => x"80",
          5760 => x"81",
          5761 => x"43",
          5762 => x"d0",
          5763 => x"78",
          5764 => x"38",
          5765 => x"08",
          5766 => x"81",
          5767 => x"59",
          5768 => x"81",
          5769 => x"59",
          5770 => x"88",
          5771 => x"94",
          5772 => x"39",
          5773 => x"08",
          5774 => x"b7",
          5775 => x"11",
          5776 => x"05",
          5777 => x"cc",
          5778 => x"84",
          5779 => x"9b",
          5780 => x"5b",
          5781 => x"2e",
          5782 => x"59",
          5783 => x"8d",
          5784 => x"2e",
          5785 => x"a0",
          5786 => x"88",
          5787 => x"8c",
          5788 => x"c7",
          5789 => x"63",
          5790 => x"62",
          5791 => x"ef",
          5792 => x"cd",
          5793 => x"bd",
          5794 => x"fe",
          5795 => x"fe",
          5796 => x"fe",
          5797 => x"81",
          5798 => x"80",
          5799 => x"38",
          5800 => x"f0",
          5801 => x"f8",
          5802 => x"fd",
          5803 => x"d3",
          5804 => x"2e",
          5805 => x"59",
          5806 => x"05",
          5807 => x"63",
          5808 => x"b7",
          5809 => x"11",
          5810 => x"05",
          5811 => x"c4",
          5812 => x"84",
          5813 => x"f7",
          5814 => x"70",
          5815 => x"81",
          5816 => x"fe",
          5817 => x"80",
          5818 => x"51",
          5819 => x"3f",
          5820 => x"33",
          5821 => x"2e",
          5822 => x"9f",
          5823 => x"38",
          5824 => x"f0",
          5825 => x"f8",
          5826 => x"fd",
          5827 => x"d3",
          5828 => x"2e",
          5829 => x"59",
          5830 => x"05",
          5831 => x"63",
          5832 => x"ff",
          5833 => x"cd",
          5834 => x"f5",
          5835 => x"aa",
          5836 => x"fe",
          5837 => x"fe",
          5838 => x"fe",
          5839 => x"81",
          5840 => x"80",
          5841 => x"38",
          5842 => x"e4",
          5843 => x"f8",
          5844 => x"fe",
          5845 => x"d3",
          5846 => x"2e",
          5847 => x"59",
          5848 => x"22",
          5849 => x"05",
          5850 => x"41",
          5851 => x"e4",
          5852 => x"f8",
          5853 => x"fe",
          5854 => x"d3",
          5855 => x"38",
          5856 => x"60",
          5857 => x"52",
          5858 => x"51",
          5859 => x"3f",
          5860 => x"79",
          5861 => x"e1",
          5862 => x"79",
          5863 => x"ae",
          5864 => x"38",
          5865 => x"87",
          5866 => x"05",
          5867 => x"b7",
          5868 => x"11",
          5869 => x"05",
          5870 => x"ca",
          5871 => x"84",
          5872 => x"92",
          5873 => x"02",
          5874 => x"79",
          5875 => x"5b",
          5876 => x"ff",
          5877 => x"cd",
          5878 => x"f3",
          5879 => x"a3",
          5880 => x"fe",
          5881 => x"fe",
          5882 => x"fe",
          5883 => x"81",
          5884 => x"80",
          5885 => x"38",
          5886 => x"e4",
          5887 => x"f8",
          5888 => x"fd",
          5889 => x"d3",
          5890 => x"2e",
          5891 => x"60",
          5892 => x"60",
          5893 => x"b7",
          5894 => x"11",
          5895 => x"05",
          5896 => x"e2",
          5897 => x"84",
          5898 => x"f4",
          5899 => x"70",
          5900 => x"81",
          5901 => x"fe",
          5902 => x"80",
          5903 => x"51",
          5904 => x"3f",
          5905 => x"33",
          5906 => x"2e",
          5907 => x"9f",
          5908 => x"38",
          5909 => x"e4",
          5910 => x"f8",
          5911 => x"fc",
          5912 => x"d3",
          5913 => x"2e",
          5914 => x"53",
          5915 => x"cd",
          5916 => x"f8",
          5917 => x"60",
          5918 => x"60",
          5919 => x"ff",
          5920 => x"cd",
          5921 => x"f2",
          5922 => x"a2",
          5923 => x"d4",
          5924 => x"a7",
          5925 => x"fe",
          5926 => x"f3",
          5927 => x"cd",
          5928 => x"f2",
          5929 => x"51",
          5930 => x"3f",
          5931 => x"84",
          5932 => x"87",
          5933 => x"0c",
          5934 => x"0b",
          5935 => x"94",
          5936 => x"84",
          5937 => x"f3",
          5938 => x"39",
          5939 => x"51",
          5940 => x"3f",
          5941 => x"0b",
          5942 => x"84",
          5943 => x"83",
          5944 => x"94",
          5945 => x"a3",
          5946 => x"fe",
          5947 => x"fe",
          5948 => x"fe",
          5949 => x"81",
          5950 => x"80",
          5951 => x"38",
          5952 => x"ce",
          5953 => x"f7",
          5954 => x"59",
          5955 => x"3d",
          5956 => x"53",
          5957 => x"51",
          5958 => x"3f",
          5959 => x"08",
          5960 => x"e7",
          5961 => x"81",
          5962 => x"fe",
          5963 => x"63",
          5964 => x"81",
          5965 => x"5e",
          5966 => x"08",
          5967 => x"cb",
          5968 => x"84",
          5969 => x"ce",
          5970 => x"f6",
          5971 => x"bb",
          5972 => x"80",
          5973 => x"e3",
          5974 => x"a6",
          5975 => x"39",
          5976 => x"51",
          5977 => x"3f",
          5978 => x"a0",
          5979 => x"a1",
          5980 => x"39",
          5981 => x"51",
          5982 => x"2e",
          5983 => x"7b",
          5984 => x"d2",
          5985 => x"2e",
          5986 => x"b7",
          5987 => x"05",
          5988 => x"bf",
          5989 => x"b0",
          5990 => x"84",
          5991 => x"cf",
          5992 => x"53",
          5993 => x"52",
          5994 => x"52",
          5995 => x"85",
          5996 => x"80",
          5997 => x"b8",
          5998 => x"64",
          5999 => x"81",
          6000 => x"54",
          6001 => x"53",
          6002 => x"52",
          6003 => x"aa",
          6004 => x"84",
          6005 => x"81",
          6006 => x"32",
          6007 => x"8a",
          6008 => x"2e",
          6009 => x"f1",
          6010 => x"cf",
          6011 => x"f5",
          6012 => x"97",
          6013 => x"0d",
          6014 => x"d3",
          6015 => x"90",
          6016 => x"87",
          6017 => x"0c",
          6018 => x"e4",
          6019 => x"94",
          6020 => x"80",
          6021 => x"c0",
          6022 => x"8c",
          6023 => x"87",
          6024 => x"0c",
          6025 => x"81",
          6026 => x"a2",
          6027 => x"d3",
          6028 => x"e7",
          6029 => x"ed",
          6030 => x"cf",
          6031 => x"e4",
          6032 => x"cf",
          6033 => x"ee",
          6034 => x"a9",
          6035 => x"ed",
          6036 => x"51",
          6037 => x"ef",
          6038 => x"04",
          6039 => x"ff",
          6040 => x"00",
          6041 => x"ff",
          6042 => x"ff",
          6043 => x"00",
          6044 => x"00",
          6045 => x"00",
          6046 => x"00",
          6047 => x"00",
          6048 => x"00",
          6049 => x"00",
          6050 => x"00",
          6051 => x"00",
          6052 => x"00",
          6053 => x"00",
          6054 => x"00",
          6055 => x"00",
          6056 => x"00",
          6057 => x"00",
          6058 => x"00",
          6059 => x"00",
          6060 => x"00",
          6061 => x"00",
          6062 => x"00",
          6063 => x"00",
          6064 => x"00",
          6065 => x"00",
          6066 => x"00",
          6067 => x"00",
          6068 => x"64",
          6069 => x"2f",
          6070 => x"25",
          6071 => x"64",
          6072 => x"2e",
          6073 => x"64",
          6074 => x"6f",
          6075 => x"6f",
          6076 => x"67",
          6077 => x"74",
          6078 => x"00",
          6079 => x"28",
          6080 => x"6d",
          6081 => x"43",
          6082 => x"6e",
          6083 => x"29",
          6084 => x"0a",
          6085 => x"69",
          6086 => x"20",
          6087 => x"6c",
          6088 => x"6e",
          6089 => x"3a",
          6090 => x"20",
          6091 => x"4e",
          6092 => x"42",
          6093 => x"20",
          6094 => x"61",
          6095 => x"25",
          6096 => x"2c",
          6097 => x"7a",
          6098 => x"30",
          6099 => x"2e",
          6100 => x"20",
          6101 => x"52",
          6102 => x"28",
          6103 => x"72",
          6104 => x"30",
          6105 => x"20",
          6106 => x"65",
          6107 => x"38",
          6108 => x"0a",
          6109 => x"20",
          6110 => x"41",
          6111 => x"53",
          6112 => x"74",
          6113 => x"38",
          6114 => x"53",
          6115 => x"3d",
          6116 => x"58",
          6117 => x"00",
          6118 => x"20",
          6119 => x"4f",
          6120 => x"0a",
          6121 => x"20",
          6122 => x"53",
          6123 => x"00",
          6124 => x"20",
          6125 => x"50",
          6126 => x"00",
          6127 => x"20",
          6128 => x"44",
          6129 => x"72",
          6130 => x"44",
          6131 => x"63",
          6132 => x"25",
          6133 => x"29",
          6134 => x"00",
          6135 => x"20",
          6136 => x"4e",
          6137 => x"52",
          6138 => x"20",
          6139 => x"54",
          6140 => x"4c",
          6141 => x"00",
          6142 => x"20",
          6143 => x"49",
          6144 => x"31",
          6145 => x"69",
          6146 => x"73",
          6147 => x"31",
          6148 => x"0a",
          6149 => x"64",
          6150 => x"73",
          6151 => x"3a",
          6152 => x"20",
          6153 => x"50",
          6154 => x"65",
          6155 => x"20",
          6156 => x"74",
          6157 => x"41",
          6158 => x"65",
          6159 => x"3d",
          6160 => x"38",
          6161 => x"00",
          6162 => x"20",
          6163 => x"50",
          6164 => x"65",
          6165 => x"79",
          6166 => x"61",
          6167 => x"41",
          6168 => x"65",
          6169 => x"3d",
          6170 => x"38",
          6171 => x"00",
          6172 => x"20",
          6173 => x"74",
          6174 => x"20",
          6175 => x"72",
          6176 => x"64",
          6177 => x"73",
          6178 => x"20",
          6179 => x"3d",
          6180 => x"38",
          6181 => x"00",
          6182 => x"20",
          6183 => x"50",
          6184 => x"64",
          6185 => x"20",
          6186 => x"20",
          6187 => x"20",
          6188 => x"20",
          6189 => x"3d",
          6190 => x"38",
          6191 => x"00",
          6192 => x"20",
          6193 => x"79",
          6194 => x"6d",
          6195 => x"6f",
          6196 => x"46",
          6197 => x"20",
          6198 => x"20",
          6199 => x"3d",
          6200 => x"38",
          6201 => x"00",
          6202 => x"6d",
          6203 => x"00",
          6204 => x"65",
          6205 => x"6d",
          6206 => x"6c",
          6207 => x"00",
          6208 => x"56",
          6209 => x"56",
          6210 => x"6e",
          6211 => x"6e",
          6212 => x"77",
          6213 => x"44",
          6214 => x"2a",
          6215 => x"3b",
          6216 => x"3f",
          6217 => x"7f",
          6218 => x"41",
          6219 => x"41",
          6220 => x"00",
          6221 => x"fe",
          6222 => x"44",
          6223 => x"2e",
          6224 => x"4f",
          6225 => x"4d",
          6226 => x"20",
          6227 => x"54",
          6228 => x"20",
          6229 => x"4f",
          6230 => x"4d",
          6231 => x"20",
          6232 => x"54",
          6233 => x"20",
          6234 => x"00",
          6235 => x"00",
          6236 => x"00",
          6237 => x"00",
          6238 => x"9a",
          6239 => x"41",
          6240 => x"45",
          6241 => x"49",
          6242 => x"92",
          6243 => x"4f",
          6244 => x"99",
          6245 => x"9d",
          6246 => x"49",
          6247 => x"a5",
          6248 => x"a9",
          6249 => x"ad",
          6250 => x"b1",
          6251 => x"b5",
          6252 => x"b9",
          6253 => x"bd",
          6254 => x"c1",
          6255 => x"c5",
          6256 => x"c9",
          6257 => x"cd",
          6258 => x"d1",
          6259 => x"d5",
          6260 => x"d9",
          6261 => x"dd",
          6262 => x"e1",
          6263 => x"e5",
          6264 => x"e9",
          6265 => x"ed",
          6266 => x"f1",
          6267 => x"f5",
          6268 => x"f9",
          6269 => x"fd",
          6270 => x"2e",
          6271 => x"5b",
          6272 => x"22",
          6273 => x"3e",
          6274 => x"00",
          6275 => x"01",
          6276 => x"10",
          6277 => x"00",
          6278 => x"00",
          6279 => x"01",
          6280 => x"04",
          6281 => x"10",
          6282 => x"00",
          6283 => x"69",
          6284 => x"00",
          6285 => x"69",
          6286 => x"6c",
          6287 => x"69",
          6288 => x"00",
          6289 => x"6c",
          6290 => x"00",
          6291 => x"65",
          6292 => x"00",
          6293 => x"63",
          6294 => x"72",
          6295 => x"64",
          6296 => x"00",
          6297 => x"65",
          6298 => x"65",
          6299 => x"65",
          6300 => x"69",
          6301 => x"69",
          6302 => x"66",
          6303 => x"66",
          6304 => x"61",
          6305 => x"00",
          6306 => x"6d",
          6307 => x"65",
          6308 => x"72",
          6309 => x"65",
          6310 => x"00",
          6311 => x"6e",
          6312 => x"00",
          6313 => x"65",
          6314 => x"00",
          6315 => x"69",
          6316 => x"45",
          6317 => x"72",
          6318 => x"6e",
          6319 => x"6e",
          6320 => x"65",
          6321 => x"72",
          6322 => x"00",
          6323 => x"69",
          6324 => x"6e",
          6325 => x"72",
          6326 => x"79",
          6327 => x"00",
          6328 => x"6f",
          6329 => x"6c",
          6330 => x"6f",
          6331 => x"2e",
          6332 => x"6f",
          6333 => x"74",
          6334 => x"6f",
          6335 => x"2e",
          6336 => x"6e",
          6337 => x"69",
          6338 => x"69",
          6339 => x"61",
          6340 => x"0a",
          6341 => x"63",
          6342 => x"73",
          6343 => x"6e",
          6344 => x"2e",
          6345 => x"69",
          6346 => x"61",
          6347 => x"61",
          6348 => x"65",
          6349 => x"74",
          6350 => x"00",
          6351 => x"69",
          6352 => x"68",
          6353 => x"6c",
          6354 => x"6e",
          6355 => x"69",
          6356 => x"00",
          6357 => x"44",
          6358 => x"20",
          6359 => x"74",
          6360 => x"72",
          6361 => x"63",
          6362 => x"2e",
          6363 => x"72",
          6364 => x"20",
          6365 => x"62",
          6366 => x"69",
          6367 => x"6e",
          6368 => x"69",
          6369 => x"00",
          6370 => x"69",
          6371 => x"6e",
          6372 => x"65",
          6373 => x"6c",
          6374 => x"0a",
          6375 => x"6f",
          6376 => x"6d",
          6377 => x"69",
          6378 => x"20",
          6379 => x"65",
          6380 => x"74",
          6381 => x"66",
          6382 => x"64",
          6383 => x"20",
          6384 => x"6b",
          6385 => x"00",
          6386 => x"6f",
          6387 => x"74",
          6388 => x"6f",
          6389 => x"64",
          6390 => x"00",
          6391 => x"69",
          6392 => x"75",
          6393 => x"6f",
          6394 => x"61",
          6395 => x"6e",
          6396 => x"6e",
          6397 => x"6c",
          6398 => x"0a",
          6399 => x"69",
          6400 => x"69",
          6401 => x"6f",
          6402 => x"64",
          6403 => x"00",
          6404 => x"6e",
          6405 => x"66",
          6406 => x"65",
          6407 => x"6d",
          6408 => x"72",
          6409 => x"00",
          6410 => x"6f",
          6411 => x"61",
          6412 => x"6f",
          6413 => x"20",
          6414 => x"65",
          6415 => x"00",
          6416 => x"61",
          6417 => x"65",
          6418 => x"73",
          6419 => x"63",
          6420 => x"65",
          6421 => x"0a",
          6422 => x"75",
          6423 => x"73",
          6424 => x"00",
          6425 => x"6e",
          6426 => x"77",
          6427 => x"72",
          6428 => x"2e",
          6429 => x"25",
          6430 => x"62",
          6431 => x"73",
          6432 => x"20",
          6433 => x"25",
          6434 => x"62",
          6435 => x"73",
          6436 => x"63",
          6437 => x"00",
          6438 => x"30",
          6439 => x"00",
          6440 => x"20",
          6441 => x"30",
          6442 => x"00",
          6443 => x"20",
          6444 => x"20",
          6445 => x"00",
          6446 => x"30",
          6447 => x"00",
          6448 => x"20",
          6449 => x"7c",
          6450 => x"0d",
          6451 => x"65",
          6452 => x"00",
          6453 => x"50",
          6454 => x"00",
          6455 => x"2a",
          6456 => x"73",
          6457 => x"00",
          6458 => x"38",
          6459 => x"2f",
          6460 => x"39",
          6461 => x"31",
          6462 => x"00",
          6463 => x"5a",
          6464 => x"20",
          6465 => x"20",
          6466 => x"78",
          6467 => x"73",
          6468 => x"20",
          6469 => x"0a",
          6470 => x"50",
          6471 => x"20",
          6472 => x"65",
          6473 => x"70",
          6474 => x"61",
          6475 => x"65",
          6476 => x"00",
          6477 => x"69",
          6478 => x"20",
          6479 => x"65",
          6480 => x"70",
          6481 => x"00",
          6482 => x"53",
          6483 => x"6e",
          6484 => x"72",
          6485 => x"0a",
          6486 => x"4f",
          6487 => x"20",
          6488 => x"69",
          6489 => x"72",
          6490 => x"74",
          6491 => x"4f",
          6492 => x"20",
          6493 => x"69",
          6494 => x"72",
          6495 => x"74",
          6496 => x"41",
          6497 => x"20",
          6498 => x"69",
          6499 => x"72",
          6500 => x"74",
          6501 => x"41",
          6502 => x"20",
          6503 => x"69",
          6504 => x"72",
          6505 => x"74",
          6506 => x"41",
          6507 => x"20",
          6508 => x"69",
          6509 => x"72",
          6510 => x"74",
          6511 => x"41",
          6512 => x"20",
          6513 => x"69",
          6514 => x"72",
          6515 => x"74",
          6516 => x"65",
          6517 => x"6e",
          6518 => x"70",
          6519 => x"6d",
          6520 => x"2e",
          6521 => x"00",
          6522 => x"6e",
          6523 => x"69",
          6524 => x"74",
          6525 => x"72",
          6526 => x"0a",
          6527 => x"3a",
          6528 => x"61",
          6529 => x"64",
          6530 => x"20",
          6531 => x"74",
          6532 => x"69",
          6533 => x"73",
          6534 => x"61",
          6535 => x"30",
          6536 => x"6c",
          6537 => x"65",
          6538 => x"69",
          6539 => x"61",
          6540 => x"6c",
          6541 => x"0a",
          6542 => x"20",
          6543 => x"61",
          6544 => x"69",
          6545 => x"69",
          6546 => x"00",
          6547 => x"6e",
          6548 => x"61",
          6549 => x"65",
          6550 => x"00",
          6551 => x"61",
          6552 => x"64",
          6553 => x"20",
          6554 => x"74",
          6555 => x"69",
          6556 => x"0a",
          6557 => x"63",
          6558 => x"0a",
          6559 => x"75",
          6560 => x"6c",
          6561 => x"69",
          6562 => x"2e",
          6563 => x"75",
          6564 => x"4d",
          6565 => x"72",
          6566 => x"00",
          6567 => x"43",
          6568 => x"6c",
          6569 => x"2e",
          6570 => x"30",
          6571 => x"25",
          6572 => x"2d",
          6573 => x"3f",
          6574 => x"00",
          6575 => x"30",
          6576 => x"25",
          6577 => x"2d",
          6578 => x"30",
          6579 => x"25",
          6580 => x"2d",
          6581 => x"69",
          6582 => x"6c",
          6583 => x"20",
          6584 => x"65",
          6585 => x"70",
          6586 => x"00",
          6587 => x"6e",
          6588 => x"69",
          6589 => x"69",
          6590 => x"72",
          6591 => x"74",
          6592 => x"00",
          6593 => x"69",
          6594 => x"6c",
          6595 => x"75",
          6596 => x"20",
          6597 => x"6f",
          6598 => x"6e",
          6599 => x"69",
          6600 => x"75",
          6601 => x"20",
          6602 => x"6f",
          6603 => x"78",
          6604 => x"74",
          6605 => x"20",
          6606 => x"65",
          6607 => x"25",
          6608 => x"20",
          6609 => x"0a",
          6610 => x"61",
          6611 => x"6e",
          6612 => x"6f",
          6613 => x"40",
          6614 => x"38",
          6615 => x"2e",
          6616 => x"00",
          6617 => x"61",
          6618 => x"72",
          6619 => x"72",
          6620 => x"20",
          6621 => x"65",
          6622 => x"64",
          6623 => x"00",
          6624 => x"65",
          6625 => x"72",
          6626 => x"67",
          6627 => x"70",
          6628 => x"61",
          6629 => x"6e",
          6630 => x"0a",
          6631 => x"6f",
          6632 => x"72",
          6633 => x"6f",
          6634 => x"67",
          6635 => x"0a",
          6636 => x"50",
          6637 => x"69",
          6638 => x"64",
          6639 => x"73",
          6640 => x"2e",
          6641 => x"00",
          6642 => x"61",
          6643 => x"6f",
          6644 => x"6e",
          6645 => x"00",
          6646 => x"75",
          6647 => x"6e",
          6648 => x"2e",
          6649 => x"6e",
          6650 => x"69",
          6651 => x"69",
          6652 => x"72",
          6653 => x"74",
          6654 => x"2e",
          6655 => x"00",
          6656 => x"00",
          6657 => x"00",
          6658 => x"00",
          6659 => x"00",
          6660 => x"01",
          6661 => x"00",
          6662 => x"00",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"f5",
          6667 => x"01",
          6668 => x"01",
          6669 => x"01",
          6670 => x"00",
          6671 => x"00",
          6672 => x"00",
          6673 => x"00",
          6674 => x"02",
          6675 => x"00",
          6676 => x"00",
          6677 => x"00",
          6678 => x"04",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"14",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"2b",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"30",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"3c",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"40",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"41",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"42",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"43",
          6711 => x"00",
          6712 => x"00",
          6713 => x"00",
          6714 => x"50",
          6715 => x"00",
          6716 => x"00",
          6717 => x"00",
          6718 => x"51",
          6719 => x"00",
          6720 => x"00",
          6721 => x"00",
          6722 => x"54",
          6723 => x"00",
          6724 => x"00",
          6725 => x"00",
          6726 => x"55",
          6727 => x"00",
          6728 => x"00",
          6729 => x"00",
          6730 => x"79",
          6731 => x"00",
          6732 => x"00",
          6733 => x"00",
          6734 => x"78",
          6735 => x"00",
          6736 => x"00",
          6737 => x"00",
          6738 => x"82",
          6739 => x"00",
          6740 => x"00",
          6741 => x"00",
          6742 => x"83",
          6743 => x"00",
          6744 => x"00",
          6745 => x"00",
          6746 => x"85",
          6747 => x"00",
          6748 => x"00",
          6749 => x"00",
          6750 => x"87",
          6751 => x"00",
          6752 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"d8",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"bc",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"dc",
           163 => x"10",
           164 => x"06",
           165 => x"92",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"dd",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"c9",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"94",
           269 => x"0b",
           270 => x"0b",
           271 => x"b2",
           272 => x"0b",
           273 => x"0b",
           274 => x"d0",
           275 => x"0b",
           276 => x"0b",
           277 => x"ee",
           278 => x"0b",
           279 => x"0b",
           280 => x"8c",
           281 => x"0b",
           282 => x"0b",
           283 => x"aa",
           284 => x"0b",
           285 => x"0b",
           286 => x"c8",
           287 => x"0b",
           288 => x"0b",
           289 => x"e6",
           290 => x"0b",
           291 => x"0b",
           292 => x"84",
           293 => x"0b",
           294 => x"0b",
           295 => x"a4",
           296 => x"0b",
           297 => x"0b",
           298 => x"c4",
           299 => x"0b",
           300 => x"0b",
           301 => x"e4",
           302 => x"0b",
           303 => x"0b",
           304 => x"84",
           305 => x"0b",
           306 => x"0b",
           307 => x"a4",
           308 => x"0b",
           309 => x"0b",
           310 => x"c4",
           311 => x"0b",
           312 => x"0b",
           313 => x"e4",
           314 => x"0b",
           315 => x"0b",
           316 => x"84",
           317 => x"0b",
           318 => x"0b",
           319 => x"a4",
           320 => x"0b",
           321 => x"0b",
           322 => x"c4",
           323 => x"0b",
           324 => x"0b",
           325 => x"e4",
           326 => x"0b",
           327 => x"0b",
           328 => x"84",
           329 => x"0b",
           330 => x"0b",
           331 => x"a3",
           332 => x"0b",
           333 => x"0b",
           334 => x"c1",
           335 => x"0b",
           336 => x"0b",
           337 => x"df",
           338 => x"0b",
           339 => x"ff",
           340 => x"ff",
           341 => x"ff",
           342 => x"ff",
           343 => x"ff",
           344 => x"ff",
           345 => x"ff",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"81",
           388 => x"82",
           389 => x"81",
           390 => x"aa",
           391 => x"d3",
           392 => x"a0",
           393 => x"d3",
           394 => x"9b",
           395 => x"90",
           396 => x"90",
           397 => x"90",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"81",
           403 => x"82",
           404 => x"81",
           405 => x"b2",
           406 => x"d3",
           407 => x"a0",
           408 => x"d3",
           409 => x"dc",
           410 => x"90",
           411 => x"90",
           412 => x"90",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"81",
           418 => x"82",
           419 => x"81",
           420 => x"b1",
           421 => x"d3",
           422 => x"a0",
           423 => x"d3",
           424 => x"b3",
           425 => x"90",
           426 => x"90",
           427 => x"90",
           428 => x"2d",
           429 => x"08",
           430 => x"04",
           431 => x"0c",
           432 => x"81",
           433 => x"82",
           434 => x"81",
           435 => x"a3",
           436 => x"d3",
           437 => x"a0",
           438 => x"d3",
           439 => x"a8",
           440 => x"90",
           441 => x"90",
           442 => x"90",
           443 => x"2d",
           444 => x"08",
           445 => x"04",
           446 => x"0c",
           447 => x"81",
           448 => x"82",
           449 => x"81",
           450 => x"80",
           451 => x"81",
           452 => x"82",
           453 => x"81",
           454 => x"80",
           455 => x"81",
           456 => x"82",
           457 => x"81",
           458 => x"80",
           459 => x"81",
           460 => x"82",
           461 => x"81",
           462 => x"80",
           463 => x"81",
           464 => x"82",
           465 => x"81",
           466 => x"80",
           467 => x"81",
           468 => x"82",
           469 => x"81",
           470 => x"81",
           471 => x"81",
           472 => x"82",
           473 => x"81",
           474 => x"80",
           475 => x"81",
           476 => x"82",
           477 => x"81",
           478 => x"80",
           479 => x"81",
           480 => x"82",
           481 => x"81",
           482 => x"80",
           483 => x"81",
           484 => x"82",
           485 => x"81",
           486 => x"80",
           487 => x"81",
           488 => x"82",
           489 => x"81",
           490 => x"81",
           491 => x"81",
           492 => x"82",
           493 => x"81",
           494 => x"81",
           495 => x"81",
           496 => x"82",
           497 => x"81",
           498 => x"81",
           499 => x"81",
           500 => x"82",
           501 => x"81",
           502 => x"80",
           503 => x"81",
           504 => x"82",
           505 => x"81",
           506 => x"81",
           507 => x"81",
           508 => x"82",
           509 => x"81",
           510 => x"81",
           511 => x"81",
           512 => x"82",
           513 => x"81",
           514 => x"80",
           515 => x"81",
           516 => x"82",
           517 => x"81",
           518 => x"80",
           519 => x"81",
           520 => x"82",
           521 => x"81",
           522 => x"80",
           523 => x"81",
           524 => x"82",
           525 => x"81",
           526 => x"80",
           527 => x"81",
           528 => x"82",
           529 => x"81",
           530 => x"81",
           531 => x"81",
           532 => x"82",
           533 => x"81",
           534 => x"81",
           535 => x"81",
           536 => x"82",
           537 => x"81",
           538 => x"81",
           539 => x"81",
           540 => x"82",
           541 => x"81",
           542 => x"80",
           543 => x"81",
           544 => x"82",
           545 => x"81",
           546 => x"81",
           547 => x"81",
           548 => x"82",
           549 => x"81",
           550 => x"b8",
           551 => x"d3",
           552 => x"a0",
           553 => x"d3",
           554 => x"fd",
           555 => x"90",
           556 => x"90",
           557 => x"90",
           558 => x"2d",
           559 => x"08",
           560 => x"04",
           561 => x"0c",
           562 => x"81",
           563 => x"82",
           564 => x"81",
           565 => x"9c",
           566 => x"d3",
           567 => x"a0",
           568 => x"d3",
           569 => x"a0",
           570 => x"90",
           571 => x"90",
           572 => x"90",
           573 => x"9f",
           574 => x"90",
           575 => x"90",
           576 => x"10",
           577 => x"10",
           578 => x"10",
           579 => x"10",
           580 => x"10",
           581 => x"10",
           582 => x"10",
           583 => x"10",
           584 => x"51",
           585 => x"73",
           586 => x"73",
           587 => x"81",
           588 => x"10",
           589 => x"07",
           590 => x"0c",
           591 => x"72",
           592 => x"81",
           593 => x"09",
           594 => x"71",
           595 => x"0a",
           596 => x"72",
           597 => x"51",
           598 => x"81",
           599 => x"81",
           600 => x"8e",
           601 => x"70",
           602 => x"0c",
           603 => x"92",
           604 => x"81",
           605 => x"f3",
           606 => x"d3",
           607 => x"81",
           608 => x"fd",
           609 => x"53",
           610 => x"08",
           611 => x"52",
           612 => x"08",
           613 => x"51",
           614 => x"81",
           615 => x"70",
           616 => x"0c",
           617 => x"0d",
           618 => x"0c",
           619 => x"90",
           620 => x"d3",
           621 => x"3d",
           622 => x"81",
           623 => x"8c",
           624 => x"81",
           625 => x"88",
           626 => x"83",
           627 => x"d3",
           628 => x"81",
           629 => x"54",
           630 => x"81",
           631 => x"04",
           632 => x"08",
           633 => x"90",
           634 => x"0d",
           635 => x"d3",
           636 => x"05",
           637 => x"90",
           638 => x"08",
           639 => x"38",
           640 => x"08",
           641 => x"30",
           642 => x"08",
           643 => x"80",
           644 => x"90",
           645 => x"0c",
           646 => x"08",
           647 => x"8a",
           648 => x"81",
           649 => x"f4",
           650 => x"d3",
           651 => x"05",
           652 => x"90",
           653 => x"0c",
           654 => x"08",
           655 => x"80",
           656 => x"81",
           657 => x"8c",
           658 => x"81",
           659 => x"8c",
           660 => x"0b",
           661 => x"08",
           662 => x"81",
           663 => x"fc",
           664 => x"38",
           665 => x"d3",
           666 => x"05",
           667 => x"90",
           668 => x"08",
           669 => x"08",
           670 => x"80",
           671 => x"90",
           672 => x"08",
           673 => x"90",
           674 => x"08",
           675 => x"3f",
           676 => x"08",
           677 => x"90",
           678 => x"0c",
           679 => x"90",
           680 => x"08",
           681 => x"38",
           682 => x"08",
           683 => x"30",
           684 => x"08",
           685 => x"81",
           686 => x"f8",
           687 => x"81",
           688 => x"54",
           689 => x"81",
           690 => x"04",
           691 => x"08",
           692 => x"90",
           693 => x"0d",
           694 => x"d3",
           695 => x"05",
           696 => x"90",
           697 => x"08",
           698 => x"38",
           699 => x"08",
           700 => x"30",
           701 => x"08",
           702 => x"81",
           703 => x"90",
           704 => x"0c",
           705 => x"08",
           706 => x"80",
           707 => x"81",
           708 => x"8c",
           709 => x"81",
           710 => x"8c",
           711 => x"53",
           712 => x"08",
           713 => x"52",
           714 => x"08",
           715 => x"51",
           716 => x"d3",
           717 => x"81",
           718 => x"f8",
           719 => x"81",
           720 => x"fc",
           721 => x"2e",
           722 => x"d3",
           723 => x"05",
           724 => x"d3",
           725 => x"05",
           726 => x"90",
           727 => x"08",
           728 => x"84",
           729 => x"3d",
           730 => x"90",
           731 => x"d3",
           732 => x"81",
           733 => x"fd",
           734 => x"0b",
           735 => x"08",
           736 => x"80",
           737 => x"90",
           738 => x"0c",
           739 => x"08",
           740 => x"81",
           741 => x"88",
           742 => x"b9",
           743 => x"90",
           744 => x"08",
           745 => x"38",
           746 => x"d3",
           747 => x"05",
           748 => x"38",
           749 => x"08",
           750 => x"10",
           751 => x"08",
           752 => x"81",
           753 => x"fc",
           754 => x"81",
           755 => x"fc",
           756 => x"b8",
           757 => x"90",
           758 => x"08",
           759 => x"e1",
           760 => x"90",
           761 => x"08",
           762 => x"08",
           763 => x"26",
           764 => x"d3",
           765 => x"05",
           766 => x"90",
           767 => x"08",
           768 => x"90",
           769 => x"0c",
           770 => x"08",
           771 => x"81",
           772 => x"fc",
           773 => x"81",
           774 => x"f8",
           775 => x"d3",
           776 => x"05",
           777 => x"81",
           778 => x"fc",
           779 => x"d3",
           780 => x"05",
           781 => x"81",
           782 => x"8c",
           783 => x"95",
           784 => x"90",
           785 => x"08",
           786 => x"38",
           787 => x"08",
           788 => x"70",
           789 => x"08",
           790 => x"51",
           791 => x"d3",
           792 => x"05",
           793 => x"d3",
           794 => x"05",
           795 => x"d3",
           796 => x"05",
           797 => x"84",
           798 => x"0d",
           799 => x"0c",
           800 => x"0d",
           801 => x"02",
           802 => x"05",
           803 => x"53",
           804 => x"27",
           805 => x"83",
           806 => x"80",
           807 => x"ff",
           808 => x"ff",
           809 => x"73",
           810 => x"05",
           811 => x"12",
           812 => x"2e",
           813 => x"ef",
           814 => x"d3",
           815 => x"3d",
           816 => x"74",
           817 => x"07",
           818 => x"2b",
           819 => x"51",
           820 => x"a5",
           821 => x"70",
           822 => x"0c",
           823 => x"84",
           824 => x"72",
           825 => x"05",
           826 => x"71",
           827 => x"53",
           828 => x"52",
           829 => x"dd",
           830 => x"27",
           831 => x"71",
           832 => x"53",
           833 => x"52",
           834 => x"f2",
           835 => x"ff",
           836 => x"3d",
           837 => x"70",
           838 => x"06",
           839 => x"70",
           840 => x"73",
           841 => x"56",
           842 => x"08",
           843 => x"38",
           844 => x"52",
           845 => x"81",
           846 => x"54",
           847 => x"9d",
           848 => x"55",
           849 => x"09",
           850 => x"38",
           851 => x"14",
           852 => x"81",
           853 => x"56",
           854 => x"e5",
           855 => x"55",
           856 => x"06",
           857 => x"06",
           858 => x"81",
           859 => x"52",
           860 => x"0d",
           861 => x"70",
           862 => x"ff",
           863 => x"f8",
           864 => x"80",
           865 => x"51",
           866 => x"84",
           867 => x"71",
           868 => x"54",
           869 => x"2e",
           870 => x"75",
           871 => x"94",
           872 => x"81",
           873 => x"87",
           874 => x"fe",
           875 => x"52",
           876 => x"88",
           877 => x"86",
           878 => x"84",
           879 => x"06",
           880 => x"14",
           881 => x"80",
           882 => x"71",
           883 => x"0c",
           884 => x"04",
           885 => x"77",
           886 => x"53",
           887 => x"80",
           888 => x"38",
           889 => x"70",
           890 => x"81",
           891 => x"81",
           892 => x"39",
           893 => x"39",
           894 => x"80",
           895 => x"81",
           896 => x"55",
           897 => x"2e",
           898 => x"55",
           899 => x"84",
           900 => x"38",
           901 => x"06",
           902 => x"2e",
           903 => x"88",
           904 => x"70",
           905 => x"34",
           906 => x"71",
           907 => x"d3",
           908 => x"3d",
           909 => x"3d",
           910 => x"72",
           911 => x"91",
           912 => x"fc",
           913 => x"51",
           914 => x"81",
           915 => x"85",
           916 => x"83",
           917 => x"72",
           918 => x"0c",
           919 => x"04",
           920 => x"76",
           921 => x"ff",
           922 => x"81",
           923 => x"26",
           924 => x"83",
           925 => x"05",
           926 => x"70",
           927 => x"8a",
           928 => x"33",
           929 => x"70",
           930 => x"fe",
           931 => x"33",
           932 => x"70",
           933 => x"f2",
           934 => x"33",
           935 => x"70",
           936 => x"e6",
           937 => x"22",
           938 => x"74",
           939 => x"80",
           940 => x"13",
           941 => x"52",
           942 => x"26",
           943 => x"81",
           944 => x"98",
           945 => x"22",
           946 => x"bc",
           947 => x"33",
           948 => x"b8",
           949 => x"33",
           950 => x"b4",
           951 => x"33",
           952 => x"b0",
           953 => x"33",
           954 => x"ac",
           955 => x"33",
           956 => x"a8",
           957 => x"c0",
           958 => x"73",
           959 => x"a0",
           960 => x"87",
           961 => x"0c",
           962 => x"81",
           963 => x"86",
           964 => x"f3",
           965 => x"5b",
           966 => x"9c",
           967 => x"0c",
           968 => x"bc",
           969 => x"7b",
           970 => x"98",
           971 => x"79",
           972 => x"87",
           973 => x"08",
           974 => x"1c",
           975 => x"98",
           976 => x"79",
           977 => x"87",
           978 => x"08",
           979 => x"1c",
           980 => x"98",
           981 => x"79",
           982 => x"87",
           983 => x"08",
           984 => x"1c",
           985 => x"98",
           986 => x"79",
           987 => x"80",
           988 => x"83",
           989 => x"59",
           990 => x"ff",
           991 => x"1b",
           992 => x"1b",
           993 => x"1b",
           994 => x"1b",
           995 => x"1b",
           996 => x"83",
           997 => x"52",
           998 => x"51",
           999 => x"8f",
          1000 => x"ff",
          1001 => x"8f",
          1002 => x"30",
          1003 => x"51",
          1004 => x"0b",
          1005 => x"fc",
          1006 => x"0d",
          1007 => x"0d",
          1008 => x"81",
          1009 => x"70",
          1010 => x"57",
          1011 => x"c0",
          1012 => x"74",
          1013 => x"38",
          1014 => x"94",
          1015 => x"70",
          1016 => x"81",
          1017 => x"52",
          1018 => x"8c",
          1019 => x"2a",
          1020 => x"51",
          1021 => x"38",
          1022 => x"70",
          1023 => x"51",
          1024 => x"8d",
          1025 => x"2a",
          1026 => x"51",
          1027 => x"be",
          1028 => x"ff",
          1029 => x"c0",
          1030 => x"70",
          1031 => x"38",
          1032 => x"90",
          1033 => x"0c",
          1034 => x"84",
          1035 => x"0d",
          1036 => x"0d",
          1037 => x"33",
          1038 => x"cf",
          1039 => x"81",
          1040 => x"55",
          1041 => x"94",
          1042 => x"80",
          1043 => x"87",
          1044 => x"51",
          1045 => x"96",
          1046 => x"06",
          1047 => x"70",
          1048 => x"38",
          1049 => x"70",
          1050 => x"51",
          1051 => x"72",
          1052 => x"81",
          1053 => x"70",
          1054 => x"38",
          1055 => x"70",
          1056 => x"51",
          1057 => x"38",
          1058 => x"06",
          1059 => x"94",
          1060 => x"80",
          1061 => x"87",
          1062 => x"52",
          1063 => x"87",
          1064 => x"f9",
          1065 => x"54",
          1066 => x"70",
          1067 => x"53",
          1068 => x"77",
          1069 => x"38",
          1070 => x"06",
          1071 => x"0b",
          1072 => x"33",
          1073 => x"06",
          1074 => x"58",
          1075 => x"84",
          1076 => x"2e",
          1077 => x"c0",
          1078 => x"70",
          1079 => x"2a",
          1080 => x"53",
          1081 => x"80",
          1082 => x"71",
          1083 => x"81",
          1084 => x"70",
          1085 => x"81",
          1086 => x"06",
          1087 => x"80",
          1088 => x"71",
          1089 => x"81",
          1090 => x"70",
          1091 => x"74",
          1092 => x"51",
          1093 => x"80",
          1094 => x"2e",
          1095 => x"c0",
          1096 => x"77",
          1097 => x"17",
          1098 => x"81",
          1099 => x"53",
          1100 => x"84",
          1101 => x"d3",
          1102 => x"3d",
          1103 => x"3d",
          1104 => x"81",
          1105 => x"70",
          1106 => x"54",
          1107 => x"94",
          1108 => x"80",
          1109 => x"87",
          1110 => x"51",
          1111 => x"82",
          1112 => x"06",
          1113 => x"70",
          1114 => x"38",
          1115 => x"06",
          1116 => x"94",
          1117 => x"80",
          1118 => x"87",
          1119 => x"52",
          1120 => x"81",
          1121 => x"d3",
          1122 => x"84",
          1123 => x"fe",
          1124 => x"0b",
          1125 => x"33",
          1126 => x"06",
          1127 => x"c0",
          1128 => x"70",
          1129 => x"38",
          1130 => x"94",
          1131 => x"70",
          1132 => x"81",
          1133 => x"51",
          1134 => x"80",
          1135 => x"72",
          1136 => x"51",
          1137 => x"80",
          1138 => x"2e",
          1139 => x"c0",
          1140 => x"71",
          1141 => x"2b",
          1142 => x"51",
          1143 => x"81",
          1144 => x"84",
          1145 => x"ff",
          1146 => x"c0",
          1147 => x"70",
          1148 => x"06",
          1149 => x"80",
          1150 => x"38",
          1151 => x"9c",
          1152 => x"80",
          1153 => x"9e",
          1154 => x"d0",
          1155 => x"c0",
          1156 => x"81",
          1157 => x"87",
          1158 => x"08",
          1159 => x"0c",
          1160 => x"94",
          1161 => x"90",
          1162 => x"9e",
          1163 => x"d0",
          1164 => x"c0",
          1165 => x"81",
          1166 => x"87",
          1167 => x"08",
          1168 => x"0c",
          1169 => x"ac",
          1170 => x"a0",
          1171 => x"9e",
          1172 => x"70",
          1173 => x"23",
          1174 => x"84",
          1175 => x"a8",
          1176 => x"81",
          1177 => x"80",
          1178 => x"9e",
          1179 => x"a0",
          1180 => x"52",
          1181 => x"2e",
          1182 => x"52",
          1183 => x"ad",
          1184 => x"87",
          1185 => x"08",
          1186 => x"80",
          1187 => x"52",
          1188 => x"83",
          1189 => x"71",
          1190 => x"34",
          1191 => x"c0",
          1192 => x"70",
          1193 => x"06",
          1194 => x"70",
          1195 => x"38",
          1196 => x"81",
          1197 => x"80",
          1198 => x"9e",
          1199 => x"90",
          1200 => x"52",
          1201 => x"2e",
          1202 => x"52",
          1203 => x"b0",
          1204 => x"87",
          1205 => x"08",
          1206 => x"06",
          1207 => x"70",
          1208 => x"38",
          1209 => x"81",
          1210 => x"80",
          1211 => x"9e",
          1212 => x"84",
          1213 => x"52",
          1214 => x"2e",
          1215 => x"52",
          1216 => x"b2",
          1217 => x"87",
          1218 => x"08",
          1219 => x"06",
          1220 => x"70",
          1221 => x"38",
          1222 => x"81",
          1223 => x"80",
          1224 => x"9e",
          1225 => x"81",
          1226 => x"52",
          1227 => x"2e",
          1228 => x"52",
          1229 => x"b4",
          1230 => x"9e",
          1231 => x"80",
          1232 => x"86",
          1233 => x"51",
          1234 => x"b5",
          1235 => x"87",
          1236 => x"08",
          1237 => x"51",
          1238 => x"80",
          1239 => x"81",
          1240 => x"d0",
          1241 => x"0b",
          1242 => x"88",
          1243 => x"06",
          1244 => x"70",
          1245 => x"38",
          1246 => x"81",
          1247 => x"87",
          1248 => x"08",
          1249 => x"51",
          1250 => x"d0",
          1251 => x"3d",
          1252 => x"3d",
          1253 => x"e8",
          1254 => x"3f",
          1255 => x"33",
          1256 => x"2e",
          1257 => x"bd",
          1258 => x"90",
          1259 => x"90",
          1260 => x"3f",
          1261 => x"33",
          1262 => x"2e",
          1263 => x"d0",
          1264 => x"81",
          1265 => x"52",
          1266 => x"51",
          1267 => x"81",
          1268 => x"54",
          1269 => x"92",
          1270 => x"8c",
          1271 => x"d0",
          1272 => x"81",
          1273 => x"89",
          1274 => x"d0",
          1275 => x"73",
          1276 => x"d0",
          1277 => x"73",
          1278 => x"38",
          1279 => x"08",
          1280 => x"90",
          1281 => x"be",
          1282 => x"94",
          1283 => x"b1",
          1284 => x"80",
          1285 => x"81",
          1286 => x"83",
          1287 => x"d0",
          1288 => x"73",
          1289 => x"38",
          1290 => x"51",
          1291 => x"81",
          1292 => x"54",
          1293 => x"88",
          1294 => x"b0",
          1295 => x"3f",
          1296 => x"33",
          1297 => x"2e",
          1298 => x"d0",
          1299 => x"81",
          1300 => x"88",
          1301 => x"d0",
          1302 => x"73",
          1303 => x"38",
          1304 => x"51",
          1305 => x"81",
          1306 => x"54",
          1307 => x"8d",
          1308 => x"b8",
          1309 => x"bf",
          1310 => x"a4",
          1311 => x"94",
          1312 => x"3f",
          1313 => x"08",
          1314 => x"a0",
          1315 => x"3f",
          1316 => x"08",
          1317 => x"c8",
          1318 => x"3f",
          1319 => x"08",
          1320 => x"f0",
          1321 => x"3f",
          1322 => x"22",
          1323 => x"98",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"c0",
          1327 => x"3f",
          1328 => x"04",
          1329 => x"02",
          1330 => x"ff",
          1331 => x"84",
          1332 => x"71",
          1333 => x"bc",
          1334 => x"71",
          1335 => x"c1",
          1336 => x"39",
          1337 => x"51",
          1338 => x"c1",
          1339 => x"39",
          1340 => x"51",
          1341 => x"c2",
          1342 => x"39",
          1343 => x"51",
          1344 => x"84",
          1345 => x"71",
          1346 => x"04",
          1347 => x"c0",
          1348 => x"04",
          1349 => x"87",
          1350 => x"70",
          1351 => x"80",
          1352 => x"74",
          1353 => x"d0",
          1354 => x"0c",
          1355 => x"04",
          1356 => x"87",
          1357 => x"70",
          1358 => x"bc",
          1359 => x"72",
          1360 => x"70",
          1361 => x"08",
          1362 => x"d0",
          1363 => x"0c",
          1364 => x"0d",
          1365 => x"bc",
          1366 => x"96",
          1367 => x"fe",
          1368 => x"93",
          1369 => x"72",
          1370 => x"81",
          1371 => x"8d",
          1372 => x"81",
          1373 => x"52",
          1374 => x"90",
          1375 => x"34",
          1376 => x"08",
          1377 => x"d3",
          1378 => x"39",
          1379 => x"08",
          1380 => x"2e",
          1381 => x"51",
          1382 => x"3d",
          1383 => x"3d",
          1384 => x"05",
          1385 => x"94",
          1386 => x"d3",
          1387 => x"51",
          1388 => x"72",
          1389 => x"0c",
          1390 => x"04",
          1391 => x"75",
          1392 => x"70",
          1393 => x"53",
          1394 => x"2e",
          1395 => x"81",
          1396 => x"81",
          1397 => x"87",
          1398 => x"85",
          1399 => x"fc",
          1400 => x"81",
          1401 => x"78",
          1402 => x"0c",
          1403 => x"33",
          1404 => x"06",
          1405 => x"80",
          1406 => x"72",
          1407 => x"51",
          1408 => x"fe",
          1409 => x"39",
          1410 => x"94",
          1411 => x"0d",
          1412 => x"0d",
          1413 => x"59",
          1414 => x"05",
          1415 => x"75",
          1416 => x"f8",
          1417 => x"2e",
          1418 => x"82",
          1419 => x"70",
          1420 => x"05",
          1421 => x"5b",
          1422 => x"2e",
          1423 => x"85",
          1424 => x"8b",
          1425 => x"2e",
          1426 => x"8a",
          1427 => x"78",
          1428 => x"5a",
          1429 => x"aa",
          1430 => x"06",
          1431 => x"84",
          1432 => x"7b",
          1433 => x"5d",
          1434 => x"59",
          1435 => x"d0",
          1436 => x"89",
          1437 => x"7a",
          1438 => x"10",
          1439 => x"d0",
          1440 => x"81",
          1441 => x"57",
          1442 => x"75",
          1443 => x"70",
          1444 => x"07",
          1445 => x"80",
          1446 => x"30",
          1447 => x"80",
          1448 => x"53",
          1449 => x"55",
          1450 => x"2e",
          1451 => x"84",
          1452 => x"81",
          1453 => x"57",
          1454 => x"2e",
          1455 => x"75",
          1456 => x"76",
          1457 => x"e0",
          1458 => x"ff",
          1459 => x"73",
          1460 => x"81",
          1461 => x"80",
          1462 => x"38",
          1463 => x"2e",
          1464 => x"73",
          1465 => x"8b",
          1466 => x"c2",
          1467 => x"38",
          1468 => x"73",
          1469 => x"81",
          1470 => x"8f",
          1471 => x"d5",
          1472 => x"38",
          1473 => x"24",
          1474 => x"80",
          1475 => x"38",
          1476 => x"73",
          1477 => x"80",
          1478 => x"ef",
          1479 => x"19",
          1480 => x"59",
          1481 => x"33",
          1482 => x"75",
          1483 => x"81",
          1484 => x"70",
          1485 => x"55",
          1486 => x"79",
          1487 => x"90",
          1488 => x"16",
          1489 => x"7b",
          1490 => x"a0",
          1491 => x"3f",
          1492 => x"53",
          1493 => x"e9",
          1494 => x"fc",
          1495 => x"81",
          1496 => x"72",
          1497 => x"b0",
          1498 => x"fb",
          1499 => x"39",
          1500 => x"83",
          1501 => x"59",
          1502 => x"82",
          1503 => x"88",
          1504 => x"8a",
          1505 => x"90",
          1506 => x"75",
          1507 => x"3f",
          1508 => x"79",
          1509 => x"81",
          1510 => x"72",
          1511 => x"38",
          1512 => x"59",
          1513 => x"84",
          1514 => x"58",
          1515 => x"80",
          1516 => x"30",
          1517 => x"80",
          1518 => x"55",
          1519 => x"25",
          1520 => x"80",
          1521 => x"74",
          1522 => x"07",
          1523 => x"0b",
          1524 => x"57",
          1525 => x"51",
          1526 => x"81",
          1527 => x"81",
          1528 => x"53",
          1529 => x"e3",
          1530 => x"d3",
          1531 => x"89",
          1532 => x"38",
          1533 => x"75",
          1534 => x"84",
          1535 => x"53",
          1536 => x"06",
          1537 => x"53",
          1538 => x"81",
          1539 => x"81",
          1540 => x"70",
          1541 => x"2a",
          1542 => x"76",
          1543 => x"38",
          1544 => x"38",
          1545 => x"70",
          1546 => x"53",
          1547 => x"8e",
          1548 => x"77",
          1549 => x"53",
          1550 => x"81",
          1551 => x"7a",
          1552 => x"55",
          1553 => x"83",
          1554 => x"79",
          1555 => x"81",
          1556 => x"72",
          1557 => x"17",
          1558 => x"27",
          1559 => x"51",
          1560 => x"75",
          1561 => x"72",
          1562 => x"81",
          1563 => x"7a",
          1564 => x"38",
          1565 => x"05",
          1566 => x"ff",
          1567 => x"70",
          1568 => x"57",
          1569 => x"76",
          1570 => x"81",
          1571 => x"72",
          1572 => x"84",
          1573 => x"f9",
          1574 => x"39",
          1575 => x"04",
          1576 => x"86",
          1577 => x"84",
          1578 => x"55",
          1579 => x"fa",
          1580 => x"3d",
          1581 => x"3d",
          1582 => x"d3",
          1583 => x"3d",
          1584 => x"75",
          1585 => x"3f",
          1586 => x"08",
          1587 => x"34",
          1588 => x"d3",
          1589 => x"3d",
          1590 => x"3d",
          1591 => x"94",
          1592 => x"d3",
          1593 => x"3d",
          1594 => x"77",
          1595 => x"a1",
          1596 => x"d3",
          1597 => x"3d",
          1598 => x"3d",
          1599 => x"81",
          1600 => x"70",
          1601 => x"55",
          1602 => x"80",
          1603 => x"38",
          1604 => x"08",
          1605 => x"81",
          1606 => x"81",
          1607 => x"72",
          1608 => x"cb",
          1609 => x"2e",
          1610 => x"88",
          1611 => x"70",
          1612 => x"51",
          1613 => x"2e",
          1614 => x"80",
          1615 => x"ff",
          1616 => x"39",
          1617 => x"c8",
          1618 => x"52",
          1619 => x"c0",
          1620 => x"52",
          1621 => x"81",
          1622 => x"51",
          1623 => x"ff",
          1624 => x"15",
          1625 => x"34",
          1626 => x"f3",
          1627 => x"72",
          1628 => x"0c",
          1629 => x"04",
          1630 => x"81",
          1631 => x"75",
          1632 => x"0c",
          1633 => x"52",
          1634 => x"3f",
          1635 => x"98",
          1636 => x"0d",
          1637 => x"0d",
          1638 => x"56",
          1639 => x"0c",
          1640 => x"70",
          1641 => x"73",
          1642 => x"81",
          1643 => x"81",
          1644 => x"ed",
          1645 => x"2e",
          1646 => x"8e",
          1647 => x"08",
          1648 => x"76",
          1649 => x"56",
          1650 => x"b0",
          1651 => x"06",
          1652 => x"75",
          1653 => x"76",
          1654 => x"70",
          1655 => x"73",
          1656 => x"8b",
          1657 => x"73",
          1658 => x"85",
          1659 => x"82",
          1660 => x"76",
          1661 => x"70",
          1662 => x"ac",
          1663 => x"a0",
          1664 => x"fa",
          1665 => x"53",
          1666 => x"57",
          1667 => x"98",
          1668 => x"39",
          1669 => x"80",
          1670 => x"26",
          1671 => x"86",
          1672 => x"80",
          1673 => x"57",
          1674 => x"74",
          1675 => x"38",
          1676 => x"27",
          1677 => x"14",
          1678 => x"06",
          1679 => x"14",
          1680 => x"06",
          1681 => x"74",
          1682 => x"f9",
          1683 => x"ff",
          1684 => x"89",
          1685 => x"38",
          1686 => x"c5",
          1687 => x"29",
          1688 => x"81",
          1689 => x"76",
          1690 => x"56",
          1691 => x"ba",
          1692 => x"2e",
          1693 => x"30",
          1694 => x"0c",
          1695 => x"81",
          1696 => x"8a",
          1697 => x"f8",
          1698 => x"7c",
          1699 => x"70",
          1700 => x"75",
          1701 => x"55",
          1702 => x"2e",
          1703 => x"87",
          1704 => x"76",
          1705 => x"73",
          1706 => x"81",
          1707 => x"81",
          1708 => x"77",
          1709 => x"70",
          1710 => x"58",
          1711 => x"09",
          1712 => x"c2",
          1713 => x"81",
          1714 => x"75",
          1715 => x"55",
          1716 => x"e2",
          1717 => x"90",
          1718 => x"f8",
          1719 => x"8f",
          1720 => x"81",
          1721 => x"75",
          1722 => x"55",
          1723 => x"81",
          1724 => x"27",
          1725 => x"d0",
          1726 => x"55",
          1727 => x"73",
          1728 => x"80",
          1729 => x"14",
          1730 => x"72",
          1731 => x"e0",
          1732 => x"80",
          1733 => x"39",
          1734 => x"55",
          1735 => x"80",
          1736 => x"e0",
          1737 => x"38",
          1738 => x"81",
          1739 => x"53",
          1740 => x"81",
          1741 => x"53",
          1742 => x"8e",
          1743 => x"70",
          1744 => x"55",
          1745 => x"27",
          1746 => x"77",
          1747 => x"74",
          1748 => x"76",
          1749 => x"77",
          1750 => x"70",
          1751 => x"55",
          1752 => x"77",
          1753 => x"38",
          1754 => x"74",
          1755 => x"55",
          1756 => x"84",
          1757 => x"0d",
          1758 => x"0d",
          1759 => x"33",
          1760 => x"70",
          1761 => x"38",
          1762 => x"11",
          1763 => x"81",
          1764 => x"83",
          1765 => x"fc",
          1766 => x"9b",
          1767 => x"84",
          1768 => x"33",
          1769 => x"51",
          1770 => x"80",
          1771 => x"84",
          1772 => x"92",
          1773 => x"51",
          1774 => x"80",
          1775 => x"81",
          1776 => x"72",
          1777 => x"92",
          1778 => x"81",
          1779 => x"0b",
          1780 => x"8c",
          1781 => x"71",
          1782 => x"06",
          1783 => x"80",
          1784 => x"87",
          1785 => x"08",
          1786 => x"38",
          1787 => x"80",
          1788 => x"71",
          1789 => x"c0",
          1790 => x"51",
          1791 => x"87",
          1792 => x"d0",
          1793 => x"81",
          1794 => x"33",
          1795 => x"d3",
          1796 => x"3d",
          1797 => x"3d",
          1798 => x"64",
          1799 => x"bf",
          1800 => x"40",
          1801 => x"74",
          1802 => x"cd",
          1803 => x"84",
          1804 => x"7a",
          1805 => x"81",
          1806 => x"72",
          1807 => x"87",
          1808 => x"11",
          1809 => x"8c",
          1810 => x"92",
          1811 => x"5a",
          1812 => x"58",
          1813 => x"c0",
          1814 => x"76",
          1815 => x"76",
          1816 => x"70",
          1817 => x"81",
          1818 => x"54",
          1819 => x"8e",
          1820 => x"52",
          1821 => x"81",
          1822 => x"81",
          1823 => x"74",
          1824 => x"53",
          1825 => x"83",
          1826 => x"78",
          1827 => x"8f",
          1828 => x"2e",
          1829 => x"c0",
          1830 => x"52",
          1831 => x"87",
          1832 => x"08",
          1833 => x"2e",
          1834 => x"84",
          1835 => x"38",
          1836 => x"87",
          1837 => x"15",
          1838 => x"70",
          1839 => x"52",
          1840 => x"ff",
          1841 => x"39",
          1842 => x"81",
          1843 => x"ff",
          1844 => x"57",
          1845 => x"90",
          1846 => x"80",
          1847 => x"71",
          1848 => x"78",
          1849 => x"38",
          1850 => x"80",
          1851 => x"80",
          1852 => x"81",
          1853 => x"72",
          1854 => x"0c",
          1855 => x"04",
          1856 => x"60",
          1857 => x"8c",
          1858 => x"33",
          1859 => x"5b",
          1860 => x"74",
          1861 => x"e1",
          1862 => x"84",
          1863 => x"79",
          1864 => x"78",
          1865 => x"06",
          1866 => x"77",
          1867 => x"87",
          1868 => x"11",
          1869 => x"8c",
          1870 => x"92",
          1871 => x"59",
          1872 => x"85",
          1873 => x"98",
          1874 => x"7d",
          1875 => x"0c",
          1876 => x"08",
          1877 => x"70",
          1878 => x"53",
          1879 => x"2e",
          1880 => x"70",
          1881 => x"33",
          1882 => x"18",
          1883 => x"2a",
          1884 => x"51",
          1885 => x"2e",
          1886 => x"c0",
          1887 => x"52",
          1888 => x"87",
          1889 => x"08",
          1890 => x"2e",
          1891 => x"84",
          1892 => x"38",
          1893 => x"87",
          1894 => x"15",
          1895 => x"70",
          1896 => x"52",
          1897 => x"ff",
          1898 => x"39",
          1899 => x"81",
          1900 => x"80",
          1901 => x"52",
          1902 => x"90",
          1903 => x"80",
          1904 => x"71",
          1905 => x"7a",
          1906 => x"38",
          1907 => x"80",
          1908 => x"80",
          1909 => x"81",
          1910 => x"72",
          1911 => x"0c",
          1912 => x"04",
          1913 => x"7e",
          1914 => x"b3",
          1915 => x"88",
          1916 => x"33",
          1917 => x"56",
          1918 => x"3f",
          1919 => x"08",
          1920 => x"83",
          1921 => x"fe",
          1922 => x"87",
          1923 => x"0c",
          1924 => x"76",
          1925 => x"38",
          1926 => x"93",
          1927 => x"2b",
          1928 => x"8c",
          1929 => x"71",
          1930 => x"38",
          1931 => x"71",
          1932 => x"c6",
          1933 => x"39",
          1934 => x"81",
          1935 => x"06",
          1936 => x"71",
          1937 => x"38",
          1938 => x"8c",
          1939 => x"e8",
          1940 => x"98",
          1941 => x"71",
          1942 => x"73",
          1943 => x"92",
          1944 => x"72",
          1945 => x"06",
          1946 => x"f7",
          1947 => x"80",
          1948 => x"88",
          1949 => x"0c",
          1950 => x"80",
          1951 => x"56",
          1952 => x"56",
          1953 => x"81",
          1954 => x"8c",
          1955 => x"fe",
          1956 => x"81",
          1957 => x"33",
          1958 => x"07",
          1959 => x"0c",
          1960 => x"3d",
          1961 => x"3d",
          1962 => x"11",
          1963 => x"33",
          1964 => x"71",
          1965 => x"81",
          1966 => x"72",
          1967 => x"75",
          1968 => x"81",
          1969 => x"52",
          1970 => x"54",
          1971 => x"0d",
          1972 => x"0d",
          1973 => x"05",
          1974 => x"52",
          1975 => x"70",
          1976 => x"34",
          1977 => x"51",
          1978 => x"83",
          1979 => x"ff",
          1980 => x"75",
          1981 => x"72",
          1982 => x"54",
          1983 => x"2a",
          1984 => x"70",
          1985 => x"34",
          1986 => x"51",
          1987 => x"81",
          1988 => x"70",
          1989 => x"70",
          1990 => x"3d",
          1991 => x"3d",
          1992 => x"77",
          1993 => x"70",
          1994 => x"38",
          1995 => x"05",
          1996 => x"70",
          1997 => x"34",
          1998 => x"eb",
          1999 => x"0d",
          2000 => x"0d",
          2001 => x"54",
          2002 => x"72",
          2003 => x"54",
          2004 => x"51",
          2005 => x"84",
          2006 => x"fc",
          2007 => x"77",
          2008 => x"53",
          2009 => x"05",
          2010 => x"70",
          2011 => x"33",
          2012 => x"ff",
          2013 => x"52",
          2014 => x"2e",
          2015 => x"80",
          2016 => x"71",
          2017 => x"0c",
          2018 => x"04",
          2019 => x"74",
          2020 => x"89",
          2021 => x"2e",
          2022 => x"11",
          2023 => x"52",
          2024 => x"70",
          2025 => x"84",
          2026 => x"0d",
          2027 => x"81",
          2028 => x"04",
          2029 => x"d3",
          2030 => x"f7",
          2031 => x"56",
          2032 => x"17",
          2033 => x"74",
          2034 => x"d6",
          2035 => x"b0",
          2036 => x"b4",
          2037 => x"81",
          2038 => x"59",
          2039 => x"81",
          2040 => x"7a",
          2041 => x"06",
          2042 => x"d3",
          2043 => x"17",
          2044 => x"08",
          2045 => x"08",
          2046 => x"08",
          2047 => x"74",
          2048 => x"38",
          2049 => x"55",
          2050 => x"09",
          2051 => x"38",
          2052 => x"18",
          2053 => x"81",
          2054 => x"f9",
          2055 => x"39",
          2056 => x"81",
          2057 => x"8b",
          2058 => x"fa",
          2059 => x"7a",
          2060 => x"57",
          2061 => x"08",
          2062 => x"75",
          2063 => x"3f",
          2064 => x"08",
          2065 => x"84",
          2066 => x"81",
          2067 => x"b4",
          2068 => x"16",
          2069 => x"be",
          2070 => x"84",
          2071 => x"85",
          2072 => x"81",
          2073 => x"17",
          2074 => x"d3",
          2075 => x"3d",
          2076 => x"3d",
          2077 => x"52",
          2078 => x"3f",
          2079 => x"08",
          2080 => x"84",
          2081 => x"38",
          2082 => x"74",
          2083 => x"81",
          2084 => x"38",
          2085 => x"59",
          2086 => x"09",
          2087 => x"e3",
          2088 => x"53",
          2089 => x"08",
          2090 => x"70",
          2091 => x"91",
          2092 => x"d5",
          2093 => x"17",
          2094 => x"3f",
          2095 => x"a4",
          2096 => x"51",
          2097 => x"86",
          2098 => x"f2",
          2099 => x"17",
          2100 => x"3f",
          2101 => x"52",
          2102 => x"51",
          2103 => x"8c",
          2104 => x"84",
          2105 => x"fc",
          2106 => x"17",
          2107 => x"70",
          2108 => x"79",
          2109 => x"52",
          2110 => x"51",
          2111 => x"77",
          2112 => x"80",
          2113 => x"81",
          2114 => x"f9",
          2115 => x"d3",
          2116 => x"2e",
          2117 => x"58",
          2118 => x"84",
          2119 => x"0d",
          2120 => x"0d",
          2121 => x"98",
          2122 => x"05",
          2123 => x"80",
          2124 => x"27",
          2125 => x"14",
          2126 => x"29",
          2127 => x"05",
          2128 => x"81",
          2129 => x"87",
          2130 => x"f9",
          2131 => x"7a",
          2132 => x"54",
          2133 => x"27",
          2134 => x"76",
          2135 => x"27",
          2136 => x"ff",
          2137 => x"58",
          2138 => x"80",
          2139 => x"82",
          2140 => x"72",
          2141 => x"38",
          2142 => x"72",
          2143 => x"8e",
          2144 => x"39",
          2145 => x"17",
          2146 => x"a4",
          2147 => x"53",
          2148 => x"fd",
          2149 => x"d3",
          2150 => x"9f",
          2151 => x"ff",
          2152 => x"11",
          2153 => x"70",
          2154 => x"18",
          2155 => x"76",
          2156 => x"53",
          2157 => x"81",
          2158 => x"80",
          2159 => x"83",
          2160 => x"b4",
          2161 => x"88",
          2162 => x"79",
          2163 => x"84",
          2164 => x"58",
          2165 => x"80",
          2166 => x"9f",
          2167 => x"80",
          2168 => x"88",
          2169 => x"08",
          2170 => x"51",
          2171 => x"81",
          2172 => x"80",
          2173 => x"10",
          2174 => x"74",
          2175 => x"51",
          2176 => x"81",
          2177 => x"83",
          2178 => x"58",
          2179 => x"87",
          2180 => x"08",
          2181 => x"51",
          2182 => x"81",
          2183 => x"9b",
          2184 => x"2b",
          2185 => x"74",
          2186 => x"51",
          2187 => x"81",
          2188 => x"f0",
          2189 => x"83",
          2190 => x"77",
          2191 => x"0c",
          2192 => x"04",
          2193 => x"7a",
          2194 => x"58",
          2195 => x"81",
          2196 => x"9e",
          2197 => x"17",
          2198 => x"96",
          2199 => x"53",
          2200 => x"81",
          2201 => x"79",
          2202 => x"72",
          2203 => x"38",
          2204 => x"72",
          2205 => x"b8",
          2206 => x"39",
          2207 => x"17",
          2208 => x"a4",
          2209 => x"53",
          2210 => x"fb",
          2211 => x"d3",
          2212 => x"81",
          2213 => x"81",
          2214 => x"83",
          2215 => x"b4",
          2216 => x"78",
          2217 => x"56",
          2218 => x"76",
          2219 => x"38",
          2220 => x"9f",
          2221 => x"33",
          2222 => x"07",
          2223 => x"74",
          2224 => x"83",
          2225 => x"89",
          2226 => x"08",
          2227 => x"51",
          2228 => x"81",
          2229 => x"59",
          2230 => x"08",
          2231 => x"74",
          2232 => x"16",
          2233 => x"84",
          2234 => x"76",
          2235 => x"88",
          2236 => x"81",
          2237 => x"8f",
          2238 => x"53",
          2239 => x"80",
          2240 => x"88",
          2241 => x"08",
          2242 => x"51",
          2243 => x"81",
          2244 => x"59",
          2245 => x"08",
          2246 => x"77",
          2247 => x"06",
          2248 => x"83",
          2249 => x"05",
          2250 => x"f7",
          2251 => x"39",
          2252 => x"a4",
          2253 => x"52",
          2254 => x"ef",
          2255 => x"84",
          2256 => x"d3",
          2257 => x"38",
          2258 => x"06",
          2259 => x"83",
          2260 => x"18",
          2261 => x"54",
          2262 => x"f6",
          2263 => x"d3",
          2264 => x"0a",
          2265 => x"52",
          2266 => x"83",
          2267 => x"83",
          2268 => x"81",
          2269 => x"8a",
          2270 => x"f8",
          2271 => x"7c",
          2272 => x"59",
          2273 => x"81",
          2274 => x"38",
          2275 => x"08",
          2276 => x"73",
          2277 => x"38",
          2278 => x"52",
          2279 => x"a4",
          2280 => x"84",
          2281 => x"d3",
          2282 => x"f2",
          2283 => x"82",
          2284 => x"39",
          2285 => x"e6",
          2286 => x"84",
          2287 => x"de",
          2288 => x"78",
          2289 => x"3f",
          2290 => x"08",
          2291 => x"84",
          2292 => x"80",
          2293 => x"d3",
          2294 => x"2e",
          2295 => x"d3",
          2296 => x"2e",
          2297 => x"53",
          2298 => x"51",
          2299 => x"81",
          2300 => x"c5",
          2301 => x"08",
          2302 => x"18",
          2303 => x"57",
          2304 => x"90",
          2305 => x"90",
          2306 => x"16",
          2307 => x"54",
          2308 => x"34",
          2309 => x"78",
          2310 => x"38",
          2311 => x"81",
          2312 => x"8a",
          2313 => x"f6",
          2314 => x"7e",
          2315 => x"5b",
          2316 => x"38",
          2317 => x"58",
          2318 => x"88",
          2319 => x"08",
          2320 => x"38",
          2321 => x"39",
          2322 => x"51",
          2323 => x"81",
          2324 => x"d3",
          2325 => x"82",
          2326 => x"d3",
          2327 => x"81",
          2328 => x"ff",
          2329 => x"38",
          2330 => x"81",
          2331 => x"26",
          2332 => x"79",
          2333 => x"08",
          2334 => x"73",
          2335 => x"b9",
          2336 => x"2e",
          2337 => x"80",
          2338 => x"1a",
          2339 => x"08",
          2340 => x"38",
          2341 => x"52",
          2342 => x"af",
          2343 => x"81",
          2344 => x"81",
          2345 => x"06",
          2346 => x"d3",
          2347 => x"81",
          2348 => x"09",
          2349 => x"72",
          2350 => x"70",
          2351 => x"d3",
          2352 => x"51",
          2353 => x"73",
          2354 => x"81",
          2355 => x"80",
          2356 => x"8c",
          2357 => x"81",
          2358 => x"38",
          2359 => x"08",
          2360 => x"73",
          2361 => x"75",
          2362 => x"77",
          2363 => x"56",
          2364 => x"76",
          2365 => x"82",
          2366 => x"26",
          2367 => x"75",
          2368 => x"f8",
          2369 => x"d3",
          2370 => x"2e",
          2371 => x"59",
          2372 => x"08",
          2373 => x"81",
          2374 => x"81",
          2375 => x"59",
          2376 => x"08",
          2377 => x"70",
          2378 => x"25",
          2379 => x"51",
          2380 => x"73",
          2381 => x"75",
          2382 => x"81",
          2383 => x"38",
          2384 => x"f5",
          2385 => x"75",
          2386 => x"f9",
          2387 => x"d3",
          2388 => x"d3",
          2389 => x"70",
          2390 => x"08",
          2391 => x"51",
          2392 => x"80",
          2393 => x"73",
          2394 => x"38",
          2395 => x"52",
          2396 => x"d0",
          2397 => x"84",
          2398 => x"a5",
          2399 => x"18",
          2400 => x"08",
          2401 => x"18",
          2402 => x"74",
          2403 => x"38",
          2404 => x"18",
          2405 => x"33",
          2406 => x"73",
          2407 => x"97",
          2408 => x"74",
          2409 => x"38",
          2410 => x"55",
          2411 => x"d3",
          2412 => x"85",
          2413 => x"75",
          2414 => x"d3",
          2415 => x"3d",
          2416 => x"3d",
          2417 => x"52",
          2418 => x"3f",
          2419 => x"08",
          2420 => x"81",
          2421 => x"80",
          2422 => x"52",
          2423 => x"c1",
          2424 => x"84",
          2425 => x"84",
          2426 => x"0c",
          2427 => x"53",
          2428 => x"15",
          2429 => x"f2",
          2430 => x"56",
          2431 => x"16",
          2432 => x"22",
          2433 => x"27",
          2434 => x"54",
          2435 => x"76",
          2436 => x"33",
          2437 => x"3f",
          2438 => x"08",
          2439 => x"38",
          2440 => x"76",
          2441 => x"70",
          2442 => x"9f",
          2443 => x"56",
          2444 => x"d3",
          2445 => x"3d",
          2446 => x"3d",
          2447 => x"71",
          2448 => x"57",
          2449 => x"0a",
          2450 => x"38",
          2451 => x"53",
          2452 => x"38",
          2453 => x"0c",
          2454 => x"54",
          2455 => x"75",
          2456 => x"73",
          2457 => x"a8",
          2458 => x"73",
          2459 => x"85",
          2460 => x"0b",
          2461 => x"5a",
          2462 => x"27",
          2463 => x"a8",
          2464 => x"18",
          2465 => x"39",
          2466 => x"70",
          2467 => x"58",
          2468 => x"b2",
          2469 => x"76",
          2470 => x"3f",
          2471 => x"08",
          2472 => x"84",
          2473 => x"bd",
          2474 => x"81",
          2475 => x"27",
          2476 => x"16",
          2477 => x"84",
          2478 => x"38",
          2479 => x"39",
          2480 => x"55",
          2481 => x"52",
          2482 => x"d5",
          2483 => x"84",
          2484 => x"0c",
          2485 => x"0c",
          2486 => x"53",
          2487 => x"80",
          2488 => x"85",
          2489 => x"94",
          2490 => x"2a",
          2491 => x"0c",
          2492 => x"06",
          2493 => x"9c",
          2494 => x"58",
          2495 => x"84",
          2496 => x"0d",
          2497 => x"0d",
          2498 => x"90",
          2499 => x"05",
          2500 => x"f0",
          2501 => x"27",
          2502 => x"0b",
          2503 => x"98",
          2504 => x"84",
          2505 => x"2e",
          2506 => x"76",
          2507 => x"58",
          2508 => x"38",
          2509 => x"15",
          2510 => x"08",
          2511 => x"38",
          2512 => x"88",
          2513 => x"53",
          2514 => x"81",
          2515 => x"c0",
          2516 => x"22",
          2517 => x"89",
          2518 => x"72",
          2519 => x"74",
          2520 => x"f3",
          2521 => x"d3",
          2522 => x"82",
          2523 => x"81",
          2524 => x"27",
          2525 => x"81",
          2526 => x"84",
          2527 => x"80",
          2528 => x"16",
          2529 => x"84",
          2530 => x"ca",
          2531 => x"38",
          2532 => x"0c",
          2533 => x"dd",
          2534 => x"08",
          2535 => x"f9",
          2536 => x"d3",
          2537 => x"87",
          2538 => x"84",
          2539 => x"80",
          2540 => x"55",
          2541 => x"08",
          2542 => x"38",
          2543 => x"d3",
          2544 => x"2e",
          2545 => x"d3",
          2546 => x"75",
          2547 => x"3f",
          2548 => x"08",
          2549 => x"94",
          2550 => x"52",
          2551 => x"c1",
          2552 => x"84",
          2553 => x"0c",
          2554 => x"0c",
          2555 => x"05",
          2556 => x"80",
          2557 => x"d3",
          2558 => x"3d",
          2559 => x"3d",
          2560 => x"71",
          2561 => x"57",
          2562 => x"51",
          2563 => x"81",
          2564 => x"54",
          2565 => x"08",
          2566 => x"81",
          2567 => x"56",
          2568 => x"52",
          2569 => x"83",
          2570 => x"84",
          2571 => x"d3",
          2572 => x"d2",
          2573 => x"84",
          2574 => x"08",
          2575 => x"54",
          2576 => x"e5",
          2577 => x"06",
          2578 => x"58",
          2579 => x"08",
          2580 => x"38",
          2581 => x"75",
          2582 => x"80",
          2583 => x"81",
          2584 => x"7a",
          2585 => x"06",
          2586 => x"39",
          2587 => x"08",
          2588 => x"76",
          2589 => x"3f",
          2590 => x"08",
          2591 => x"84",
          2592 => x"ff",
          2593 => x"84",
          2594 => x"06",
          2595 => x"54",
          2596 => x"84",
          2597 => x"0d",
          2598 => x"0d",
          2599 => x"52",
          2600 => x"3f",
          2601 => x"08",
          2602 => x"06",
          2603 => x"51",
          2604 => x"83",
          2605 => x"06",
          2606 => x"14",
          2607 => x"3f",
          2608 => x"08",
          2609 => x"07",
          2610 => x"d3",
          2611 => x"3d",
          2612 => x"3d",
          2613 => x"70",
          2614 => x"06",
          2615 => x"53",
          2616 => x"ed",
          2617 => x"33",
          2618 => x"83",
          2619 => x"06",
          2620 => x"90",
          2621 => x"15",
          2622 => x"3f",
          2623 => x"04",
          2624 => x"7b",
          2625 => x"84",
          2626 => x"58",
          2627 => x"80",
          2628 => x"38",
          2629 => x"52",
          2630 => x"8f",
          2631 => x"84",
          2632 => x"d3",
          2633 => x"f5",
          2634 => x"08",
          2635 => x"53",
          2636 => x"84",
          2637 => x"39",
          2638 => x"70",
          2639 => x"81",
          2640 => x"51",
          2641 => x"16",
          2642 => x"84",
          2643 => x"81",
          2644 => x"38",
          2645 => x"ae",
          2646 => x"81",
          2647 => x"54",
          2648 => x"2e",
          2649 => x"8f",
          2650 => x"81",
          2651 => x"76",
          2652 => x"54",
          2653 => x"09",
          2654 => x"38",
          2655 => x"7a",
          2656 => x"80",
          2657 => x"fa",
          2658 => x"d3",
          2659 => x"81",
          2660 => x"89",
          2661 => x"08",
          2662 => x"86",
          2663 => x"98",
          2664 => x"81",
          2665 => x"8b",
          2666 => x"fb",
          2667 => x"70",
          2668 => x"81",
          2669 => x"fc",
          2670 => x"d3",
          2671 => x"81",
          2672 => x"b4",
          2673 => x"08",
          2674 => x"ec",
          2675 => x"d3",
          2676 => x"81",
          2677 => x"a0",
          2678 => x"81",
          2679 => x"52",
          2680 => x"51",
          2681 => x"8b",
          2682 => x"52",
          2683 => x"51",
          2684 => x"81",
          2685 => x"34",
          2686 => x"84",
          2687 => x"0d",
          2688 => x"0d",
          2689 => x"98",
          2690 => x"70",
          2691 => x"ec",
          2692 => x"d3",
          2693 => x"38",
          2694 => x"53",
          2695 => x"81",
          2696 => x"34",
          2697 => x"04",
          2698 => x"78",
          2699 => x"80",
          2700 => x"34",
          2701 => x"80",
          2702 => x"38",
          2703 => x"18",
          2704 => x"9c",
          2705 => x"70",
          2706 => x"56",
          2707 => x"a0",
          2708 => x"71",
          2709 => x"81",
          2710 => x"81",
          2711 => x"89",
          2712 => x"06",
          2713 => x"73",
          2714 => x"55",
          2715 => x"55",
          2716 => x"81",
          2717 => x"81",
          2718 => x"74",
          2719 => x"75",
          2720 => x"52",
          2721 => x"13",
          2722 => x"08",
          2723 => x"33",
          2724 => x"9c",
          2725 => x"11",
          2726 => x"8a",
          2727 => x"84",
          2728 => x"96",
          2729 => x"e7",
          2730 => x"84",
          2731 => x"23",
          2732 => x"e7",
          2733 => x"d3",
          2734 => x"17",
          2735 => x"0d",
          2736 => x"0d",
          2737 => x"5e",
          2738 => x"70",
          2739 => x"55",
          2740 => x"83",
          2741 => x"73",
          2742 => x"91",
          2743 => x"2e",
          2744 => x"1d",
          2745 => x"0c",
          2746 => x"15",
          2747 => x"70",
          2748 => x"56",
          2749 => x"09",
          2750 => x"38",
          2751 => x"80",
          2752 => x"30",
          2753 => x"78",
          2754 => x"54",
          2755 => x"73",
          2756 => x"60",
          2757 => x"54",
          2758 => x"96",
          2759 => x"0b",
          2760 => x"80",
          2761 => x"f6",
          2762 => x"d3",
          2763 => x"85",
          2764 => x"3d",
          2765 => x"5c",
          2766 => x"53",
          2767 => x"51",
          2768 => x"80",
          2769 => x"88",
          2770 => x"5c",
          2771 => x"09",
          2772 => x"d4",
          2773 => x"70",
          2774 => x"71",
          2775 => x"30",
          2776 => x"73",
          2777 => x"51",
          2778 => x"57",
          2779 => x"38",
          2780 => x"75",
          2781 => x"17",
          2782 => x"75",
          2783 => x"30",
          2784 => x"51",
          2785 => x"80",
          2786 => x"38",
          2787 => x"87",
          2788 => x"26",
          2789 => x"77",
          2790 => x"a4",
          2791 => x"27",
          2792 => x"a0",
          2793 => x"39",
          2794 => x"33",
          2795 => x"57",
          2796 => x"27",
          2797 => x"75",
          2798 => x"30",
          2799 => x"32",
          2800 => x"80",
          2801 => x"25",
          2802 => x"56",
          2803 => x"80",
          2804 => x"84",
          2805 => x"58",
          2806 => x"70",
          2807 => x"55",
          2808 => x"09",
          2809 => x"38",
          2810 => x"80",
          2811 => x"30",
          2812 => x"77",
          2813 => x"54",
          2814 => x"81",
          2815 => x"ae",
          2816 => x"06",
          2817 => x"54",
          2818 => x"74",
          2819 => x"80",
          2820 => x"7b",
          2821 => x"30",
          2822 => x"70",
          2823 => x"25",
          2824 => x"07",
          2825 => x"51",
          2826 => x"a7",
          2827 => x"8b",
          2828 => x"39",
          2829 => x"54",
          2830 => x"8c",
          2831 => x"ff",
          2832 => x"f8",
          2833 => x"54",
          2834 => x"e1",
          2835 => x"84",
          2836 => x"b2",
          2837 => x"70",
          2838 => x"71",
          2839 => x"54",
          2840 => x"81",
          2841 => x"80",
          2842 => x"38",
          2843 => x"76",
          2844 => x"df",
          2845 => x"54",
          2846 => x"81",
          2847 => x"55",
          2848 => x"34",
          2849 => x"52",
          2850 => x"51",
          2851 => x"81",
          2852 => x"bf",
          2853 => x"16",
          2854 => x"26",
          2855 => x"16",
          2856 => x"06",
          2857 => x"17",
          2858 => x"34",
          2859 => x"fd",
          2860 => x"19",
          2861 => x"80",
          2862 => x"79",
          2863 => x"81",
          2864 => x"81",
          2865 => x"85",
          2866 => x"54",
          2867 => x"8f",
          2868 => x"86",
          2869 => x"39",
          2870 => x"f3",
          2871 => x"73",
          2872 => x"80",
          2873 => x"52",
          2874 => x"ce",
          2875 => x"84",
          2876 => x"d3",
          2877 => x"d7",
          2878 => x"08",
          2879 => x"e6",
          2880 => x"d3",
          2881 => x"81",
          2882 => x"80",
          2883 => x"1b",
          2884 => x"55",
          2885 => x"2e",
          2886 => x"8b",
          2887 => x"06",
          2888 => x"1c",
          2889 => x"33",
          2890 => x"70",
          2891 => x"55",
          2892 => x"38",
          2893 => x"52",
          2894 => x"9f",
          2895 => x"84",
          2896 => x"8b",
          2897 => x"7a",
          2898 => x"3f",
          2899 => x"75",
          2900 => x"57",
          2901 => x"2e",
          2902 => x"84",
          2903 => x"06",
          2904 => x"75",
          2905 => x"81",
          2906 => x"2a",
          2907 => x"73",
          2908 => x"38",
          2909 => x"54",
          2910 => x"fb",
          2911 => x"80",
          2912 => x"34",
          2913 => x"c1",
          2914 => x"06",
          2915 => x"38",
          2916 => x"39",
          2917 => x"70",
          2918 => x"54",
          2919 => x"86",
          2920 => x"84",
          2921 => x"06",
          2922 => x"73",
          2923 => x"38",
          2924 => x"83",
          2925 => x"b4",
          2926 => x"51",
          2927 => x"81",
          2928 => x"88",
          2929 => x"ea",
          2930 => x"d3",
          2931 => x"3d",
          2932 => x"3d",
          2933 => x"ff",
          2934 => x"71",
          2935 => x"5c",
          2936 => x"80",
          2937 => x"38",
          2938 => x"05",
          2939 => x"a0",
          2940 => x"71",
          2941 => x"38",
          2942 => x"71",
          2943 => x"81",
          2944 => x"38",
          2945 => x"11",
          2946 => x"06",
          2947 => x"70",
          2948 => x"38",
          2949 => x"81",
          2950 => x"05",
          2951 => x"76",
          2952 => x"38",
          2953 => x"c2",
          2954 => x"77",
          2955 => x"57",
          2956 => x"05",
          2957 => x"70",
          2958 => x"33",
          2959 => x"53",
          2960 => x"99",
          2961 => x"e0",
          2962 => x"ff",
          2963 => x"ff",
          2964 => x"70",
          2965 => x"38",
          2966 => x"81",
          2967 => x"51",
          2968 => x"9f",
          2969 => x"72",
          2970 => x"81",
          2971 => x"70",
          2972 => x"72",
          2973 => x"32",
          2974 => x"72",
          2975 => x"73",
          2976 => x"53",
          2977 => x"70",
          2978 => x"38",
          2979 => x"19",
          2980 => x"75",
          2981 => x"38",
          2982 => x"83",
          2983 => x"74",
          2984 => x"59",
          2985 => x"39",
          2986 => x"33",
          2987 => x"d3",
          2988 => x"3d",
          2989 => x"3d",
          2990 => x"80",
          2991 => x"34",
          2992 => x"17",
          2993 => x"75",
          2994 => x"3f",
          2995 => x"d3",
          2996 => x"80",
          2997 => x"16",
          2998 => x"3f",
          2999 => x"08",
          3000 => x"06",
          3001 => x"73",
          3002 => x"2e",
          3003 => x"80",
          3004 => x"0b",
          3005 => x"56",
          3006 => x"e9",
          3007 => x"06",
          3008 => x"57",
          3009 => x"32",
          3010 => x"80",
          3011 => x"51",
          3012 => x"8a",
          3013 => x"e8",
          3014 => x"06",
          3015 => x"53",
          3016 => x"52",
          3017 => x"51",
          3018 => x"81",
          3019 => x"55",
          3020 => x"08",
          3021 => x"38",
          3022 => x"c2",
          3023 => x"86",
          3024 => x"97",
          3025 => x"84",
          3026 => x"d3",
          3027 => x"2e",
          3028 => x"55",
          3029 => x"84",
          3030 => x"0d",
          3031 => x"0d",
          3032 => x"05",
          3033 => x"33",
          3034 => x"75",
          3035 => x"fc",
          3036 => x"d3",
          3037 => x"8b",
          3038 => x"81",
          3039 => x"24",
          3040 => x"81",
          3041 => x"84",
          3042 => x"a0",
          3043 => x"55",
          3044 => x"73",
          3045 => x"e6",
          3046 => x"0c",
          3047 => x"06",
          3048 => x"57",
          3049 => x"ae",
          3050 => x"33",
          3051 => x"3f",
          3052 => x"08",
          3053 => x"70",
          3054 => x"55",
          3055 => x"76",
          3056 => x"b8",
          3057 => x"2a",
          3058 => x"51",
          3059 => x"72",
          3060 => x"86",
          3061 => x"74",
          3062 => x"15",
          3063 => x"81",
          3064 => x"d7",
          3065 => x"d3",
          3066 => x"ff",
          3067 => x"06",
          3068 => x"56",
          3069 => x"38",
          3070 => x"8f",
          3071 => x"2a",
          3072 => x"51",
          3073 => x"72",
          3074 => x"80",
          3075 => x"52",
          3076 => x"3f",
          3077 => x"08",
          3078 => x"57",
          3079 => x"09",
          3080 => x"e2",
          3081 => x"74",
          3082 => x"56",
          3083 => x"33",
          3084 => x"72",
          3085 => x"38",
          3086 => x"51",
          3087 => x"81",
          3088 => x"57",
          3089 => x"84",
          3090 => x"ff",
          3091 => x"56",
          3092 => x"25",
          3093 => x"0b",
          3094 => x"56",
          3095 => x"05",
          3096 => x"83",
          3097 => x"2e",
          3098 => x"52",
          3099 => x"c6",
          3100 => x"84",
          3101 => x"06",
          3102 => x"27",
          3103 => x"16",
          3104 => x"27",
          3105 => x"56",
          3106 => x"84",
          3107 => x"56",
          3108 => x"84",
          3109 => x"14",
          3110 => x"3f",
          3111 => x"08",
          3112 => x"06",
          3113 => x"80",
          3114 => x"06",
          3115 => x"80",
          3116 => x"db",
          3117 => x"d3",
          3118 => x"ff",
          3119 => x"77",
          3120 => x"d8",
          3121 => x"de",
          3122 => x"84",
          3123 => x"9c",
          3124 => x"c4",
          3125 => x"15",
          3126 => x"14",
          3127 => x"70",
          3128 => x"51",
          3129 => x"56",
          3130 => x"84",
          3131 => x"81",
          3132 => x"71",
          3133 => x"16",
          3134 => x"53",
          3135 => x"23",
          3136 => x"8b",
          3137 => x"73",
          3138 => x"80",
          3139 => x"8d",
          3140 => x"39",
          3141 => x"51",
          3142 => x"81",
          3143 => x"53",
          3144 => x"08",
          3145 => x"72",
          3146 => x"8d",
          3147 => x"ce",
          3148 => x"14",
          3149 => x"3f",
          3150 => x"08",
          3151 => x"06",
          3152 => x"38",
          3153 => x"51",
          3154 => x"81",
          3155 => x"55",
          3156 => x"51",
          3157 => x"81",
          3158 => x"83",
          3159 => x"53",
          3160 => x"80",
          3161 => x"38",
          3162 => x"78",
          3163 => x"2a",
          3164 => x"78",
          3165 => x"86",
          3166 => x"22",
          3167 => x"31",
          3168 => x"f6",
          3169 => x"84",
          3170 => x"d3",
          3171 => x"2e",
          3172 => x"81",
          3173 => x"80",
          3174 => x"f5",
          3175 => x"83",
          3176 => x"ff",
          3177 => x"38",
          3178 => x"9f",
          3179 => x"38",
          3180 => x"39",
          3181 => x"80",
          3182 => x"38",
          3183 => x"98",
          3184 => x"a0",
          3185 => x"1c",
          3186 => x"0c",
          3187 => x"17",
          3188 => x"76",
          3189 => x"81",
          3190 => x"80",
          3191 => x"d9",
          3192 => x"d3",
          3193 => x"ff",
          3194 => x"8d",
          3195 => x"8e",
          3196 => x"8a",
          3197 => x"14",
          3198 => x"3f",
          3199 => x"08",
          3200 => x"74",
          3201 => x"a2",
          3202 => x"79",
          3203 => x"ee",
          3204 => x"a8",
          3205 => x"15",
          3206 => x"2e",
          3207 => x"10",
          3208 => x"2a",
          3209 => x"05",
          3210 => x"ff",
          3211 => x"53",
          3212 => x"9c",
          3213 => x"81",
          3214 => x"0b",
          3215 => x"ff",
          3216 => x"0c",
          3217 => x"84",
          3218 => x"83",
          3219 => x"06",
          3220 => x"80",
          3221 => x"d8",
          3222 => x"d3",
          3223 => x"ff",
          3224 => x"72",
          3225 => x"81",
          3226 => x"38",
          3227 => x"73",
          3228 => x"3f",
          3229 => x"08",
          3230 => x"81",
          3231 => x"84",
          3232 => x"b2",
          3233 => x"87",
          3234 => x"84",
          3235 => x"ff",
          3236 => x"82",
          3237 => x"09",
          3238 => x"c8",
          3239 => x"51",
          3240 => x"81",
          3241 => x"84",
          3242 => x"d2",
          3243 => x"06",
          3244 => x"98",
          3245 => x"ee",
          3246 => x"84",
          3247 => x"85",
          3248 => x"09",
          3249 => x"38",
          3250 => x"51",
          3251 => x"81",
          3252 => x"90",
          3253 => x"a0",
          3254 => x"ca",
          3255 => x"84",
          3256 => x"0c",
          3257 => x"81",
          3258 => x"81",
          3259 => x"81",
          3260 => x"72",
          3261 => x"80",
          3262 => x"0c",
          3263 => x"81",
          3264 => x"90",
          3265 => x"fb",
          3266 => x"54",
          3267 => x"80",
          3268 => x"73",
          3269 => x"80",
          3270 => x"72",
          3271 => x"80",
          3272 => x"86",
          3273 => x"15",
          3274 => x"71",
          3275 => x"81",
          3276 => x"81",
          3277 => x"d0",
          3278 => x"d3",
          3279 => x"06",
          3280 => x"38",
          3281 => x"54",
          3282 => x"80",
          3283 => x"71",
          3284 => x"81",
          3285 => x"87",
          3286 => x"fa",
          3287 => x"ab",
          3288 => x"58",
          3289 => x"05",
          3290 => x"e6",
          3291 => x"80",
          3292 => x"84",
          3293 => x"38",
          3294 => x"08",
          3295 => x"d3",
          3296 => x"08",
          3297 => x"80",
          3298 => x"80",
          3299 => x"54",
          3300 => x"84",
          3301 => x"34",
          3302 => x"75",
          3303 => x"2e",
          3304 => x"53",
          3305 => x"53",
          3306 => x"f7",
          3307 => x"d3",
          3308 => x"73",
          3309 => x"0c",
          3310 => x"04",
          3311 => x"67",
          3312 => x"80",
          3313 => x"59",
          3314 => x"78",
          3315 => x"c8",
          3316 => x"06",
          3317 => x"3d",
          3318 => x"99",
          3319 => x"52",
          3320 => x"3f",
          3321 => x"08",
          3322 => x"84",
          3323 => x"38",
          3324 => x"52",
          3325 => x"52",
          3326 => x"3f",
          3327 => x"08",
          3328 => x"84",
          3329 => x"02",
          3330 => x"33",
          3331 => x"55",
          3332 => x"25",
          3333 => x"55",
          3334 => x"54",
          3335 => x"81",
          3336 => x"80",
          3337 => x"74",
          3338 => x"81",
          3339 => x"75",
          3340 => x"3f",
          3341 => x"08",
          3342 => x"02",
          3343 => x"91",
          3344 => x"81",
          3345 => x"82",
          3346 => x"06",
          3347 => x"80",
          3348 => x"88",
          3349 => x"39",
          3350 => x"58",
          3351 => x"38",
          3352 => x"70",
          3353 => x"54",
          3354 => x"81",
          3355 => x"52",
          3356 => x"a5",
          3357 => x"84",
          3358 => x"88",
          3359 => x"62",
          3360 => x"d4",
          3361 => x"54",
          3362 => x"15",
          3363 => x"62",
          3364 => x"e8",
          3365 => x"52",
          3366 => x"51",
          3367 => x"7a",
          3368 => x"83",
          3369 => x"80",
          3370 => x"38",
          3371 => x"08",
          3372 => x"53",
          3373 => x"3d",
          3374 => x"dd",
          3375 => x"d3",
          3376 => x"81",
          3377 => x"82",
          3378 => x"39",
          3379 => x"38",
          3380 => x"33",
          3381 => x"70",
          3382 => x"55",
          3383 => x"2e",
          3384 => x"55",
          3385 => x"77",
          3386 => x"81",
          3387 => x"73",
          3388 => x"38",
          3389 => x"54",
          3390 => x"a0",
          3391 => x"82",
          3392 => x"52",
          3393 => x"a3",
          3394 => x"84",
          3395 => x"18",
          3396 => x"55",
          3397 => x"84",
          3398 => x"38",
          3399 => x"70",
          3400 => x"54",
          3401 => x"86",
          3402 => x"c0",
          3403 => x"b0",
          3404 => x"1b",
          3405 => x"1b",
          3406 => x"70",
          3407 => x"d9",
          3408 => x"84",
          3409 => x"84",
          3410 => x"0c",
          3411 => x"52",
          3412 => x"3f",
          3413 => x"08",
          3414 => x"08",
          3415 => x"77",
          3416 => x"86",
          3417 => x"1a",
          3418 => x"1a",
          3419 => x"91",
          3420 => x"0b",
          3421 => x"80",
          3422 => x"0c",
          3423 => x"70",
          3424 => x"54",
          3425 => x"81",
          3426 => x"d3",
          3427 => x"2e",
          3428 => x"81",
          3429 => x"94",
          3430 => x"17",
          3431 => x"2b",
          3432 => x"57",
          3433 => x"52",
          3434 => x"9f",
          3435 => x"84",
          3436 => x"d3",
          3437 => x"26",
          3438 => x"55",
          3439 => x"08",
          3440 => x"81",
          3441 => x"79",
          3442 => x"31",
          3443 => x"70",
          3444 => x"25",
          3445 => x"76",
          3446 => x"81",
          3447 => x"55",
          3448 => x"38",
          3449 => x"0c",
          3450 => x"75",
          3451 => x"54",
          3452 => x"a2",
          3453 => x"7a",
          3454 => x"3f",
          3455 => x"08",
          3456 => x"55",
          3457 => x"89",
          3458 => x"84",
          3459 => x"1a",
          3460 => x"80",
          3461 => x"54",
          3462 => x"84",
          3463 => x"0d",
          3464 => x"0d",
          3465 => x"64",
          3466 => x"59",
          3467 => x"90",
          3468 => x"52",
          3469 => x"cf",
          3470 => x"84",
          3471 => x"d3",
          3472 => x"38",
          3473 => x"55",
          3474 => x"86",
          3475 => x"82",
          3476 => x"19",
          3477 => x"55",
          3478 => x"80",
          3479 => x"38",
          3480 => x"0b",
          3481 => x"82",
          3482 => x"39",
          3483 => x"1a",
          3484 => x"82",
          3485 => x"19",
          3486 => x"08",
          3487 => x"7c",
          3488 => x"74",
          3489 => x"2e",
          3490 => x"94",
          3491 => x"83",
          3492 => x"56",
          3493 => x"38",
          3494 => x"22",
          3495 => x"89",
          3496 => x"55",
          3497 => x"75",
          3498 => x"19",
          3499 => x"39",
          3500 => x"52",
          3501 => x"93",
          3502 => x"84",
          3503 => x"75",
          3504 => x"38",
          3505 => x"ff",
          3506 => x"98",
          3507 => x"19",
          3508 => x"51",
          3509 => x"81",
          3510 => x"80",
          3511 => x"38",
          3512 => x"08",
          3513 => x"2a",
          3514 => x"80",
          3515 => x"38",
          3516 => x"8a",
          3517 => x"5c",
          3518 => x"27",
          3519 => x"7a",
          3520 => x"54",
          3521 => x"52",
          3522 => x"51",
          3523 => x"81",
          3524 => x"fe",
          3525 => x"83",
          3526 => x"56",
          3527 => x"9f",
          3528 => x"08",
          3529 => x"74",
          3530 => x"38",
          3531 => x"b4",
          3532 => x"16",
          3533 => x"89",
          3534 => x"51",
          3535 => x"77",
          3536 => x"b9",
          3537 => x"1a",
          3538 => x"08",
          3539 => x"84",
          3540 => x"57",
          3541 => x"27",
          3542 => x"56",
          3543 => x"52",
          3544 => x"c7",
          3545 => x"84",
          3546 => x"38",
          3547 => x"19",
          3548 => x"06",
          3549 => x"52",
          3550 => x"a2",
          3551 => x"31",
          3552 => x"7f",
          3553 => x"94",
          3554 => x"94",
          3555 => x"5c",
          3556 => x"80",
          3557 => x"d3",
          3558 => x"3d",
          3559 => x"3d",
          3560 => x"65",
          3561 => x"5d",
          3562 => x"0c",
          3563 => x"05",
          3564 => x"f6",
          3565 => x"d3",
          3566 => x"81",
          3567 => x"8a",
          3568 => x"33",
          3569 => x"2e",
          3570 => x"56",
          3571 => x"90",
          3572 => x"81",
          3573 => x"06",
          3574 => x"87",
          3575 => x"2e",
          3576 => x"95",
          3577 => x"91",
          3578 => x"56",
          3579 => x"81",
          3580 => x"34",
          3581 => x"8e",
          3582 => x"08",
          3583 => x"56",
          3584 => x"84",
          3585 => x"5c",
          3586 => x"82",
          3587 => x"18",
          3588 => x"ff",
          3589 => x"74",
          3590 => x"7e",
          3591 => x"ff",
          3592 => x"2a",
          3593 => x"7a",
          3594 => x"8c",
          3595 => x"08",
          3596 => x"38",
          3597 => x"39",
          3598 => x"52",
          3599 => x"e7",
          3600 => x"84",
          3601 => x"d3",
          3602 => x"2e",
          3603 => x"74",
          3604 => x"91",
          3605 => x"2e",
          3606 => x"74",
          3607 => x"88",
          3608 => x"38",
          3609 => x"0c",
          3610 => x"15",
          3611 => x"08",
          3612 => x"06",
          3613 => x"51",
          3614 => x"81",
          3615 => x"fe",
          3616 => x"18",
          3617 => x"51",
          3618 => x"81",
          3619 => x"80",
          3620 => x"38",
          3621 => x"08",
          3622 => x"2a",
          3623 => x"80",
          3624 => x"38",
          3625 => x"8a",
          3626 => x"5b",
          3627 => x"27",
          3628 => x"7b",
          3629 => x"54",
          3630 => x"52",
          3631 => x"51",
          3632 => x"81",
          3633 => x"fe",
          3634 => x"b0",
          3635 => x"31",
          3636 => x"79",
          3637 => x"84",
          3638 => x"16",
          3639 => x"89",
          3640 => x"52",
          3641 => x"cc",
          3642 => x"55",
          3643 => x"16",
          3644 => x"2b",
          3645 => x"39",
          3646 => x"94",
          3647 => x"93",
          3648 => x"cd",
          3649 => x"d3",
          3650 => x"e3",
          3651 => x"b0",
          3652 => x"76",
          3653 => x"94",
          3654 => x"ff",
          3655 => x"71",
          3656 => x"7b",
          3657 => x"38",
          3658 => x"18",
          3659 => x"51",
          3660 => x"81",
          3661 => x"fd",
          3662 => x"53",
          3663 => x"18",
          3664 => x"06",
          3665 => x"51",
          3666 => x"7e",
          3667 => x"83",
          3668 => x"76",
          3669 => x"17",
          3670 => x"1e",
          3671 => x"18",
          3672 => x"0c",
          3673 => x"58",
          3674 => x"74",
          3675 => x"38",
          3676 => x"8c",
          3677 => x"90",
          3678 => x"33",
          3679 => x"55",
          3680 => x"34",
          3681 => x"81",
          3682 => x"90",
          3683 => x"f8",
          3684 => x"8b",
          3685 => x"53",
          3686 => x"f2",
          3687 => x"d3",
          3688 => x"81",
          3689 => x"80",
          3690 => x"16",
          3691 => x"2a",
          3692 => x"51",
          3693 => x"80",
          3694 => x"38",
          3695 => x"52",
          3696 => x"e7",
          3697 => x"84",
          3698 => x"d3",
          3699 => x"d4",
          3700 => x"08",
          3701 => x"a0",
          3702 => x"73",
          3703 => x"88",
          3704 => x"74",
          3705 => x"51",
          3706 => x"8c",
          3707 => x"9c",
          3708 => x"fb",
          3709 => x"b2",
          3710 => x"15",
          3711 => x"3f",
          3712 => x"15",
          3713 => x"3f",
          3714 => x"0b",
          3715 => x"78",
          3716 => x"3f",
          3717 => x"08",
          3718 => x"81",
          3719 => x"57",
          3720 => x"34",
          3721 => x"84",
          3722 => x"0d",
          3723 => x"0d",
          3724 => x"54",
          3725 => x"81",
          3726 => x"53",
          3727 => x"08",
          3728 => x"3d",
          3729 => x"73",
          3730 => x"3f",
          3731 => x"08",
          3732 => x"84",
          3733 => x"81",
          3734 => x"74",
          3735 => x"d3",
          3736 => x"3d",
          3737 => x"3d",
          3738 => x"51",
          3739 => x"8b",
          3740 => x"81",
          3741 => x"24",
          3742 => x"d3",
          3743 => x"d3",
          3744 => x"52",
          3745 => x"84",
          3746 => x"0d",
          3747 => x"0d",
          3748 => x"3d",
          3749 => x"94",
          3750 => x"c1",
          3751 => x"84",
          3752 => x"d3",
          3753 => x"e0",
          3754 => x"63",
          3755 => x"d4",
          3756 => x"8d",
          3757 => x"84",
          3758 => x"d3",
          3759 => x"38",
          3760 => x"05",
          3761 => x"2b",
          3762 => x"80",
          3763 => x"76",
          3764 => x"0c",
          3765 => x"02",
          3766 => x"70",
          3767 => x"81",
          3768 => x"56",
          3769 => x"9e",
          3770 => x"53",
          3771 => x"db",
          3772 => x"d3",
          3773 => x"15",
          3774 => x"81",
          3775 => x"84",
          3776 => x"06",
          3777 => x"55",
          3778 => x"84",
          3779 => x"0d",
          3780 => x"0d",
          3781 => x"5b",
          3782 => x"80",
          3783 => x"ff",
          3784 => x"9f",
          3785 => x"b5",
          3786 => x"84",
          3787 => x"d3",
          3788 => x"fc",
          3789 => x"7a",
          3790 => x"08",
          3791 => x"64",
          3792 => x"2e",
          3793 => x"a0",
          3794 => x"70",
          3795 => x"ea",
          3796 => x"84",
          3797 => x"d3",
          3798 => x"d4",
          3799 => x"7b",
          3800 => x"3f",
          3801 => x"08",
          3802 => x"84",
          3803 => x"38",
          3804 => x"51",
          3805 => x"81",
          3806 => x"45",
          3807 => x"51",
          3808 => x"81",
          3809 => x"57",
          3810 => x"08",
          3811 => x"80",
          3812 => x"da",
          3813 => x"d3",
          3814 => x"81",
          3815 => x"a4",
          3816 => x"7b",
          3817 => x"3f",
          3818 => x"84",
          3819 => x"38",
          3820 => x"51",
          3821 => x"81",
          3822 => x"57",
          3823 => x"08",
          3824 => x"38",
          3825 => x"09",
          3826 => x"38",
          3827 => x"e0",
          3828 => x"dc",
          3829 => x"ff",
          3830 => x"74",
          3831 => x"3f",
          3832 => x"78",
          3833 => x"33",
          3834 => x"56",
          3835 => x"91",
          3836 => x"05",
          3837 => x"81",
          3838 => x"56",
          3839 => x"f5",
          3840 => x"54",
          3841 => x"81",
          3842 => x"80",
          3843 => x"78",
          3844 => x"55",
          3845 => x"11",
          3846 => x"18",
          3847 => x"58",
          3848 => x"34",
          3849 => x"ff",
          3850 => x"55",
          3851 => x"34",
          3852 => x"77",
          3853 => x"81",
          3854 => x"ff",
          3855 => x"55",
          3856 => x"34",
          3857 => x"d3",
          3858 => x"84",
          3859 => x"e8",
          3860 => x"70",
          3861 => x"56",
          3862 => x"76",
          3863 => x"81",
          3864 => x"70",
          3865 => x"56",
          3866 => x"82",
          3867 => x"78",
          3868 => x"80",
          3869 => x"27",
          3870 => x"19",
          3871 => x"7a",
          3872 => x"5c",
          3873 => x"55",
          3874 => x"7a",
          3875 => x"5c",
          3876 => x"2e",
          3877 => x"85",
          3878 => x"94",
          3879 => x"81",
          3880 => x"73",
          3881 => x"81",
          3882 => x"7a",
          3883 => x"38",
          3884 => x"76",
          3885 => x"0c",
          3886 => x"04",
          3887 => x"7b",
          3888 => x"fc",
          3889 => x"53",
          3890 => x"bb",
          3891 => x"84",
          3892 => x"d3",
          3893 => x"fa",
          3894 => x"33",
          3895 => x"f2",
          3896 => x"08",
          3897 => x"27",
          3898 => x"15",
          3899 => x"2a",
          3900 => x"51",
          3901 => x"83",
          3902 => x"94",
          3903 => x"80",
          3904 => x"0c",
          3905 => x"2e",
          3906 => x"79",
          3907 => x"70",
          3908 => x"51",
          3909 => x"2e",
          3910 => x"52",
          3911 => x"ff",
          3912 => x"81",
          3913 => x"ff",
          3914 => x"70",
          3915 => x"ff",
          3916 => x"81",
          3917 => x"73",
          3918 => x"76",
          3919 => x"06",
          3920 => x"0c",
          3921 => x"98",
          3922 => x"58",
          3923 => x"39",
          3924 => x"54",
          3925 => x"73",
          3926 => x"cd",
          3927 => x"d3",
          3928 => x"81",
          3929 => x"81",
          3930 => x"38",
          3931 => x"08",
          3932 => x"9b",
          3933 => x"84",
          3934 => x"0c",
          3935 => x"0c",
          3936 => x"81",
          3937 => x"76",
          3938 => x"38",
          3939 => x"94",
          3940 => x"94",
          3941 => x"16",
          3942 => x"2a",
          3943 => x"51",
          3944 => x"72",
          3945 => x"38",
          3946 => x"51",
          3947 => x"81",
          3948 => x"54",
          3949 => x"08",
          3950 => x"d3",
          3951 => x"a7",
          3952 => x"74",
          3953 => x"3f",
          3954 => x"08",
          3955 => x"2e",
          3956 => x"74",
          3957 => x"79",
          3958 => x"14",
          3959 => x"38",
          3960 => x"0c",
          3961 => x"94",
          3962 => x"94",
          3963 => x"83",
          3964 => x"72",
          3965 => x"38",
          3966 => x"51",
          3967 => x"81",
          3968 => x"94",
          3969 => x"91",
          3970 => x"53",
          3971 => x"81",
          3972 => x"34",
          3973 => x"39",
          3974 => x"81",
          3975 => x"05",
          3976 => x"08",
          3977 => x"08",
          3978 => x"38",
          3979 => x"0c",
          3980 => x"80",
          3981 => x"72",
          3982 => x"73",
          3983 => x"53",
          3984 => x"8c",
          3985 => x"16",
          3986 => x"38",
          3987 => x"0c",
          3988 => x"81",
          3989 => x"8b",
          3990 => x"f9",
          3991 => x"56",
          3992 => x"80",
          3993 => x"38",
          3994 => x"3d",
          3995 => x"8a",
          3996 => x"51",
          3997 => x"81",
          3998 => x"55",
          3999 => x"08",
          4000 => x"77",
          4001 => x"52",
          4002 => x"b5",
          4003 => x"84",
          4004 => x"d3",
          4005 => x"c3",
          4006 => x"33",
          4007 => x"55",
          4008 => x"24",
          4009 => x"16",
          4010 => x"2a",
          4011 => x"51",
          4012 => x"80",
          4013 => x"9c",
          4014 => x"77",
          4015 => x"3f",
          4016 => x"08",
          4017 => x"77",
          4018 => x"22",
          4019 => x"74",
          4020 => x"ce",
          4021 => x"d3",
          4022 => x"74",
          4023 => x"81",
          4024 => x"85",
          4025 => x"74",
          4026 => x"38",
          4027 => x"74",
          4028 => x"d3",
          4029 => x"3d",
          4030 => x"3d",
          4031 => x"3d",
          4032 => x"70",
          4033 => x"ff",
          4034 => x"84",
          4035 => x"81",
          4036 => x"73",
          4037 => x"0d",
          4038 => x"0d",
          4039 => x"3d",
          4040 => x"71",
          4041 => x"e7",
          4042 => x"d3",
          4043 => x"81",
          4044 => x"80",
          4045 => x"93",
          4046 => x"84",
          4047 => x"51",
          4048 => x"81",
          4049 => x"53",
          4050 => x"81",
          4051 => x"52",
          4052 => x"ac",
          4053 => x"84",
          4054 => x"d3",
          4055 => x"2e",
          4056 => x"85",
          4057 => x"87",
          4058 => x"84",
          4059 => x"74",
          4060 => x"d5",
          4061 => x"52",
          4062 => x"89",
          4063 => x"84",
          4064 => x"70",
          4065 => x"07",
          4066 => x"81",
          4067 => x"06",
          4068 => x"54",
          4069 => x"84",
          4070 => x"0d",
          4071 => x"0d",
          4072 => x"53",
          4073 => x"53",
          4074 => x"56",
          4075 => x"81",
          4076 => x"55",
          4077 => x"08",
          4078 => x"52",
          4079 => x"81",
          4080 => x"84",
          4081 => x"d3",
          4082 => x"38",
          4083 => x"05",
          4084 => x"2b",
          4085 => x"80",
          4086 => x"86",
          4087 => x"76",
          4088 => x"38",
          4089 => x"51",
          4090 => x"74",
          4091 => x"0c",
          4092 => x"04",
          4093 => x"63",
          4094 => x"80",
          4095 => x"ec",
          4096 => x"3d",
          4097 => x"3f",
          4098 => x"08",
          4099 => x"84",
          4100 => x"38",
          4101 => x"73",
          4102 => x"08",
          4103 => x"13",
          4104 => x"58",
          4105 => x"26",
          4106 => x"7c",
          4107 => x"39",
          4108 => x"cc",
          4109 => x"81",
          4110 => x"d3",
          4111 => x"33",
          4112 => x"81",
          4113 => x"06",
          4114 => x"75",
          4115 => x"52",
          4116 => x"05",
          4117 => x"3f",
          4118 => x"08",
          4119 => x"38",
          4120 => x"08",
          4121 => x"38",
          4122 => x"08",
          4123 => x"d3",
          4124 => x"80",
          4125 => x"81",
          4126 => x"59",
          4127 => x"14",
          4128 => x"ca",
          4129 => x"39",
          4130 => x"81",
          4131 => x"57",
          4132 => x"38",
          4133 => x"18",
          4134 => x"ff",
          4135 => x"81",
          4136 => x"5b",
          4137 => x"08",
          4138 => x"7c",
          4139 => x"12",
          4140 => x"52",
          4141 => x"82",
          4142 => x"06",
          4143 => x"14",
          4144 => x"cb",
          4145 => x"84",
          4146 => x"ff",
          4147 => x"70",
          4148 => x"82",
          4149 => x"51",
          4150 => x"b4",
          4151 => x"bb",
          4152 => x"d3",
          4153 => x"0a",
          4154 => x"70",
          4155 => x"84",
          4156 => x"51",
          4157 => x"ff",
          4158 => x"56",
          4159 => x"38",
          4160 => x"7c",
          4161 => x"0c",
          4162 => x"81",
          4163 => x"74",
          4164 => x"7a",
          4165 => x"0c",
          4166 => x"04",
          4167 => x"79",
          4168 => x"05",
          4169 => x"57",
          4170 => x"81",
          4171 => x"56",
          4172 => x"08",
          4173 => x"91",
          4174 => x"75",
          4175 => x"90",
          4176 => x"81",
          4177 => x"06",
          4178 => x"87",
          4179 => x"2e",
          4180 => x"94",
          4181 => x"73",
          4182 => x"27",
          4183 => x"73",
          4184 => x"d3",
          4185 => x"88",
          4186 => x"76",
          4187 => x"3f",
          4188 => x"08",
          4189 => x"0c",
          4190 => x"39",
          4191 => x"52",
          4192 => x"bf",
          4193 => x"d3",
          4194 => x"2e",
          4195 => x"83",
          4196 => x"81",
          4197 => x"81",
          4198 => x"06",
          4199 => x"56",
          4200 => x"a0",
          4201 => x"81",
          4202 => x"98",
          4203 => x"94",
          4204 => x"08",
          4205 => x"84",
          4206 => x"51",
          4207 => x"81",
          4208 => x"56",
          4209 => x"8c",
          4210 => x"17",
          4211 => x"07",
          4212 => x"18",
          4213 => x"2e",
          4214 => x"91",
          4215 => x"55",
          4216 => x"84",
          4217 => x"0d",
          4218 => x"0d",
          4219 => x"3d",
          4220 => x"52",
          4221 => x"da",
          4222 => x"d3",
          4223 => x"81",
          4224 => x"81",
          4225 => x"45",
          4226 => x"52",
          4227 => x"52",
          4228 => x"3f",
          4229 => x"08",
          4230 => x"84",
          4231 => x"38",
          4232 => x"05",
          4233 => x"2a",
          4234 => x"51",
          4235 => x"55",
          4236 => x"38",
          4237 => x"54",
          4238 => x"81",
          4239 => x"80",
          4240 => x"70",
          4241 => x"54",
          4242 => x"81",
          4243 => x"52",
          4244 => x"c5",
          4245 => x"84",
          4246 => x"2a",
          4247 => x"51",
          4248 => x"80",
          4249 => x"38",
          4250 => x"d3",
          4251 => x"15",
          4252 => x"86",
          4253 => x"81",
          4254 => x"5c",
          4255 => x"3d",
          4256 => x"c7",
          4257 => x"d3",
          4258 => x"81",
          4259 => x"80",
          4260 => x"d3",
          4261 => x"73",
          4262 => x"3f",
          4263 => x"08",
          4264 => x"84",
          4265 => x"87",
          4266 => x"39",
          4267 => x"08",
          4268 => x"38",
          4269 => x"08",
          4270 => x"77",
          4271 => x"3f",
          4272 => x"08",
          4273 => x"08",
          4274 => x"d3",
          4275 => x"80",
          4276 => x"55",
          4277 => x"94",
          4278 => x"2e",
          4279 => x"53",
          4280 => x"51",
          4281 => x"81",
          4282 => x"55",
          4283 => x"78",
          4284 => x"fe",
          4285 => x"84",
          4286 => x"81",
          4287 => x"a0",
          4288 => x"e9",
          4289 => x"53",
          4290 => x"05",
          4291 => x"51",
          4292 => x"81",
          4293 => x"54",
          4294 => x"08",
          4295 => x"78",
          4296 => x"8e",
          4297 => x"58",
          4298 => x"81",
          4299 => x"54",
          4300 => x"08",
          4301 => x"54",
          4302 => x"81",
          4303 => x"84",
          4304 => x"06",
          4305 => x"02",
          4306 => x"33",
          4307 => x"81",
          4308 => x"86",
          4309 => x"f6",
          4310 => x"74",
          4311 => x"70",
          4312 => x"c3",
          4313 => x"84",
          4314 => x"56",
          4315 => x"08",
          4316 => x"54",
          4317 => x"08",
          4318 => x"81",
          4319 => x"82",
          4320 => x"84",
          4321 => x"09",
          4322 => x"38",
          4323 => x"b4",
          4324 => x"b0",
          4325 => x"84",
          4326 => x"51",
          4327 => x"81",
          4328 => x"54",
          4329 => x"08",
          4330 => x"8b",
          4331 => x"b4",
          4332 => x"b7",
          4333 => x"54",
          4334 => x"15",
          4335 => x"90",
          4336 => x"34",
          4337 => x"0a",
          4338 => x"19",
          4339 => x"9f",
          4340 => x"78",
          4341 => x"51",
          4342 => x"a0",
          4343 => x"11",
          4344 => x"05",
          4345 => x"b6",
          4346 => x"ae",
          4347 => x"15",
          4348 => x"78",
          4349 => x"53",
          4350 => x"3f",
          4351 => x"0b",
          4352 => x"77",
          4353 => x"3f",
          4354 => x"08",
          4355 => x"84",
          4356 => x"82",
          4357 => x"52",
          4358 => x"51",
          4359 => x"3f",
          4360 => x"52",
          4361 => x"aa",
          4362 => x"90",
          4363 => x"34",
          4364 => x"0b",
          4365 => x"78",
          4366 => x"b6",
          4367 => x"84",
          4368 => x"39",
          4369 => x"52",
          4370 => x"be",
          4371 => x"81",
          4372 => x"99",
          4373 => x"da",
          4374 => x"3d",
          4375 => x"d2",
          4376 => x"53",
          4377 => x"84",
          4378 => x"3d",
          4379 => x"3f",
          4380 => x"08",
          4381 => x"84",
          4382 => x"38",
          4383 => x"3d",
          4384 => x"3d",
          4385 => x"cc",
          4386 => x"d3",
          4387 => x"81",
          4388 => x"82",
          4389 => x"81",
          4390 => x"81",
          4391 => x"86",
          4392 => x"aa",
          4393 => x"a4",
          4394 => x"a8",
          4395 => x"05",
          4396 => x"ea",
          4397 => x"77",
          4398 => x"70",
          4399 => x"b4",
          4400 => x"3d",
          4401 => x"51",
          4402 => x"81",
          4403 => x"55",
          4404 => x"08",
          4405 => x"6f",
          4406 => x"06",
          4407 => x"a2",
          4408 => x"92",
          4409 => x"81",
          4410 => x"d3",
          4411 => x"2e",
          4412 => x"81",
          4413 => x"51",
          4414 => x"81",
          4415 => x"55",
          4416 => x"08",
          4417 => x"68",
          4418 => x"a8",
          4419 => x"05",
          4420 => x"51",
          4421 => x"3f",
          4422 => x"33",
          4423 => x"8b",
          4424 => x"84",
          4425 => x"06",
          4426 => x"73",
          4427 => x"a0",
          4428 => x"8b",
          4429 => x"54",
          4430 => x"15",
          4431 => x"33",
          4432 => x"70",
          4433 => x"55",
          4434 => x"2e",
          4435 => x"6e",
          4436 => x"df",
          4437 => x"78",
          4438 => x"3f",
          4439 => x"08",
          4440 => x"ff",
          4441 => x"82",
          4442 => x"84",
          4443 => x"80",
          4444 => x"d3",
          4445 => x"78",
          4446 => x"af",
          4447 => x"84",
          4448 => x"d4",
          4449 => x"55",
          4450 => x"08",
          4451 => x"81",
          4452 => x"73",
          4453 => x"81",
          4454 => x"63",
          4455 => x"76",
          4456 => x"3f",
          4457 => x"0b",
          4458 => x"87",
          4459 => x"84",
          4460 => x"77",
          4461 => x"3f",
          4462 => x"08",
          4463 => x"84",
          4464 => x"78",
          4465 => x"aa",
          4466 => x"84",
          4467 => x"81",
          4468 => x"a8",
          4469 => x"ed",
          4470 => x"80",
          4471 => x"02",
          4472 => x"df",
          4473 => x"57",
          4474 => x"3d",
          4475 => x"96",
          4476 => x"e9",
          4477 => x"84",
          4478 => x"d3",
          4479 => x"cf",
          4480 => x"65",
          4481 => x"d4",
          4482 => x"b5",
          4483 => x"84",
          4484 => x"d3",
          4485 => x"38",
          4486 => x"05",
          4487 => x"06",
          4488 => x"73",
          4489 => x"a7",
          4490 => x"09",
          4491 => x"71",
          4492 => x"06",
          4493 => x"55",
          4494 => x"15",
          4495 => x"81",
          4496 => x"34",
          4497 => x"b4",
          4498 => x"d3",
          4499 => x"74",
          4500 => x"0c",
          4501 => x"04",
          4502 => x"64",
          4503 => x"93",
          4504 => x"52",
          4505 => x"d1",
          4506 => x"d3",
          4507 => x"81",
          4508 => x"80",
          4509 => x"58",
          4510 => x"3d",
          4511 => x"c8",
          4512 => x"d3",
          4513 => x"81",
          4514 => x"b4",
          4515 => x"c7",
          4516 => x"a0",
          4517 => x"55",
          4518 => x"84",
          4519 => x"17",
          4520 => x"2b",
          4521 => x"96",
          4522 => x"b0",
          4523 => x"54",
          4524 => x"15",
          4525 => x"ff",
          4526 => x"81",
          4527 => x"55",
          4528 => x"84",
          4529 => x"0d",
          4530 => x"0d",
          4531 => x"5a",
          4532 => x"3d",
          4533 => x"99",
          4534 => x"81",
          4535 => x"84",
          4536 => x"84",
          4537 => x"81",
          4538 => x"07",
          4539 => x"55",
          4540 => x"2e",
          4541 => x"81",
          4542 => x"55",
          4543 => x"2e",
          4544 => x"7b",
          4545 => x"80",
          4546 => x"70",
          4547 => x"be",
          4548 => x"d3",
          4549 => x"81",
          4550 => x"80",
          4551 => x"52",
          4552 => x"dc",
          4553 => x"84",
          4554 => x"d3",
          4555 => x"38",
          4556 => x"08",
          4557 => x"08",
          4558 => x"56",
          4559 => x"19",
          4560 => x"59",
          4561 => x"74",
          4562 => x"56",
          4563 => x"ec",
          4564 => x"75",
          4565 => x"74",
          4566 => x"2e",
          4567 => x"16",
          4568 => x"33",
          4569 => x"73",
          4570 => x"38",
          4571 => x"84",
          4572 => x"06",
          4573 => x"7a",
          4574 => x"76",
          4575 => x"07",
          4576 => x"54",
          4577 => x"80",
          4578 => x"80",
          4579 => x"7b",
          4580 => x"53",
          4581 => x"93",
          4582 => x"84",
          4583 => x"d3",
          4584 => x"38",
          4585 => x"55",
          4586 => x"56",
          4587 => x"8b",
          4588 => x"56",
          4589 => x"83",
          4590 => x"75",
          4591 => x"51",
          4592 => x"3f",
          4593 => x"08",
          4594 => x"81",
          4595 => x"98",
          4596 => x"e6",
          4597 => x"53",
          4598 => x"b8",
          4599 => x"3d",
          4600 => x"3f",
          4601 => x"08",
          4602 => x"08",
          4603 => x"d3",
          4604 => x"98",
          4605 => x"a0",
          4606 => x"70",
          4607 => x"ae",
          4608 => x"6d",
          4609 => x"81",
          4610 => x"57",
          4611 => x"74",
          4612 => x"38",
          4613 => x"81",
          4614 => x"81",
          4615 => x"52",
          4616 => x"89",
          4617 => x"84",
          4618 => x"a5",
          4619 => x"33",
          4620 => x"54",
          4621 => x"3f",
          4622 => x"08",
          4623 => x"38",
          4624 => x"76",
          4625 => x"05",
          4626 => x"39",
          4627 => x"08",
          4628 => x"15",
          4629 => x"ff",
          4630 => x"73",
          4631 => x"38",
          4632 => x"83",
          4633 => x"56",
          4634 => x"75",
          4635 => x"81",
          4636 => x"33",
          4637 => x"2e",
          4638 => x"52",
          4639 => x"51",
          4640 => x"3f",
          4641 => x"08",
          4642 => x"ff",
          4643 => x"38",
          4644 => x"88",
          4645 => x"8a",
          4646 => x"38",
          4647 => x"ec",
          4648 => x"75",
          4649 => x"74",
          4650 => x"73",
          4651 => x"05",
          4652 => x"17",
          4653 => x"70",
          4654 => x"34",
          4655 => x"70",
          4656 => x"ff",
          4657 => x"55",
          4658 => x"26",
          4659 => x"8b",
          4660 => x"86",
          4661 => x"e5",
          4662 => x"38",
          4663 => x"99",
          4664 => x"05",
          4665 => x"70",
          4666 => x"73",
          4667 => x"81",
          4668 => x"ff",
          4669 => x"ed",
          4670 => x"80",
          4671 => x"91",
          4672 => x"55",
          4673 => x"3f",
          4674 => x"08",
          4675 => x"84",
          4676 => x"38",
          4677 => x"51",
          4678 => x"3f",
          4679 => x"08",
          4680 => x"84",
          4681 => x"76",
          4682 => x"67",
          4683 => x"34",
          4684 => x"81",
          4685 => x"84",
          4686 => x"06",
          4687 => x"80",
          4688 => x"2e",
          4689 => x"81",
          4690 => x"ff",
          4691 => x"81",
          4692 => x"54",
          4693 => x"08",
          4694 => x"53",
          4695 => x"08",
          4696 => x"ff",
          4697 => x"67",
          4698 => x"8b",
          4699 => x"53",
          4700 => x"51",
          4701 => x"3f",
          4702 => x"0b",
          4703 => x"79",
          4704 => x"ee",
          4705 => x"84",
          4706 => x"55",
          4707 => x"84",
          4708 => x"0d",
          4709 => x"0d",
          4710 => x"88",
          4711 => x"05",
          4712 => x"fc",
          4713 => x"54",
          4714 => x"d2",
          4715 => x"d3",
          4716 => x"81",
          4717 => x"82",
          4718 => x"1a",
          4719 => x"82",
          4720 => x"80",
          4721 => x"8c",
          4722 => x"78",
          4723 => x"1a",
          4724 => x"2a",
          4725 => x"51",
          4726 => x"90",
          4727 => x"82",
          4728 => x"58",
          4729 => x"81",
          4730 => x"39",
          4731 => x"22",
          4732 => x"70",
          4733 => x"56",
          4734 => x"fe",
          4735 => x"14",
          4736 => x"30",
          4737 => x"9f",
          4738 => x"84",
          4739 => x"19",
          4740 => x"5a",
          4741 => x"81",
          4742 => x"38",
          4743 => x"77",
          4744 => x"82",
          4745 => x"56",
          4746 => x"74",
          4747 => x"ff",
          4748 => x"81",
          4749 => x"55",
          4750 => x"75",
          4751 => x"82",
          4752 => x"84",
          4753 => x"ff",
          4754 => x"d3",
          4755 => x"2e",
          4756 => x"81",
          4757 => x"8e",
          4758 => x"56",
          4759 => x"09",
          4760 => x"38",
          4761 => x"59",
          4762 => x"77",
          4763 => x"06",
          4764 => x"87",
          4765 => x"39",
          4766 => x"ba",
          4767 => x"55",
          4768 => x"2e",
          4769 => x"15",
          4770 => x"2e",
          4771 => x"83",
          4772 => x"75",
          4773 => x"7e",
          4774 => x"a8",
          4775 => x"84",
          4776 => x"d3",
          4777 => x"ce",
          4778 => x"16",
          4779 => x"56",
          4780 => x"38",
          4781 => x"19",
          4782 => x"8c",
          4783 => x"7d",
          4784 => x"38",
          4785 => x"0c",
          4786 => x"0c",
          4787 => x"80",
          4788 => x"73",
          4789 => x"98",
          4790 => x"05",
          4791 => x"57",
          4792 => x"26",
          4793 => x"7b",
          4794 => x"0c",
          4795 => x"81",
          4796 => x"84",
          4797 => x"54",
          4798 => x"84",
          4799 => x"0d",
          4800 => x"0d",
          4801 => x"88",
          4802 => x"05",
          4803 => x"54",
          4804 => x"c5",
          4805 => x"56",
          4806 => x"d3",
          4807 => x"8b",
          4808 => x"d3",
          4809 => x"29",
          4810 => x"05",
          4811 => x"55",
          4812 => x"84",
          4813 => x"34",
          4814 => x"08",
          4815 => x"5f",
          4816 => x"51",
          4817 => x"3f",
          4818 => x"08",
          4819 => x"70",
          4820 => x"57",
          4821 => x"8b",
          4822 => x"82",
          4823 => x"06",
          4824 => x"56",
          4825 => x"38",
          4826 => x"05",
          4827 => x"7e",
          4828 => x"f0",
          4829 => x"84",
          4830 => x"67",
          4831 => x"2e",
          4832 => x"82",
          4833 => x"8b",
          4834 => x"75",
          4835 => x"80",
          4836 => x"81",
          4837 => x"2e",
          4838 => x"80",
          4839 => x"38",
          4840 => x"0a",
          4841 => x"ff",
          4842 => x"55",
          4843 => x"86",
          4844 => x"8a",
          4845 => x"89",
          4846 => x"2a",
          4847 => x"77",
          4848 => x"59",
          4849 => x"81",
          4850 => x"70",
          4851 => x"07",
          4852 => x"56",
          4853 => x"38",
          4854 => x"05",
          4855 => x"7e",
          4856 => x"80",
          4857 => x"81",
          4858 => x"8a",
          4859 => x"83",
          4860 => x"06",
          4861 => x"08",
          4862 => x"74",
          4863 => x"41",
          4864 => x"56",
          4865 => x"8a",
          4866 => x"61",
          4867 => x"55",
          4868 => x"27",
          4869 => x"93",
          4870 => x"80",
          4871 => x"38",
          4872 => x"70",
          4873 => x"43",
          4874 => x"95",
          4875 => x"06",
          4876 => x"2e",
          4877 => x"77",
          4878 => x"74",
          4879 => x"83",
          4880 => x"06",
          4881 => x"82",
          4882 => x"2e",
          4883 => x"78",
          4884 => x"2e",
          4885 => x"80",
          4886 => x"ae",
          4887 => x"2a",
          4888 => x"81",
          4889 => x"56",
          4890 => x"2e",
          4891 => x"77",
          4892 => x"81",
          4893 => x"79",
          4894 => x"70",
          4895 => x"5a",
          4896 => x"86",
          4897 => x"27",
          4898 => x"52",
          4899 => x"f9",
          4900 => x"d3",
          4901 => x"29",
          4902 => x"70",
          4903 => x"55",
          4904 => x"0b",
          4905 => x"08",
          4906 => x"05",
          4907 => x"ff",
          4908 => x"27",
          4909 => x"88",
          4910 => x"ae",
          4911 => x"2a",
          4912 => x"81",
          4913 => x"56",
          4914 => x"2e",
          4915 => x"77",
          4916 => x"81",
          4917 => x"79",
          4918 => x"70",
          4919 => x"5a",
          4920 => x"86",
          4921 => x"27",
          4922 => x"52",
          4923 => x"f9",
          4924 => x"d3",
          4925 => x"84",
          4926 => x"d3",
          4927 => x"f5",
          4928 => x"81",
          4929 => x"84",
          4930 => x"d3",
          4931 => x"71",
          4932 => x"83",
          4933 => x"5e",
          4934 => x"89",
          4935 => x"5c",
          4936 => x"1c",
          4937 => x"05",
          4938 => x"ff",
          4939 => x"70",
          4940 => x"31",
          4941 => x"57",
          4942 => x"83",
          4943 => x"06",
          4944 => x"1c",
          4945 => x"5c",
          4946 => x"1d",
          4947 => x"29",
          4948 => x"31",
          4949 => x"55",
          4950 => x"87",
          4951 => x"7c",
          4952 => x"7a",
          4953 => x"31",
          4954 => x"f8",
          4955 => x"d3",
          4956 => x"7d",
          4957 => x"81",
          4958 => x"81",
          4959 => x"83",
          4960 => x"80",
          4961 => x"87",
          4962 => x"81",
          4963 => x"fd",
          4964 => x"f8",
          4965 => x"2e",
          4966 => x"80",
          4967 => x"ff",
          4968 => x"d3",
          4969 => x"a0",
          4970 => x"38",
          4971 => x"74",
          4972 => x"86",
          4973 => x"fd",
          4974 => x"81",
          4975 => x"80",
          4976 => x"83",
          4977 => x"39",
          4978 => x"08",
          4979 => x"92",
          4980 => x"b8",
          4981 => x"59",
          4982 => x"27",
          4983 => x"86",
          4984 => x"55",
          4985 => x"09",
          4986 => x"38",
          4987 => x"f5",
          4988 => x"38",
          4989 => x"55",
          4990 => x"86",
          4991 => x"80",
          4992 => x"7a",
          4993 => x"b9",
          4994 => x"81",
          4995 => x"7a",
          4996 => x"8a",
          4997 => x"52",
          4998 => x"ff",
          4999 => x"79",
          5000 => x"7b",
          5001 => x"06",
          5002 => x"51",
          5003 => x"3f",
          5004 => x"1c",
          5005 => x"32",
          5006 => x"96",
          5007 => x"06",
          5008 => x"91",
          5009 => x"a1",
          5010 => x"55",
          5011 => x"ff",
          5012 => x"74",
          5013 => x"06",
          5014 => x"51",
          5015 => x"3f",
          5016 => x"52",
          5017 => x"ff",
          5018 => x"f8",
          5019 => x"34",
          5020 => x"1b",
          5021 => x"d9",
          5022 => x"52",
          5023 => x"ff",
          5024 => x"60",
          5025 => x"51",
          5026 => x"3f",
          5027 => x"09",
          5028 => x"cb",
          5029 => x"b2",
          5030 => x"c3",
          5031 => x"a0",
          5032 => x"52",
          5033 => x"ff",
          5034 => x"82",
          5035 => x"51",
          5036 => x"3f",
          5037 => x"1b",
          5038 => x"95",
          5039 => x"b2",
          5040 => x"a0",
          5041 => x"80",
          5042 => x"1c",
          5043 => x"80",
          5044 => x"93",
          5045 => x"c0",
          5046 => x"1b",
          5047 => x"82",
          5048 => x"52",
          5049 => x"ff",
          5050 => x"7c",
          5051 => x"06",
          5052 => x"51",
          5053 => x"3f",
          5054 => x"a4",
          5055 => x"0b",
          5056 => x"93",
          5057 => x"d4",
          5058 => x"51",
          5059 => x"3f",
          5060 => x"52",
          5061 => x"70",
          5062 => x"9f",
          5063 => x"54",
          5064 => x"52",
          5065 => x"9b",
          5066 => x"56",
          5067 => x"08",
          5068 => x"7d",
          5069 => x"81",
          5070 => x"38",
          5071 => x"86",
          5072 => x"52",
          5073 => x"9b",
          5074 => x"80",
          5075 => x"7a",
          5076 => x"ed",
          5077 => x"85",
          5078 => x"7a",
          5079 => x"8f",
          5080 => x"85",
          5081 => x"83",
          5082 => x"ff",
          5083 => x"ff",
          5084 => x"e8",
          5085 => x"9e",
          5086 => x"52",
          5087 => x"51",
          5088 => x"3f",
          5089 => x"52",
          5090 => x"9e",
          5091 => x"54",
          5092 => x"53",
          5093 => x"51",
          5094 => x"3f",
          5095 => x"16",
          5096 => x"7e",
          5097 => x"d8",
          5098 => x"80",
          5099 => x"ff",
          5100 => x"7f",
          5101 => x"7d",
          5102 => x"81",
          5103 => x"f8",
          5104 => x"ff",
          5105 => x"ff",
          5106 => x"51",
          5107 => x"3f",
          5108 => x"88",
          5109 => x"39",
          5110 => x"f8",
          5111 => x"2e",
          5112 => x"55",
          5113 => x"51",
          5114 => x"3f",
          5115 => x"57",
          5116 => x"83",
          5117 => x"76",
          5118 => x"7a",
          5119 => x"ff",
          5120 => x"81",
          5121 => x"82",
          5122 => x"80",
          5123 => x"84",
          5124 => x"51",
          5125 => x"3f",
          5126 => x"78",
          5127 => x"74",
          5128 => x"18",
          5129 => x"2e",
          5130 => x"79",
          5131 => x"2e",
          5132 => x"55",
          5133 => x"62",
          5134 => x"74",
          5135 => x"75",
          5136 => x"7e",
          5137 => x"b8",
          5138 => x"84",
          5139 => x"38",
          5140 => x"78",
          5141 => x"74",
          5142 => x"56",
          5143 => x"93",
          5144 => x"66",
          5145 => x"26",
          5146 => x"56",
          5147 => x"83",
          5148 => x"64",
          5149 => x"77",
          5150 => x"84",
          5151 => x"52",
          5152 => x"9d",
          5153 => x"d4",
          5154 => x"51",
          5155 => x"3f",
          5156 => x"55",
          5157 => x"81",
          5158 => x"34",
          5159 => x"16",
          5160 => x"16",
          5161 => x"16",
          5162 => x"05",
          5163 => x"c1",
          5164 => x"fe",
          5165 => x"fe",
          5166 => x"34",
          5167 => x"08",
          5168 => x"07",
          5169 => x"16",
          5170 => x"84",
          5171 => x"34",
          5172 => x"c6",
          5173 => x"9c",
          5174 => x"52",
          5175 => x"51",
          5176 => x"3f",
          5177 => x"53",
          5178 => x"51",
          5179 => x"3f",
          5180 => x"d3",
          5181 => x"38",
          5182 => x"52",
          5183 => x"99",
          5184 => x"56",
          5185 => x"08",
          5186 => x"39",
          5187 => x"39",
          5188 => x"39",
          5189 => x"08",
          5190 => x"d3",
          5191 => x"3d",
          5192 => x"3d",
          5193 => x"71",
          5194 => x"8e",
          5195 => x"29",
          5196 => x"05",
          5197 => x"04",
          5198 => x"51",
          5199 => x"81",
          5200 => x"80",
          5201 => x"c5",
          5202 => x"f2",
          5203 => x"e0",
          5204 => x"39",
          5205 => x"51",
          5206 => x"81",
          5207 => x"80",
          5208 => x"c6",
          5209 => x"d6",
          5210 => x"a4",
          5211 => x"39",
          5212 => x"51",
          5213 => x"81",
          5214 => x"80",
          5215 => x"c6",
          5216 => x"39",
          5217 => x"51",
          5218 => x"c7",
          5219 => x"39",
          5220 => x"51",
          5221 => x"c7",
          5222 => x"39",
          5223 => x"51",
          5224 => x"c8",
          5225 => x"39",
          5226 => x"51",
          5227 => x"c8",
          5228 => x"39",
          5229 => x"51",
          5230 => x"c8",
          5231 => x"87",
          5232 => x"3d",
          5233 => x"3d",
          5234 => x"56",
          5235 => x"e7",
          5236 => x"74",
          5237 => x"e8",
          5238 => x"39",
          5239 => x"74",
          5240 => x"96",
          5241 => x"84",
          5242 => x"51",
          5243 => x"3f",
          5244 => x"08",
          5245 => x"75",
          5246 => x"f4",
          5247 => x"a0",
          5248 => x"0d",
          5249 => x"0d",
          5250 => x"02",
          5251 => x"c7",
          5252 => x"73",
          5253 => x"5d",
          5254 => x"5c",
          5255 => x"81",
          5256 => x"ff",
          5257 => x"81",
          5258 => x"ff",
          5259 => x"80",
          5260 => x"27",
          5261 => x"79",
          5262 => x"38",
          5263 => x"a7",
          5264 => x"39",
          5265 => x"72",
          5266 => x"38",
          5267 => x"81",
          5268 => x"ff",
          5269 => x"89",
          5270 => x"b0",
          5271 => x"dc",
          5272 => x"55",
          5273 => x"74",
          5274 => x"78",
          5275 => x"72",
          5276 => x"c9",
          5277 => x"8c",
          5278 => x"39",
          5279 => x"51",
          5280 => x"3f",
          5281 => x"a1",
          5282 => x"53",
          5283 => x"8e",
          5284 => x"52",
          5285 => x"51",
          5286 => x"3f",
          5287 => x"c9",
          5288 => x"86",
          5289 => x"15",
          5290 => x"fe",
          5291 => x"ff",
          5292 => x"c9",
          5293 => x"86",
          5294 => x"55",
          5295 => x"aa",
          5296 => x"70",
          5297 => x"26",
          5298 => x"9f",
          5299 => x"38",
          5300 => x"8b",
          5301 => x"fe",
          5302 => x"73",
          5303 => x"a0",
          5304 => x"d9",
          5305 => x"55",
          5306 => x"c9",
          5307 => x"85",
          5308 => x"16",
          5309 => x"56",
          5310 => x"3f",
          5311 => x"08",
          5312 => x"98",
          5313 => x"74",
          5314 => x"81",
          5315 => x"fe",
          5316 => x"81",
          5317 => x"98",
          5318 => x"2c",
          5319 => x"70",
          5320 => x"07",
          5321 => x"56",
          5322 => x"74",
          5323 => x"38",
          5324 => x"74",
          5325 => x"81",
          5326 => x"80",
          5327 => x"7a",
          5328 => x"76",
          5329 => x"38",
          5330 => x"81",
          5331 => x"8d",
          5332 => x"ec",
          5333 => x"02",
          5334 => x"e3",
          5335 => x"72",
          5336 => x"07",
          5337 => x"87",
          5338 => x"07",
          5339 => x"5a",
          5340 => x"57",
          5341 => x"38",
          5342 => x"52",
          5343 => x"52",
          5344 => x"3f",
          5345 => x"08",
          5346 => x"84",
          5347 => x"81",
          5348 => x"87",
          5349 => x"0c",
          5350 => x"08",
          5351 => x"d4",
          5352 => x"80",
          5353 => x"76",
          5354 => x"3f",
          5355 => x"08",
          5356 => x"84",
          5357 => x"7a",
          5358 => x"2e",
          5359 => x"19",
          5360 => x"59",
          5361 => x"3d",
          5362 => x"cc",
          5363 => x"30",
          5364 => x"80",
          5365 => x"79",
          5366 => x"38",
          5367 => x"90",
          5368 => x"cc",
          5369 => x"98",
          5370 => x"78",
          5371 => x"3f",
          5372 => x"81",
          5373 => x"96",
          5374 => x"f9",
          5375 => x"02",
          5376 => x"05",
          5377 => x"ff",
          5378 => x"7a",
          5379 => x"fe",
          5380 => x"d3",
          5381 => x"38",
          5382 => x"88",
          5383 => x"2e",
          5384 => x"39",
          5385 => x"54",
          5386 => x"53",
          5387 => x"51",
          5388 => x"d3",
          5389 => x"83",
          5390 => x"76",
          5391 => x"0c",
          5392 => x"04",
          5393 => x"02",
          5394 => x"81",
          5395 => x"81",
          5396 => x"55",
          5397 => x"3f",
          5398 => x"22",
          5399 => x"e4",
          5400 => x"e8",
          5401 => x"f4",
          5402 => x"a5",
          5403 => x"c9",
          5404 => x"88",
          5405 => x"80",
          5406 => x"fe",
          5407 => x"86",
          5408 => x"fe",
          5409 => x"c0",
          5410 => x"53",
          5411 => x"3f",
          5412 => x"f6",
          5413 => x"ca",
          5414 => x"f8",
          5415 => x"51",
          5416 => x"3f",
          5417 => x"70",
          5418 => x"52",
          5419 => x"95",
          5420 => x"fe",
          5421 => x"81",
          5422 => x"fe",
          5423 => x"80",
          5424 => x"df",
          5425 => x"2a",
          5426 => x"51",
          5427 => x"2e",
          5428 => x"51",
          5429 => x"3f",
          5430 => x"51",
          5431 => x"3f",
          5432 => x"f5",
          5433 => x"83",
          5434 => x"06",
          5435 => x"80",
          5436 => x"81",
          5437 => x"ab",
          5438 => x"d8",
          5439 => x"a3",
          5440 => x"fe",
          5441 => x"72",
          5442 => x"81",
          5443 => x"71",
          5444 => x"38",
          5445 => x"f5",
          5446 => x"ca",
          5447 => x"f7",
          5448 => x"51",
          5449 => x"3f",
          5450 => x"70",
          5451 => x"52",
          5452 => x"95",
          5453 => x"fe",
          5454 => x"81",
          5455 => x"fe",
          5456 => x"80",
          5457 => x"db",
          5458 => x"2a",
          5459 => x"51",
          5460 => x"2e",
          5461 => x"51",
          5462 => x"3f",
          5463 => x"51",
          5464 => x"3f",
          5465 => x"f4",
          5466 => x"87",
          5467 => x"06",
          5468 => x"80",
          5469 => x"81",
          5470 => x"a7",
          5471 => x"a8",
          5472 => x"9f",
          5473 => x"fe",
          5474 => x"72",
          5475 => x"81",
          5476 => x"71",
          5477 => x"38",
          5478 => x"f4",
          5479 => x"cb",
          5480 => x"f5",
          5481 => x"51",
          5482 => x"3f",
          5483 => x"3f",
          5484 => x"04",
          5485 => x"78",
          5486 => x"55",
          5487 => x"80",
          5488 => x"38",
          5489 => x"77",
          5490 => x"33",
          5491 => x"39",
          5492 => x"80",
          5493 => x"81",
          5494 => x"57",
          5495 => x"2e",
          5496 => x"53",
          5497 => x"84",
          5498 => x"38",
          5499 => x"06",
          5500 => x"2e",
          5501 => x"88",
          5502 => x"70",
          5503 => x"34",
          5504 => x"90",
          5505 => x"c4",
          5506 => x"53",
          5507 => x"55",
          5508 => x"3f",
          5509 => x"08",
          5510 => x"15",
          5511 => x"81",
          5512 => x"38",
          5513 => x"81",
          5514 => x"53",
          5515 => x"d2",
          5516 => x"72",
          5517 => x"0c",
          5518 => x"04",
          5519 => x"80",
          5520 => x"ea",
          5521 => x"5c",
          5522 => x"51",
          5523 => x"3f",
          5524 => x"08",
          5525 => x"59",
          5526 => x"09",
          5527 => x"38",
          5528 => x"52",
          5529 => x"52",
          5530 => x"ca",
          5531 => x"78",
          5532 => x"b4",
          5533 => x"e3",
          5534 => x"84",
          5535 => x"88",
          5536 => x"80",
          5537 => x"39",
          5538 => x"5c",
          5539 => x"51",
          5540 => x"3f",
          5541 => x"46",
          5542 => x"53",
          5543 => x"51",
          5544 => x"3f",
          5545 => x"64",
          5546 => x"ce",
          5547 => x"fe",
          5548 => x"fd",
          5549 => x"d3",
          5550 => x"2b",
          5551 => x"51",
          5552 => x"c3",
          5553 => x"38",
          5554 => x"24",
          5555 => x"78",
          5556 => x"bc",
          5557 => x"24",
          5558 => x"82",
          5559 => x"38",
          5560 => x"8a",
          5561 => x"2e",
          5562 => x"8d",
          5563 => x"84",
          5564 => x"38",
          5565 => x"82",
          5566 => x"f9",
          5567 => x"c0",
          5568 => x"38",
          5569 => x"24",
          5570 => x"b0",
          5571 => x"38",
          5572 => x"84",
          5573 => x"dd",
          5574 => x"c1",
          5575 => x"38",
          5576 => x"2e",
          5577 => x"8c",
          5578 => x"80",
          5579 => x"ba",
          5580 => x"f8",
          5581 => x"78",
          5582 => x"8a",
          5583 => x"80",
          5584 => x"38",
          5585 => x"2e",
          5586 => x"8c",
          5587 => x"80",
          5588 => x"dc",
          5589 => x"d5",
          5590 => x"38",
          5591 => x"78",
          5592 => x"8b",
          5593 => x"81",
          5594 => x"38",
          5595 => x"2e",
          5596 => x"78",
          5597 => x"8b",
          5598 => x"f9",
          5599 => x"85",
          5600 => x"38",
          5601 => x"2e",
          5602 => x"8b",
          5603 => x"3d",
          5604 => x"53",
          5605 => x"51",
          5606 => x"3f",
          5607 => x"08",
          5608 => x"cc",
          5609 => x"c7",
          5610 => x"fe",
          5611 => x"fe",
          5612 => x"ff",
          5613 => x"81",
          5614 => x"80",
          5615 => x"81",
          5616 => x"38",
          5617 => x"80",
          5618 => x"52",
          5619 => x"05",
          5620 => x"87",
          5621 => x"d3",
          5622 => x"ff",
          5623 => x"8e",
          5624 => x"cc",
          5625 => x"d4",
          5626 => x"fd",
          5627 => x"cc",
          5628 => x"d2",
          5629 => x"fe",
          5630 => x"fe",
          5631 => x"ff",
          5632 => x"81",
          5633 => x"80",
          5634 => x"38",
          5635 => x"52",
          5636 => x"05",
          5637 => x"8b",
          5638 => x"d3",
          5639 => x"81",
          5640 => x"8a",
          5641 => x"3d",
          5642 => x"53",
          5643 => x"51",
          5644 => x"3f",
          5645 => x"08",
          5646 => x"38",
          5647 => x"fc",
          5648 => x"3d",
          5649 => x"53",
          5650 => x"51",
          5651 => x"3f",
          5652 => x"08",
          5653 => x"d3",
          5654 => x"63",
          5655 => x"fc",
          5656 => x"ff",
          5657 => x"02",
          5658 => x"33",
          5659 => x"63",
          5660 => x"81",
          5661 => x"51",
          5662 => x"3f",
          5663 => x"08",
          5664 => x"81",
          5665 => x"fe",
          5666 => x"81",
          5667 => x"39",
          5668 => x"f8",
          5669 => x"ea",
          5670 => x"d3",
          5671 => x"3d",
          5672 => x"52",
          5673 => x"8e",
          5674 => x"81",
          5675 => x"52",
          5676 => x"9f",
          5677 => x"39",
          5678 => x"f8",
          5679 => x"ea",
          5680 => x"d3",
          5681 => x"3d",
          5682 => x"52",
          5683 => x"e6",
          5684 => x"84",
          5685 => x"fe",
          5686 => x"5a",
          5687 => x"3f",
          5688 => x"08",
          5689 => x"f8",
          5690 => x"fe",
          5691 => x"81",
          5692 => x"81",
          5693 => x"80",
          5694 => x"81",
          5695 => x"81",
          5696 => x"78",
          5697 => x"7a",
          5698 => x"3f",
          5699 => x"08",
          5700 => x"f8",
          5701 => x"84",
          5702 => x"86",
          5703 => x"39",
          5704 => x"f4",
          5705 => x"f8",
          5706 => x"80",
          5707 => x"d3",
          5708 => x"2e",
          5709 => x"b7",
          5710 => x"11",
          5711 => x"05",
          5712 => x"d1",
          5713 => x"84",
          5714 => x"fa",
          5715 => x"3d",
          5716 => x"53",
          5717 => x"51",
          5718 => x"3f",
          5719 => x"08",
          5720 => x"d3",
          5721 => x"81",
          5722 => x"fe",
          5723 => x"63",
          5724 => x"79",
          5725 => x"38",
          5726 => x"7a",
          5727 => x"5c",
          5728 => x"26",
          5729 => x"cc",
          5730 => x"ba",
          5731 => x"fe",
          5732 => x"fe",
          5733 => x"fe",
          5734 => x"81",
          5735 => x"80",
          5736 => x"d0",
          5737 => x"78",
          5738 => x"38",
          5739 => x"08",
          5740 => x"81",
          5741 => x"59",
          5742 => x"88",
          5743 => x"88",
          5744 => x"39",
          5745 => x"33",
          5746 => x"38",
          5747 => x"33",
          5748 => x"2e",
          5749 => x"d0",
          5750 => x"89",
          5751 => x"a0",
          5752 => x"05",
          5753 => x"fe",
          5754 => x"fe",
          5755 => x"fe",
          5756 => x"81",
          5757 => x"80",
          5758 => x"d0",
          5759 => x"78",
          5760 => x"38",
          5761 => x"08",
          5762 => x"81",
          5763 => x"59",
          5764 => x"88",
          5765 => x"8c",
          5766 => x"39",
          5767 => x"33",
          5768 => x"38",
          5769 => x"33",
          5770 => x"2e",
          5771 => x"d0",
          5772 => x"88",
          5773 => x"a0",
          5774 => x"43",
          5775 => x"ec",
          5776 => x"f8",
          5777 => x"fe",
          5778 => x"d3",
          5779 => x"2e",
          5780 => x"62",
          5781 => x"88",
          5782 => x"81",
          5783 => x"2e",
          5784 => x"80",
          5785 => x"79",
          5786 => x"38",
          5787 => x"cd",
          5788 => x"f6",
          5789 => x"55",
          5790 => x"53",
          5791 => x"51",
          5792 => x"81",
          5793 => x"84",
          5794 => x"3d",
          5795 => x"53",
          5796 => x"51",
          5797 => x"3f",
          5798 => x"08",
          5799 => x"ec",
          5800 => x"fe",
          5801 => x"fe",
          5802 => x"fe",
          5803 => x"81",
          5804 => x"80",
          5805 => x"63",
          5806 => x"cb",
          5807 => x"34",
          5808 => x"44",
          5809 => x"f0",
          5810 => x"f8",
          5811 => x"fd",
          5812 => x"d3",
          5813 => x"38",
          5814 => x"63",
          5815 => x"52",
          5816 => x"51",
          5817 => x"3f",
          5818 => x"79",
          5819 => x"8a",
          5820 => x"79",
          5821 => x"ae",
          5822 => x"38",
          5823 => x"a0",
          5824 => x"fe",
          5825 => x"fe",
          5826 => x"fe",
          5827 => x"81",
          5828 => x"80",
          5829 => x"63",
          5830 => x"cb",
          5831 => x"34",
          5832 => x"44",
          5833 => x"81",
          5834 => x"fe",
          5835 => x"ff",
          5836 => x"3d",
          5837 => x"53",
          5838 => x"51",
          5839 => x"3f",
          5840 => x"08",
          5841 => x"c4",
          5842 => x"fe",
          5843 => x"fe",
          5844 => x"fe",
          5845 => x"81",
          5846 => x"80",
          5847 => x"60",
          5848 => x"05",
          5849 => x"82",
          5850 => x"78",
          5851 => x"fe",
          5852 => x"fe",
          5853 => x"fe",
          5854 => x"81",
          5855 => x"df",
          5856 => x"39",
          5857 => x"54",
          5858 => x"bc",
          5859 => x"90",
          5860 => x"52",
          5861 => x"fa",
          5862 => x"45",
          5863 => x"78",
          5864 => x"e8",
          5865 => x"26",
          5866 => x"84",
          5867 => x"39",
          5868 => x"e4",
          5869 => x"f8",
          5870 => x"fd",
          5871 => x"d3",
          5872 => x"2e",
          5873 => x"59",
          5874 => x"22",
          5875 => x"05",
          5876 => x"41",
          5877 => x"81",
          5878 => x"fe",
          5879 => x"ff",
          5880 => x"3d",
          5881 => x"53",
          5882 => x"51",
          5883 => x"3f",
          5884 => x"08",
          5885 => x"94",
          5886 => x"fe",
          5887 => x"fe",
          5888 => x"fe",
          5889 => x"81",
          5890 => x"80",
          5891 => x"60",
          5892 => x"59",
          5893 => x"41",
          5894 => x"e4",
          5895 => x"f8",
          5896 => x"fc",
          5897 => x"d3",
          5898 => x"38",
          5899 => x"60",
          5900 => x"52",
          5901 => x"51",
          5902 => x"3f",
          5903 => x"79",
          5904 => x"b6",
          5905 => x"79",
          5906 => x"ae",
          5907 => x"38",
          5908 => x"a8",
          5909 => x"fe",
          5910 => x"fe",
          5911 => x"fe",
          5912 => x"81",
          5913 => x"80",
          5914 => x"7f",
          5915 => x"81",
          5916 => x"fe",
          5917 => x"60",
          5918 => x"59",
          5919 => x"41",
          5920 => x"81",
          5921 => x"fe",
          5922 => x"ff",
          5923 => x"cd",
          5924 => x"f2",
          5925 => x"51",
          5926 => x"3f",
          5927 => x"81",
          5928 => x"fe",
          5929 => x"a2",
          5930 => x"e8",
          5931 => x"39",
          5932 => x"0b",
          5933 => x"84",
          5934 => x"81",
          5935 => x"94",
          5936 => x"ce",
          5937 => x"f1",
          5938 => x"c0",
          5939 => x"98",
          5940 => x"e8",
          5941 => x"83",
          5942 => x"94",
          5943 => x"80",
          5944 => x"c0",
          5945 => x"f3",
          5946 => x"3d",
          5947 => x"53",
          5948 => x"51",
          5949 => x"3f",
          5950 => x"08",
          5951 => x"8c",
          5952 => x"81",
          5953 => x"fe",
          5954 => x"63",
          5955 => x"b7",
          5956 => x"11",
          5957 => x"05",
          5958 => x"f9",
          5959 => x"84",
          5960 => x"f2",
          5961 => x"52",
          5962 => x"51",
          5963 => x"3f",
          5964 => x"2d",
          5965 => x"08",
          5966 => x"84",
          5967 => x"f2",
          5968 => x"d3",
          5969 => x"81",
          5970 => x"fe",
          5971 => x"f2",
          5972 => x"cf",
          5973 => x"f0",
          5974 => x"c5",
          5975 => x"ac",
          5976 => x"9c",
          5977 => x"d4",
          5978 => x"ff",
          5979 => x"ec",
          5980 => x"98",
          5981 => x"33",
          5982 => x"80",
          5983 => x"38",
          5984 => x"80",
          5985 => x"80",
          5986 => x"38",
          5987 => x"f8",
          5988 => x"e0",
          5989 => x"cf",
          5990 => x"d3",
          5991 => x"81",
          5992 => x"80",
          5993 => x"b8",
          5994 => x"70",
          5995 => x"f6",
          5996 => x"d0",
          5997 => x"d3",
          5998 => x"56",
          5999 => x"46",
          6000 => x"80",
          6001 => x"80",
          6002 => x"80",
          6003 => x"ec",
          6004 => x"d3",
          6005 => x"7c",
          6006 => x"81",
          6007 => x"78",
          6008 => x"ff",
          6009 => x"06",
          6010 => x"81",
          6011 => x"fe",
          6012 => x"f1",
          6013 => x"3d",
          6014 => x"81",
          6015 => x"9b",
          6016 => x"0b",
          6017 => x"8c",
          6018 => x"86",
          6019 => x"c0",
          6020 => x"8c",
          6021 => x"87",
          6022 => x"0c",
          6023 => x"0b",
          6024 => x"94",
          6025 => x"0b",
          6026 => x"0c",
          6027 => x"81",
          6028 => x"fe",
          6029 => x"fe",
          6030 => x"81",
          6031 => x"fe",
          6032 => x"81",
          6033 => x"fe",
          6034 => x"81",
          6035 => x"fe",
          6036 => x"81",
          6037 => x"3f",
          6038 => x"80",
          6039 => x"00",
          6040 => x"ff",
          6041 => x"ff",
          6042 => x"ff",
          6043 => x"00",
          6044 => x"00",
          6045 => x"00",
          6046 => x"00",
          6047 => x"00",
          6048 => x"00",
          6049 => x"00",
          6050 => x"00",
          6051 => x"00",
          6052 => x"00",
          6053 => x"00",
          6054 => x"00",
          6055 => x"00",
          6056 => x"00",
          6057 => x"00",
          6058 => x"00",
          6059 => x"00",
          6060 => x"00",
          6061 => x"00",
          6062 => x"00",
          6063 => x"00",
          6064 => x"00",
          6065 => x"00",
          6066 => x"00",
          6067 => x"00",
          6068 => x"25",
          6069 => x"64",
          6070 => x"20",
          6071 => x"25",
          6072 => x"64",
          6073 => x"25",
          6074 => x"53",
          6075 => x"43",
          6076 => x"69",
          6077 => x"61",
          6078 => x"6e",
          6079 => x"20",
          6080 => x"6f",
          6081 => x"6f",
          6082 => x"6f",
          6083 => x"67",
          6084 => x"3a",
          6085 => x"76",
          6086 => x"73",
          6087 => x"70",
          6088 => x"65",
          6089 => x"64",
          6090 => x"20",
          6091 => x"49",
          6092 => x"20",
          6093 => x"4d",
          6094 => x"74",
          6095 => x"3d",
          6096 => x"58",
          6097 => x"69",
          6098 => x"25",
          6099 => x"29",
          6100 => x"20",
          6101 => x"42",
          6102 => x"20",
          6103 => x"61",
          6104 => x"25",
          6105 => x"2c",
          6106 => x"7a",
          6107 => x"30",
          6108 => x"2e",
          6109 => x"20",
          6110 => x"52",
          6111 => x"28",
          6112 => x"72",
          6113 => x"30",
          6114 => x"20",
          6115 => x"65",
          6116 => x"38",
          6117 => x"0a",
          6118 => x"20",
          6119 => x"49",
          6120 => x"4c",
          6121 => x"20",
          6122 => x"50",
          6123 => x"00",
          6124 => x"20",
          6125 => x"53",
          6126 => x"00",
          6127 => x"20",
          6128 => x"53",
          6129 => x"61",
          6130 => x"28",
          6131 => x"69",
          6132 => x"3d",
          6133 => x"58",
          6134 => x"00",
          6135 => x"20",
          6136 => x"49",
          6137 => x"52",
          6138 => x"54",
          6139 => x"4e",
          6140 => x"4c",
          6141 => x"0a",
          6142 => x"20",
          6143 => x"54",
          6144 => x"52",
          6145 => x"54",
          6146 => x"72",
          6147 => x"30",
          6148 => x"2e",
          6149 => x"41",
          6150 => x"65",
          6151 => x"73",
          6152 => x"20",
          6153 => x"43",
          6154 => x"52",
          6155 => x"74",
          6156 => x"63",
          6157 => x"20",
          6158 => x"72",
          6159 => x"20",
          6160 => x"30",
          6161 => x"00",
          6162 => x"20",
          6163 => x"43",
          6164 => x"4d",
          6165 => x"72",
          6166 => x"74",
          6167 => x"20",
          6168 => x"72",
          6169 => x"20",
          6170 => x"30",
          6171 => x"00",
          6172 => x"20",
          6173 => x"53",
          6174 => x"6b",
          6175 => x"61",
          6176 => x"41",
          6177 => x"65",
          6178 => x"20",
          6179 => x"20",
          6180 => x"30",
          6181 => x"00",
          6182 => x"20",
          6183 => x"5a",
          6184 => x"49",
          6185 => x"20",
          6186 => x"20",
          6187 => x"20",
          6188 => x"20",
          6189 => x"20",
          6190 => x"30",
          6191 => x"00",
          6192 => x"20",
          6193 => x"53",
          6194 => x"65",
          6195 => x"6c",
          6196 => x"20",
          6197 => x"71",
          6198 => x"20",
          6199 => x"20",
          6200 => x"30",
          6201 => x"00",
          6202 => x"53",
          6203 => x"6c",
          6204 => x"4d",
          6205 => x"75",
          6206 => x"46",
          6207 => x"00",
          6208 => x"45",
          6209 => x"45",
          6210 => x"69",
          6211 => x"55",
          6212 => x"6f",
          6213 => x"53",
          6214 => x"22",
          6215 => x"3a",
          6216 => x"3e",
          6217 => x"7c",
          6218 => x"46",
          6219 => x"46",
          6220 => x"32",
          6221 => x"eb",
          6222 => x"53",
          6223 => x"35",
          6224 => x"4e",
          6225 => x"41",
          6226 => x"20",
          6227 => x"41",
          6228 => x"20",
          6229 => x"4e",
          6230 => x"41",
          6231 => x"20",
          6232 => x"41",
          6233 => x"20",
          6234 => x"00",
          6235 => x"00",
          6236 => x"00",
          6237 => x"00",
          6238 => x"80",
          6239 => x"8e",
          6240 => x"45",
          6241 => x"49",
          6242 => x"90",
          6243 => x"99",
          6244 => x"59",
          6245 => x"9c",
          6246 => x"41",
          6247 => x"a5",
          6248 => x"a8",
          6249 => x"ac",
          6250 => x"b0",
          6251 => x"b4",
          6252 => x"b8",
          6253 => x"bc",
          6254 => x"c0",
          6255 => x"c4",
          6256 => x"c8",
          6257 => x"cc",
          6258 => x"d0",
          6259 => x"d4",
          6260 => x"d8",
          6261 => x"dc",
          6262 => x"e0",
          6263 => x"e4",
          6264 => x"e8",
          6265 => x"ec",
          6266 => x"f0",
          6267 => x"f4",
          6268 => x"f8",
          6269 => x"fc",
          6270 => x"2b",
          6271 => x"3d",
          6272 => x"5c",
          6273 => x"3c",
          6274 => x"7f",
          6275 => x"00",
          6276 => x"00",
          6277 => x"01",
          6278 => x"00",
          6279 => x"00",
          6280 => x"00",
          6281 => x"00",
          6282 => x"00",
          6283 => x"64",
          6284 => x"74",
          6285 => x"64",
          6286 => x"74",
          6287 => x"66",
          6288 => x"74",
          6289 => x"66",
          6290 => x"64",
          6291 => x"66",
          6292 => x"63",
          6293 => x"6d",
          6294 => x"61",
          6295 => x"6d",
          6296 => x"70",
          6297 => x"6d",
          6298 => x"6d",
          6299 => x"6d",
          6300 => x"68",
          6301 => x"68",
          6302 => x"68",
          6303 => x"68",
          6304 => x"63",
          6305 => x"00",
          6306 => x"6a",
          6307 => x"72",
          6308 => x"61",
          6309 => x"72",
          6310 => x"74",
          6311 => x"69",
          6312 => x"00",
          6313 => x"74",
          6314 => x"00",
          6315 => x"44",
          6316 => x"20",
          6317 => x"6f",
          6318 => x"49",
          6319 => x"72",
          6320 => x"20",
          6321 => x"6f",
          6322 => x"00",
          6323 => x"44",
          6324 => x"20",
          6325 => x"20",
          6326 => x"64",
          6327 => x"00",
          6328 => x"4e",
          6329 => x"69",
          6330 => x"66",
          6331 => x"64",
          6332 => x"4e",
          6333 => x"61",
          6334 => x"66",
          6335 => x"64",
          6336 => x"49",
          6337 => x"6c",
          6338 => x"66",
          6339 => x"6e",
          6340 => x"2e",
          6341 => x"41",
          6342 => x"73",
          6343 => x"65",
          6344 => x"64",
          6345 => x"46",
          6346 => x"20",
          6347 => x"65",
          6348 => x"20",
          6349 => x"73",
          6350 => x"0a",
          6351 => x"46",
          6352 => x"20",
          6353 => x"64",
          6354 => x"69",
          6355 => x"6c",
          6356 => x"0a",
          6357 => x"53",
          6358 => x"73",
          6359 => x"69",
          6360 => x"70",
          6361 => x"65",
          6362 => x"64",
          6363 => x"44",
          6364 => x"65",
          6365 => x"6d",
          6366 => x"20",
          6367 => x"69",
          6368 => x"6c",
          6369 => x"0a",
          6370 => x"44",
          6371 => x"20",
          6372 => x"20",
          6373 => x"62",
          6374 => x"2e",
          6375 => x"4e",
          6376 => x"6f",
          6377 => x"74",
          6378 => x"65",
          6379 => x"6c",
          6380 => x"73",
          6381 => x"20",
          6382 => x"6e",
          6383 => x"6e",
          6384 => x"73",
          6385 => x"00",
          6386 => x"46",
          6387 => x"61",
          6388 => x"62",
          6389 => x"65",
          6390 => x"00",
          6391 => x"54",
          6392 => x"6f",
          6393 => x"20",
          6394 => x"72",
          6395 => x"6f",
          6396 => x"61",
          6397 => x"6c",
          6398 => x"2e",
          6399 => x"46",
          6400 => x"20",
          6401 => x"6c",
          6402 => x"65",
          6403 => x"00",
          6404 => x"49",
          6405 => x"66",
          6406 => x"69",
          6407 => x"20",
          6408 => x"6f",
          6409 => x"0a",
          6410 => x"54",
          6411 => x"6d",
          6412 => x"20",
          6413 => x"6e",
          6414 => x"6c",
          6415 => x"0a",
          6416 => x"50",
          6417 => x"6d",
          6418 => x"72",
          6419 => x"6e",
          6420 => x"72",
          6421 => x"2e",
          6422 => x"53",
          6423 => x"65",
          6424 => x"0a",
          6425 => x"55",
          6426 => x"6f",
          6427 => x"65",
          6428 => x"72",
          6429 => x"0a",
          6430 => x"20",
          6431 => x"65",
          6432 => x"73",
          6433 => x"20",
          6434 => x"20",
          6435 => x"65",
          6436 => x"65",
          6437 => x"00",
          6438 => x"25",
          6439 => x"00",
          6440 => x"3a",
          6441 => x"25",
          6442 => x"00",
          6443 => x"20",
          6444 => x"20",
          6445 => x"00",
          6446 => x"25",
          6447 => x"00",
          6448 => x"20",
          6449 => x"20",
          6450 => x"7c",
          6451 => x"72",
          6452 => x"00",
          6453 => x"5a",
          6454 => x"41",
          6455 => x"0a",
          6456 => x"25",
          6457 => x"00",
          6458 => x"31",
          6459 => x"37",
          6460 => x"31",
          6461 => x"76",
          6462 => x"00",
          6463 => x"20",
          6464 => x"2c",
          6465 => x"76",
          6466 => x"32",
          6467 => x"25",
          6468 => x"73",
          6469 => x"0a",
          6470 => x"5a",
          6471 => x"41",
          6472 => x"74",
          6473 => x"75",
          6474 => x"48",
          6475 => x"6c",
          6476 => x"00",
          6477 => x"54",
          6478 => x"72",
          6479 => x"74",
          6480 => x"75",
          6481 => x"00",
          6482 => x"50",
          6483 => x"69",
          6484 => x"72",
          6485 => x"74",
          6486 => x"49",
          6487 => x"4c",
          6488 => x"20",
          6489 => x"65",
          6490 => x"70",
          6491 => x"49",
          6492 => x"4c",
          6493 => x"20",
          6494 => x"65",
          6495 => x"70",
          6496 => x"55",
          6497 => x"30",
          6498 => x"20",
          6499 => x"65",
          6500 => x"70",
          6501 => x"55",
          6502 => x"30",
          6503 => x"20",
          6504 => x"65",
          6505 => x"70",
          6506 => x"55",
          6507 => x"31",
          6508 => x"20",
          6509 => x"65",
          6510 => x"70",
          6511 => x"55",
          6512 => x"31",
          6513 => x"20",
          6514 => x"65",
          6515 => x"70",
          6516 => x"53",
          6517 => x"69",
          6518 => x"75",
          6519 => x"69",
          6520 => x"2e",
          6521 => x"00",
          6522 => x"45",
          6523 => x"6c",
          6524 => x"20",
          6525 => x"65",
          6526 => x"2e",
          6527 => x"30",
          6528 => x"46",
          6529 => x"65",
          6530 => x"6f",
          6531 => x"69",
          6532 => x"6c",
          6533 => x"20",
          6534 => x"63",
          6535 => x"20",
          6536 => x"70",
          6537 => x"73",
          6538 => x"6e",
          6539 => x"6d",
          6540 => x"61",
          6541 => x"2e",
          6542 => x"2a",
          6543 => x"42",
          6544 => x"64",
          6545 => x"20",
          6546 => x"0a",
          6547 => x"49",
          6548 => x"69",
          6549 => x"73",
          6550 => x"0a",
          6551 => x"46",
          6552 => x"65",
          6553 => x"6f",
          6554 => x"69",
          6555 => x"6c",
          6556 => x"2e",
          6557 => x"72",
          6558 => x"64",
          6559 => x"25",
          6560 => x"43",
          6561 => x"72",
          6562 => x"2e",
          6563 => x"44",
          6564 => x"20",
          6565 => x"6f",
          6566 => x"00",
          6567 => x"0a",
          6568 => x"70",
          6569 => x"65",
          6570 => x"25",
          6571 => x"20",
          6572 => x"58",
          6573 => x"3f",
          6574 => x"00",
          6575 => x"25",
          6576 => x"20",
          6577 => x"58",
          6578 => x"25",
          6579 => x"20",
          6580 => x"58",
          6581 => x"44",
          6582 => x"62",
          6583 => x"67",
          6584 => x"74",
          6585 => x"75",
          6586 => x"0a",
          6587 => x"45",
          6588 => x"6c",
          6589 => x"20",
          6590 => x"65",
          6591 => x"70",
          6592 => x"00",
          6593 => x"44",
          6594 => x"62",
          6595 => x"20",
          6596 => x"74",
          6597 => x"66",
          6598 => x"45",
          6599 => x"6c",
          6600 => x"20",
          6601 => x"74",
          6602 => x"66",
          6603 => x"45",
          6604 => x"75",
          6605 => x"67",
          6606 => x"64",
          6607 => x"20",
          6608 => x"78",
          6609 => x"2e",
          6610 => x"43",
          6611 => x"69",
          6612 => x"63",
          6613 => x"20",
          6614 => x"30",
          6615 => x"2e",
          6616 => x"00",
          6617 => x"43",
          6618 => x"20",
          6619 => x"75",
          6620 => x"64",
          6621 => x"64",
          6622 => x"25",
          6623 => x"0a",
          6624 => x"52",
          6625 => x"61",
          6626 => x"6e",
          6627 => x"70",
          6628 => x"63",
          6629 => x"6f",
          6630 => x"2e",
          6631 => x"43",
          6632 => x"20",
          6633 => x"6f",
          6634 => x"6e",
          6635 => x"2e",
          6636 => x"5a",
          6637 => x"62",
          6638 => x"25",
          6639 => x"25",
          6640 => x"73",
          6641 => x"00",
          6642 => x"42",
          6643 => x"63",
          6644 => x"61",
          6645 => x"0a",
          6646 => x"52",
          6647 => x"69",
          6648 => x"2e",
          6649 => x"45",
          6650 => x"6c",
          6651 => x"20",
          6652 => x"65",
          6653 => x"70",
          6654 => x"2e",
          6655 => x"00",
          6656 => x"00",
          6657 => x"00",
          6658 => x"00",
          6659 => x"00",
          6660 => x"00",
          6661 => x"00",
          6662 => x"00",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"05",
          6667 => x"00",
          6668 => x"01",
          6669 => x"80",
          6670 => x"01",
          6671 => x"00",
          6672 => x"01",
          6673 => x"00",
          6674 => x"01",
          6675 => x"00",
          6676 => x"00",
          6677 => x"00",
          6678 => x"01",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"01",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"01",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"01",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"01",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"01",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"01",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"01",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"01",
          6711 => x"00",
          6712 => x"00",
          6713 => x"00",
          6714 => x"01",
          6715 => x"00",
          6716 => x"00",
          6717 => x"00",
          6718 => x"01",
          6719 => x"00",
          6720 => x"00",
          6721 => x"00",
          6722 => x"01",
          6723 => x"00",
          6724 => x"00",
          6725 => x"00",
          6726 => x"01",
          6727 => x"00",
          6728 => x"00",
          6729 => x"00",
          6730 => x"01",
          6731 => x"00",
          6732 => x"00",
          6733 => x"00",
          6734 => x"01",
          6735 => x"00",
          6736 => x"00",
          6737 => x"00",
          6738 => x"01",
          6739 => x"00",
          6740 => x"00",
          6741 => x"00",
          6742 => x"01",
          6743 => x"00",
          6744 => x"00",
          6745 => x"00",
          6746 => x"01",
          6747 => x"00",
          6748 => x"00",
          6749 => x"00",
          6750 => x"01",
          6751 => x"00",
          6752 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
