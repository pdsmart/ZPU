-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"ff",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"ae",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c3",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c5",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"d4",
           386 => x"b3",
           387 => x"d4",
           388 => x"90",
           389 => x"d4",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"84",
           396 => x"82",
           397 => x"af",
           398 => x"d8",
           399 => x"80",
           400 => x"d8",
           401 => x"ad",
           402 => x"d4",
           403 => x"90",
           404 => x"d4",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"84",
           419 => x"82",
           420 => x"96",
           421 => x"d8",
           422 => x"80",
           423 => x"d8",
           424 => x"cd",
           425 => x"d4",
           426 => x"90",
           427 => x"d4",
           428 => x"dd",
           429 => x"d4",
           430 => x"90",
           431 => x"d4",
           432 => x"bb",
           433 => x"d4",
           434 => x"90",
           435 => x"d4",
           436 => x"f8",
           437 => x"d4",
           438 => x"90",
           439 => x"d4",
           440 => x"ef",
           441 => x"d4",
           442 => x"90",
           443 => x"d4",
           444 => x"a2",
           445 => x"d4",
           446 => x"90",
           447 => x"d4",
           448 => x"c7",
           449 => x"d4",
           450 => x"90",
           451 => x"d4",
           452 => x"c6",
           453 => x"d4",
           454 => x"90",
           455 => x"d4",
           456 => x"ac",
           457 => x"d4",
           458 => x"90",
           459 => x"d4",
           460 => x"ac",
           461 => x"d4",
           462 => x"90",
           463 => x"d4",
           464 => x"84",
           465 => x"d4",
           466 => x"90",
           467 => x"d4",
           468 => x"ed",
           469 => x"d4",
           470 => x"90",
           471 => x"d4",
           472 => x"a3",
           473 => x"d4",
           474 => x"90",
           475 => x"d4",
           476 => x"a7",
           477 => x"d4",
           478 => x"90",
           479 => x"d4",
           480 => x"c7",
           481 => x"d4",
           482 => x"90",
           483 => x"d4",
           484 => x"e6",
           485 => x"d4",
           486 => x"90",
           487 => x"d4",
           488 => x"da",
           489 => x"d4",
           490 => x"90",
           491 => x"d4",
           492 => x"bc",
           493 => x"d4",
           494 => x"90",
           495 => x"d4",
           496 => x"b6",
           497 => x"d4",
           498 => x"90",
           499 => x"d4",
           500 => x"ec",
           501 => x"d4",
           502 => x"90",
           503 => x"d4",
           504 => x"bb",
           505 => x"d4",
           506 => x"90",
           507 => x"d4",
           508 => x"bc",
           509 => x"d4",
           510 => x"90",
           511 => x"d4",
           512 => x"a6",
           513 => x"d4",
           514 => x"90",
           515 => x"d4",
           516 => x"ff",
           517 => x"d4",
           518 => x"90",
           519 => x"d4",
           520 => x"aa",
           521 => x"d4",
           522 => x"90",
           523 => x"d4",
           524 => x"c3",
           525 => x"d4",
           526 => x"90",
           527 => x"d4",
           528 => x"ad",
           529 => x"d4",
           530 => x"90",
           531 => x"d4",
           532 => x"b8",
           533 => x"d4",
           534 => x"90",
           535 => x"d4",
           536 => x"bf",
           537 => x"d4",
           538 => x"90",
           539 => x"d4",
           540 => x"e6",
           541 => x"d4",
           542 => x"90",
           543 => x"d4",
           544 => x"ab",
           545 => x"d4",
           546 => x"90",
           547 => x"d4",
           548 => x"e0",
           549 => x"d4",
           550 => x"90",
           551 => x"d4",
           552 => x"cc",
           553 => x"d4",
           554 => x"90",
           555 => x"d4",
           556 => x"ee",
           557 => x"d4",
           558 => x"90",
           559 => x"d4",
           560 => x"d8",
           561 => x"d4",
           562 => x"90",
           563 => x"d4",
           564 => x"bc",
           565 => x"d4",
           566 => x"90",
           567 => x"d4",
           568 => x"a1",
           569 => x"d4",
           570 => x"90",
           571 => x"d4",
           572 => x"c5",
           573 => x"d4",
           574 => x"90",
           575 => x"d4",
           576 => x"a8",
           577 => x"d4",
           578 => x"90",
           579 => x"d4",
           580 => x"98",
           581 => x"d4",
           582 => x"90",
           583 => x"d4",
           584 => x"82",
           585 => x"d4",
           586 => x"90",
           587 => x"d4",
           588 => x"aa",
           589 => x"d4",
           590 => x"90",
           591 => x"d4",
           592 => x"a2",
           593 => x"d4",
           594 => x"90",
           595 => x"d4",
           596 => x"ec",
           597 => x"d4",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"c8",
           623 => x"b4",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"d4",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"d8",
           637 => x"05",
           638 => x"d8",
           639 => x"05",
           640 => x"f4",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"d4",
           652 => x"d8",
           653 => x"3d",
           654 => x"d4",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"d8",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"d8",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"d8",
           675 => x"05",
           676 => x"d4",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"d8",
           683 => x"05",
           684 => x"90",
           685 => x"c8",
           686 => x"d8",
           687 => x"05",
           688 => x"d8",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"d8",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"d8",
           709 => x"05",
           710 => x"72",
           711 => x"d4",
           712 => x"08",
           713 => x"d4",
           714 => x"0c",
           715 => x"d4",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"d4",
           722 => x"0d",
           723 => x"d8",
           724 => x"05",
           725 => x"d4",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"d8",
           730 => x"05",
           731 => x"d4",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"d4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"d4",
           756 => x"d8",
           757 => x"3d",
           758 => x"d4",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"d8",
           769 => x"82",
           770 => x"f8",
           771 => x"d8",
           772 => x"05",
           773 => x"d8",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"d4",
           779 => x"0d",
           780 => x"d8",
           781 => x"05",
           782 => x"d4",
           783 => x"08",
           784 => x"8c",
           785 => x"d8",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"d4",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"d4",
           804 => x"08",
           805 => x"d8",
           806 => x"05",
           807 => x"d4",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"d4",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"d8",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"d4",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"d8",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"d8",
           863 => x"05",
           864 => x"d4",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"d4",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"d8",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"d4",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"d8",
           889 => x"05",
           890 => x"d4",
           891 => x"33",
           892 => x"d8",
           893 => x"05",
           894 => x"d8",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"d4",
           901 => x"51",
           902 => x"72",
           903 => x"d4",
           904 => x"22",
           905 => x"51",
           906 => x"d8",
           907 => x"05",
           908 => x"d4",
           909 => x"22",
           910 => x"51",
           911 => x"d8",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"d8",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"d8",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"d4",
           930 => x"23",
           931 => x"d8",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"d4",
           938 => x"23",
           939 => x"bf",
           940 => x"d4",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"d8",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"d4",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"d4",
           969 => x"0c",
           970 => x"d8",
           971 => x"05",
           972 => x"d4",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"d8",
           982 => x"05",
           983 => x"a2",
           984 => x"d8",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"d4",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"d8",
           993 => x"05",
           994 => x"d4",
           995 => x"22",
           996 => x"d4",
           997 => x"22",
           998 => x"54",
           999 => x"d8",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"d4",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"d8",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"d4",
          1020 => x"08",
          1021 => x"c1",
          1022 => x"c8",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"d4",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"d4",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"d4",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"d8",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"d8",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"d4",
          1069 => x"22",
          1070 => x"51",
          1071 => x"d8",
          1072 => x"05",
          1073 => x"d4",
          1074 => x"08",
          1075 => x"d4",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"d8",
          1081 => x"05",
          1082 => x"39",
          1083 => x"d8",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"d4",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"d4",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"d8",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"d8",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"d8",
          1127 => x"d8",
          1128 => x"05",
          1129 => x"d4",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"d8",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"d8",
          1147 => x"05",
          1148 => x"33",
          1149 => x"d4",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"d4",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"d4",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"d4",
          1172 => x"08",
          1173 => x"ab",
          1174 => x"c8",
          1175 => x"d8",
          1176 => x"05",
          1177 => x"d8",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"d4",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"d4",
          1193 => x"22",
          1194 => x"53",
          1195 => x"d4",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"d8",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"d8",
          1225 => x"05",
          1226 => x"d4",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"d8",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"d4",
          1247 => x"33",
          1248 => x"d4",
          1249 => x"33",
          1250 => x"54",
          1251 => x"d8",
          1252 => x"05",
          1253 => x"d4",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"d8",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"d4",
          1269 => x"23",
          1270 => x"d8",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"d4",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"d4",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"d4",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"d8",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"d8",
          1381 => x"05",
          1382 => x"54",
          1383 => x"d8",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"d8",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"d4",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"d8",
          1397 => x"05",
          1398 => x"d8",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"d8",
          1407 => x"05",
          1408 => x"51",
          1409 => x"d8",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"d4",
          1420 => x"08",
          1421 => x"d8",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"d8",
          1430 => x"05",
          1431 => x"51",
          1432 => x"d8",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"d4",
          1444 => x"08",
          1445 => x"d8",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"d4",
          1452 => x"08",
          1453 => x"d4",
          1454 => x"08",
          1455 => x"d8",
          1456 => x"05",
          1457 => x"d4",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"d4",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"d8",
          1479 => x"05",
          1480 => x"d8",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"d4",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"d4",
          1496 => x"34",
          1497 => x"d8",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"d8",
          1506 => x"05",
          1507 => x"08",
          1508 => x"d4",
          1509 => x"0c",
          1510 => x"d8",
          1511 => x"05",
          1512 => x"c8",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"d4",
          1516 => x"d8",
          1517 => x"3d",
          1518 => x"a8",
          1519 => x"d8",
          1520 => x"05",
          1521 => x"d8",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"c8",
          1525 => x"d8",
          1526 => x"85",
          1527 => x"d8",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"d4",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"d8",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"d4",
          1549 => x"0c",
          1550 => x"d8",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"f4",
          1567 => x"f4",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"d8",
          1582 => x"3d",
          1583 => x"d4",
          1584 => x"d8",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"d8",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"d8",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"d4",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"d8",
          1625 => x"05",
          1626 => x"d8",
          1627 => x"05",
          1628 => x"d8",
          1629 => x"05",
          1630 => x"c8",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"d4",
          1634 => x"d8",
          1635 => x"3d",
          1636 => x"ac",
          1637 => x"d8",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"c8",
          1642 => x"3d",
          1643 => x"d4",
          1644 => x"d8",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"d8",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"d4",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"d4",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"d8",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"d8",
          1689 => x"05",
          1690 => x"d8",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"d8",
          1696 => x"72",
          1697 => x"d8",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"d4",
          1702 => x"08",
          1703 => x"d4",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"d8",
          1707 => x"05",
          1708 => x"d4",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"d4",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"d4",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"d8",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"d8",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"d4",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"d4",
          1761 => x"08",
          1762 => x"d8",
          1763 => x"05",
          1764 => x"d4",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"d8",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"d8",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"c8",
          1783 => x"d8",
          1784 => x"05",
          1785 => x"d8",
          1786 => x"05",
          1787 => x"80",
          1788 => x"d8",
          1789 => x"05",
          1790 => x"d4",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"d8",
          1795 => x"05",
          1796 => x"d8",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"d8",
          1810 => x"05",
          1811 => x"d8",
          1812 => x"05",
          1813 => x"34",
          1814 => x"d8",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"d8",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"d8",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"d8",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"d8",
          1836 => x"05",
          1837 => x"d4",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"d8",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"d4",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"d4",
          1853 => x"08",
          1854 => x"90",
          1855 => x"d4",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"d8",
          1863 => x"05",
          1864 => x"d8",
          1865 => x"05",
          1866 => x"d4",
          1867 => x"08",
          1868 => x"d8",
          1869 => x"05",
          1870 => x"d4",
          1871 => x"08",
          1872 => x"d8",
          1873 => x"05",
          1874 => x"d4",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"d4",
          1878 => x"08",
          1879 => x"d8",
          1880 => x"05",
          1881 => x"d4",
          1882 => x"08",
          1883 => x"d8",
          1884 => x"05",
          1885 => x"d4",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"d4",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"d4",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"d4",
          1905 => x"08",
          1906 => x"d8",
          1907 => x"05",
          1908 => x"d4",
          1909 => x"08",
          1910 => x"71",
          1911 => x"d4",
          1912 => x"08",
          1913 => x"d8",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"d4",
          1922 => x"d8",
          1923 => x"3d",
          1924 => x"d4",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"d4",
          1931 => x"08",
          1932 => x"d8",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"d8",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"d8",
          1942 => x"05",
          1943 => x"d4",
          1944 => x"08",
          1945 => x"d8",
          1946 => x"84",
          1947 => x"d8",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"d8",
          1954 => x"05",
          1955 => x"d4",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"d4",
          1978 => x"d8",
          1979 => x"3d",
          1980 => x"d4",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"d8",
          1986 => x"05",
          1987 => x"d4",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"d4",
          1991 => x"08",
          1992 => x"d8",
          1993 => x"05",
          1994 => x"d4",
          1995 => x"08",
          1996 => x"d8",
          1997 => x"05",
          1998 => x"d4",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"d8",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"d8",
          2008 => x"05",
          2009 => x"71",
          2010 => x"d8",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"d4",
          2016 => x"08",
          2017 => x"c8",
          2018 => x"3d",
          2019 => x"d4",
          2020 => x"d8",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"d8",
          2024 => x"05",
          2025 => x"81",
          2026 => x"d8",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"d4",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"d4",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"d8",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"d4",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"d8",
          2059 => x"05",
          2060 => x"80",
          2061 => x"d8",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"d8",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"d4",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"d4",
          2079 => x"08",
          2080 => x"d8",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"d8",
          2090 => x"05",
          2091 => x"c8",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"d4",
          2095 => x"d8",
          2096 => x"3d",
          2097 => x"d4",
          2098 => x"08",
          2099 => x"08",
          2100 => x"82",
          2101 => x"8c",
          2102 => x"38",
          2103 => x"d8",
          2104 => x"05",
          2105 => x"39",
          2106 => x"08",
          2107 => x"52",
          2108 => x"d8",
          2109 => x"05",
          2110 => x"82",
          2111 => x"f8",
          2112 => x"81",
          2113 => x"51",
          2114 => x"9f",
          2115 => x"d4",
          2116 => x"08",
          2117 => x"d8",
          2118 => x"05",
          2119 => x"d4",
          2120 => x"08",
          2121 => x"38",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"05",
          2125 => x"08",
          2126 => x"82",
          2127 => x"f8",
          2128 => x"d8",
          2129 => x"05",
          2130 => x"82",
          2131 => x"fc",
          2132 => x"82",
          2133 => x"fc",
          2134 => x"d8",
          2135 => x"3d",
          2136 => x"d4",
          2137 => x"d8",
          2138 => x"82",
          2139 => x"fe",
          2140 => x"d8",
          2141 => x"05",
          2142 => x"d4",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"80",
          2146 => x"38",
          2147 => x"08",
          2148 => x"81",
          2149 => x"d4",
          2150 => x"0c",
          2151 => x"08",
          2152 => x"ff",
          2153 => x"d4",
          2154 => x"0c",
          2155 => x"08",
          2156 => x"80",
          2157 => x"82",
          2158 => x"8c",
          2159 => x"70",
          2160 => x"08",
          2161 => x"52",
          2162 => x"34",
          2163 => x"08",
          2164 => x"81",
          2165 => x"d4",
          2166 => x"0c",
          2167 => x"82",
          2168 => x"88",
          2169 => x"82",
          2170 => x"51",
          2171 => x"82",
          2172 => x"04",
          2173 => x"08",
          2174 => x"d4",
          2175 => x"0d",
          2176 => x"d8",
          2177 => x"05",
          2178 => x"d4",
          2179 => x"08",
          2180 => x"38",
          2181 => x"08",
          2182 => x"30",
          2183 => x"08",
          2184 => x"80",
          2185 => x"d4",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"8a",
          2189 => x"82",
          2190 => x"f4",
          2191 => x"d8",
          2192 => x"05",
          2193 => x"d4",
          2194 => x"0c",
          2195 => x"08",
          2196 => x"80",
          2197 => x"82",
          2198 => x"8c",
          2199 => x"82",
          2200 => x"8c",
          2201 => x"0b",
          2202 => x"08",
          2203 => x"82",
          2204 => x"fc",
          2205 => x"38",
          2206 => x"d8",
          2207 => x"05",
          2208 => x"d4",
          2209 => x"08",
          2210 => x"08",
          2211 => x"80",
          2212 => x"d4",
          2213 => x"08",
          2214 => x"d4",
          2215 => x"08",
          2216 => x"3f",
          2217 => x"08",
          2218 => x"d4",
          2219 => x"0c",
          2220 => x"d4",
          2221 => x"08",
          2222 => x"38",
          2223 => x"08",
          2224 => x"30",
          2225 => x"08",
          2226 => x"82",
          2227 => x"f8",
          2228 => x"82",
          2229 => x"54",
          2230 => x"82",
          2231 => x"04",
          2232 => x"08",
          2233 => x"d4",
          2234 => x"0d",
          2235 => x"d8",
          2236 => x"05",
          2237 => x"d4",
          2238 => x"08",
          2239 => x"38",
          2240 => x"08",
          2241 => x"30",
          2242 => x"08",
          2243 => x"81",
          2244 => x"d4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"80",
          2248 => x"82",
          2249 => x"8c",
          2250 => x"82",
          2251 => x"8c",
          2252 => x"53",
          2253 => x"08",
          2254 => x"52",
          2255 => x"08",
          2256 => x"51",
          2257 => x"82",
          2258 => x"70",
          2259 => x"08",
          2260 => x"54",
          2261 => x"08",
          2262 => x"80",
          2263 => x"82",
          2264 => x"f8",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"d8",
          2268 => x"05",
          2269 => x"d8",
          2270 => x"87",
          2271 => x"d8",
          2272 => x"82",
          2273 => x"02",
          2274 => x"0c",
          2275 => x"80",
          2276 => x"d4",
          2277 => x"08",
          2278 => x"d4",
          2279 => x"08",
          2280 => x"3f",
          2281 => x"08",
          2282 => x"c8",
          2283 => x"3d",
          2284 => x"d4",
          2285 => x"d8",
          2286 => x"82",
          2287 => x"fd",
          2288 => x"53",
          2289 => x"08",
          2290 => x"52",
          2291 => x"08",
          2292 => x"51",
          2293 => x"d8",
          2294 => x"82",
          2295 => x"54",
          2296 => x"82",
          2297 => x"04",
          2298 => x"08",
          2299 => x"d4",
          2300 => x"0d",
          2301 => x"d8",
          2302 => x"05",
          2303 => x"82",
          2304 => x"f8",
          2305 => x"d8",
          2306 => x"05",
          2307 => x"d4",
          2308 => x"08",
          2309 => x"82",
          2310 => x"fc",
          2311 => x"2e",
          2312 => x"0b",
          2313 => x"08",
          2314 => x"24",
          2315 => x"d8",
          2316 => x"05",
          2317 => x"d8",
          2318 => x"05",
          2319 => x"d4",
          2320 => x"08",
          2321 => x"d4",
          2322 => x"0c",
          2323 => x"82",
          2324 => x"fc",
          2325 => x"2e",
          2326 => x"82",
          2327 => x"8c",
          2328 => x"d8",
          2329 => x"05",
          2330 => x"38",
          2331 => x"08",
          2332 => x"82",
          2333 => x"8c",
          2334 => x"82",
          2335 => x"88",
          2336 => x"d8",
          2337 => x"05",
          2338 => x"d4",
          2339 => x"08",
          2340 => x"d4",
          2341 => x"0c",
          2342 => x"08",
          2343 => x"81",
          2344 => x"d4",
          2345 => x"0c",
          2346 => x"08",
          2347 => x"81",
          2348 => x"d4",
          2349 => x"0c",
          2350 => x"82",
          2351 => x"90",
          2352 => x"2e",
          2353 => x"d8",
          2354 => x"05",
          2355 => x"d8",
          2356 => x"05",
          2357 => x"39",
          2358 => x"08",
          2359 => x"70",
          2360 => x"08",
          2361 => x"51",
          2362 => x"08",
          2363 => x"82",
          2364 => x"85",
          2365 => x"d8",
          2366 => x"82",
          2367 => x"02",
          2368 => x"0c",
          2369 => x"80",
          2370 => x"d4",
          2371 => x"34",
          2372 => x"08",
          2373 => x"53",
          2374 => x"82",
          2375 => x"88",
          2376 => x"08",
          2377 => x"33",
          2378 => x"d8",
          2379 => x"05",
          2380 => x"ff",
          2381 => x"a0",
          2382 => x"06",
          2383 => x"d8",
          2384 => x"05",
          2385 => x"81",
          2386 => x"53",
          2387 => x"d8",
          2388 => x"05",
          2389 => x"ad",
          2390 => x"06",
          2391 => x"0b",
          2392 => x"08",
          2393 => x"82",
          2394 => x"88",
          2395 => x"08",
          2396 => x"0c",
          2397 => x"53",
          2398 => x"d8",
          2399 => x"05",
          2400 => x"d4",
          2401 => x"33",
          2402 => x"2e",
          2403 => x"81",
          2404 => x"d8",
          2405 => x"05",
          2406 => x"81",
          2407 => x"70",
          2408 => x"72",
          2409 => x"d4",
          2410 => x"34",
          2411 => x"08",
          2412 => x"82",
          2413 => x"e8",
          2414 => x"d8",
          2415 => x"05",
          2416 => x"2e",
          2417 => x"d8",
          2418 => x"05",
          2419 => x"2e",
          2420 => x"cd",
          2421 => x"82",
          2422 => x"f4",
          2423 => x"d8",
          2424 => x"05",
          2425 => x"81",
          2426 => x"70",
          2427 => x"72",
          2428 => x"d4",
          2429 => x"34",
          2430 => x"82",
          2431 => x"d4",
          2432 => x"34",
          2433 => x"08",
          2434 => x"70",
          2435 => x"71",
          2436 => x"51",
          2437 => x"82",
          2438 => x"f8",
          2439 => x"fe",
          2440 => x"d4",
          2441 => x"33",
          2442 => x"26",
          2443 => x"0b",
          2444 => x"08",
          2445 => x"83",
          2446 => x"d8",
          2447 => x"05",
          2448 => x"73",
          2449 => x"82",
          2450 => x"f8",
          2451 => x"72",
          2452 => x"38",
          2453 => x"0b",
          2454 => x"08",
          2455 => x"82",
          2456 => x"0b",
          2457 => x"08",
          2458 => x"b2",
          2459 => x"d4",
          2460 => x"33",
          2461 => x"27",
          2462 => x"d8",
          2463 => x"05",
          2464 => x"b9",
          2465 => x"8d",
          2466 => x"82",
          2467 => x"ec",
          2468 => x"a5",
          2469 => x"82",
          2470 => x"f4",
          2471 => x"0b",
          2472 => x"08",
          2473 => x"82",
          2474 => x"f8",
          2475 => x"a0",
          2476 => x"cf",
          2477 => x"d4",
          2478 => x"33",
          2479 => x"73",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"11",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"d8",
          2486 => x"05",
          2487 => x"51",
          2488 => x"d8",
          2489 => x"05",
          2490 => x"d4",
          2491 => x"33",
          2492 => x"27",
          2493 => x"d8",
          2494 => x"05",
          2495 => x"51",
          2496 => x"d8",
          2497 => x"05",
          2498 => x"d4",
          2499 => x"33",
          2500 => x"26",
          2501 => x"0b",
          2502 => x"08",
          2503 => x"81",
          2504 => x"d8",
          2505 => x"05",
          2506 => x"d4",
          2507 => x"33",
          2508 => x"74",
          2509 => x"80",
          2510 => x"d4",
          2511 => x"0c",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"12",
          2519 => x"08",
          2520 => x"82",
          2521 => x"88",
          2522 => x"08",
          2523 => x"0c",
          2524 => x"51",
          2525 => x"72",
          2526 => x"d4",
          2527 => x"34",
          2528 => x"82",
          2529 => x"f0",
          2530 => x"72",
          2531 => x"38",
          2532 => x"08",
          2533 => x"30",
          2534 => x"08",
          2535 => x"82",
          2536 => x"8c",
          2537 => x"d8",
          2538 => x"05",
          2539 => x"53",
          2540 => x"d8",
          2541 => x"05",
          2542 => x"d4",
          2543 => x"08",
          2544 => x"0c",
          2545 => x"82",
          2546 => x"04",
          2547 => x"08",
          2548 => x"d4",
          2549 => x"0d",
          2550 => x"d8",
          2551 => x"05",
          2552 => x"d4",
          2553 => x"08",
          2554 => x"0c",
          2555 => x"08",
          2556 => x"70",
          2557 => x"72",
          2558 => x"82",
          2559 => x"f8",
          2560 => x"81",
          2561 => x"72",
          2562 => x"81",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"82",
          2568 => x"f8",
          2569 => x"72",
          2570 => x"81",
          2571 => x"81",
          2572 => x"d4",
          2573 => x"34",
          2574 => x"08",
          2575 => x"70",
          2576 => x"71",
          2577 => x"51",
          2578 => x"82",
          2579 => x"f8",
          2580 => x"d8",
          2581 => x"05",
          2582 => x"b0",
          2583 => x"06",
          2584 => x"82",
          2585 => x"88",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"53",
          2589 => x"d8",
          2590 => x"05",
          2591 => x"d4",
          2592 => x"33",
          2593 => x"08",
          2594 => x"82",
          2595 => x"e8",
          2596 => x"e2",
          2597 => x"82",
          2598 => x"e8",
          2599 => x"f8",
          2600 => x"80",
          2601 => x"0b",
          2602 => x"08",
          2603 => x"82",
          2604 => x"88",
          2605 => x"08",
          2606 => x"0c",
          2607 => x"53",
          2608 => x"d8",
          2609 => x"05",
          2610 => x"39",
          2611 => x"d8",
          2612 => x"05",
          2613 => x"d4",
          2614 => x"08",
          2615 => x"05",
          2616 => x"08",
          2617 => x"33",
          2618 => x"08",
          2619 => x"80",
          2620 => x"d8",
          2621 => x"05",
          2622 => x"a0",
          2623 => x"81",
          2624 => x"d4",
          2625 => x"0c",
          2626 => x"82",
          2627 => x"f8",
          2628 => x"af",
          2629 => x"38",
          2630 => x"08",
          2631 => x"53",
          2632 => x"83",
          2633 => x"80",
          2634 => x"d4",
          2635 => x"0c",
          2636 => x"88",
          2637 => x"d4",
          2638 => x"34",
          2639 => x"d8",
          2640 => x"05",
          2641 => x"73",
          2642 => x"82",
          2643 => x"f8",
          2644 => x"72",
          2645 => x"38",
          2646 => x"0b",
          2647 => x"08",
          2648 => x"82",
          2649 => x"0b",
          2650 => x"08",
          2651 => x"80",
          2652 => x"d4",
          2653 => x"0c",
          2654 => x"08",
          2655 => x"53",
          2656 => x"81",
          2657 => x"d8",
          2658 => x"05",
          2659 => x"e0",
          2660 => x"38",
          2661 => x"08",
          2662 => x"e0",
          2663 => x"72",
          2664 => x"08",
          2665 => x"82",
          2666 => x"f8",
          2667 => x"11",
          2668 => x"82",
          2669 => x"f8",
          2670 => x"d8",
          2671 => x"05",
          2672 => x"73",
          2673 => x"82",
          2674 => x"f8",
          2675 => x"11",
          2676 => x"82",
          2677 => x"f8",
          2678 => x"d8",
          2679 => x"05",
          2680 => x"89",
          2681 => x"80",
          2682 => x"d4",
          2683 => x"0c",
          2684 => x"82",
          2685 => x"f8",
          2686 => x"d8",
          2687 => x"05",
          2688 => x"72",
          2689 => x"38",
          2690 => x"d8",
          2691 => x"05",
          2692 => x"39",
          2693 => x"08",
          2694 => x"70",
          2695 => x"08",
          2696 => x"29",
          2697 => x"08",
          2698 => x"70",
          2699 => x"d4",
          2700 => x"0c",
          2701 => x"08",
          2702 => x"70",
          2703 => x"71",
          2704 => x"51",
          2705 => x"53",
          2706 => x"d8",
          2707 => x"05",
          2708 => x"39",
          2709 => x"08",
          2710 => x"53",
          2711 => x"90",
          2712 => x"d4",
          2713 => x"08",
          2714 => x"d4",
          2715 => x"0c",
          2716 => x"08",
          2717 => x"82",
          2718 => x"fc",
          2719 => x"0c",
          2720 => x"82",
          2721 => x"ec",
          2722 => x"d8",
          2723 => x"05",
          2724 => x"c8",
          2725 => x"0d",
          2726 => x"0c",
          2727 => x"0d",
          2728 => x"70",
          2729 => x"74",
          2730 => x"e3",
          2731 => x"75",
          2732 => x"d1",
          2733 => x"c8",
          2734 => x"0c",
          2735 => x"54",
          2736 => x"74",
          2737 => x"a0",
          2738 => x"06",
          2739 => x"15",
          2740 => x"80",
          2741 => x"29",
          2742 => x"05",
          2743 => x"56",
          2744 => x"82",
          2745 => x"53",
          2746 => x"08",
          2747 => x"3f",
          2748 => x"08",
          2749 => x"16",
          2750 => x"81",
          2751 => x"38",
          2752 => x"81",
          2753 => x"54",
          2754 => x"c9",
          2755 => x"73",
          2756 => x"0c",
          2757 => x"04",
          2758 => x"73",
          2759 => x"26",
          2760 => x"71",
          2761 => x"ae",
          2762 => x"71",
          2763 => x"b4",
          2764 => x"80",
          2765 => x"f0",
          2766 => x"39",
          2767 => x"51",
          2768 => x"82",
          2769 => x"80",
          2770 => x"b5",
          2771 => x"e4",
          2772 => x"b0",
          2773 => x"39",
          2774 => x"51",
          2775 => x"82",
          2776 => x"80",
          2777 => x"b5",
          2778 => x"c8",
          2779 => x"84",
          2780 => x"39",
          2781 => x"51",
          2782 => x"b6",
          2783 => x"39",
          2784 => x"51",
          2785 => x"b6",
          2786 => x"39",
          2787 => x"51",
          2788 => x"b7",
          2789 => x"39",
          2790 => x"51",
          2791 => x"b7",
          2792 => x"39",
          2793 => x"51",
          2794 => x"b7",
          2795 => x"39",
          2796 => x"51",
          2797 => x"83",
          2798 => x"fb",
          2799 => x"79",
          2800 => x"87",
          2801 => x"38",
          2802 => x"87",
          2803 => x"90",
          2804 => x"52",
          2805 => x"ab",
          2806 => x"c8",
          2807 => x"51",
          2808 => x"82",
          2809 => x"54",
          2810 => x"52",
          2811 => x"51",
          2812 => x"3f",
          2813 => x"04",
          2814 => x"66",
          2815 => x"80",
          2816 => x"5b",
          2817 => x"78",
          2818 => x"07",
          2819 => x"57",
          2820 => x"56",
          2821 => x"26",
          2822 => x"56",
          2823 => x"70",
          2824 => x"51",
          2825 => x"74",
          2826 => x"81",
          2827 => x"8c",
          2828 => x"56",
          2829 => x"3f",
          2830 => x"08",
          2831 => x"c8",
          2832 => x"82",
          2833 => x"87",
          2834 => x"0c",
          2835 => x"08",
          2836 => x"d4",
          2837 => x"80",
          2838 => x"75",
          2839 => x"cc",
          2840 => x"c8",
          2841 => x"d8",
          2842 => x"38",
          2843 => x"80",
          2844 => x"74",
          2845 => x"59",
          2846 => x"96",
          2847 => x"51",
          2848 => x"3f",
          2849 => x"78",
          2850 => x"7b",
          2851 => x"2a",
          2852 => x"57",
          2853 => x"80",
          2854 => x"82",
          2855 => x"87",
          2856 => x"08",
          2857 => x"fe",
          2858 => x"56",
          2859 => x"c8",
          2860 => x"0d",
          2861 => x"0d",
          2862 => x"05",
          2863 => x"59",
          2864 => x"80",
          2865 => x"7b",
          2866 => x"3f",
          2867 => x"08",
          2868 => x"77",
          2869 => x"38",
          2870 => x"bf",
          2871 => x"82",
          2872 => x"82",
          2873 => x"82",
          2874 => x"82",
          2875 => x"54",
          2876 => x"08",
          2877 => x"a8",
          2878 => x"b8",
          2879 => x"b9",
          2880 => x"f4",
          2881 => x"55",
          2882 => x"d8",
          2883 => x"52",
          2884 => x"2d",
          2885 => x"08",
          2886 => x"79",
          2887 => x"d8",
          2888 => x"3d",
          2889 => x"3d",
          2890 => x"63",
          2891 => x"80",
          2892 => x"73",
          2893 => x"41",
          2894 => x"5e",
          2895 => x"52",
          2896 => x"51",
          2897 => x"3f",
          2898 => x"51",
          2899 => x"3f",
          2900 => x"79",
          2901 => x"38",
          2902 => x"89",
          2903 => x"2e",
          2904 => x"c6",
          2905 => x"53",
          2906 => x"8e",
          2907 => x"52",
          2908 => x"51",
          2909 => x"3f",
          2910 => x"b9",
          2911 => x"b8",
          2912 => x"15",
          2913 => x"39",
          2914 => x"72",
          2915 => x"38",
          2916 => x"82",
          2917 => x"ff",
          2918 => x"89",
          2919 => x"8c",
          2920 => x"b4",
          2921 => x"55",
          2922 => x"18",
          2923 => x"27",
          2924 => x"33",
          2925 => x"98",
          2926 => x"9c",
          2927 => x"82",
          2928 => x"ff",
          2929 => x"81",
          2930 => x"f4",
          2931 => x"a0",
          2932 => x"3f",
          2933 => x"82",
          2934 => x"ff",
          2935 => x"80",
          2936 => x"27",
          2937 => x"74",
          2938 => x"55",
          2939 => x"72",
          2940 => x"38",
          2941 => x"53",
          2942 => x"83",
          2943 => x"75",
          2944 => x"81",
          2945 => x"53",
          2946 => x"90",
          2947 => x"fe",
          2948 => x"82",
          2949 => x"52",
          2950 => x"39",
          2951 => x"08",
          2952 => x"d7",
          2953 => x"15",
          2954 => x"39",
          2955 => x"51",
          2956 => x"78",
          2957 => x"5c",
          2958 => x"3f",
          2959 => x"08",
          2960 => x"98",
          2961 => x"76",
          2962 => x"81",
          2963 => x"a0",
          2964 => x"d8",
          2965 => x"2b",
          2966 => x"70",
          2967 => x"30",
          2968 => x"70",
          2969 => x"07",
          2970 => x"06",
          2971 => x"59",
          2972 => x"80",
          2973 => x"38",
          2974 => x"09",
          2975 => x"38",
          2976 => x"39",
          2977 => x"72",
          2978 => x"b2",
          2979 => x"72",
          2980 => x"0c",
          2981 => x"04",
          2982 => x"02",
          2983 => x"82",
          2984 => x"82",
          2985 => x"55",
          2986 => x"3f",
          2987 => x"22",
          2988 => x"3f",
          2989 => x"54",
          2990 => x"53",
          2991 => x"33",
          2992 => x"d4",
          2993 => x"90",
          2994 => x"2e",
          2995 => x"8d",
          2996 => x"0d",
          2997 => x"0d",
          2998 => x"80",
          2999 => x"b6",
          3000 => x"9c",
          3001 => x"b9",
          3002 => x"d8",
          3003 => x"9c",
          3004 => x"81",
          3005 => x"06",
          3006 => x"80",
          3007 => x"81",
          3008 => x"3f",
          3009 => x"51",
          3010 => x"80",
          3011 => x"3f",
          3012 => x"70",
          3013 => x"52",
          3014 => x"92",
          3015 => x"9c",
          3016 => x"ba",
          3017 => x"9c",
          3018 => x"9b",
          3019 => x"83",
          3020 => x"06",
          3021 => x"80",
          3022 => x"81",
          3023 => x"3f",
          3024 => x"51",
          3025 => x"80",
          3026 => x"3f",
          3027 => x"70",
          3028 => x"52",
          3029 => x"92",
          3030 => x"9b",
          3031 => x"ba",
          3032 => x"e0",
          3033 => x"9b",
          3034 => x"85",
          3035 => x"06",
          3036 => x"80",
          3037 => x"81",
          3038 => x"3f",
          3039 => x"51",
          3040 => x"80",
          3041 => x"3f",
          3042 => x"70",
          3043 => x"52",
          3044 => x"92",
          3045 => x"9b",
          3046 => x"ba",
          3047 => x"a4",
          3048 => x"9b",
          3049 => x"87",
          3050 => x"06",
          3051 => x"80",
          3052 => x"81",
          3053 => x"3f",
          3054 => x"51",
          3055 => x"80",
          3056 => x"3f",
          3057 => x"70",
          3058 => x"52",
          3059 => x"92",
          3060 => x"9a",
          3061 => x"bb",
          3062 => x"e8",
          3063 => x"9a",
          3064 => x"ba",
          3065 => x"0d",
          3066 => x"0d",
          3067 => x"05",
          3068 => x"70",
          3069 => x"80",
          3070 => x"e2",
          3071 => x"0b",
          3072 => x"33",
          3073 => x"38",
          3074 => x"bb",
          3075 => x"ef",
          3076 => x"8e",
          3077 => x"d8",
          3078 => x"70",
          3079 => x"08",
          3080 => x"82",
          3081 => x"51",
          3082 => x"0b",
          3083 => x"34",
          3084 => x"d3",
          3085 => x"73",
          3086 => x"81",
          3087 => x"82",
          3088 => x"74",
          3089 => x"81",
          3090 => x"82",
          3091 => x"80",
          3092 => x"82",
          3093 => x"51",
          3094 => x"91",
          3095 => x"d8",
          3096 => x"e2",
          3097 => x"0b",
          3098 => x"c4",
          3099 => x"82",
          3100 => x"54",
          3101 => x"09",
          3102 => x"38",
          3103 => x"53",
          3104 => x"51",
          3105 => x"80",
          3106 => x"c8",
          3107 => x"0d",
          3108 => x"0d",
          3109 => x"82",
          3110 => x"5f",
          3111 => x"7c",
          3112 => x"cb",
          3113 => x"c8",
          3114 => x"06",
          3115 => x"2e",
          3116 => x"a3",
          3117 => x"59",
          3118 => x"bb",
          3119 => x"51",
          3120 => x"7c",
          3121 => x"82",
          3122 => x"81",
          3123 => x"82",
          3124 => x"7d",
          3125 => x"82",
          3126 => x"91",
          3127 => x"70",
          3128 => x"bc",
          3129 => x"b1",
          3130 => x"3d",
          3131 => x"80",
          3132 => x"51",
          3133 => x"b4",
          3134 => x"05",
          3135 => x"3f",
          3136 => x"08",
          3137 => x"90",
          3138 => x"78",
          3139 => x"89",
          3140 => x"80",
          3141 => x"d9",
          3142 => x"2e",
          3143 => x"78",
          3144 => x"38",
          3145 => x"81",
          3146 => x"82",
          3147 => x"78",
          3148 => x"ae",
          3149 => x"39",
          3150 => x"82",
          3151 => x"94",
          3152 => x"38",
          3153 => x"78",
          3154 => x"fc",
          3155 => x"24",
          3156 => x"b0",
          3157 => x"38",
          3158 => x"84",
          3159 => x"d9",
          3160 => x"2e",
          3161 => x"78",
          3162 => x"86",
          3163 => x"c9",
          3164 => x"d5",
          3165 => x"38",
          3166 => x"24",
          3167 => x"80",
          3168 => x"d9",
          3169 => x"d0",
          3170 => x"78",
          3171 => x"89",
          3172 => x"80",
          3173 => x"a5",
          3174 => x"39",
          3175 => x"2e",
          3176 => x"78",
          3177 => x"8c",
          3178 => x"8d",
          3179 => x"82",
          3180 => x"38",
          3181 => x"24",
          3182 => x"80",
          3183 => x"f6",
          3184 => x"f9",
          3185 => x"38",
          3186 => x"78",
          3187 => x"8d",
          3188 => x"81",
          3189 => x"db",
          3190 => x"39",
          3191 => x"80",
          3192 => x"84",
          3193 => x"e4",
          3194 => x"c8",
          3195 => x"82",
          3196 => x"8f",
          3197 => x"3d",
          3198 => x"53",
          3199 => x"51",
          3200 => x"82",
          3201 => x"80",
          3202 => x"81",
          3203 => x"38",
          3204 => x"80",
          3205 => x"52",
          3206 => x"05",
          3207 => x"c8",
          3208 => x"d8",
          3209 => x"ff",
          3210 => x"8d",
          3211 => x"b4",
          3212 => x"3f",
          3213 => x"aa",
          3214 => x"c4",
          3215 => x"39",
          3216 => x"80",
          3217 => x"84",
          3218 => x"80",
          3219 => x"c8",
          3220 => x"fd",
          3221 => x"53",
          3222 => x"80",
          3223 => x"51",
          3224 => x"3f",
          3225 => x"08",
          3226 => x"dc",
          3227 => x"39",
          3228 => x"80",
          3229 => x"84",
          3230 => x"d0",
          3231 => x"c8",
          3232 => x"87",
          3233 => x"26",
          3234 => x"b4",
          3235 => x"11",
          3236 => x"05",
          3237 => x"3f",
          3238 => x"08",
          3239 => x"d8",
          3240 => x"63",
          3241 => x"e4",
          3242 => x"ff",
          3243 => x"02",
          3244 => x"33",
          3245 => x"63",
          3246 => x"82",
          3247 => x"51",
          3248 => x"3f",
          3249 => x"08",
          3250 => x"82",
          3251 => x"ca",
          3252 => x"5d",
          3253 => x"b4",
          3254 => x"05",
          3255 => x"3f",
          3256 => x"08",
          3257 => x"84",
          3258 => x"90",
          3259 => x"53",
          3260 => x"08",
          3261 => x"f1",
          3262 => x"d1",
          3263 => x"ff",
          3264 => x"8f",
          3265 => x"d8",
          3266 => x"3d",
          3267 => x"52",
          3268 => x"3f",
          3269 => x"08",
          3270 => x"84",
          3271 => x"90",
          3272 => x"d8",
          3273 => x"3d",
          3274 => x"52",
          3275 => x"3f",
          3276 => x"58",
          3277 => x"57",
          3278 => x"55",
          3279 => x"08",
          3280 => x"54",
          3281 => x"52",
          3282 => x"e9",
          3283 => x"c8",
          3284 => x"fb",
          3285 => x"d8",
          3286 => x"ef",
          3287 => x"82",
          3288 => x"ff",
          3289 => x"ff",
          3290 => x"e8",
          3291 => x"d8",
          3292 => x"2e",
          3293 => x"b4",
          3294 => x"11",
          3295 => x"05",
          3296 => x"3f",
          3297 => x"08",
          3298 => x"d6",
          3299 => x"fe",
          3300 => x"ff",
          3301 => x"e8",
          3302 => x"d8",
          3303 => x"38",
          3304 => x"08",
          3305 => x"e8",
          3306 => x"ac",
          3307 => x"5c",
          3308 => x"27",
          3309 => x"61",
          3310 => x"70",
          3311 => x"0c",
          3312 => x"f5",
          3313 => x"39",
          3314 => x"80",
          3315 => x"84",
          3316 => x"f8",
          3317 => x"c8",
          3318 => x"fa",
          3319 => x"3d",
          3320 => x"53",
          3321 => x"51",
          3322 => x"82",
          3323 => x"80",
          3324 => x"38",
          3325 => x"f8",
          3326 => x"84",
          3327 => x"cc",
          3328 => x"c8",
          3329 => x"f9",
          3330 => x"bc",
          3331 => x"ab",
          3332 => x"5a",
          3333 => x"81",
          3334 => x"59",
          3335 => x"05",
          3336 => x"34",
          3337 => x"42",
          3338 => x"3d",
          3339 => x"53",
          3340 => x"51",
          3341 => x"82",
          3342 => x"80",
          3343 => x"38",
          3344 => x"fc",
          3345 => x"84",
          3346 => x"80",
          3347 => x"c8",
          3348 => x"f9",
          3349 => x"3d",
          3350 => x"53",
          3351 => x"51",
          3352 => x"82",
          3353 => x"80",
          3354 => x"38",
          3355 => x"51",
          3356 => x"3f",
          3357 => x"63",
          3358 => x"61",
          3359 => x"33",
          3360 => x"78",
          3361 => x"38",
          3362 => x"54",
          3363 => x"79",
          3364 => x"94",
          3365 => x"c0",
          3366 => x"62",
          3367 => x"5a",
          3368 => x"51",
          3369 => x"f8",
          3370 => x"3d",
          3371 => x"53",
          3372 => x"51",
          3373 => x"82",
          3374 => x"80",
          3375 => x"d7",
          3376 => x"78",
          3377 => x"38",
          3378 => x"08",
          3379 => x"39",
          3380 => x"33",
          3381 => x"2e",
          3382 => x"d6",
          3383 => x"bc",
          3384 => x"b6",
          3385 => x"80",
          3386 => x"82",
          3387 => x"44",
          3388 => x"d7",
          3389 => x"78",
          3390 => x"38",
          3391 => x"08",
          3392 => x"82",
          3393 => x"59",
          3394 => x"88",
          3395 => x"8c",
          3396 => x"39",
          3397 => x"08",
          3398 => x"44",
          3399 => x"fc",
          3400 => x"84",
          3401 => x"a4",
          3402 => x"c8",
          3403 => x"38",
          3404 => x"33",
          3405 => x"2e",
          3406 => x"d6",
          3407 => x"80",
          3408 => x"d7",
          3409 => x"78",
          3410 => x"38",
          3411 => x"08",
          3412 => x"82",
          3413 => x"59",
          3414 => x"88",
          3415 => x"80",
          3416 => x"39",
          3417 => x"33",
          3418 => x"2e",
          3419 => x"d7",
          3420 => x"99",
          3421 => x"b2",
          3422 => x"80",
          3423 => x"82",
          3424 => x"43",
          3425 => x"d7",
          3426 => x"05",
          3427 => x"fe",
          3428 => x"ff",
          3429 => x"e4",
          3430 => x"d8",
          3431 => x"2e",
          3432 => x"62",
          3433 => x"88",
          3434 => x"81",
          3435 => x"32",
          3436 => x"72",
          3437 => x"70",
          3438 => x"51",
          3439 => x"80",
          3440 => x"7a",
          3441 => x"38",
          3442 => x"bd",
          3443 => x"93",
          3444 => x"63",
          3445 => x"62",
          3446 => x"ee",
          3447 => x"bd",
          3448 => x"d0",
          3449 => x"ff",
          3450 => x"ff",
          3451 => x"e3",
          3452 => x"d8",
          3453 => x"2e",
          3454 => x"b4",
          3455 => x"11",
          3456 => x"05",
          3457 => x"3f",
          3458 => x"08",
          3459 => x"38",
          3460 => x"80",
          3461 => x"79",
          3462 => x"05",
          3463 => x"fe",
          3464 => x"ff",
          3465 => x"e3",
          3466 => x"d8",
          3467 => x"38",
          3468 => x"63",
          3469 => x"52",
          3470 => x"51",
          3471 => x"3f",
          3472 => x"08",
          3473 => x"52",
          3474 => x"a7",
          3475 => x"45",
          3476 => x"78",
          3477 => x"8a",
          3478 => x"27",
          3479 => x"3d",
          3480 => x"53",
          3481 => x"51",
          3482 => x"82",
          3483 => x"80",
          3484 => x"63",
          3485 => x"cb",
          3486 => x"34",
          3487 => x"44",
          3488 => x"82",
          3489 => x"c2",
          3490 => x"a7",
          3491 => x"fe",
          3492 => x"ff",
          3493 => x"dc",
          3494 => x"d8",
          3495 => x"2e",
          3496 => x"b4",
          3497 => x"11",
          3498 => x"05",
          3499 => x"3f",
          3500 => x"08",
          3501 => x"38",
          3502 => x"be",
          3503 => x"70",
          3504 => x"23",
          3505 => x"3d",
          3506 => x"53",
          3507 => x"51",
          3508 => x"82",
          3509 => x"e0",
          3510 => x"39",
          3511 => x"54",
          3512 => x"d8",
          3513 => x"f0",
          3514 => x"a8",
          3515 => x"f8",
          3516 => x"ff",
          3517 => x"79",
          3518 => x"59",
          3519 => x"f3",
          3520 => x"9f",
          3521 => x"60",
          3522 => x"d0",
          3523 => x"fe",
          3524 => x"ff",
          3525 => x"db",
          3526 => x"d8",
          3527 => x"2e",
          3528 => x"59",
          3529 => x"22",
          3530 => x"05",
          3531 => x"41",
          3532 => x"82",
          3533 => x"c1",
          3534 => x"a0",
          3535 => x"fe",
          3536 => x"ff",
          3537 => x"db",
          3538 => x"d8",
          3539 => x"2e",
          3540 => x"b4",
          3541 => x"11",
          3542 => x"05",
          3543 => x"3f",
          3544 => x"08",
          3545 => x"38",
          3546 => x"0c",
          3547 => x"05",
          3548 => x"fe",
          3549 => x"ff",
          3550 => x"da",
          3551 => x"d8",
          3552 => x"38",
          3553 => x"60",
          3554 => x"52",
          3555 => x"51",
          3556 => x"3f",
          3557 => x"08",
          3558 => x"52",
          3559 => x"a5",
          3560 => x"45",
          3561 => x"78",
          3562 => x"b6",
          3563 => x"27",
          3564 => x"3d",
          3565 => x"53",
          3566 => x"51",
          3567 => x"82",
          3568 => x"80",
          3569 => x"60",
          3570 => x"59",
          3571 => x"41",
          3572 => x"82",
          3573 => x"c0",
          3574 => x"ab",
          3575 => x"f4",
          3576 => x"3f",
          3577 => x"89",
          3578 => x"39",
          3579 => x"51",
          3580 => x"3f",
          3581 => x"dd",
          3582 => x"39",
          3583 => x"51",
          3584 => x"3f",
          3585 => x"0b",
          3586 => x"84",
          3587 => x"81",
          3588 => x"94",
          3589 => x"ca",
          3590 => x"b4",
          3591 => x"c3",
          3592 => x"83",
          3593 => x"94",
          3594 => x"80",
          3595 => x"c0",
          3596 => x"f1",
          3597 => x"3d",
          3598 => x"53",
          3599 => x"51",
          3600 => x"82",
          3601 => x"80",
          3602 => x"38",
          3603 => x"be",
          3604 => x"a3",
          3605 => x"59",
          3606 => x"3d",
          3607 => x"53",
          3608 => x"51",
          3609 => x"82",
          3610 => x"80",
          3611 => x"38",
          3612 => x"be",
          3613 => x"a2",
          3614 => x"59",
          3615 => x"d8",
          3616 => x"2e",
          3617 => x"82",
          3618 => x"52",
          3619 => x"51",
          3620 => x"3f",
          3621 => x"82",
          3622 => x"ff",
          3623 => x"ff",
          3624 => x"f0",
          3625 => x"bf",
          3626 => x"be",
          3627 => x"59",
          3628 => x"91",
          3629 => x"aa",
          3630 => x"79",
          3631 => x"80",
          3632 => x"38",
          3633 => x"59",
          3634 => x"81",
          3635 => x"3d",
          3636 => x"51",
          3637 => x"82",
          3638 => x"5b",
          3639 => x"82",
          3640 => x"7b",
          3641 => x"38",
          3642 => x"8c",
          3643 => x"39",
          3644 => x"ad",
          3645 => x"39",
          3646 => x"56",
          3647 => x"bf",
          3648 => x"53",
          3649 => x"52",
          3650 => x"b0",
          3651 => x"a4",
          3652 => x"39",
          3653 => x"3d",
          3654 => x"51",
          3655 => x"ab",
          3656 => x"82",
          3657 => x"80",
          3658 => x"e4",
          3659 => x"ff",
          3660 => x"ff",
          3661 => x"93",
          3662 => x"80",
          3663 => x"f0",
          3664 => x"ff",
          3665 => x"ff",
          3666 => x"82",
          3667 => x"82",
          3668 => x"80",
          3669 => x"80",
          3670 => x"80",
          3671 => x"80",
          3672 => x"ff",
          3673 => x"e6",
          3674 => x"d8",
          3675 => x"d8",
          3676 => x"70",
          3677 => x"07",
          3678 => x"5b",
          3679 => x"5a",
          3680 => x"83",
          3681 => x"78",
          3682 => x"78",
          3683 => x"38",
          3684 => x"81",
          3685 => x"59",
          3686 => x"38",
          3687 => x"7d",
          3688 => x"59",
          3689 => x"7e",
          3690 => x"81",
          3691 => x"38",
          3692 => x"51",
          3693 => x"3f",
          3694 => x"f5",
          3695 => x"0b",
          3696 => x"34",
          3697 => x"8c",
          3698 => x"55",
          3699 => x"52",
          3700 => x"af",
          3701 => x"c8",
          3702 => x"75",
          3703 => x"87",
          3704 => x"73",
          3705 => x"3f",
          3706 => x"c8",
          3707 => x"0c",
          3708 => x"9c",
          3709 => x"55",
          3710 => x"52",
          3711 => x"83",
          3712 => x"c8",
          3713 => x"75",
          3714 => x"87",
          3715 => x"73",
          3716 => x"3f",
          3717 => x"c8",
          3718 => x"0c",
          3719 => x"0b",
          3720 => x"84",
          3721 => x"83",
          3722 => x"94",
          3723 => x"fa",
          3724 => x"fd",
          3725 => x"02",
          3726 => x"05",
          3727 => x"82",
          3728 => x"87",
          3729 => x"13",
          3730 => x"0c",
          3731 => x"0c",
          3732 => x"3f",
          3733 => x"82",
          3734 => x"ff",
          3735 => x"82",
          3736 => x"ff",
          3737 => x"80",
          3738 => x"92",
          3739 => x"51",
          3740 => x"ec",
          3741 => x"04",
          3742 => x"80",
          3743 => x"71",
          3744 => x"87",
          3745 => x"d8",
          3746 => x"ff",
          3747 => x"ff",
          3748 => x"72",
          3749 => x"38",
          3750 => x"c8",
          3751 => x"0d",
          3752 => x"0d",
          3753 => x"54",
          3754 => x"52",
          3755 => x"2e",
          3756 => x"72",
          3757 => x"a0",
          3758 => x"06",
          3759 => x"13",
          3760 => x"72",
          3761 => x"a2",
          3762 => x"06",
          3763 => x"13",
          3764 => x"72",
          3765 => x"2e",
          3766 => x"9f",
          3767 => x"81",
          3768 => x"72",
          3769 => x"70",
          3770 => x"38",
          3771 => x"80",
          3772 => x"73",
          3773 => x"39",
          3774 => x"80",
          3775 => x"54",
          3776 => x"83",
          3777 => x"70",
          3778 => x"38",
          3779 => x"80",
          3780 => x"54",
          3781 => x"09",
          3782 => x"38",
          3783 => x"a2",
          3784 => x"70",
          3785 => x"07",
          3786 => x"70",
          3787 => x"38",
          3788 => x"81",
          3789 => x"71",
          3790 => x"51",
          3791 => x"c8",
          3792 => x"0d",
          3793 => x"0d",
          3794 => x"08",
          3795 => x"38",
          3796 => x"05",
          3797 => x"d3",
          3798 => x"d8",
          3799 => x"38",
          3800 => x"39",
          3801 => x"82",
          3802 => x"86",
          3803 => x"fc",
          3804 => x"82",
          3805 => x"05",
          3806 => x"52",
          3807 => x"81",
          3808 => x"13",
          3809 => x"51",
          3810 => x"9e",
          3811 => x"38",
          3812 => x"51",
          3813 => x"97",
          3814 => x"38",
          3815 => x"51",
          3816 => x"bb",
          3817 => x"38",
          3818 => x"51",
          3819 => x"bb",
          3820 => x"38",
          3821 => x"55",
          3822 => x"87",
          3823 => x"d9",
          3824 => x"22",
          3825 => x"73",
          3826 => x"80",
          3827 => x"0b",
          3828 => x"9c",
          3829 => x"87",
          3830 => x"0c",
          3831 => x"87",
          3832 => x"0c",
          3833 => x"87",
          3834 => x"0c",
          3835 => x"87",
          3836 => x"0c",
          3837 => x"87",
          3838 => x"0c",
          3839 => x"87",
          3840 => x"0c",
          3841 => x"98",
          3842 => x"87",
          3843 => x"0c",
          3844 => x"c0",
          3845 => x"80",
          3846 => x"d8",
          3847 => x"3d",
          3848 => x"3d",
          3849 => x"87",
          3850 => x"5d",
          3851 => x"87",
          3852 => x"08",
          3853 => x"23",
          3854 => x"b8",
          3855 => x"82",
          3856 => x"c0",
          3857 => x"5a",
          3858 => x"34",
          3859 => x"b0",
          3860 => x"84",
          3861 => x"c0",
          3862 => x"5a",
          3863 => x"34",
          3864 => x"a8",
          3865 => x"86",
          3866 => x"c0",
          3867 => x"5c",
          3868 => x"23",
          3869 => x"a0",
          3870 => x"8a",
          3871 => x"7d",
          3872 => x"ff",
          3873 => x"7b",
          3874 => x"06",
          3875 => x"33",
          3876 => x"33",
          3877 => x"33",
          3878 => x"33",
          3879 => x"33",
          3880 => x"ff",
          3881 => x"82",
          3882 => x"ff",
          3883 => x"8f",
          3884 => x"fb",
          3885 => x"9f",
          3886 => x"d6",
          3887 => x"81",
          3888 => x"55",
          3889 => x"94",
          3890 => x"80",
          3891 => x"87",
          3892 => x"51",
          3893 => x"96",
          3894 => x"06",
          3895 => x"70",
          3896 => x"38",
          3897 => x"70",
          3898 => x"51",
          3899 => x"72",
          3900 => x"81",
          3901 => x"70",
          3902 => x"38",
          3903 => x"70",
          3904 => x"51",
          3905 => x"38",
          3906 => x"06",
          3907 => x"94",
          3908 => x"80",
          3909 => x"87",
          3910 => x"52",
          3911 => x"74",
          3912 => x"0c",
          3913 => x"04",
          3914 => x"02",
          3915 => x"70",
          3916 => x"2a",
          3917 => x"70",
          3918 => x"34",
          3919 => x"04",
          3920 => x"02",
          3921 => x"58",
          3922 => x"09",
          3923 => x"38",
          3924 => x"51",
          3925 => x"d6",
          3926 => x"81",
          3927 => x"56",
          3928 => x"84",
          3929 => x"2e",
          3930 => x"c0",
          3931 => x"72",
          3932 => x"2a",
          3933 => x"55",
          3934 => x"80",
          3935 => x"73",
          3936 => x"81",
          3937 => x"72",
          3938 => x"81",
          3939 => x"06",
          3940 => x"80",
          3941 => x"73",
          3942 => x"81",
          3943 => x"72",
          3944 => x"75",
          3945 => x"53",
          3946 => x"80",
          3947 => x"2e",
          3948 => x"c0",
          3949 => x"77",
          3950 => x"0b",
          3951 => x"0c",
          3952 => x"04",
          3953 => x"79",
          3954 => x"33",
          3955 => x"06",
          3956 => x"70",
          3957 => x"fc",
          3958 => x"ff",
          3959 => x"82",
          3960 => x"70",
          3961 => x"59",
          3962 => x"87",
          3963 => x"51",
          3964 => x"86",
          3965 => x"94",
          3966 => x"08",
          3967 => x"70",
          3968 => x"54",
          3969 => x"2e",
          3970 => x"91",
          3971 => x"06",
          3972 => x"d7",
          3973 => x"32",
          3974 => x"51",
          3975 => x"2e",
          3976 => x"93",
          3977 => x"06",
          3978 => x"ff",
          3979 => x"81",
          3980 => x"87",
          3981 => x"52",
          3982 => x"86",
          3983 => x"94",
          3984 => x"72",
          3985 => x"74",
          3986 => x"ff",
          3987 => x"57",
          3988 => x"38",
          3989 => x"c8",
          3990 => x"0d",
          3991 => x"0d",
          3992 => x"33",
          3993 => x"06",
          3994 => x"c0",
          3995 => x"72",
          3996 => x"38",
          3997 => x"94",
          3998 => x"70",
          3999 => x"81",
          4000 => x"51",
          4001 => x"e2",
          4002 => x"ff",
          4003 => x"c0",
          4004 => x"70",
          4005 => x"38",
          4006 => x"90",
          4007 => x"70",
          4008 => x"82",
          4009 => x"51",
          4010 => x"04",
          4011 => x"82",
          4012 => x"81",
          4013 => x"d8",
          4014 => x"fe",
          4015 => x"d6",
          4016 => x"81",
          4017 => x"53",
          4018 => x"84",
          4019 => x"2e",
          4020 => x"c0",
          4021 => x"71",
          4022 => x"2a",
          4023 => x"51",
          4024 => x"52",
          4025 => x"a0",
          4026 => x"ff",
          4027 => x"c0",
          4028 => x"70",
          4029 => x"38",
          4030 => x"90",
          4031 => x"70",
          4032 => x"98",
          4033 => x"51",
          4034 => x"c8",
          4035 => x"0d",
          4036 => x"0d",
          4037 => x"80",
          4038 => x"2a",
          4039 => x"51",
          4040 => x"84",
          4041 => x"c0",
          4042 => x"82",
          4043 => x"87",
          4044 => x"08",
          4045 => x"0c",
          4046 => x"94",
          4047 => x"f4",
          4048 => x"9e",
          4049 => x"d6",
          4050 => x"c0",
          4051 => x"82",
          4052 => x"87",
          4053 => x"08",
          4054 => x"0c",
          4055 => x"ac",
          4056 => x"84",
          4057 => x"9e",
          4058 => x"d7",
          4059 => x"c0",
          4060 => x"82",
          4061 => x"87",
          4062 => x"08",
          4063 => x"0c",
          4064 => x"bc",
          4065 => x"94",
          4066 => x"9e",
          4067 => x"d7",
          4068 => x"c0",
          4069 => x"82",
          4070 => x"87",
          4071 => x"08",
          4072 => x"d7",
          4073 => x"c0",
          4074 => x"82",
          4075 => x"87",
          4076 => x"08",
          4077 => x"0c",
          4078 => x"8c",
          4079 => x"ac",
          4080 => x"82",
          4081 => x"80",
          4082 => x"9e",
          4083 => x"84",
          4084 => x"51",
          4085 => x"80",
          4086 => x"81",
          4087 => x"d7",
          4088 => x"0b",
          4089 => x"90",
          4090 => x"80",
          4091 => x"52",
          4092 => x"2e",
          4093 => x"52",
          4094 => x"b2",
          4095 => x"87",
          4096 => x"08",
          4097 => x"0a",
          4098 => x"52",
          4099 => x"83",
          4100 => x"71",
          4101 => x"34",
          4102 => x"c0",
          4103 => x"70",
          4104 => x"06",
          4105 => x"70",
          4106 => x"38",
          4107 => x"82",
          4108 => x"80",
          4109 => x"9e",
          4110 => x"a0",
          4111 => x"51",
          4112 => x"80",
          4113 => x"81",
          4114 => x"d7",
          4115 => x"0b",
          4116 => x"90",
          4117 => x"80",
          4118 => x"52",
          4119 => x"2e",
          4120 => x"52",
          4121 => x"b6",
          4122 => x"87",
          4123 => x"08",
          4124 => x"80",
          4125 => x"52",
          4126 => x"83",
          4127 => x"71",
          4128 => x"34",
          4129 => x"c0",
          4130 => x"70",
          4131 => x"06",
          4132 => x"70",
          4133 => x"38",
          4134 => x"82",
          4135 => x"80",
          4136 => x"9e",
          4137 => x"81",
          4138 => x"51",
          4139 => x"80",
          4140 => x"81",
          4141 => x"d7",
          4142 => x"0b",
          4143 => x"90",
          4144 => x"c0",
          4145 => x"52",
          4146 => x"2e",
          4147 => x"52",
          4148 => x"ba",
          4149 => x"87",
          4150 => x"08",
          4151 => x"06",
          4152 => x"70",
          4153 => x"38",
          4154 => x"82",
          4155 => x"87",
          4156 => x"08",
          4157 => x"06",
          4158 => x"51",
          4159 => x"82",
          4160 => x"80",
          4161 => x"9e",
          4162 => x"84",
          4163 => x"52",
          4164 => x"2e",
          4165 => x"52",
          4166 => x"bd",
          4167 => x"9e",
          4168 => x"83",
          4169 => x"84",
          4170 => x"51",
          4171 => x"be",
          4172 => x"87",
          4173 => x"08",
          4174 => x"51",
          4175 => x"80",
          4176 => x"81",
          4177 => x"d7",
          4178 => x"c0",
          4179 => x"70",
          4180 => x"51",
          4181 => x"c0",
          4182 => x"0d",
          4183 => x"0d",
          4184 => x"51",
          4185 => x"3f",
          4186 => x"33",
          4187 => x"2e",
          4188 => x"c0",
          4189 => x"90",
          4190 => x"c0",
          4191 => x"ac",
          4192 => x"d7",
          4193 => x"73",
          4194 => x"38",
          4195 => x"08",
          4196 => x"08",
          4197 => x"82",
          4198 => x"ff",
          4199 => x"82",
          4200 => x"54",
          4201 => x"94",
          4202 => x"84",
          4203 => x"88",
          4204 => x"52",
          4205 => x"51",
          4206 => x"3f",
          4207 => x"33",
          4208 => x"2e",
          4209 => x"d6",
          4210 => x"d6",
          4211 => x"54",
          4212 => x"bc",
          4213 => x"80",
          4214 => x"b5",
          4215 => x"80",
          4216 => x"82",
          4217 => x"82",
          4218 => x"11",
          4219 => x"c1",
          4220 => x"8f",
          4221 => x"d7",
          4222 => x"73",
          4223 => x"38",
          4224 => x"08",
          4225 => x"08",
          4226 => x"82",
          4227 => x"ff",
          4228 => x"82",
          4229 => x"54",
          4230 => x"8e",
          4231 => x"bc",
          4232 => x"c2",
          4233 => x"8f",
          4234 => x"d7",
          4235 => x"73",
          4236 => x"38",
          4237 => x"33",
          4238 => x"b0",
          4239 => x"98",
          4240 => x"bd",
          4241 => x"80",
          4242 => x"82",
          4243 => x"52",
          4244 => x"51",
          4245 => x"3f",
          4246 => x"33",
          4247 => x"2e",
          4248 => x"c2",
          4249 => x"aa",
          4250 => x"d7",
          4251 => x"73",
          4252 => x"38",
          4253 => x"51",
          4254 => x"3f",
          4255 => x"33",
          4256 => x"2e",
          4257 => x"c3",
          4258 => x"aa",
          4259 => x"d7",
          4260 => x"73",
          4261 => x"38",
          4262 => x"51",
          4263 => x"3f",
          4264 => x"33",
          4265 => x"2e",
          4266 => x"c3",
          4267 => x"aa",
          4268 => x"c3",
          4269 => x"aa",
          4270 => x"d7",
          4271 => x"82",
          4272 => x"ff",
          4273 => x"82",
          4274 => x"52",
          4275 => x"51",
          4276 => x"3f",
          4277 => x"08",
          4278 => x"88",
          4279 => x"f8",
          4280 => x"b0",
          4281 => x"fb",
          4282 => x"a0",
          4283 => x"c4",
          4284 => x"8d",
          4285 => x"d7",
          4286 => x"bd",
          4287 => x"75",
          4288 => x"3f",
          4289 => x"08",
          4290 => x"29",
          4291 => x"54",
          4292 => x"c8",
          4293 => x"c4",
          4294 => x"8d",
          4295 => x"d7",
          4296 => x"73",
          4297 => x"38",
          4298 => x"08",
          4299 => x"c0",
          4300 => x"c0",
          4301 => x"d8",
          4302 => x"84",
          4303 => x"71",
          4304 => x"82",
          4305 => x"52",
          4306 => x"51",
          4307 => x"3f",
          4308 => x"33",
          4309 => x"2e",
          4310 => x"d7",
          4311 => x"bd",
          4312 => x"75",
          4313 => x"3f",
          4314 => x"08",
          4315 => x"29",
          4316 => x"54",
          4317 => x"c8",
          4318 => x"c5",
          4319 => x"8c",
          4320 => x"51",
          4321 => x"3f",
          4322 => x"04",
          4323 => x"02",
          4324 => x"ff",
          4325 => x"84",
          4326 => x"71",
          4327 => x"af",
          4328 => x"71",
          4329 => x"c5",
          4330 => x"39",
          4331 => x"51",
          4332 => x"c5",
          4333 => x"39",
          4334 => x"51",
          4335 => x"c6",
          4336 => x"39",
          4337 => x"51",
          4338 => x"3f",
          4339 => x"04",
          4340 => x"0c",
          4341 => x"0d",
          4342 => x"84",
          4343 => x"52",
          4344 => x"70",
          4345 => x"82",
          4346 => x"72",
          4347 => x"0d",
          4348 => x"0d",
          4349 => x"84",
          4350 => x"d7",
          4351 => x"80",
          4352 => x"09",
          4353 => x"c4",
          4354 => x"82",
          4355 => x"73",
          4356 => x"3d",
          4357 => x"0b",
          4358 => x"84",
          4359 => x"d7",
          4360 => x"c0",
          4361 => x"04",
          4362 => x"76",
          4363 => x"98",
          4364 => x"2b",
          4365 => x"72",
          4366 => x"82",
          4367 => x"51",
          4368 => x"80",
          4369 => x"94",
          4370 => x"53",
          4371 => x"9c",
          4372 => x"90",
          4373 => x"02",
          4374 => x"05",
          4375 => x"52",
          4376 => x"72",
          4377 => x"06",
          4378 => x"53",
          4379 => x"c8",
          4380 => x"0d",
          4381 => x"0d",
          4382 => x"05",
          4383 => x"71",
          4384 => x"54",
          4385 => x"b1",
          4386 => x"ac",
          4387 => x"51",
          4388 => x"3f",
          4389 => x"08",
          4390 => x"ff",
          4391 => x"82",
          4392 => x"52",
          4393 => x"aa",
          4394 => x"33",
          4395 => x"72",
          4396 => x"81",
          4397 => x"cc",
          4398 => x"ff",
          4399 => x"74",
          4400 => x"3d",
          4401 => x"3d",
          4402 => x"84",
          4403 => x"33",
          4404 => x"bb",
          4405 => x"d8",
          4406 => x"84",
          4407 => x"c8",
          4408 => x"51",
          4409 => x"58",
          4410 => x"2e",
          4411 => x"51",
          4412 => x"82",
          4413 => x"70",
          4414 => x"d7",
          4415 => x"19",
          4416 => x"56",
          4417 => x"3f",
          4418 => x"08",
          4419 => x"d8",
          4420 => x"84",
          4421 => x"c8",
          4422 => x"51",
          4423 => x"80",
          4424 => x"75",
          4425 => x"74",
          4426 => x"b9",
          4427 => x"a0",
          4428 => x"55",
          4429 => x"a0",
          4430 => x"ff",
          4431 => x"75",
          4432 => x"80",
          4433 => x"a0",
          4434 => x"2e",
          4435 => x"d8",
          4436 => x"75",
          4437 => x"38",
          4438 => x"33",
          4439 => x"38",
          4440 => x"05",
          4441 => x"78",
          4442 => x"80",
          4443 => x"82",
          4444 => x"52",
          4445 => x"a0",
          4446 => x"d8",
          4447 => x"80",
          4448 => x"8c",
          4449 => x"fd",
          4450 => x"d7",
          4451 => x"54",
          4452 => x"71",
          4453 => x"38",
          4454 => x"d0",
          4455 => x"0c",
          4456 => x"14",
          4457 => x"80",
          4458 => x"80",
          4459 => x"a0",
          4460 => x"9c",
          4461 => x"80",
          4462 => x"71",
          4463 => x"86",
          4464 => x"9c",
          4465 => x"a4",
          4466 => x"82",
          4467 => x"85",
          4468 => x"dc",
          4469 => x"57",
          4470 => x"d8",
          4471 => x"80",
          4472 => x"82",
          4473 => x"80",
          4474 => x"d8",
          4475 => x"80",
          4476 => x"3d",
          4477 => x"81",
          4478 => x"82",
          4479 => x"80",
          4480 => x"75",
          4481 => x"fd",
          4482 => x"c8",
          4483 => x"0b",
          4484 => x"08",
          4485 => x"82",
          4486 => x"ff",
          4487 => x"55",
          4488 => x"34",
          4489 => x"52",
          4490 => x"c9",
          4491 => x"ff",
          4492 => x"74",
          4493 => x"81",
          4494 => x"38",
          4495 => x"04",
          4496 => x"aa",
          4497 => x"3d",
          4498 => x"81",
          4499 => x"80",
          4500 => x"9c",
          4501 => x"f4",
          4502 => x"d8",
          4503 => x"95",
          4504 => x"82",
          4505 => x"54",
          4506 => x"52",
          4507 => x"52",
          4508 => x"d8",
          4509 => x"c8",
          4510 => x"a5",
          4511 => x"ff",
          4512 => x"82",
          4513 => x"81",
          4514 => x"80",
          4515 => x"c8",
          4516 => x"38",
          4517 => x"08",
          4518 => x"17",
          4519 => x"74",
          4520 => x"70",
          4521 => x"07",
          4522 => x"55",
          4523 => x"2e",
          4524 => x"ff",
          4525 => x"d8",
          4526 => x"11",
          4527 => x"80",
          4528 => x"82",
          4529 => x"80",
          4530 => x"82",
          4531 => x"ff",
          4532 => x"78",
          4533 => x"81",
          4534 => x"75",
          4535 => x"ff",
          4536 => x"79",
          4537 => x"9d",
          4538 => x"08",
          4539 => x"c8",
          4540 => x"80",
          4541 => x"d8",
          4542 => x"3d",
          4543 => x"3d",
          4544 => x"71",
          4545 => x"33",
          4546 => x"58",
          4547 => x"09",
          4548 => x"38",
          4549 => x"05",
          4550 => x"27",
          4551 => x"17",
          4552 => x"71",
          4553 => x"55",
          4554 => x"09",
          4555 => x"38",
          4556 => x"ea",
          4557 => x"73",
          4558 => x"d8",
          4559 => x"08",
          4560 => x"ad",
          4561 => x"d8",
          4562 => x"79",
          4563 => x"51",
          4564 => x"3f",
          4565 => x"08",
          4566 => x"84",
          4567 => x"74",
          4568 => x"38",
          4569 => x"88",
          4570 => x"fc",
          4571 => x"39",
          4572 => x"8c",
          4573 => x"53",
          4574 => x"c0",
          4575 => x"d8",
          4576 => x"2e",
          4577 => x"1b",
          4578 => x"77",
          4579 => x"3f",
          4580 => x"08",
          4581 => x"55",
          4582 => x"74",
          4583 => x"81",
          4584 => x"ff",
          4585 => x"82",
          4586 => x"8b",
          4587 => x"73",
          4588 => x"0c",
          4589 => x"04",
          4590 => x"b0",
          4591 => x"3d",
          4592 => x"08",
          4593 => x"80",
          4594 => x"34",
          4595 => x"33",
          4596 => x"08",
          4597 => x"81",
          4598 => x"82",
          4599 => x"55",
          4600 => x"38",
          4601 => x"80",
          4602 => x"38",
          4603 => x"06",
          4604 => x"80",
          4605 => x"38",
          4606 => x"86",
          4607 => x"c8",
          4608 => x"9c",
          4609 => x"c8",
          4610 => x"81",
          4611 => x"53",
          4612 => x"d8",
          4613 => x"80",
          4614 => x"82",
          4615 => x"80",
          4616 => x"82",
          4617 => x"ff",
          4618 => x"80",
          4619 => x"d8",
          4620 => x"82",
          4621 => x"53",
          4622 => x"90",
          4623 => x"54",
          4624 => x"3f",
          4625 => x"08",
          4626 => x"c8",
          4627 => x"09",
          4628 => x"d0",
          4629 => x"c8",
          4630 => x"ab",
          4631 => x"d8",
          4632 => x"80",
          4633 => x"c8",
          4634 => x"38",
          4635 => x"08",
          4636 => x"17",
          4637 => x"74",
          4638 => x"74",
          4639 => x"52",
          4640 => x"c2",
          4641 => x"70",
          4642 => x"5c",
          4643 => x"27",
          4644 => x"5b",
          4645 => x"09",
          4646 => x"97",
          4647 => x"75",
          4648 => x"34",
          4649 => x"82",
          4650 => x"80",
          4651 => x"f9",
          4652 => x"3d",
          4653 => x"3f",
          4654 => x"08",
          4655 => x"98",
          4656 => x"78",
          4657 => x"38",
          4658 => x"06",
          4659 => x"33",
          4660 => x"70",
          4661 => x"f0",
          4662 => x"98",
          4663 => x"2c",
          4664 => x"05",
          4665 => x"82",
          4666 => x"70",
          4667 => x"33",
          4668 => x"51",
          4669 => x"59",
          4670 => x"56",
          4671 => x"80",
          4672 => x"74",
          4673 => x"74",
          4674 => x"29",
          4675 => x"05",
          4676 => x"51",
          4677 => x"24",
          4678 => x"76",
          4679 => x"77",
          4680 => x"3f",
          4681 => x"08",
          4682 => x"54",
          4683 => x"d7",
          4684 => x"f0",
          4685 => x"56",
          4686 => x"81",
          4687 => x"81",
          4688 => x"70",
          4689 => x"81",
          4690 => x"51",
          4691 => x"26",
          4692 => x"53",
          4693 => x"51",
          4694 => x"82",
          4695 => x"81",
          4696 => x"73",
          4697 => x"39",
          4698 => x"80",
          4699 => x"38",
          4700 => x"74",
          4701 => x"34",
          4702 => x"70",
          4703 => x"f0",
          4704 => x"98",
          4705 => x"2c",
          4706 => x"70",
          4707 => x"c6",
          4708 => x"5e",
          4709 => x"57",
          4710 => x"74",
          4711 => x"81",
          4712 => x"38",
          4713 => x"14",
          4714 => x"80",
          4715 => x"84",
          4716 => x"82",
          4717 => x"92",
          4718 => x"f0",
          4719 => x"82",
          4720 => x"78",
          4721 => x"75",
          4722 => x"54",
          4723 => x"fd",
          4724 => x"84",
          4725 => x"d8",
          4726 => x"08",
          4727 => x"8c",
          4728 => x"7e",
          4729 => x"38",
          4730 => x"33",
          4731 => x"27",
          4732 => x"98",
          4733 => x"2c",
          4734 => x"75",
          4735 => x"74",
          4736 => x"33",
          4737 => x"74",
          4738 => x"29",
          4739 => x"05",
          4740 => x"82",
          4741 => x"56",
          4742 => x"39",
          4743 => x"33",
          4744 => x"54",
          4745 => x"8c",
          4746 => x"54",
          4747 => x"74",
          4748 => x"88",
          4749 => x"7e",
          4750 => x"81",
          4751 => x"82",
          4752 => x"82",
          4753 => x"70",
          4754 => x"29",
          4755 => x"05",
          4756 => x"82",
          4757 => x"5a",
          4758 => x"74",
          4759 => x"38",
          4760 => x"08",
          4761 => x"70",
          4762 => x"ff",
          4763 => x"74",
          4764 => x"29",
          4765 => x"05",
          4766 => x"82",
          4767 => x"56",
          4768 => x"75",
          4769 => x"82",
          4770 => x"70",
          4771 => x"98",
          4772 => x"88",
          4773 => x"56",
          4774 => x"25",
          4775 => x"82",
          4776 => x"52",
          4777 => x"9e",
          4778 => x"81",
          4779 => x"81",
          4780 => x"70",
          4781 => x"f0",
          4782 => x"51",
          4783 => x"24",
          4784 => x"ee",
          4785 => x"34",
          4786 => x"1b",
          4787 => x"8c",
          4788 => x"82",
          4789 => x"f3",
          4790 => x"fd",
          4791 => x"8c",
          4792 => x"ff",
          4793 => x"73",
          4794 => x"c6",
          4795 => x"88",
          4796 => x"54",
          4797 => x"88",
          4798 => x"54",
          4799 => x"8c",
          4800 => x"ac",
          4801 => x"51",
          4802 => x"3f",
          4803 => x"33",
          4804 => x"70",
          4805 => x"f0",
          4806 => x"51",
          4807 => x"74",
          4808 => x"74",
          4809 => x"14",
          4810 => x"82",
          4811 => x"52",
          4812 => x"ff",
          4813 => x"74",
          4814 => x"29",
          4815 => x"05",
          4816 => x"82",
          4817 => x"58",
          4818 => x"75",
          4819 => x"82",
          4820 => x"52",
          4821 => x"9c",
          4822 => x"f0",
          4823 => x"98",
          4824 => x"2c",
          4825 => x"33",
          4826 => x"57",
          4827 => x"fa",
          4828 => x"f4",
          4829 => x"88",
          4830 => x"b6",
          4831 => x"80",
          4832 => x"80",
          4833 => x"98",
          4834 => x"88",
          4835 => x"55",
          4836 => x"de",
          4837 => x"39",
          4838 => x"33",
          4839 => x"80",
          4840 => x"f4",
          4841 => x"8a",
          4842 => x"86",
          4843 => x"88",
          4844 => x"f6",
          4845 => x"d8",
          4846 => x"ff",
          4847 => x"96",
          4848 => x"88",
          4849 => x"80",
          4850 => x"81",
          4851 => x"79",
          4852 => x"3f",
          4853 => x"7a",
          4854 => x"82",
          4855 => x"80",
          4856 => x"88",
          4857 => x"d8",
          4858 => x"3d",
          4859 => x"f0",
          4860 => x"73",
          4861 => x"ba",
          4862 => x"ac",
          4863 => x"51",
          4864 => x"3f",
          4865 => x"33",
          4866 => x"73",
          4867 => x"34",
          4868 => x"06",
          4869 => x"82",
          4870 => x"82",
          4871 => x"55",
          4872 => x"2e",
          4873 => x"ff",
          4874 => x"82",
          4875 => x"74",
          4876 => x"98",
          4877 => x"ff",
          4878 => x"55",
          4879 => x"ad",
          4880 => x"54",
          4881 => x"74",
          4882 => x"ac",
          4883 => x"33",
          4884 => x"de",
          4885 => x"80",
          4886 => x"80",
          4887 => x"98",
          4888 => x"88",
          4889 => x"55",
          4890 => x"d5",
          4891 => x"ac",
          4892 => x"51",
          4893 => x"3f",
          4894 => x"33",
          4895 => x"70",
          4896 => x"f0",
          4897 => x"51",
          4898 => x"74",
          4899 => x"38",
          4900 => x"08",
          4901 => x"ff",
          4902 => x"74",
          4903 => x"29",
          4904 => x"05",
          4905 => x"82",
          4906 => x"58",
          4907 => x"75",
          4908 => x"f7",
          4909 => x"f0",
          4910 => x"81",
          4911 => x"f0",
          4912 => x"56",
          4913 => x"27",
          4914 => x"82",
          4915 => x"52",
          4916 => x"73",
          4917 => x"34",
          4918 => x"33",
          4919 => x"99",
          4920 => x"f0",
          4921 => x"81",
          4922 => x"f0",
          4923 => x"56",
          4924 => x"26",
          4925 => x"ba",
          4926 => x"8c",
          4927 => x"82",
          4928 => x"ee",
          4929 => x"0b",
          4930 => x"34",
          4931 => x"f0",
          4932 => x"9e",
          4933 => x"38",
          4934 => x"08",
          4935 => x"2e",
          4936 => x"51",
          4937 => x"3f",
          4938 => x"08",
          4939 => x"34",
          4940 => x"08",
          4941 => x"81",
          4942 => x"52",
          4943 => x"a3",
          4944 => x"5b",
          4945 => x"7a",
          4946 => x"d7",
          4947 => x"11",
          4948 => x"74",
          4949 => x"38",
          4950 => x"a1",
          4951 => x"d8",
          4952 => x"f0",
          4953 => x"d8",
          4954 => x"ff",
          4955 => x"53",
          4956 => x"51",
          4957 => x"3f",
          4958 => x"80",
          4959 => x"08",
          4960 => x"2e",
          4961 => x"74",
          4962 => x"f9",
          4963 => x"7a",
          4964 => x"81",
          4965 => x"82",
          4966 => x"55",
          4967 => x"a4",
          4968 => x"ff",
          4969 => x"82",
          4970 => x"82",
          4971 => x"82",
          4972 => x"81",
          4973 => x"05",
          4974 => x"79",
          4975 => x"a5",
          4976 => x"39",
          4977 => x"82",
          4978 => x"70",
          4979 => x"74",
          4980 => x"38",
          4981 => x"a0",
          4982 => x"d8",
          4983 => x"f0",
          4984 => x"d8",
          4985 => x"ff",
          4986 => x"53",
          4987 => x"51",
          4988 => x"3f",
          4989 => x"73",
          4990 => x"5b",
          4991 => x"82",
          4992 => x"74",
          4993 => x"f0",
          4994 => x"f0",
          4995 => x"79",
          4996 => x"3f",
          4997 => x"82",
          4998 => x"70",
          4999 => x"82",
          5000 => x"59",
          5001 => x"77",
          5002 => x"38",
          5003 => x"08",
          5004 => x"54",
          5005 => x"8c",
          5006 => x"70",
          5007 => x"ff",
          5008 => x"f4",
          5009 => x"f0",
          5010 => x"73",
          5011 => x"e2",
          5012 => x"ac",
          5013 => x"51",
          5014 => x"3f",
          5015 => x"33",
          5016 => x"73",
          5017 => x"34",
          5018 => x"f9",
          5019 => x"c0",
          5020 => x"d8",
          5021 => x"80",
          5022 => x"bc",
          5023 => x"53",
          5024 => x"c0",
          5025 => x"a5",
          5026 => x"d8",
          5027 => x"80",
          5028 => x"34",
          5029 => x"81",
          5030 => x"d8",
          5031 => x"77",
          5032 => x"76",
          5033 => x"82",
          5034 => x"54",
          5035 => x"34",
          5036 => x"34",
          5037 => x"08",
          5038 => x"22",
          5039 => x"80",
          5040 => x"83",
          5041 => x"70",
          5042 => x"51",
          5043 => x"88",
          5044 => x"89",
          5045 => x"d8",
          5046 => x"88",
          5047 => x"c0",
          5048 => x"11",
          5049 => x"77",
          5050 => x"76",
          5051 => x"89",
          5052 => x"ff",
          5053 => x"52",
          5054 => x"72",
          5055 => x"fb",
          5056 => x"82",
          5057 => x"ff",
          5058 => x"51",
          5059 => x"d8",
          5060 => x"3d",
          5061 => x"3d",
          5062 => x"05",
          5063 => x"05",
          5064 => x"71",
          5065 => x"c0",
          5066 => x"2b",
          5067 => x"83",
          5068 => x"70",
          5069 => x"33",
          5070 => x"07",
          5071 => x"ae",
          5072 => x"81",
          5073 => x"07",
          5074 => x"53",
          5075 => x"54",
          5076 => x"53",
          5077 => x"77",
          5078 => x"18",
          5079 => x"c0",
          5080 => x"88",
          5081 => x"70",
          5082 => x"74",
          5083 => x"82",
          5084 => x"70",
          5085 => x"81",
          5086 => x"88",
          5087 => x"83",
          5088 => x"f8",
          5089 => x"56",
          5090 => x"73",
          5091 => x"06",
          5092 => x"54",
          5093 => x"82",
          5094 => x"81",
          5095 => x"72",
          5096 => x"82",
          5097 => x"16",
          5098 => x"34",
          5099 => x"34",
          5100 => x"04",
          5101 => x"82",
          5102 => x"02",
          5103 => x"05",
          5104 => x"2b",
          5105 => x"11",
          5106 => x"33",
          5107 => x"71",
          5108 => x"58",
          5109 => x"55",
          5110 => x"84",
          5111 => x"13",
          5112 => x"2b",
          5113 => x"2a",
          5114 => x"52",
          5115 => x"34",
          5116 => x"34",
          5117 => x"08",
          5118 => x"11",
          5119 => x"33",
          5120 => x"71",
          5121 => x"56",
          5122 => x"72",
          5123 => x"33",
          5124 => x"71",
          5125 => x"70",
          5126 => x"56",
          5127 => x"86",
          5128 => x"87",
          5129 => x"d8",
          5130 => x"70",
          5131 => x"33",
          5132 => x"07",
          5133 => x"ff",
          5134 => x"2a",
          5135 => x"53",
          5136 => x"34",
          5137 => x"34",
          5138 => x"04",
          5139 => x"02",
          5140 => x"82",
          5141 => x"71",
          5142 => x"11",
          5143 => x"12",
          5144 => x"2b",
          5145 => x"29",
          5146 => x"81",
          5147 => x"98",
          5148 => x"2b",
          5149 => x"53",
          5150 => x"56",
          5151 => x"71",
          5152 => x"f6",
          5153 => x"fe",
          5154 => x"d8",
          5155 => x"16",
          5156 => x"12",
          5157 => x"2b",
          5158 => x"07",
          5159 => x"33",
          5160 => x"71",
          5161 => x"70",
          5162 => x"ff",
          5163 => x"52",
          5164 => x"5a",
          5165 => x"05",
          5166 => x"54",
          5167 => x"13",
          5168 => x"13",
          5169 => x"c0",
          5170 => x"70",
          5171 => x"33",
          5172 => x"71",
          5173 => x"56",
          5174 => x"72",
          5175 => x"81",
          5176 => x"88",
          5177 => x"81",
          5178 => x"70",
          5179 => x"51",
          5180 => x"72",
          5181 => x"81",
          5182 => x"3d",
          5183 => x"3d",
          5184 => x"c0",
          5185 => x"05",
          5186 => x"70",
          5187 => x"11",
          5188 => x"83",
          5189 => x"8b",
          5190 => x"2b",
          5191 => x"59",
          5192 => x"73",
          5193 => x"81",
          5194 => x"88",
          5195 => x"8c",
          5196 => x"22",
          5197 => x"88",
          5198 => x"53",
          5199 => x"73",
          5200 => x"14",
          5201 => x"c0",
          5202 => x"70",
          5203 => x"33",
          5204 => x"71",
          5205 => x"56",
          5206 => x"72",
          5207 => x"33",
          5208 => x"71",
          5209 => x"70",
          5210 => x"55",
          5211 => x"82",
          5212 => x"83",
          5213 => x"d8",
          5214 => x"82",
          5215 => x"12",
          5216 => x"2b",
          5217 => x"c8",
          5218 => x"87",
          5219 => x"f7",
          5220 => x"82",
          5221 => x"31",
          5222 => x"83",
          5223 => x"70",
          5224 => x"fd",
          5225 => x"d8",
          5226 => x"83",
          5227 => x"82",
          5228 => x"12",
          5229 => x"2b",
          5230 => x"07",
          5231 => x"33",
          5232 => x"71",
          5233 => x"90",
          5234 => x"42",
          5235 => x"5b",
          5236 => x"54",
          5237 => x"8d",
          5238 => x"80",
          5239 => x"fe",
          5240 => x"84",
          5241 => x"33",
          5242 => x"71",
          5243 => x"83",
          5244 => x"11",
          5245 => x"53",
          5246 => x"55",
          5247 => x"34",
          5248 => x"06",
          5249 => x"14",
          5250 => x"c0",
          5251 => x"84",
          5252 => x"13",
          5253 => x"2b",
          5254 => x"2a",
          5255 => x"56",
          5256 => x"16",
          5257 => x"16",
          5258 => x"c0",
          5259 => x"80",
          5260 => x"34",
          5261 => x"14",
          5262 => x"c0",
          5263 => x"84",
          5264 => x"85",
          5265 => x"d8",
          5266 => x"70",
          5267 => x"33",
          5268 => x"07",
          5269 => x"80",
          5270 => x"2a",
          5271 => x"56",
          5272 => x"34",
          5273 => x"34",
          5274 => x"04",
          5275 => x"73",
          5276 => x"c0",
          5277 => x"f7",
          5278 => x"80",
          5279 => x"71",
          5280 => x"3f",
          5281 => x"04",
          5282 => x"80",
          5283 => x"f8",
          5284 => x"d8",
          5285 => x"ff",
          5286 => x"d8",
          5287 => x"11",
          5288 => x"33",
          5289 => x"07",
          5290 => x"56",
          5291 => x"ff",
          5292 => x"78",
          5293 => x"38",
          5294 => x"17",
          5295 => x"12",
          5296 => x"2b",
          5297 => x"ff",
          5298 => x"31",
          5299 => x"ff",
          5300 => x"27",
          5301 => x"56",
          5302 => x"79",
          5303 => x"73",
          5304 => x"38",
          5305 => x"5b",
          5306 => x"85",
          5307 => x"88",
          5308 => x"54",
          5309 => x"78",
          5310 => x"2e",
          5311 => x"79",
          5312 => x"76",
          5313 => x"d8",
          5314 => x"70",
          5315 => x"33",
          5316 => x"07",
          5317 => x"ff",
          5318 => x"5a",
          5319 => x"73",
          5320 => x"38",
          5321 => x"54",
          5322 => x"81",
          5323 => x"54",
          5324 => x"81",
          5325 => x"7a",
          5326 => x"06",
          5327 => x"51",
          5328 => x"81",
          5329 => x"80",
          5330 => x"52",
          5331 => x"c6",
          5332 => x"c0",
          5333 => x"86",
          5334 => x"12",
          5335 => x"2b",
          5336 => x"07",
          5337 => x"55",
          5338 => x"17",
          5339 => x"ff",
          5340 => x"2a",
          5341 => x"54",
          5342 => x"34",
          5343 => x"06",
          5344 => x"15",
          5345 => x"c0",
          5346 => x"2b",
          5347 => x"1e",
          5348 => x"87",
          5349 => x"88",
          5350 => x"88",
          5351 => x"5e",
          5352 => x"54",
          5353 => x"34",
          5354 => x"34",
          5355 => x"08",
          5356 => x"11",
          5357 => x"33",
          5358 => x"71",
          5359 => x"53",
          5360 => x"74",
          5361 => x"86",
          5362 => x"87",
          5363 => x"d8",
          5364 => x"16",
          5365 => x"11",
          5366 => x"33",
          5367 => x"07",
          5368 => x"53",
          5369 => x"56",
          5370 => x"16",
          5371 => x"16",
          5372 => x"c0",
          5373 => x"05",
          5374 => x"d8",
          5375 => x"3d",
          5376 => x"3d",
          5377 => x"82",
          5378 => x"84",
          5379 => x"3f",
          5380 => x"80",
          5381 => x"71",
          5382 => x"3f",
          5383 => x"08",
          5384 => x"d8",
          5385 => x"3d",
          5386 => x"3d",
          5387 => x"40",
          5388 => x"42",
          5389 => x"c0",
          5390 => x"09",
          5391 => x"38",
          5392 => x"7b",
          5393 => x"51",
          5394 => x"82",
          5395 => x"54",
          5396 => x"7e",
          5397 => x"51",
          5398 => x"7e",
          5399 => x"39",
          5400 => x"8f",
          5401 => x"c8",
          5402 => x"ff",
          5403 => x"c0",
          5404 => x"31",
          5405 => x"83",
          5406 => x"70",
          5407 => x"11",
          5408 => x"12",
          5409 => x"2b",
          5410 => x"31",
          5411 => x"ff",
          5412 => x"29",
          5413 => x"88",
          5414 => x"33",
          5415 => x"71",
          5416 => x"70",
          5417 => x"44",
          5418 => x"41",
          5419 => x"5b",
          5420 => x"5b",
          5421 => x"25",
          5422 => x"81",
          5423 => x"75",
          5424 => x"ff",
          5425 => x"54",
          5426 => x"83",
          5427 => x"88",
          5428 => x"88",
          5429 => x"33",
          5430 => x"71",
          5431 => x"90",
          5432 => x"47",
          5433 => x"54",
          5434 => x"8b",
          5435 => x"31",
          5436 => x"ff",
          5437 => x"77",
          5438 => x"fe",
          5439 => x"54",
          5440 => x"09",
          5441 => x"38",
          5442 => x"c0",
          5443 => x"ff",
          5444 => x"81",
          5445 => x"8e",
          5446 => x"24",
          5447 => x"51",
          5448 => x"81",
          5449 => x"18",
          5450 => x"24",
          5451 => x"79",
          5452 => x"33",
          5453 => x"71",
          5454 => x"53",
          5455 => x"f4",
          5456 => x"78",
          5457 => x"3f",
          5458 => x"08",
          5459 => x"06",
          5460 => x"53",
          5461 => x"82",
          5462 => x"11",
          5463 => x"55",
          5464 => x"b7",
          5465 => x"c0",
          5466 => x"05",
          5467 => x"ff",
          5468 => x"81",
          5469 => x"15",
          5470 => x"24",
          5471 => x"78",
          5472 => x"3f",
          5473 => x"08",
          5474 => x"33",
          5475 => x"71",
          5476 => x"53",
          5477 => x"9c",
          5478 => x"78",
          5479 => x"3f",
          5480 => x"08",
          5481 => x"06",
          5482 => x"53",
          5483 => x"82",
          5484 => x"11",
          5485 => x"55",
          5486 => x"df",
          5487 => x"c0",
          5488 => x"05",
          5489 => x"19",
          5490 => x"83",
          5491 => x"58",
          5492 => x"7f",
          5493 => x"b0",
          5494 => x"c8",
          5495 => x"d8",
          5496 => x"2e",
          5497 => x"53",
          5498 => x"d8",
          5499 => x"ff",
          5500 => x"73",
          5501 => x"3f",
          5502 => x"78",
          5503 => x"80",
          5504 => x"78",
          5505 => x"3f",
          5506 => x"2b",
          5507 => x"08",
          5508 => x"51",
          5509 => x"7b",
          5510 => x"d8",
          5511 => x"3d",
          5512 => x"3d",
          5513 => x"29",
          5514 => x"fb",
          5515 => x"d8",
          5516 => x"82",
          5517 => x"80",
          5518 => x"73",
          5519 => x"82",
          5520 => x"51",
          5521 => x"3f",
          5522 => x"c8",
          5523 => x"0d",
          5524 => x"0d",
          5525 => x"33",
          5526 => x"70",
          5527 => x"38",
          5528 => x"11",
          5529 => x"82",
          5530 => x"83",
          5531 => x"fc",
          5532 => x"9b",
          5533 => x"84",
          5534 => x"33",
          5535 => x"51",
          5536 => x"80",
          5537 => x"84",
          5538 => x"92",
          5539 => x"51",
          5540 => x"80",
          5541 => x"81",
          5542 => x"72",
          5543 => x"92",
          5544 => x"81",
          5545 => x"0b",
          5546 => x"8c",
          5547 => x"71",
          5548 => x"06",
          5549 => x"80",
          5550 => x"87",
          5551 => x"08",
          5552 => x"38",
          5553 => x"80",
          5554 => x"71",
          5555 => x"c0",
          5556 => x"51",
          5557 => x"87",
          5558 => x"d8",
          5559 => x"82",
          5560 => x"33",
          5561 => x"d8",
          5562 => x"3d",
          5563 => x"3d",
          5564 => x"64",
          5565 => x"bf",
          5566 => x"40",
          5567 => x"74",
          5568 => x"cd",
          5569 => x"c8",
          5570 => x"7a",
          5571 => x"81",
          5572 => x"72",
          5573 => x"87",
          5574 => x"11",
          5575 => x"8c",
          5576 => x"92",
          5577 => x"5a",
          5578 => x"58",
          5579 => x"c0",
          5580 => x"76",
          5581 => x"76",
          5582 => x"70",
          5583 => x"81",
          5584 => x"54",
          5585 => x"8e",
          5586 => x"52",
          5587 => x"81",
          5588 => x"81",
          5589 => x"74",
          5590 => x"53",
          5591 => x"83",
          5592 => x"78",
          5593 => x"8f",
          5594 => x"2e",
          5595 => x"c0",
          5596 => x"52",
          5597 => x"87",
          5598 => x"08",
          5599 => x"2e",
          5600 => x"84",
          5601 => x"38",
          5602 => x"87",
          5603 => x"15",
          5604 => x"70",
          5605 => x"52",
          5606 => x"ff",
          5607 => x"39",
          5608 => x"81",
          5609 => x"ff",
          5610 => x"57",
          5611 => x"90",
          5612 => x"80",
          5613 => x"71",
          5614 => x"78",
          5615 => x"38",
          5616 => x"80",
          5617 => x"80",
          5618 => x"81",
          5619 => x"72",
          5620 => x"0c",
          5621 => x"04",
          5622 => x"60",
          5623 => x"8c",
          5624 => x"33",
          5625 => x"5b",
          5626 => x"74",
          5627 => x"e1",
          5628 => x"c8",
          5629 => x"79",
          5630 => x"78",
          5631 => x"06",
          5632 => x"77",
          5633 => x"87",
          5634 => x"11",
          5635 => x"8c",
          5636 => x"92",
          5637 => x"59",
          5638 => x"85",
          5639 => x"98",
          5640 => x"7d",
          5641 => x"0c",
          5642 => x"08",
          5643 => x"70",
          5644 => x"53",
          5645 => x"2e",
          5646 => x"70",
          5647 => x"33",
          5648 => x"18",
          5649 => x"2a",
          5650 => x"51",
          5651 => x"2e",
          5652 => x"c0",
          5653 => x"52",
          5654 => x"87",
          5655 => x"08",
          5656 => x"2e",
          5657 => x"84",
          5658 => x"38",
          5659 => x"87",
          5660 => x"15",
          5661 => x"70",
          5662 => x"52",
          5663 => x"ff",
          5664 => x"39",
          5665 => x"81",
          5666 => x"80",
          5667 => x"52",
          5668 => x"90",
          5669 => x"80",
          5670 => x"71",
          5671 => x"7a",
          5672 => x"38",
          5673 => x"80",
          5674 => x"80",
          5675 => x"81",
          5676 => x"72",
          5677 => x"0c",
          5678 => x"04",
          5679 => x"7a",
          5680 => x"a3",
          5681 => x"88",
          5682 => x"33",
          5683 => x"56",
          5684 => x"3f",
          5685 => x"08",
          5686 => x"83",
          5687 => x"fe",
          5688 => x"87",
          5689 => x"0c",
          5690 => x"76",
          5691 => x"38",
          5692 => x"93",
          5693 => x"2b",
          5694 => x"8c",
          5695 => x"71",
          5696 => x"38",
          5697 => x"71",
          5698 => x"c6",
          5699 => x"39",
          5700 => x"81",
          5701 => x"06",
          5702 => x"71",
          5703 => x"38",
          5704 => x"8c",
          5705 => x"e8",
          5706 => x"98",
          5707 => x"71",
          5708 => x"73",
          5709 => x"92",
          5710 => x"72",
          5711 => x"06",
          5712 => x"f7",
          5713 => x"80",
          5714 => x"88",
          5715 => x"0c",
          5716 => x"80",
          5717 => x"56",
          5718 => x"56",
          5719 => x"82",
          5720 => x"88",
          5721 => x"fe",
          5722 => x"81",
          5723 => x"33",
          5724 => x"07",
          5725 => x"0c",
          5726 => x"3d",
          5727 => x"3d",
          5728 => x"11",
          5729 => x"33",
          5730 => x"71",
          5731 => x"81",
          5732 => x"72",
          5733 => x"75",
          5734 => x"82",
          5735 => x"52",
          5736 => x"54",
          5737 => x"0d",
          5738 => x"0d",
          5739 => x"05",
          5740 => x"52",
          5741 => x"70",
          5742 => x"34",
          5743 => x"51",
          5744 => x"83",
          5745 => x"ff",
          5746 => x"75",
          5747 => x"72",
          5748 => x"54",
          5749 => x"2a",
          5750 => x"70",
          5751 => x"34",
          5752 => x"51",
          5753 => x"81",
          5754 => x"70",
          5755 => x"70",
          5756 => x"3d",
          5757 => x"3d",
          5758 => x"77",
          5759 => x"70",
          5760 => x"38",
          5761 => x"05",
          5762 => x"70",
          5763 => x"34",
          5764 => x"eb",
          5765 => x"0d",
          5766 => x"0d",
          5767 => x"54",
          5768 => x"72",
          5769 => x"54",
          5770 => x"51",
          5771 => x"84",
          5772 => x"fc",
          5773 => x"77",
          5774 => x"53",
          5775 => x"05",
          5776 => x"70",
          5777 => x"33",
          5778 => x"ff",
          5779 => x"52",
          5780 => x"2e",
          5781 => x"80",
          5782 => x"71",
          5783 => x"0c",
          5784 => x"04",
          5785 => x"74",
          5786 => x"89",
          5787 => x"2e",
          5788 => x"11",
          5789 => x"52",
          5790 => x"70",
          5791 => x"c8",
          5792 => x"0d",
          5793 => x"82",
          5794 => x"04",
          5795 => x"77",
          5796 => x"70",
          5797 => x"33",
          5798 => x"55",
          5799 => x"ff",
          5800 => x"c8",
          5801 => x"72",
          5802 => x"38",
          5803 => x"72",
          5804 => x"b6",
          5805 => x"c8",
          5806 => x"ff",
          5807 => x"80",
          5808 => x"73",
          5809 => x"55",
          5810 => x"c8",
          5811 => x"0d",
          5812 => x"0d",
          5813 => x"0b",
          5814 => x"56",
          5815 => x"2e",
          5816 => x"81",
          5817 => x"08",
          5818 => x"70",
          5819 => x"33",
          5820 => x"e4",
          5821 => x"c8",
          5822 => x"09",
          5823 => x"38",
          5824 => x"08",
          5825 => x"b4",
          5826 => x"a8",
          5827 => x"a0",
          5828 => x"56",
          5829 => x"27",
          5830 => x"16",
          5831 => x"82",
          5832 => x"06",
          5833 => x"54",
          5834 => x"78",
          5835 => x"33",
          5836 => x"3f",
          5837 => x"5a",
          5838 => x"c8",
          5839 => x"0d",
          5840 => x"0d",
          5841 => x"56",
          5842 => x"b4",
          5843 => x"af",
          5844 => x"fe",
          5845 => x"d8",
          5846 => x"82",
          5847 => x"9f",
          5848 => x"74",
          5849 => x"52",
          5850 => x"51",
          5851 => x"82",
          5852 => x"80",
          5853 => x"ff",
          5854 => x"74",
          5855 => x"76",
          5856 => x"0c",
          5857 => x"04",
          5858 => x"7a",
          5859 => x"fe",
          5860 => x"d8",
          5861 => x"82",
          5862 => x"81",
          5863 => x"33",
          5864 => x"2e",
          5865 => x"80",
          5866 => x"17",
          5867 => x"81",
          5868 => x"06",
          5869 => x"84",
          5870 => x"d8",
          5871 => x"b8",
          5872 => x"56",
          5873 => x"82",
          5874 => x"84",
          5875 => x"fb",
          5876 => x"8b",
          5877 => x"52",
          5878 => x"eb",
          5879 => x"85",
          5880 => x"84",
          5881 => x"fb",
          5882 => x"17",
          5883 => x"a0",
          5884 => x"d3",
          5885 => x"08",
          5886 => x"17",
          5887 => x"3f",
          5888 => x"81",
          5889 => x"19",
          5890 => x"53",
          5891 => x"17",
          5892 => x"c4",
          5893 => x"18",
          5894 => x"80",
          5895 => x"33",
          5896 => x"3f",
          5897 => x"08",
          5898 => x"38",
          5899 => x"82",
          5900 => x"8a",
          5901 => x"fb",
          5902 => x"fe",
          5903 => x"08",
          5904 => x"56",
          5905 => x"74",
          5906 => x"38",
          5907 => x"75",
          5908 => x"16",
          5909 => x"53",
          5910 => x"c8",
          5911 => x"0d",
          5912 => x"0d",
          5913 => x"08",
          5914 => x"81",
          5915 => x"df",
          5916 => x"15",
          5917 => x"d7",
          5918 => x"33",
          5919 => x"82",
          5920 => x"38",
          5921 => x"89",
          5922 => x"2e",
          5923 => x"bf",
          5924 => x"2e",
          5925 => x"81",
          5926 => x"81",
          5927 => x"89",
          5928 => x"08",
          5929 => x"52",
          5930 => x"3f",
          5931 => x"08",
          5932 => x"74",
          5933 => x"14",
          5934 => x"81",
          5935 => x"2a",
          5936 => x"05",
          5937 => x"57",
          5938 => x"f5",
          5939 => x"c8",
          5940 => x"38",
          5941 => x"06",
          5942 => x"33",
          5943 => x"78",
          5944 => x"06",
          5945 => x"5c",
          5946 => x"53",
          5947 => x"38",
          5948 => x"06",
          5949 => x"39",
          5950 => x"a8",
          5951 => x"52",
          5952 => x"bd",
          5953 => x"c8",
          5954 => x"38",
          5955 => x"fe",
          5956 => x"b8",
          5957 => x"cf",
          5958 => x"c8",
          5959 => x"ff",
          5960 => x"39",
          5961 => x"a8",
          5962 => x"52",
          5963 => x"91",
          5964 => x"c8",
          5965 => x"76",
          5966 => x"fc",
          5967 => x"b8",
          5968 => x"ba",
          5969 => x"c8",
          5970 => x"06",
          5971 => x"81",
          5972 => x"d8",
          5973 => x"3d",
          5974 => x"3d",
          5975 => x"7e",
          5976 => x"82",
          5977 => x"27",
          5978 => x"76",
          5979 => x"27",
          5980 => x"75",
          5981 => x"79",
          5982 => x"38",
          5983 => x"89",
          5984 => x"2e",
          5985 => x"80",
          5986 => x"2e",
          5987 => x"81",
          5988 => x"81",
          5989 => x"89",
          5990 => x"08",
          5991 => x"52",
          5992 => x"3f",
          5993 => x"08",
          5994 => x"c8",
          5995 => x"38",
          5996 => x"06",
          5997 => x"81",
          5998 => x"06",
          5999 => x"77",
          6000 => x"2e",
          6001 => x"84",
          6002 => x"06",
          6003 => x"06",
          6004 => x"53",
          6005 => x"81",
          6006 => x"34",
          6007 => x"a8",
          6008 => x"52",
          6009 => x"d9",
          6010 => x"c8",
          6011 => x"d8",
          6012 => x"94",
          6013 => x"ff",
          6014 => x"05",
          6015 => x"54",
          6016 => x"38",
          6017 => x"74",
          6018 => x"06",
          6019 => x"07",
          6020 => x"74",
          6021 => x"39",
          6022 => x"a8",
          6023 => x"52",
          6024 => x"9d",
          6025 => x"c8",
          6026 => x"d8",
          6027 => x"d8",
          6028 => x"ff",
          6029 => x"76",
          6030 => x"06",
          6031 => x"05",
          6032 => x"3f",
          6033 => x"87",
          6034 => x"08",
          6035 => x"51",
          6036 => x"82",
          6037 => x"59",
          6038 => x"08",
          6039 => x"f0",
          6040 => x"82",
          6041 => x"06",
          6042 => x"05",
          6043 => x"54",
          6044 => x"3f",
          6045 => x"08",
          6046 => x"74",
          6047 => x"51",
          6048 => x"81",
          6049 => x"34",
          6050 => x"c8",
          6051 => x"0d",
          6052 => x"0d",
          6053 => x"72",
          6054 => x"56",
          6055 => x"27",
          6056 => x"9c",
          6057 => x"9d",
          6058 => x"2e",
          6059 => x"53",
          6060 => x"51",
          6061 => x"82",
          6062 => x"54",
          6063 => x"08",
          6064 => x"93",
          6065 => x"80",
          6066 => x"54",
          6067 => x"82",
          6068 => x"54",
          6069 => x"74",
          6070 => x"fb",
          6071 => x"d8",
          6072 => x"82",
          6073 => x"80",
          6074 => x"38",
          6075 => x"08",
          6076 => x"38",
          6077 => x"08",
          6078 => x"38",
          6079 => x"52",
          6080 => x"d6",
          6081 => x"c8",
          6082 => x"9c",
          6083 => x"11",
          6084 => x"57",
          6085 => x"74",
          6086 => x"81",
          6087 => x"0c",
          6088 => x"81",
          6089 => x"84",
          6090 => x"55",
          6091 => x"ff",
          6092 => x"54",
          6093 => x"c8",
          6094 => x"0d",
          6095 => x"0d",
          6096 => x"08",
          6097 => x"79",
          6098 => x"17",
          6099 => x"80",
          6100 => x"9c",
          6101 => x"26",
          6102 => x"58",
          6103 => x"52",
          6104 => x"fd",
          6105 => x"74",
          6106 => x"08",
          6107 => x"38",
          6108 => x"08",
          6109 => x"c8",
          6110 => x"82",
          6111 => x"17",
          6112 => x"c8",
          6113 => x"c7",
          6114 => x"94",
          6115 => x"56",
          6116 => x"2e",
          6117 => x"77",
          6118 => x"81",
          6119 => x"38",
          6120 => x"9c",
          6121 => x"26",
          6122 => x"56",
          6123 => x"51",
          6124 => x"80",
          6125 => x"c8",
          6126 => x"09",
          6127 => x"38",
          6128 => x"08",
          6129 => x"c8",
          6130 => x"30",
          6131 => x"80",
          6132 => x"07",
          6133 => x"08",
          6134 => x"55",
          6135 => x"ef",
          6136 => x"c8",
          6137 => x"95",
          6138 => x"08",
          6139 => x"27",
          6140 => x"9c",
          6141 => x"89",
          6142 => x"85",
          6143 => x"db",
          6144 => x"81",
          6145 => x"17",
          6146 => x"89",
          6147 => x"75",
          6148 => x"ac",
          6149 => x"7a",
          6150 => x"3f",
          6151 => x"08",
          6152 => x"38",
          6153 => x"d8",
          6154 => x"2e",
          6155 => x"86",
          6156 => x"c8",
          6157 => x"d8",
          6158 => x"70",
          6159 => x"07",
          6160 => x"7c",
          6161 => x"55",
          6162 => x"f8",
          6163 => x"2e",
          6164 => x"ff",
          6165 => x"55",
          6166 => x"ff",
          6167 => x"76",
          6168 => x"3f",
          6169 => x"08",
          6170 => x"08",
          6171 => x"d8",
          6172 => x"80",
          6173 => x"55",
          6174 => x"94",
          6175 => x"2e",
          6176 => x"53",
          6177 => x"51",
          6178 => x"82",
          6179 => x"55",
          6180 => x"75",
          6181 => x"9c",
          6182 => x"05",
          6183 => x"56",
          6184 => x"26",
          6185 => x"15",
          6186 => x"84",
          6187 => x"07",
          6188 => x"18",
          6189 => x"ff",
          6190 => x"2e",
          6191 => x"39",
          6192 => x"39",
          6193 => x"08",
          6194 => x"81",
          6195 => x"74",
          6196 => x"0c",
          6197 => x"04",
          6198 => x"7a",
          6199 => x"f3",
          6200 => x"d8",
          6201 => x"81",
          6202 => x"c8",
          6203 => x"38",
          6204 => x"51",
          6205 => x"82",
          6206 => x"82",
          6207 => x"b4",
          6208 => x"84",
          6209 => x"52",
          6210 => x"52",
          6211 => x"3f",
          6212 => x"39",
          6213 => x"8a",
          6214 => x"75",
          6215 => x"38",
          6216 => x"19",
          6217 => x"81",
          6218 => x"ed",
          6219 => x"d8",
          6220 => x"2e",
          6221 => x"15",
          6222 => x"70",
          6223 => x"07",
          6224 => x"53",
          6225 => x"75",
          6226 => x"0c",
          6227 => x"04",
          6228 => x"7a",
          6229 => x"58",
          6230 => x"f0",
          6231 => x"80",
          6232 => x"9f",
          6233 => x"80",
          6234 => x"90",
          6235 => x"17",
          6236 => x"aa",
          6237 => x"53",
          6238 => x"88",
          6239 => x"08",
          6240 => x"38",
          6241 => x"53",
          6242 => x"17",
          6243 => x"72",
          6244 => x"fe",
          6245 => x"08",
          6246 => x"80",
          6247 => x"16",
          6248 => x"2b",
          6249 => x"75",
          6250 => x"73",
          6251 => x"f5",
          6252 => x"d8",
          6253 => x"82",
          6254 => x"ff",
          6255 => x"81",
          6256 => x"c8",
          6257 => x"38",
          6258 => x"82",
          6259 => x"26",
          6260 => x"58",
          6261 => x"73",
          6262 => x"39",
          6263 => x"51",
          6264 => x"82",
          6265 => x"98",
          6266 => x"94",
          6267 => x"17",
          6268 => x"58",
          6269 => x"9a",
          6270 => x"81",
          6271 => x"74",
          6272 => x"98",
          6273 => x"83",
          6274 => x"b8",
          6275 => x"0c",
          6276 => x"82",
          6277 => x"8a",
          6278 => x"f8",
          6279 => x"70",
          6280 => x"08",
          6281 => x"57",
          6282 => x"0a",
          6283 => x"38",
          6284 => x"15",
          6285 => x"08",
          6286 => x"72",
          6287 => x"cb",
          6288 => x"ff",
          6289 => x"81",
          6290 => x"13",
          6291 => x"94",
          6292 => x"74",
          6293 => x"85",
          6294 => x"22",
          6295 => x"73",
          6296 => x"38",
          6297 => x"8a",
          6298 => x"05",
          6299 => x"06",
          6300 => x"8a",
          6301 => x"73",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"81",
          6305 => x"c8",
          6306 => x"ff",
          6307 => x"82",
          6308 => x"ff",
          6309 => x"38",
          6310 => x"82",
          6311 => x"26",
          6312 => x"7b",
          6313 => x"98",
          6314 => x"55",
          6315 => x"94",
          6316 => x"73",
          6317 => x"3f",
          6318 => x"08",
          6319 => x"82",
          6320 => x"80",
          6321 => x"38",
          6322 => x"d8",
          6323 => x"2e",
          6324 => x"55",
          6325 => x"08",
          6326 => x"38",
          6327 => x"08",
          6328 => x"fb",
          6329 => x"d8",
          6330 => x"38",
          6331 => x"0c",
          6332 => x"51",
          6333 => x"82",
          6334 => x"98",
          6335 => x"90",
          6336 => x"16",
          6337 => x"15",
          6338 => x"74",
          6339 => x"0c",
          6340 => x"04",
          6341 => x"7b",
          6342 => x"5b",
          6343 => x"52",
          6344 => x"ac",
          6345 => x"c8",
          6346 => x"d8",
          6347 => x"ec",
          6348 => x"c8",
          6349 => x"17",
          6350 => x"51",
          6351 => x"82",
          6352 => x"54",
          6353 => x"08",
          6354 => x"82",
          6355 => x"9c",
          6356 => x"33",
          6357 => x"72",
          6358 => x"09",
          6359 => x"38",
          6360 => x"d8",
          6361 => x"72",
          6362 => x"55",
          6363 => x"53",
          6364 => x"8e",
          6365 => x"56",
          6366 => x"09",
          6367 => x"38",
          6368 => x"d8",
          6369 => x"81",
          6370 => x"fd",
          6371 => x"d8",
          6372 => x"82",
          6373 => x"80",
          6374 => x"38",
          6375 => x"09",
          6376 => x"38",
          6377 => x"82",
          6378 => x"8b",
          6379 => x"fd",
          6380 => x"9a",
          6381 => x"eb",
          6382 => x"d8",
          6383 => x"ff",
          6384 => x"70",
          6385 => x"53",
          6386 => x"09",
          6387 => x"38",
          6388 => x"eb",
          6389 => x"d8",
          6390 => x"2b",
          6391 => x"72",
          6392 => x"0c",
          6393 => x"04",
          6394 => x"77",
          6395 => x"ff",
          6396 => x"9a",
          6397 => x"55",
          6398 => x"76",
          6399 => x"53",
          6400 => x"09",
          6401 => x"38",
          6402 => x"52",
          6403 => x"eb",
          6404 => x"3d",
          6405 => x"3d",
          6406 => x"80",
          6407 => x"70",
          6408 => x"81",
          6409 => x"74",
          6410 => x"56",
          6411 => x"70",
          6412 => x"ff",
          6413 => x"51",
          6414 => x"38",
          6415 => x"c8",
          6416 => x"0d",
          6417 => x"0d",
          6418 => x"59",
          6419 => x"5f",
          6420 => x"70",
          6421 => x"19",
          6422 => x"83",
          6423 => x"19",
          6424 => x"51",
          6425 => x"82",
          6426 => x"5b",
          6427 => x"08",
          6428 => x"9c",
          6429 => x"33",
          6430 => x"86",
          6431 => x"82",
          6432 => x"15",
          6433 => x"70",
          6434 => x"58",
          6435 => x"1a",
          6436 => x"c8",
          6437 => x"81",
          6438 => x"81",
          6439 => x"81",
          6440 => x"c8",
          6441 => x"ae",
          6442 => x"06",
          6443 => x"53",
          6444 => x"53",
          6445 => x"82",
          6446 => x"77",
          6447 => x"56",
          6448 => x"09",
          6449 => x"38",
          6450 => x"7f",
          6451 => x"81",
          6452 => x"ef",
          6453 => x"2e",
          6454 => x"81",
          6455 => x"86",
          6456 => x"06",
          6457 => x"80",
          6458 => x"8d",
          6459 => x"81",
          6460 => x"90",
          6461 => x"1d",
          6462 => x"5d",
          6463 => x"09",
          6464 => x"9c",
          6465 => x"33",
          6466 => x"2e",
          6467 => x"81",
          6468 => x"1e",
          6469 => x"52",
          6470 => x"3f",
          6471 => x"08",
          6472 => x"06",
          6473 => x"f8",
          6474 => x"70",
          6475 => x"8d",
          6476 => x"51",
          6477 => x"58",
          6478 => x"d0",
          6479 => x"05",
          6480 => x"3f",
          6481 => x"08",
          6482 => x"06",
          6483 => x"2e",
          6484 => x"81",
          6485 => x"c8",
          6486 => x"1a",
          6487 => x"75",
          6488 => x"14",
          6489 => x"75",
          6490 => x"2e",
          6491 => x"b0",
          6492 => x"57",
          6493 => x"c1",
          6494 => x"70",
          6495 => x"81",
          6496 => x"55",
          6497 => x"8e",
          6498 => x"fe",
          6499 => x"73",
          6500 => x"80",
          6501 => x"1c",
          6502 => x"06",
          6503 => x"39",
          6504 => x"72",
          6505 => x"7b",
          6506 => x"51",
          6507 => x"82",
          6508 => x"81",
          6509 => x"72",
          6510 => x"38",
          6511 => x"1a",
          6512 => x"80",
          6513 => x"f8",
          6514 => x"d8",
          6515 => x"82",
          6516 => x"89",
          6517 => x"08",
          6518 => x"86",
          6519 => x"98",
          6520 => x"82",
          6521 => x"90",
          6522 => x"f2",
          6523 => x"70",
          6524 => x"80",
          6525 => x"f6",
          6526 => x"d8",
          6527 => x"82",
          6528 => x"83",
          6529 => x"ff",
          6530 => x"ff",
          6531 => x"0c",
          6532 => x"52",
          6533 => x"a9",
          6534 => x"c8",
          6535 => x"d8",
          6536 => x"85",
          6537 => x"08",
          6538 => x"57",
          6539 => x"84",
          6540 => x"39",
          6541 => x"bf",
          6542 => x"ff",
          6543 => x"73",
          6544 => x"75",
          6545 => x"82",
          6546 => x"83",
          6547 => x"06",
          6548 => x"8f",
          6549 => x"73",
          6550 => x"74",
          6551 => x"81",
          6552 => x"38",
          6553 => x"70",
          6554 => x"81",
          6555 => x"55",
          6556 => x"38",
          6557 => x"70",
          6558 => x"54",
          6559 => x"92",
          6560 => x"33",
          6561 => x"06",
          6562 => x"08",
          6563 => x"58",
          6564 => x"7c",
          6565 => x"06",
          6566 => x"8d",
          6567 => x"7d",
          6568 => x"81",
          6569 => x"38",
          6570 => x"9a",
          6571 => x"e5",
          6572 => x"d8",
          6573 => x"ff",
          6574 => x"74",
          6575 => x"76",
          6576 => x"06",
          6577 => x"05",
          6578 => x"75",
          6579 => x"ca",
          6580 => x"77",
          6581 => x"8f",
          6582 => x"c8",
          6583 => x"ff",
          6584 => x"80",
          6585 => x"77",
          6586 => x"80",
          6587 => x"51",
          6588 => x"3f",
          6589 => x"08",
          6590 => x"70",
          6591 => x"81",
          6592 => x"80",
          6593 => x"74",
          6594 => x"08",
          6595 => x"06",
          6596 => x"75",
          6597 => x"75",
          6598 => x"2e",
          6599 => x"b3",
          6600 => x"5b",
          6601 => x"ff",
          6602 => x"33",
          6603 => x"70",
          6604 => x"55",
          6605 => x"2e",
          6606 => x"80",
          6607 => x"77",
          6608 => x"22",
          6609 => x"8b",
          6610 => x"70",
          6611 => x"51",
          6612 => x"81",
          6613 => x"5c",
          6614 => x"93",
          6615 => x"f9",
          6616 => x"d8",
          6617 => x"ff",
          6618 => x"7e",
          6619 => x"ab",
          6620 => x"06",
          6621 => x"38",
          6622 => x"19",
          6623 => x"08",
          6624 => x"3f",
          6625 => x"08",
          6626 => x"38",
          6627 => x"ff",
          6628 => x"0c",
          6629 => x"51",
          6630 => x"82",
          6631 => x"58",
          6632 => x"08",
          6633 => x"e8",
          6634 => x"d8",
          6635 => x"3d",
          6636 => x"3d",
          6637 => x"08",
          6638 => x"81",
          6639 => x"5d",
          6640 => x"73",
          6641 => x"73",
          6642 => x"70",
          6643 => x"5d",
          6644 => x"8d",
          6645 => x"70",
          6646 => x"22",
          6647 => x"f0",
          6648 => x"a0",
          6649 => x"92",
          6650 => x"5f",
          6651 => x"3f",
          6652 => x"05",
          6653 => x"54",
          6654 => x"82",
          6655 => x"c0",
          6656 => x"34",
          6657 => x"1c",
          6658 => x"58",
          6659 => x"52",
          6660 => x"e2",
          6661 => x"27",
          6662 => x"7a",
          6663 => x"70",
          6664 => x"06",
          6665 => x"80",
          6666 => x"74",
          6667 => x"06",
          6668 => x"55",
          6669 => x"81",
          6670 => x"07",
          6671 => x"71",
          6672 => x"81",
          6673 => x"56",
          6674 => x"2e",
          6675 => x"84",
          6676 => x"56",
          6677 => x"76",
          6678 => x"38",
          6679 => x"55",
          6680 => x"05",
          6681 => x"57",
          6682 => x"bf",
          6683 => x"74",
          6684 => x"87",
          6685 => x"76",
          6686 => x"ff",
          6687 => x"2a",
          6688 => x"74",
          6689 => x"3d",
          6690 => x"54",
          6691 => x"34",
          6692 => x"b5",
          6693 => x"54",
          6694 => x"ad",
          6695 => x"70",
          6696 => x"e3",
          6697 => x"d8",
          6698 => x"2e",
          6699 => x"17",
          6700 => x"2e",
          6701 => x"15",
          6702 => x"55",
          6703 => x"89",
          6704 => x"70",
          6705 => x"d0",
          6706 => x"77",
          6707 => x"54",
          6708 => x"16",
          6709 => x"56",
          6710 => x"8a",
          6711 => x"81",
          6712 => x"58",
          6713 => x"78",
          6714 => x"27",
          6715 => x"51",
          6716 => x"82",
          6717 => x"8b",
          6718 => x"5b",
          6719 => x"27",
          6720 => x"87",
          6721 => x"e4",
          6722 => x"38",
          6723 => x"08",
          6724 => x"c8",
          6725 => x"09",
          6726 => x"df",
          6727 => x"cb",
          6728 => x"1b",
          6729 => x"cb",
          6730 => x"81",
          6731 => x"06",
          6732 => x"81",
          6733 => x"2e",
          6734 => x"52",
          6735 => x"fe",
          6736 => x"82",
          6737 => x"19",
          6738 => x"79",
          6739 => x"3f",
          6740 => x"08",
          6741 => x"c8",
          6742 => x"38",
          6743 => x"78",
          6744 => x"d4",
          6745 => x"2b",
          6746 => x"71",
          6747 => x"79",
          6748 => x"3f",
          6749 => x"08",
          6750 => x"c8",
          6751 => x"38",
          6752 => x"f5",
          6753 => x"d8",
          6754 => x"ff",
          6755 => x"1a",
          6756 => x"51",
          6757 => x"82",
          6758 => x"57",
          6759 => x"08",
          6760 => x"8c",
          6761 => x"1b",
          6762 => x"ff",
          6763 => x"5b",
          6764 => x"34",
          6765 => x"17",
          6766 => x"c8",
          6767 => x"34",
          6768 => x"08",
          6769 => x"51",
          6770 => x"77",
          6771 => x"05",
          6772 => x"73",
          6773 => x"2e",
          6774 => x"10",
          6775 => x"81",
          6776 => x"54",
          6777 => x"ca",
          6778 => x"76",
          6779 => x"b9",
          6780 => x"38",
          6781 => x"54",
          6782 => x"8c",
          6783 => x"38",
          6784 => x"ff",
          6785 => x"74",
          6786 => x"22",
          6787 => x"86",
          6788 => x"c0",
          6789 => x"76",
          6790 => x"83",
          6791 => x"52",
          6792 => x"f7",
          6793 => x"c8",
          6794 => x"d8",
          6795 => x"c9",
          6796 => x"59",
          6797 => x"38",
          6798 => x"52",
          6799 => x"81",
          6800 => x"c8",
          6801 => x"d8",
          6802 => x"38",
          6803 => x"d8",
          6804 => x"9c",
          6805 => x"df",
          6806 => x"53",
          6807 => x"9c",
          6808 => x"df",
          6809 => x"1a",
          6810 => x"33",
          6811 => x"55",
          6812 => x"34",
          6813 => x"1d",
          6814 => x"74",
          6815 => x"0c",
          6816 => x"04",
          6817 => x"78",
          6818 => x"12",
          6819 => x"08",
          6820 => x"55",
          6821 => x"94",
          6822 => x"74",
          6823 => x"3f",
          6824 => x"08",
          6825 => x"c8",
          6826 => x"38",
          6827 => x"52",
          6828 => x"8d",
          6829 => x"c8",
          6830 => x"d8",
          6831 => x"38",
          6832 => x"53",
          6833 => x"81",
          6834 => x"34",
          6835 => x"77",
          6836 => x"82",
          6837 => x"52",
          6838 => x"bf",
          6839 => x"c8",
          6840 => x"d8",
          6841 => x"2e",
          6842 => x"84",
          6843 => x"06",
          6844 => x"54",
          6845 => x"c8",
          6846 => x"0d",
          6847 => x"0d",
          6848 => x"08",
          6849 => x"80",
          6850 => x"34",
          6851 => x"80",
          6852 => x"38",
          6853 => x"ff",
          6854 => x"38",
          6855 => x"7f",
          6856 => x"70",
          6857 => x"5b",
          6858 => x"77",
          6859 => x"38",
          6860 => x"70",
          6861 => x"5b",
          6862 => x"97",
          6863 => x"80",
          6864 => x"ff",
          6865 => x"53",
          6866 => x"26",
          6867 => x"5b",
          6868 => x"76",
          6869 => x"81",
          6870 => x"58",
          6871 => x"b5",
          6872 => x"2b",
          6873 => x"80",
          6874 => x"82",
          6875 => x"83",
          6876 => x"55",
          6877 => x"27",
          6878 => x"76",
          6879 => x"74",
          6880 => x"72",
          6881 => x"97",
          6882 => x"55",
          6883 => x"30",
          6884 => x"78",
          6885 => x"72",
          6886 => x"52",
          6887 => x"80",
          6888 => x"80",
          6889 => x"74",
          6890 => x"55",
          6891 => x"80",
          6892 => x"08",
          6893 => x"70",
          6894 => x"54",
          6895 => x"38",
          6896 => x"80",
          6897 => x"79",
          6898 => x"53",
          6899 => x"05",
          6900 => x"82",
          6901 => x"70",
          6902 => x"5a",
          6903 => x"08",
          6904 => x"81",
          6905 => x"53",
          6906 => x"b7",
          6907 => x"2e",
          6908 => x"84",
          6909 => x"55",
          6910 => x"70",
          6911 => x"07",
          6912 => x"54",
          6913 => x"26",
          6914 => x"80",
          6915 => x"ae",
          6916 => x"05",
          6917 => x"17",
          6918 => x"70",
          6919 => x"34",
          6920 => x"8a",
          6921 => x"b5",
          6922 => x"88",
          6923 => x"0b",
          6924 => x"96",
          6925 => x"72",
          6926 => x"76",
          6927 => x"0b",
          6928 => x"81",
          6929 => x"39",
          6930 => x"1a",
          6931 => x"57",
          6932 => x"80",
          6933 => x"18",
          6934 => x"56",
          6935 => x"bf",
          6936 => x"72",
          6937 => x"38",
          6938 => x"8c",
          6939 => x"53",
          6940 => x"87",
          6941 => x"2a",
          6942 => x"72",
          6943 => x"72",
          6944 => x"72",
          6945 => x"38",
          6946 => x"83",
          6947 => x"56",
          6948 => x"70",
          6949 => x"34",
          6950 => x"15",
          6951 => x"33",
          6952 => x"59",
          6953 => x"38",
          6954 => x"05",
          6955 => x"82",
          6956 => x"1c",
          6957 => x"33",
          6958 => x"85",
          6959 => x"19",
          6960 => x"08",
          6961 => x"33",
          6962 => x"9c",
          6963 => x"11",
          6964 => x"aa",
          6965 => x"c8",
          6966 => x"96",
          6967 => x"87",
          6968 => x"c8",
          6969 => x"23",
          6970 => x"d8",
          6971 => x"d8",
          6972 => x"19",
          6973 => x"0d",
          6974 => x"0d",
          6975 => x"41",
          6976 => x"70",
          6977 => x"55",
          6978 => x"83",
          6979 => x"73",
          6980 => x"92",
          6981 => x"2e",
          6982 => x"98",
          6983 => x"1f",
          6984 => x"81",
          6985 => x"64",
          6986 => x"56",
          6987 => x"2e",
          6988 => x"83",
          6989 => x"73",
          6990 => x"70",
          6991 => x"25",
          6992 => x"51",
          6993 => x"38",
          6994 => x"0c",
          6995 => x"51",
          6996 => x"26",
          6997 => x"80",
          6998 => x"34",
          6999 => x"51",
          7000 => x"82",
          7001 => x"56",
          7002 => x"63",
          7003 => x"8c",
          7004 => x"54",
          7005 => x"3d",
          7006 => x"da",
          7007 => x"d8",
          7008 => x"2e",
          7009 => x"83",
          7010 => x"82",
          7011 => x"27",
          7012 => x"10",
          7013 => x"c8",
          7014 => x"55",
          7015 => x"23",
          7016 => x"82",
          7017 => x"83",
          7018 => x"70",
          7019 => x"30",
          7020 => x"71",
          7021 => x"51",
          7022 => x"73",
          7023 => x"80",
          7024 => x"38",
          7025 => x"26",
          7026 => x"52",
          7027 => x"51",
          7028 => x"82",
          7029 => x"81",
          7030 => x"81",
          7031 => x"d7",
          7032 => x"1a",
          7033 => x"23",
          7034 => x"ff",
          7035 => x"15",
          7036 => x"70",
          7037 => x"57",
          7038 => x"09",
          7039 => x"38",
          7040 => x"80",
          7041 => x"30",
          7042 => x"79",
          7043 => x"54",
          7044 => x"74",
          7045 => x"27",
          7046 => x"78",
          7047 => x"81",
          7048 => x"79",
          7049 => x"ae",
          7050 => x"80",
          7051 => x"82",
          7052 => x"06",
          7053 => x"82",
          7054 => x"73",
          7055 => x"81",
          7056 => x"38",
          7057 => x"73",
          7058 => x"81",
          7059 => x"78",
          7060 => x"80",
          7061 => x"0b",
          7062 => x"58",
          7063 => x"78",
          7064 => x"a0",
          7065 => x"70",
          7066 => x"34",
          7067 => x"8a",
          7068 => x"38",
          7069 => x"54",
          7070 => x"34",
          7071 => x"78",
          7072 => x"38",
          7073 => x"fe",
          7074 => x"22",
          7075 => x"72",
          7076 => x"30",
          7077 => x"51",
          7078 => x"56",
          7079 => x"2e",
          7080 => x"87",
          7081 => x"59",
          7082 => x"78",
          7083 => x"55",
          7084 => x"23",
          7085 => x"86",
          7086 => x"39",
          7087 => x"57",
          7088 => x"80",
          7089 => x"83",
          7090 => x"56",
          7091 => x"a0",
          7092 => x"06",
          7093 => x"1d",
          7094 => x"70",
          7095 => x"5d",
          7096 => x"f2",
          7097 => x"38",
          7098 => x"ff",
          7099 => x"ae",
          7100 => x"06",
          7101 => x"83",
          7102 => x"80",
          7103 => x"79",
          7104 => x"70",
          7105 => x"73",
          7106 => x"38",
          7107 => x"fe",
          7108 => x"19",
          7109 => x"2e",
          7110 => x"15",
          7111 => x"55",
          7112 => x"09",
          7113 => x"38",
          7114 => x"52",
          7115 => x"d5",
          7116 => x"70",
          7117 => x"5f",
          7118 => x"70",
          7119 => x"5f",
          7120 => x"80",
          7121 => x"38",
          7122 => x"96",
          7123 => x"32",
          7124 => x"80",
          7125 => x"54",
          7126 => x"8c",
          7127 => x"2e",
          7128 => x"83",
          7129 => x"39",
          7130 => x"5b",
          7131 => x"83",
          7132 => x"7c",
          7133 => x"30",
          7134 => x"80",
          7135 => x"07",
          7136 => x"55",
          7137 => x"a6",
          7138 => x"2e",
          7139 => x"7c",
          7140 => x"38",
          7141 => x"57",
          7142 => x"81",
          7143 => x"5d",
          7144 => x"7c",
          7145 => x"fc",
          7146 => x"ff",
          7147 => x"ff",
          7148 => x"38",
          7149 => x"57",
          7150 => x"75",
          7151 => x"c2",
          7152 => x"c8",
          7153 => x"ff",
          7154 => x"2a",
          7155 => x"51",
          7156 => x"80",
          7157 => x"75",
          7158 => x"82",
          7159 => x"33",
          7160 => x"ff",
          7161 => x"38",
          7162 => x"73",
          7163 => x"38",
          7164 => x"7f",
          7165 => x"c0",
          7166 => x"a0",
          7167 => x"2a",
          7168 => x"75",
          7169 => x"58",
          7170 => x"75",
          7171 => x"38",
          7172 => x"c9",
          7173 => x"cc",
          7174 => x"c8",
          7175 => x"8a",
          7176 => x"77",
          7177 => x"56",
          7178 => x"bf",
          7179 => x"99",
          7180 => x"7b",
          7181 => x"ff",
          7182 => x"73",
          7183 => x"38",
          7184 => x"e0",
          7185 => x"ff",
          7186 => x"55",
          7187 => x"a0",
          7188 => x"74",
          7189 => x"58",
          7190 => x"a0",
          7191 => x"73",
          7192 => x"09",
          7193 => x"38",
          7194 => x"1f",
          7195 => x"2e",
          7196 => x"88",
          7197 => x"2b",
          7198 => x"5c",
          7199 => x"54",
          7200 => x"8d",
          7201 => x"06",
          7202 => x"2e",
          7203 => x"85",
          7204 => x"07",
          7205 => x"2a",
          7206 => x"51",
          7207 => x"38",
          7208 => x"54",
          7209 => x"85",
          7210 => x"07",
          7211 => x"2a",
          7212 => x"51",
          7213 => x"2e",
          7214 => x"88",
          7215 => x"ab",
          7216 => x"51",
          7217 => x"82",
          7218 => x"ab",
          7219 => x"56",
          7220 => x"08",
          7221 => x"38",
          7222 => x"08",
          7223 => x"81",
          7224 => x"38",
          7225 => x"70",
          7226 => x"82",
          7227 => x"54",
          7228 => x"96",
          7229 => x"06",
          7230 => x"2e",
          7231 => x"ff",
          7232 => x"1f",
          7233 => x"80",
          7234 => x"81",
          7235 => x"bb",
          7236 => x"b7",
          7237 => x"2a",
          7238 => x"51",
          7239 => x"38",
          7240 => x"70",
          7241 => x"81",
          7242 => x"55",
          7243 => x"e1",
          7244 => x"08",
          7245 => x"60",
          7246 => x"52",
          7247 => x"ef",
          7248 => x"c8",
          7249 => x"0c",
          7250 => x"75",
          7251 => x"0c",
          7252 => x"04",
          7253 => x"7c",
          7254 => x"08",
          7255 => x"55",
          7256 => x"59",
          7257 => x"81",
          7258 => x"70",
          7259 => x"33",
          7260 => x"52",
          7261 => x"2e",
          7262 => x"ee",
          7263 => x"2e",
          7264 => x"81",
          7265 => x"33",
          7266 => x"81",
          7267 => x"52",
          7268 => x"26",
          7269 => x"14",
          7270 => x"06",
          7271 => x"52",
          7272 => x"80",
          7273 => x"0b",
          7274 => x"59",
          7275 => x"7a",
          7276 => x"70",
          7277 => x"33",
          7278 => x"05",
          7279 => x"9f",
          7280 => x"53",
          7281 => x"89",
          7282 => x"70",
          7283 => x"54",
          7284 => x"12",
          7285 => x"26",
          7286 => x"12",
          7287 => x"06",
          7288 => x"30",
          7289 => x"51",
          7290 => x"2e",
          7291 => x"85",
          7292 => x"be",
          7293 => x"74",
          7294 => x"30",
          7295 => x"9f",
          7296 => x"2a",
          7297 => x"54",
          7298 => x"2e",
          7299 => x"15",
          7300 => x"55",
          7301 => x"ff",
          7302 => x"39",
          7303 => x"86",
          7304 => x"7c",
          7305 => x"51",
          7306 => x"f0",
          7307 => x"70",
          7308 => x"0c",
          7309 => x"04",
          7310 => x"78",
          7311 => x"83",
          7312 => x"0b",
          7313 => x"79",
          7314 => x"d1",
          7315 => x"55",
          7316 => x"08",
          7317 => x"84",
          7318 => x"ce",
          7319 => x"d8",
          7320 => x"ff",
          7321 => x"83",
          7322 => x"d4",
          7323 => x"81",
          7324 => x"38",
          7325 => x"17",
          7326 => x"74",
          7327 => x"09",
          7328 => x"38",
          7329 => x"81",
          7330 => x"30",
          7331 => x"79",
          7332 => x"54",
          7333 => x"74",
          7334 => x"09",
          7335 => x"38",
          7336 => x"ca",
          7337 => x"ee",
          7338 => x"87",
          7339 => x"c8",
          7340 => x"d8",
          7341 => x"2e",
          7342 => x"53",
          7343 => x"52",
          7344 => x"51",
          7345 => x"82",
          7346 => x"55",
          7347 => x"08",
          7348 => x"38",
          7349 => x"82",
          7350 => x"88",
          7351 => x"f2",
          7352 => x"02",
          7353 => x"cb",
          7354 => x"55",
          7355 => x"60",
          7356 => x"3f",
          7357 => x"08",
          7358 => x"80",
          7359 => x"c8",
          7360 => x"84",
          7361 => x"c8",
          7362 => x"82",
          7363 => x"70",
          7364 => x"8c",
          7365 => x"2e",
          7366 => x"73",
          7367 => x"81",
          7368 => x"33",
          7369 => x"80",
          7370 => x"81",
          7371 => x"c6",
          7372 => x"d8",
          7373 => x"ff",
          7374 => x"06",
          7375 => x"98",
          7376 => x"2e",
          7377 => x"74",
          7378 => x"81",
          7379 => x"8a",
          7380 => x"b4",
          7381 => x"39",
          7382 => x"77",
          7383 => x"81",
          7384 => x"33",
          7385 => x"3f",
          7386 => x"08",
          7387 => x"70",
          7388 => x"55",
          7389 => x"86",
          7390 => x"80",
          7391 => x"74",
          7392 => x"81",
          7393 => x"8a",
          7394 => x"fc",
          7395 => x"53",
          7396 => x"fd",
          7397 => x"d8",
          7398 => x"ff",
          7399 => x"82",
          7400 => x"06",
          7401 => x"8c",
          7402 => x"58",
          7403 => x"fa",
          7404 => x"58",
          7405 => x"2e",
          7406 => x"fe",
          7407 => x"be",
          7408 => x"c8",
          7409 => x"78",
          7410 => x"5a",
          7411 => x"90",
          7412 => x"75",
          7413 => x"38",
          7414 => x"3d",
          7415 => x"70",
          7416 => x"08",
          7417 => x"7a",
          7418 => x"38",
          7419 => x"51",
          7420 => x"82",
          7421 => x"81",
          7422 => x"81",
          7423 => x"38",
          7424 => x"83",
          7425 => x"38",
          7426 => x"84",
          7427 => x"38",
          7428 => x"81",
          7429 => x"38",
          7430 => x"51",
          7431 => x"82",
          7432 => x"83",
          7433 => x"53",
          7434 => x"2e",
          7435 => x"84",
          7436 => x"ce",
          7437 => x"af",
          7438 => x"c8",
          7439 => x"ff",
          7440 => x"8d",
          7441 => x"14",
          7442 => x"3f",
          7443 => x"08",
          7444 => x"15",
          7445 => x"14",
          7446 => x"34",
          7447 => x"33",
          7448 => x"81",
          7449 => x"54",
          7450 => x"72",
          7451 => x"98",
          7452 => x"ff",
          7453 => x"29",
          7454 => x"33",
          7455 => x"72",
          7456 => x"72",
          7457 => x"38",
          7458 => x"06",
          7459 => x"2e",
          7460 => x"56",
          7461 => x"80",
          7462 => x"c9",
          7463 => x"d8",
          7464 => x"82",
          7465 => x"88",
          7466 => x"8f",
          7467 => x"56",
          7468 => x"38",
          7469 => x"51",
          7470 => x"82",
          7471 => x"83",
          7472 => x"55",
          7473 => x"80",
          7474 => x"c9",
          7475 => x"d8",
          7476 => x"80",
          7477 => x"c9",
          7478 => x"d8",
          7479 => x"ff",
          7480 => x"8d",
          7481 => x"2e",
          7482 => x"88",
          7483 => x"14",
          7484 => x"05",
          7485 => x"75",
          7486 => x"38",
          7487 => x"52",
          7488 => x"51",
          7489 => x"3f",
          7490 => x"08",
          7491 => x"c8",
          7492 => x"82",
          7493 => x"d8",
          7494 => x"ff",
          7495 => x"26",
          7496 => x"57",
          7497 => x"f5",
          7498 => x"82",
          7499 => x"f5",
          7500 => x"81",
          7501 => x"8d",
          7502 => x"2e",
          7503 => x"82",
          7504 => x"16",
          7505 => x"16",
          7506 => x"70",
          7507 => x"7a",
          7508 => x"0c",
          7509 => x"83",
          7510 => x"06",
          7511 => x"e2",
          7512 => x"83",
          7513 => x"c8",
          7514 => x"ff",
          7515 => x"56",
          7516 => x"38",
          7517 => x"38",
          7518 => x"51",
          7519 => x"82",
          7520 => x"ac",
          7521 => x"82",
          7522 => x"39",
          7523 => x"80",
          7524 => x"38",
          7525 => x"15",
          7526 => x"53",
          7527 => x"8d",
          7528 => x"15",
          7529 => x"76",
          7530 => x"51",
          7531 => x"13",
          7532 => x"8d",
          7533 => x"15",
          7534 => x"cc",
          7535 => x"94",
          7536 => x"0b",
          7537 => x"ff",
          7538 => x"15",
          7539 => x"2e",
          7540 => x"81",
          7541 => x"e8",
          7542 => x"8b",
          7543 => x"c8",
          7544 => x"ff",
          7545 => x"81",
          7546 => x"06",
          7547 => x"81",
          7548 => x"51",
          7549 => x"82",
          7550 => x"80",
          7551 => x"d8",
          7552 => x"15",
          7553 => x"14",
          7554 => x"3f",
          7555 => x"08",
          7556 => x"06",
          7557 => x"d4",
          7558 => x"81",
          7559 => x"38",
          7560 => x"c6",
          7561 => x"d8",
          7562 => x"8b",
          7563 => x"2e",
          7564 => x"b3",
          7565 => x"14",
          7566 => x"3f",
          7567 => x"08",
          7568 => x"e4",
          7569 => x"81",
          7570 => x"84",
          7571 => x"c6",
          7572 => x"d8",
          7573 => x"15",
          7574 => x"14",
          7575 => x"3f",
          7576 => x"08",
          7577 => x"76",
          7578 => x"f0",
          7579 => x"05",
          7580 => x"f0",
          7581 => x"86",
          7582 => x"f0",
          7583 => x"15",
          7584 => x"98",
          7585 => x"56",
          7586 => x"c8",
          7587 => x"0d",
          7588 => x"0d",
          7589 => x"55",
          7590 => x"ba",
          7591 => x"53",
          7592 => x"b2",
          7593 => x"52",
          7594 => x"aa",
          7595 => x"22",
          7596 => x"57",
          7597 => x"2e",
          7598 => x"9a",
          7599 => x"33",
          7600 => x"8d",
          7601 => x"c8",
          7602 => x"52",
          7603 => x"71",
          7604 => x"55",
          7605 => x"53",
          7606 => x"0c",
          7607 => x"d8",
          7608 => x"3d",
          7609 => x"3d",
          7610 => x"05",
          7611 => x"89",
          7612 => x"52",
          7613 => x"3f",
          7614 => x"0b",
          7615 => x"08",
          7616 => x"82",
          7617 => x"84",
          7618 => x"90",
          7619 => x"55",
          7620 => x"2e",
          7621 => x"74",
          7622 => x"73",
          7623 => x"38",
          7624 => x"78",
          7625 => x"54",
          7626 => x"92",
          7627 => x"89",
          7628 => x"84",
          7629 => x"a7",
          7630 => x"c8",
          7631 => x"82",
          7632 => x"88",
          7633 => x"ea",
          7634 => x"02",
          7635 => x"eb",
          7636 => x"59",
          7637 => x"80",
          7638 => x"38",
          7639 => x"70",
          7640 => x"cc",
          7641 => x"3d",
          7642 => x"58",
          7643 => x"82",
          7644 => x"55",
          7645 => x"08",
          7646 => x"7a",
          7647 => x"8c",
          7648 => x"56",
          7649 => x"82",
          7650 => x"55",
          7651 => x"08",
          7652 => x"80",
          7653 => x"70",
          7654 => x"57",
          7655 => x"83",
          7656 => x"77",
          7657 => x"73",
          7658 => x"ab",
          7659 => x"2e",
          7660 => x"84",
          7661 => x"06",
          7662 => x"51",
          7663 => x"82",
          7664 => x"55",
          7665 => x"b2",
          7666 => x"06",
          7667 => x"b8",
          7668 => x"2a",
          7669 => x"51",
          7670 => x"2e",
          7671 => x"55",
          7672 => x"77",
          7673 => x"74",
          7674 => x"77",
          7675 => x"81",
          7676 => x"73",
          7677 => x"af",
          7678 => x"7a",
          7679 => x"3f",
          7680 => x"08",
          7681 => x"b2",
          7682 => x"8e",
          7683 => x"b7",
          7684 => x"a0",
          7685 => x"34",
          7686 => x"52",
          7687 => x"c8",
          7688 => x"62",
          7689 => x"c3",
          7690 => x"54",
          7691 => x"15",
          7692 => x"2e",
          7693 => x"7a",
          7694 => x"51",
          7695 => x"75",
          7696 => x"d0",
          7697 => x"c9",
          7698 => x"c8",
          7699 => x"d8",
          7700 => x"ca",
          7701 => x"74",
          7702 => x"02",
          7703 => x"70",
          7704 => x"81",
          7705 => x"56",
          7706 => x"86",
          7707 => x"82",
          7708 => x"81",
          7709 => x"06",
          7710 => x"80",
          7711 => x"75",
          7712 => x"73",
          7713 => x"38",
          7714 => x"92",
          7715 => x"7a",
          7716 => x"3f",
          7717 => x"08",
          7718 => x"90",
          7719 => x"55",
          7720 => x"08",
          7721 => x"77",
          7722 => x"81",
          7723 => x"73",
          7724 => x"38",
          7725 => x"07",
          7726 => x"11",
          7727 => x"0c",
          7728 => x"0c",
          7729 => x"52",
          7730 => x"3f",
          7731 => x"08",
          7732 => x"08",
          7733 => x"63",
          7734 => x"5a",
          7735 => x"82",
          7736 => x"82",
          7737 => x"8c",
          7738 => x"7a",
          7739 => x"17",
          7740 => x"23",
          7741 => x"34",
          7742 => x"1a",
          7743 => x"9c",
          7744 => x"0b",
          7745 => x"77",
          7746 => x"81",
          7747 => x"73",
          7748 => x"8d",
          7749 => x"c8",
          7750 => x"81",
          7751 => x"d8",
          7752 => x"1a",
          7753 => x"22",
          7754 => x"7b",
          7755 => x"a8",
          7756 => x"78",
          7757 => x"3f",
          7758 => x"08",
          7759 => x"c8",
          7760 => x"83",
          7761 => x"82",
          7762 => x"ff",
          7763 => x"06",
          7764 => x"55",
          7765 => x"56",
          7766 => x"76",
          7767 => x"51",
          7768 => x"27",
          7769 => x"70",
          7770 => x"5a",
          7771 => x"76",
          7772 => x"74",
          7773 => x"83",
          7774 => x"73",
          7775 => x"38",
          7776 => x"51",
          7777 => x"82",
          7778 => x"85",
          7779 => x"8e",
          7780 => x"2a",
          7781 => x"08",
          7782 => x"0c",
          7783 => x"79",
          7784 => x"73",
          7785 => x"0c",
          7786 => x"04",
          7787 => x"60",
          7788 => x"40",
          7789 => x"80",
          7790 => x"3d",
          7791 => x"78",
          7792 => x"3f",
          7793 => x"08",
          7794 => x"c8",
          7795 => x"91",
          7796 => x"74",
          7797 => x"38",
          7798 => x"c7",
          7799 => x"33",
          7800 => x"87",
          7801 => x"2e",
          7802 => x"95",
          7803 => x"91",
          7804 => x"56",
          7805 => x"81",
          7806 => x"34",
          7807 => x"a3",
          7808 => x"08",
          7809 => x"31",
          7810 => x"27",
          7811 => x"5c",
          7812 => x"82",
          7813 => x"19",
          7814 => x"ff",
          7815 => x"74",
          7816 => x"7e",
          7817 => x"ff",
          7818 => x"2a",
          7819 => x"79",
          7820 => x"87",
          7821 => x"08",
          7822 => x"98",
          7823 => x"78",
          7824 => x"3f",
          7825 => x"08",
          7826 => x"27",
          7827 => x"74",
          7828 => x"a3",
          7829 => x"1a",
          7830 => x"08",
          7831 => x"c3",
          7832 => x"d8",
          7833 => x"2e",
          7834 => x"82",
          7835 => x"1a",
          7836 => x"59",
          7837 => x"2e",
          7838 => x"77",
          7839 => x"11",
          7840 => x"55",
          7841 => x"85",
          7842 => x"31",
          7843 => x"76",
          7844 => x"81",
          7845 => x"ff",
          7846 => x"82",
          7847 => x"fe",
          7848 => x"83",
          7849 => x"56",
          7850 => x"a0",
          7851 => x"08",
          7852 => x"74",
          7853 => x"38",
          7854 => x"b8",
          7855 => x"16",
          7856 => x"89",
          7857 => x"51",
          7858 => x"3f",
          7859 => x"56",
          7860 => x"9c",
          7861 => x"19",
          7862 => x"06",
          7863 => x"31",
          7864 => x"76",
          7865 => x"7b",
          7866 => x"08",
          7867 => x"c0",
          7868 => x"d8",
          7869 => x"ff",
          7870 => x"94",
          7871 => x"ff",
          7872 => x"05",
          7873 => x"ff",
          7874 => x"7b",
          7875 => x"08",
          7876 => x"76",
          7877 => x"08",
          7878 => x"0c",
          7879 => x"f0",
          7880 => x"75",
          7881 => x"0c",
          7882 => x"04",
          7883 => x"60",
          7884 => x"40",
          7885 => x"80",
          7886 => x"3d",
          7887 => x"77",
          7888 => x"3f",
          7889 => x"08",
          7890 => x"c8",
          7891 => x"91",
          7892 => x"74",
          7893 => x"38",
          7894 => x"be",
          7895 => x"33",
          7896 => x"70",
          7897 => x"56",
          7898 => x"74",
          7899 => x"aa",
          7900 => x"82",
          7901 => x"34",
          7902 => x"9e",
          7903 => x"91",
          7904 => x"56",
          7905 => x"94",
          7906 => x"11",
          7907 => x"76",
          7908 => x"75",
          7909 => x"80",
          7910 => x"38",
          7911 => x"70",
          7912 => x"56",
          7913 => x"81",
          7914 => x"11",
          7915 => x"77",
          7916 => x"5c",
          7917 => x"38",
          7918 => x"88",
          7919 => x"74",
          7920 => x"52",
          7921 => x"18",
          7922 => x"51",
          7923 => x"82",
          7924 => x"55",
          7925 => x"08",
          7926 => x"b1",
          7927 => x"2e",
          7928 => x"74",
          7929 => x"95",
          7930 => x"19",
          7931 => x"08",
          7932 => x"88",
          7933 => x"55",
          7934 => x"9c",
          7935 => x"09",
          7936 => x"38",
          7937 => x"bd",
          7938 => x"d8",
          7939 => x"ed",
          7940 => x"08",
          7941 => x"c0",
          7942 => x"d8",
          7943 => x"2e",
          7944 => x"82",
          7945 => x"1b",
          7946 => x"5a",
          7947 => x"2e",
          7948 => x"78",
          7949 => x"11",
          7950 => x"55",
          7951 => x"85",
          7952 => x"31",
          7953 => x"76",
          7954 => x"81",
          7955 => x"ff",
          7956 => x"82",
          7957 => x"fe",
          7958 => x"b4",
          7959 => x"31",
          7960 => x"79",
          7961 => x"84",
          7962 => x"16",
          7963 => x"89",
          7964 => x"52",
          7965 => x"ff",
          7966 => x"7e",
          7967 => x"83",
          7968 => x"89",
          7969 => x"de",
          7970 => x"08",
          7971 => x"26",
          7972 => x"51",
          7973 => x"3f",
          7974 => x"08",
          7975 => x"7e",
          7976 => x"0c",
          7977 => x"19",
          7978 => x"08",
          7979 => x"84",
          7980 => x"57",
          7981 => x"27",
          7982 => x"56",
          7983 => x"52",
          7984 => x"bc",
          7985 => x"d8",
          7986 => x"b1",
          7987 => x"7c",
          7988 => x"08",
          7989 => x"1f",
          7990 => x"ff",
          7991 => x"7e",
          7992 => x"83",
          7993 => x"76",
          7994 => x"17",
          7995 => x"1e",
          7996 => x"18",
          7997 => x"0c",
          7998 => x"58",
          7999 => x"74",
          8000 => x"38",
          8001 => x"8c",
          8002 => x"8a",
          8003 => x"33",
          8004 => x"55",
          8005 => x"34",
          8006 => x"82",
          8007 => x"90",
          8008 => x"f8",
          8009 => x"8b",
          8010 => x"53",
          8011 => x"f2",
          8012 => x"d8",
          8013 => x"82",
          8014 => x"81",
          8015 => x"16",
          8016 => x"2a",
          8017 => x"51",
          8018 => x"80",
          8019 => x"38",
          8020 => x"52",
          8021 => x"bb",
          8022 => x"d8",
          8023 => x"82",
          8024 => x"80",
          8025 => x"16",
          8026 => x"33",
          8027 => x"55",
          8028 => x"34",
          8029 => x"53",
          8030 => x"08",
          8031 => x"3f",
          8032 => x"52",
          8033 => x"ff",
          8034 => x"82",
          8035 => x"52",
          8036 => x"ff",
          8037 => x"76",
          8038 => x"51",
          8039 => x"3f",
          8040 => x"0b",
          8041 => x"78",
          8042 => x"dc",
          8043 => x"c8",
          8044 => x"33",
          8045 => x"55",
          8046 => x"17",
          8047 => x"d8",
          8048 => x"3d",
          8049 => x"3d",
          8050 => x"52",
          8051 => x"3f",
          8052 => x"08",
          8053 => x"c8",
          8054 => x"86",
          8055 => x"52",
          8056 => x"ad",
          8057 => x"c8",
          8058 => x"d8",
          8059 => x"38",
          8060 => x"08",
          8061 => x"82",
          8062 => x"86",
          8063 => x"ff",
          8064 => x"3d",
          8065 => x"3f",
          8066 => x"0b",
          8067 => x"08",
          8068 => x"82",
          8069 => x"82",
          8070 => x"80",
          8071 => x"d8",
          8072 => x"3d",
          8073 => x"3d",
          8074 => x"94",
          8075 => x"52",
          8076 => x"e9",
          8077 => x"d8",
          8078 => x"82",
          8079 => x"80",
          8080 => x"58",
          8081 => x"3d",
          8082 => x"dd",
          8083 => x"d8",
          8084 => x"82",
          8085 => x"bc",
          8086 => x"c7",
          8087 => x"98",
          8088 => x"73",
          8089 => x"38",
          8090 => x"12",
          8091 => x"39",
          8092 => x"33",
          8093 => x"70",
          8094 => x"55",
          8095 => x"2e",
          8096 => x"7f",
          8097 => x"54",
          8098 => x"82",
          8099 => x"98",
          8100 => x"39",
          8101 => x"08",
          8102 => x"81",
          8103 => x"85",
          8104 => x"d8",
          8105 => x"3d",
          8106 => x"a3",
          8107 => x"e1",
          8108 => x"e1",
          8109 => x"5b",
          8110 => x"80",
          8111 => x"3d",
          8112 => x"52",
          8113 => x"51",
          8114 => x"82",
          8115 => x"57",
          8116 => x"08",
          8117 => x"7b",
          8118 => x"0c",
          8119 => x"11",
          8120 => x"3d",
          8121 => x"80",
          8122 => x"54",
          8123 => x"82",
          8124 => x"52",
          8125 => x"70",
          8126 => x"d4",
          8127 => x"c8",
          8128 => x"d8",
          8129 => x"ef",
          8130 => x"3d",
          8131 => x"51",
          8132 => x"3f",
          8133 => x"08",
          8134 => x"c8",
          8135 => x"38",
          8136 => x"08",
          8137 => x"c9",
          8138 => x"d8",
          8139 => x"d6",
          8140 => x"52",
          8141 => x"98",
          8142 => x"c8",
          8143 => x"d8",
          8144 => x"b3",
          8145 => x"74",
          8146 => x"3f",
          8147 => x"08",
          8148 => x"c8",
          8149 => x"80",
          8150 => x"52",
          8151 => x"cf",
          8152 => x"d8",
          8153 => x"a6",
          8154 => x"74",
          8155 => x"3f",
          8156 => x"08",
          8157 => x"c8",
          8158 => x"c9",
          8159 => x"2e",
          8160 => x"86",
          8161 => x"81",
          8162 => x"81",
          8163 => x"df",
          8164 => x"05",
          8165 => x"d6",
          8166 => x"93",
          8167 => x"82",
          8168 => x"56",
          8169 => x"80",
          8170 => x"02",
          8171 => x"55",
          8172 => x"16",
          8173 => x"56",
          8174 => x"38",
          8175 => x"73",
          8176 => x"99",
          8177 => x"2e",
          8178 => x"16",
          8179 => x"ff",
          8180 => x"3d",
          8181 => x"18",
          8182 => x"58",
          8183 => x"33",
          8184 => x"eb",
          8185 => x"80",
          8186 => x"11",
          8187 => x"74",
          8188 => x"39",
          8189 => x"09",
          8190 => x"38",
          8191 => x"e1",
          8192 => x"55",
          8193 => x"34",
          8194 => x"f0",
          8195 => x"84",
          8196 => x"c0",
          8197 => x"70",
          8198 => x"56",
          8199 => x"76",
          8200 => x"81",
          8201 => x"70",
          8202 => x"56",
          8203 => x"82",
          8204 => x"78",
          8205 => x"80",
          8206 => x"27",
          8207 => x"19",
          8208 => x"7a",
          8209 => x"5c",
          8210 => x"55",
          8211 => x"7a",
          8212 => x"5c",
          8213 => x"2e",
          8214 => x"85",
          8215 => x"97",
          8216 => x"3d",
          8217 => x"19",
          8218 => x"33",
          8219 => x"05",
          8220 => x"78",
          8221 => x"80",
          8222 => x"82",
          8223 => x"80",
          8224 => x"04",
          8225 => x"7b",
          8226 => x"fc",
          8227 => x"53",
          8228 => x"fd",
          8229 => x"c8",
          8230 => x"d8",
          8231 => x"fe",
          8232 => x"33",
          8233 => x"f6",
          8234 => x"08",
          8235 => x"27",
          8236 => x"15",
          8237 => x"2a",
          8238 => x"51",
          8239 => x"83",
          8240 => x"94",
          8241 => x"80",
          8242 => x"0c",
          8243 => x"2e",
          8244 => x"79",
          8245 => x"70",
          8246 => x"51",
          8247 => x"2e",
          8248 => x"52",
          8249 => x"fe",
          8250 => x"82",
          8251 => x"ff",
          8252 => x"70",
          8253 => x"fe",
          8254 => x"82",
          8255 => x"73",
          8256 => x"76",
          8257 => x"06",
          8258 => x"0c",
          8259 => x"98",
          8260 => x"58",
          8261 => x"39",
          8262 => x"54",
          8263 => x"73",
          8264 => x"ff",
          8265 => x"82",
          8266 => x"54",
          8267 => x"08",
          8268 => x"9d",
          8269 => x"c8",
          8270 => x"81",
          8271 => x"d8",
          8272 => x"16",
          8273 => x"16",
          8274 => x"2e",
          8275 => x"76",
          8276 => x"de",
          8277 => x"31",
          8278 => x"18",
          8279 => x"90",
          8280 => x"81",
          8281 => x"06",
          8282 => x"56",
          8283 => x"9b",
          8284 => x"74",
          8285 => x"c5",
          8286 => x"c8",
          8287 => x"d8",
          8288 => x"38",
          8289 => x"08",
          8290 => x"73",
          8291 => x"ff",
          8292 => x"82",
          8293 => x"54",
          8294 => x"bf",
          8295 => x"27",
          8296 => x"53",
          8297 => x"08",
          8298 => x"73",
          8299 => x"ff",
          8300 => x"15",
          8301 => x"16",
          8302 => x"ff",
          8303 => x"80",
          8304 => x"73",
          8305 => x"ff",
          8306 => x"82",
          8307 => x"94",
          8308 => x"91",
          8309 => x"53",
          8310 => x"81",
          8311 => x"34",
          8312 => x"39",
          8313 => x"82",
          8314 => x"05",
          8315 => x"08",
          8316 => x"08",
          8317 => x"38",
          8318 => x"0c",
          8319 => x"80",
          8320 => x"72",
          8321 => x"73",
          8322 => x"53",
          8323 => x"8c",
          8324 => x"16",
          8325 => x"38",
          8326 => x"0c",
          8327 => x"82",
          8328 => x"8b",
          8329 => x"f9",
          8330 => x"56",
          8331 => x"80",
          8332 => x"38",
          8333 => x"3d",
          8334 => x"8a",
          8335 => x"51",
          8336 => x"82",
          8337 => x"55",
          8338 => x"08",
          8339 => x"77",
          8340 => x"52",
          8341 => x"a1",
          8342 => x"c8",
          8343 => x"d8",
          8344 => x"c4",
          8345 => x"33",
          8346 => x"55",
          8347 => x"24",
          8348 => x"16",
          8349 => x"2a",
          8350 => x"51",
          8351 => x"80",
          8352 => x"9c",
          8353 => x"77",
          8354 => x"3f",
          8355 => x"08",
          8356 => x"77",
          8357 => x"22",
          8358 => x"74",
          8359 => x"ff",
          8360 => x"82",
          8361 => x"55",
          8362 => x"09",
          8363 => x"38",
          8364 => x"39",
          8365 => x"84",
          8366 => x"0c",
          8367 => x"82",
          8368 => x"89",
          8369 => x"fc",
          8370 => x"87",
          8371 => x"53",
          8372 => x"e7",
          8373 => x"d8",
          8374 => x"38",
          8375 => x"08",
          8376 => x"3d",
          8377 => x"3d",
          8378 => x"89",
          8379 => x"54",
          8380 => x"54",
          8381 => x"82",
          8382 => x"53",
          8383 => x"08",
          8384 => x"74",
          8385 => x"d8",
          8386 => x"73",
          8387 => x"c0",
          8388 => x"c8",
          8389 => x"cb",
          8390 => x"c8",
          8391 => x"51",
          8392 => x"82",
          8393 => x"53",
          8394 => x"08",
          8395 => x"81",
          8396 => x"80",
          8397 => x"82",
          8398 => x"a7",
          8399 => x"73",
          8400 => x"3f",
          8401 => x"51",
          8402 => x"3f",
          8403 => x"08",
          8404 => x"30",
          8405 => x"9f",
          8406 => x"d8",
          8407 => x"51",
          8408 => x"72",
          8409 => x"0c",
          8410 => x"04",
          8411 => x"66",
          8412 => x"89",
          8413 => x"97",
          8414 => x"de",
          8415 => x"d8",
          8416 => x"82",
          8417 => x"b2",
          8418 => x"75",
          8419 => x"3f",
          8420 => x"08",
          8421 => x"c8",
          8422 => x"02",
          8423 => x"33",
          8424 => x"55",
          8425 => x"25",
          8426 => x"55",
          8427 => x"80",
          8428 => x"76",
          8429 => x"ce",
          8430 => x"82",
          8431 => x"95",
          8432 => x"f0",
          8433 => x"65",
          8434 => x"53",
          8435 => x"05",
          8436 => x"51",
          8437 => x"82",
          8438 => x"5b",
          8439 => x"08",
          8440 => x"7c",
          8441 => x"08",
          8442 => x"fe",
          8443 => x"08",
          8444 => x"55",
          8445 => x"91",
          8446 => x"0c",
          8447 => x"81",
          8448 => x"39",
          8449 => x"c9",
          8450 => x"c8",
          8451 => x"55",
          8452 => x"2e",
          8453 => x"80",
          8454 => x"75",
          8455 => x"52",
          8456 => x"05",
          8457 => x"b9",
          8458 => x"c8",
          8459 => x"cf",
          8460 => x"c8",
          8461 => x"cc",
          8462 => x"c8",
          8463 => x"82",
          8464 => x"07",
          8465 => x"05",
          8466 => x"53",
          8467 => x"9c",
          8468 => x"26",
          8469 => x"f9",
          8470 => x"08",
          8471 => x"08",
          8472 => x"98",
          8473 => x"81",
          8474 => x"58",
          8475 => x"3f",
          8476 => x"08",
          8477 => x"c8",
          8478 => x"38",
          8479 => x"77",
          8480 => x"5d",
          8481 => x"74",
          8482 => x"81",
          8483 => x"b8",
          8484 => x"a9",
          8485 => x"d8",
          8486 => x"ff",
          8487 => x"30",
          8488 => x"1b",
          8489 => x"5b",
          8490 => x"39",
          8491 => x"ff",
          8492 => x"82",
          8493 => x"f0",
          8494 => x"30",
          8495 => x"1b",
          8496 => x"5b",
          8497 => x"83",
          8498 => x"58",
          8499 => x"92",
          8500 => x"0c",
          8501 => x"12",
          8502 => x"33",
          8503 => x"54",
          8504 => x"34",
          8505 => x"c8",
          8506 => x"0d",
          8507 => x"0d",
          8508 => x"fc",
          8509 => x"52",
          8510 => x"3f",
          8511 => x"08",
          8512 => x"c8",
          8513 => x"38",
          8514 => x"56",
          8515 => x"38",
          8516 => x"70",
          8517 => x"81",
          8518 => x"55",
          8519 => x"80",
          8520 => x"38",
          8521 => x"54",
          8522 => x"08",
          8523 => x"38",
          8524 => x"82",
          8525 => x"53",
          8526 => x"52",
          8527 => x"b2",
          8528 => x"d8",
          8529 => x"88",
          8530 => x"80",
          8531 => x"17",
          8532 => x"51",
          8533 => x"3f",
          8534 => x"08",
          8535 => x"81",
          8536 => x"81",
          8537 => x"c8",
          8538 => x"09",
          8539 => x"38",
          8540 => x"39",
          8541 => x"77",
          8542 => x"c8",
          8543 => x"08",
          8544 => x"98",
          8545 => x"82",
          8546 => x"52",
          8547 => x"b2",
          8548 => x"d8",
          8549 => x"94",
          8550 => x"18",
          8551 => x"33",
          8552 => x"54",
          8553 => x"34",
          8554 => x"85",
          8555 => x"18",
          8556 => x"74",
          8557 => x"0c",
          8558 => x"04",
          8559 => x"82",
          8560 => x"ff",
          8561 => x"a3",
          8562 => x"93",
          8563 => x"c8",
          8564 => x"d8",
          8565 => x"f9",
          8566 => x"a3",
          8567 => x"96",
          8568 => x"58",
          8569 => x"82",
          8570 => x"55",
          8571 => x"08",
          8572 => x"02",
          8573 => x"33",
          8574 => x"70",
          8575 => x"55",
          8576 => x"73",
          8577 => x"75",
          8578 => x"80",
          8579 => x"c1",
          8580 => x"da",
          8581 => x"81",
          8582 => x"87",
          8583 => x"b1",
          8584 => x"78",
          8585 => x"87",
          8586 => x"c8",
          8587 => x"2a",
          8588 => x"51",
          8589 => x"80",
          8590 => x"38",
          8591 => x"d8",
          8592 => x"15",
          8593 => x"89",
          8594 => x"82",
          8595 => x"5c",
          8596 => x"3d",
          8597 => x"ff",
          8598 => x"82",
          8599 => x"55",
          8600 => x"08",
          8601 => x"82",
          8602 => x"52",
          8603 => x"bb",
          8604 => x"d8",
          8605 => x"82",
          8606 => x"86",
          8607 => x"80",
          8608 => x"d8",
          8609 => x"2e",
          8610 => x"d8",
          8611 => x"c1",
          8612 => x"c7",
          8613 => x"d8",
          8614 => x"d8",
          8615 => x"70",
          8616 => x"08",
          8617 => x"51",
          8618 => x"80",
          8619 => x"73",
          8620 => x"38",
          8621 => x"52",
          8622 => x"af",
          8623 => x"d8",
          8624 => x"74",
          8625 => x"51",
          8626 => x"3f",
          8627 => x"08",
          8628 => x"d8",
          8629 => x"3d",
          8630 => x"3d",
          8631 => x"9a",
          8632 => x"05",
          8633 => x"51",
          8634 => x"82",
          8635 => x"54",
          8636 => x"08",
          8637 => x"78",
          8638 => x"8e",
          8639 => x"58",
          8640 => x"82",
          8641 => x"54",
          8642 => x"08",
          8643 => x"54",
          8644 => x"82",
          8645 => x"84",
          8646 => x"06",
          8647 => x"02",
          8648 => x"33",
          8649 => x"81",
          8650 => x"86",
          8651 => x"fd",
          8652 => x"74",
          8653 => x"70",
          8654 => x"b0",
          8655 => x"d8",
          8656 => x"55",
          8657 => x"c8",
          8658 => x"87",
          8659 => x"c8",
          8660 => x"09",
          8661 => x"38",
          8662 => x"d8",
          8663 => x"2e",
          8664 => x"86",
          8665 => x"81",
          8666 => x"81",
          8667 => x"d8",
          8668 => x"78",
          8669 => x"e0",
          8670 => x"c8",
          8671 => x"d8",
          8672 => x"9f",
          8673 => x"a0",
          8674 => x"51",
          8675 => x"3f",
          8676 => x"0b",
          8677 => x"78",
          8678 => x"80",
          8679 => x"82",
          8680 => x"52",
          8681 => x"51",
          8682 => x"3f",
          8683 => x"b8",
          8684 => x"ff",
          8685 => x"a0",
          8686 => x"11",
          8687 => x"05",
          8688 => x"b2",
          8689 => x"ae",
          8690 => x"15",
          8691 => x"78",
          8692 => x"53",
          8693 => x"90",
          8694 => x"81",
          8695 => x"34",
          8696 => x"bf",
          8697 => x"d8",
          8698 => x"82",
          8699 => x"b3",
          8700 => x"b2",
          8701 => x"96",
          8702 => x"a3",
          8703 => x"53",
          8704 => x"51",
          8705 => x"3f",
          8706 => x"0b",
          8707 => x"78",
          8708 => x"83",
          8709 => x"51",
          8710 => x"3f",
          8711 => x"08",
          8712 => x"80",
          8713 => x"76",
          8714 => x"e5",
          8715 => x"d8",
          8716 => x"3d",
          8717 => x"3d",
          8718 => x"84",
          8719 => x"94",
          8720 => x"aa",
          8721 => x"05",
          8722 => x"51",
          8723 => x"82",
          8724 => x"55",
          8725 => x"08",
          8726 => x"78",
          8727 => x"08",
          8728 => x"70",
          8729 => x"91",
          8730 => x"c8",
          8731 => x"d8",
          8732 => x"be",
          8733 => x"9f",
          8734 => x"a0",
          8735 => x"55",
          8736 => x"38",
          8737 => x"3d",
          8738 => x"3d",
          8739 => x"51",
          8740 => x"3f",
          8741 => x"52",
          8742 => x"52",
          8743 => x"d6",
          8744 => x"08",
          8745 => x"c8",
          8746 => x"d8",
          8747 => x"82",
          8748 => x"97",
          8749 => x"3d",
          8750 => x"81",
          8751 => x"65",
          8752 => x"2e",
          8753 => x"55",
          8754 => x"82",
          8755 => x"84",
          8756 => x"06",
          8757 => x"73",
          8758 => x"d6",
          8759 => x"c8",
          8760 => x"d8",
          8761 => x"ca",
          8762 => x"93",
          8763 => x"ff",
          8764 => x"8d",
          8765 => x"a1",
          8766 => x"af",
          8767 => x"17",
          8768 => x"33",
          8769 => x"70",
          8770 => x"55",
          8771 => x"38",
          8772 => x"54",
          8773 => x"34",
          8774 => x"0b",
          8775 => x"8b",
          8776 => x"84",
          8777 => x"06",
          8778 => x"73",
          8779 => x"e7",
          8780 => x"2e",
          8781 => x"75",
          8782 => x"ff",
          8783 => x"82",
          8784 => x"52",
          8785 => x"a5",
          8786 => x"55",
          8787 => x"08",
          8788 => x"de",
          8789 => x"c8",
          8790 => x"51",
          8791 => x"3f",
          8792 => x"08",
          8793 => x"11",
          8794 => x"82",
          8795 => x"80",
          8796 => x"16",
          8797 => x"ae",
          8798 => x"06",
          8799 => x"53",
          8800 => x"51",
          8801 => x"3f",
          8802 => x"0b",
          8803 => x"87",
          8804 => x"c8",
          8805 => x"77",
          8806 => x"3f",
          8807 => x"08",
          8808 => x"c8",
          8809 => x"78",
          8810 => x"dc",
          8811 => x"c8",
          8812 => x"82",
          8813 => x"aa",
          8814 => x"ec",
          8815 => x"80",
          8816 => x"02",
          8817 => x"e3",
          8818 => x"57",
          8819 => x"3d",
          8820 => x"97",
          8821 => x"87",
          8822 => x"c8",
          8823 => x"d8",
          8824 => x"cf",
          8825 => x"66",
          8826 => x"d0",
          8827 => x"89",
          8828 => x"c8",
          8829 => x"d8",
          8830 => x"38",
          8831 => x"05",
          8832 => x"06",
          8833 => x"73",
          8834 => x"a7",
          8835 => x"09",
          8836 => x"71",
          8837 => x"06",
          8838 => x"55",
          8839 => x"15",
          8840 => x"81",
          8841 => x"34",
          8842 => x"a2",
          8843 => x"d8",
          8844 => x"74",
          8845 => x"0c",
          8846 => x"04",
          8847 => x"65",
          8848 => x"94",
          8849 => x"52",
          8850 => x"d1",
          8851 => x"d8",
          8852 => x"82",
          8853 => x"80",
          8854 => x"58",
          8855 => x"3d",
          8856 => x"c5",
          8857 => x"d8",
          8858 => x"82",
          8859 => x"b4",
          8860 => x"c7",
          8861 => x"a0",
          8862 => x"55",
          8863 => x"84",
          8864 => x"17",
          8865 => x"2b",
          8866 => x"96",
          8867 => x"9e",
          8868 => x"54",
          8869 => x"15",
          8870 => x"ff",
          8871 => x"82",
          8872 => x"55",
          8873 => x"c8",
          8874 => x"0d",
          8875 => x"0d",
          8876 => x"5a",
          8877 => x"3d",
          8878 => x"9a",
          8879 => x"9f",
          8880 => x"c8",
          8881 => x"c8",
          8882 => x"82",
          8883 => x"07",
          8884 => x"55",
          8885 => x"2e",
          8886 => x"81",
          8887 => x"55",
          8888 => x"2e",
          8889 => x"7b",
          8890 => x"80",
          8891 => x"70",
          8892 => x"ac",
          8893 => x"d8",
          8894 => x"82",
          8895 => x"80",
          8896 => x"52",
          8897 => x"b2",
          8898 => x"d8",
          8899 => x"82",
          8900 => x"bf",
          8901 => x"c8",
          8902 => x"c8",
          8903 => x"59",
          8904 => x"81",
          8905 => x"56",
          8906 => x"33",
          8907 => x"16",
          8908 => x"27",
          8909 => x"56",
          8910 => x"80",
          8911 => x"80",
          8912 => x"ff",
          8913 => x"70",
          8914 => x"56",
          8915 => x"e8",
          8916 => x"76",
          8917 => x"81",
          8918 => x"80",
          8919 => x"57",
          8920 => x"78",
          8921 => x"51",
          8922 => x"2e",
          8923 => x"73",
          8924 => x"38",
          8925 => x"08",
          8926 => x"9f",
          8927 => x"d8",
          8928 => x"82",
          8929 => x"a7",
          8930 => x"33",
          8931 => x"c3",
          8932 => x"2e",
          8933 => x"e4",
          8934 => x"2e",
          8935 => x"56",
          8936 => x"05",
          8937 => x"d6",
          8938 => x"c8",
          8939 => x"76",
          8940 => x"0c",
          8941 => x"04",
          8942 => x"82",
          8943 => x"ff",
          8944 => x"9d",
          8945 => x"97",
          8946 => x"c8",
          8947 => x"c8",
          8948 => x"82",
          8949 => x"82",
          8950 => x"53",
          8951 => x"3d",
          8952 => x"ff",
          8953 => x"73",
          8954 => x"51",
          8955 => x"74",
          8956 => x"38",
          8957 => x"3d",
          8958 => x"90",
          8959 => x"c8",
          8960 => x"ff",
          8961 => x"38",
          8962 => x"08",
          8963 => x"3f",
          8964 => x"82",
          8965 => x"51",
          8966 => x"82",
          8967 => x"83",
          8968 => x"55",
          8969 => x"a3",
          8970 => x"82",
          8971 => x"ff",
          8972 => x"82",
          8973 => x"93",
          8974 => x"75",
          8975 => x"75",
          8976 => x"38",
          8977 => x"76",
          8978 => x"86",
          8979 => x"39",
          8980 => x"27",
          8981 => x"88",
          8982 => x"77",
          8983 => x"59",
          8984 => x"56",
          8985 => x"81",
          8986 => x"81",
          8987 => x"33",
          8988 => x"73",
          8989 => x"fe",
          8990 => x"33",
          8991 => x"73",
          8992 => x"81",
          8993 => x"80",
          8994 => x"02",
          8995 => x"75",
          8996 => x"51",
          8997 => x"2e",
          8998 => x"87",
          8999 => x"56",
          9000 => x"78",
          9001 => x"80",
          9002 => x"70",
          9003 => x"a9",
          9004 => x"d8",
          9005 => x"82",
          9006 => x"80",
          9007 => x"52",
          9008 => x"af",
          9009 => x"d8",
          9010 => x"82",
          9011 => x"8d",
          9012 => x"c4",
          9013 => x"e5",
          9014 => x"c6",
          9015 => x"c8",
          9016 => x"09",
          9017 => x"cc",
          9018 => x"75",
          9019 => x"c4",
          9020 => x"74",
          9021 => x"9c",
          9022 => x"c8",
          9023 => x"d8",
          9024 => x"38",
          9025 => x"d8",
          9026 => x"66",
          9027 => x"89",
          9028 => x"88",
          9029 => x"34",
          9030 => x"52",
          9031 => x"99",
          9032 => x"54",
          9033 => x"15",
          9034 => x"ff",
          9035 => x"82",
          9036 => x"54",
          9037 => x"82",
          9038 => x"9c",
          9039 => x"f2",
          9040 => x"62",
          9041 => x"80",
          9042 => x"93",
          9043 => x"55",
          9044 => x"5e",
          9045 => x"3f",
          9046 => x"08",
          9047 => x"c8",
          9048 => x"38",
          9049 => x"58",
          9050 => x"38",
          9051 => x"97",
          9052 => x"08",
          9053 => x"38",
          9054 => x"70",
          9055 => x"81",
          9056 => x"55",
          9057 => x"87",
          9058 => x"39",
          9059 => x"90",
          9060 => x"82",
          9061 => x"8a",
          9062 => x"89",
          9063 => x"7f",
          9064 => x"56",
          9065 => x"3f",
          9066 => x"06",
          9067 => x"72",
          9068 => x"82",
          9069 => x"05",
          9070 => x"7c",
          9071 => x"55",
          9072 => x"27",
          9073 => x"16",
          9074 => x"83",
          9075 => x"76",
          9076 => x"80",
          9077 => x"79",
          9078 => x"85",
          9079 => x"7f",
          9080 => x"14",
          9081 => x"83",
          9082 => x"82",
          9083 => x"81",
          9084 => x"38",
          9085 => x"08",
          9086 => x"95",
          9087 => x"c8",
          9088 => x"81",
          9089 => x"7b",
          9090 => x"06",
          9091 => x"39",
          9092 => x"56",
          9093 => x"09",
          9094 => x"b9",
          9095 => x"80",
          9096 => x"80",
          9097 => x"78",
          9098 => x"7a",
          9099 => x"38",
          9100 => x"73",
          9101 => x"81",
          9102 => x"ff",
          9103 => x"74",
          9104 => x"ff",
          9105 => x"82",
          9106 => x"58",
          9107 => x"08",
          9108 => x"74",
          9109 => x"16",
          9110 => x"73",
          9111 => x"39",
          9112 => x"7e",
          9113 => x"0c",
          9114 => x"2e",
          9115 => x"88",
          9116 => x"8c",
          9117 => x"1a",
          9118 => x"07",
          9119 => x"1b",
          9120 => x"08",
          9121 => x"16",
          9122 => x"75",
          9123 => x"38",
          9124 => x"94",
          9125 => x"15",
          9126 => x"54",
          9127 => x"34",
          9128 => x"82",
          9129 => x"90",
          9130 => x"e9",
          9131 => x"6d",
          9132 => x"80",
          9133 => x"9d",
          9134 => x"5c",
          9135 => x"3f",
          9136 => x"0b",
          9137 => x"08",
          9138 => x"38",
          9139 => x"08",
          9140 => x"f0",
          9141 => x"08",
          9142 => x"80",
          9143 => x"80",
          9144 => x"d8",
          9145 => x"ff",
          9146 => x"52",
          9147 => x"8e",
          9148 => x"d8",
          9149 => x"ff",
          9150 => x"06",
          9151 => x"56",
          9152 => x"38",
          9153 => x"70",
          9154 => x"55",
          9155 => x"8b",
          9156 => x"3d",
          9157 => x"83",
          9158 => x"ff",
          9159 => x"82",
          9160 => x"99",
          9161 => x"74",
          9162 => x"38",
          9163 => x"80",
          9164 => x"ff",
          9165 => x"55",
          9166 => x"83",
          9167 => x"78",
          9168 => x"38",
          9169 => x"26",
          9170 => x"81",
          9171 => x"8b",
          9172 => x"79",
          9173 => x"80",
          9174 => x"93",
          9175 => x"39",
          9176 => x"6e",
          9177 => x"89",
          9178 => x"48",
          9179 => x"83",
          9180 => x"61",
          9181 => x"25",
          9182 => x"55",
          9183 => x"8a",
          9184 => x"3d",
          9185 => x"81",
          9186 => x"ff",
          9187 => x"81",
          9188 => x"c8",
          9189 => x"38",
          9190 => x"70",
          9191 => x"d8",
          9192 => x"56",
          9193 => x"38",
          9194 => x"55",
          9195 => x"75",
          9196 => x"38",
          9197 => x"70",
          9198 => x"ff",
          9199 => x"83",
          9200 => x"78",
          9201 => x"89",
          9202 => x"81",
          9203 => x"06",
          9204 => x"80",
          9205 => x"77",
          9206 => x"74",
          9207 => x"8d",
          9208 => x"06",
          9209 => x"2e",
          9210 => x"77",
          9211 => x"93",
          9212 => x"74",
          9213 => x"cb",
          9214 => x"7d",
          9215 => x"81",
          9216 => x"38",
          9217 => x"66",
          9218 => x"81",
          9219 => x"84",
          9220 => x"74",
          9221 => x"38",
          9222 => x"98",
          9223 => x"84",
          9224 => x"82",
          9225 => x"57",
          9226 => x"80",
          9227 => x"76",
          9228 => x"38",
          9229 => x"51",
          9230 => x"3f",
          9231 => x"08",
          9232 => x"87",
          9233 => x"2a",
          9234 => x"5c",
          9235 => x"d8",
          9236 => x"80",
          9237 => x"44",
          9238 => x"0a",
          9239 => x"ec",
          9240 => x"39",
          9241 => x"66",
          9242 => x"81",
          9243 => x"f4",
          9244 => x"74",
          9245 => x"38",
          9246 => x"98",
          9247 => x"f4",
          9248 => x"82",
          9249 => x"57",
          9250 => x"80",
          9251 => x"76",
          9252 => x"38",
          9253 => x"51",
          9254 => x"3f",
          9255 => x"08",
          9256 => x"57",
          9257 => x"08",
          9258 => x"96",
          9259 => x"82",
          9260 => x"10",
          9261 => x"08",
          9262 => x"72",
          9263 => x"59",
          9264 => x"ff",
          9265 => x"5d",
          9266 => x"44",
          9267 => x"11",
          9268 => x"70",
          9269 => x"71",
          9270 => x"06",
          9271 => x"52",
          9272 => x"40",
          9273 => x"09",
          9274 => x"38",
          9275 => x"18",
          9276 => x"39",
          9277 => x"79",
          9278 => x"70",
          9279 => x"58",
          9280 => x"76",
          9281 => x"38",
          9282 => x"7d",
          9283 => x"70",
          9284 => x"55",
          9285 => x"3f",
          9286 => x"08",
          9287 => x"2e",
          9288 => x"9b",
          9289 => x"c8",
          9290 => x"f5",
          9291 => x"38",
          9292 => x"38",
          9293 => x"59",
          9294 => x"38",
          9295 => x"7d",
          9296 => x"81",
          9297 => x"38",
          9298 => x"0b",
          9299 => x"08",
          9300 => x"78",
          9301 => x"1a",
          9302 => x"c0",
          9303 => x"74",
          9304 => x"39",
          9305 => x"55",
          9306 => x"8f",
          9307 => x"fd",
          9308 => x"d8",
          9309 => x"f5",
          9310 => x"78",
          9311 => x"79",
          9312 => x"80",
          9313 => x"f1",
          9314 => x"39",
          9315 => x"81",
          9316 => x"06",
          9317 => x"55",
          9318 => x"27",
          9319 => x"81",
          9320 => x"56",
          9321 => x"38",
          9322 => x"80",
          9323 => x"ff",
          9324 => x"8b",
          9325 => x"8c",
          9326 => x"ff",
          9327 => x"84",
          9328 => x"1b",
          9329 => x"e1",
          9330 => x"1c",
          9331 => x"ff",
          9332 => x"8e",
          9333 => x"8f",
          9334 => x"0b",
          9335 => x"7d",
          9336 => x"30",
          9337 => x"84",
          9338 => x"51",
          9339 => x"51",
          9340 => x"3f",
          9341 => x"83",
          9342 => x"90",
          9343 => x"ff",
          9344 => x"93",
          9345 => x"8f",
          9346 => x"39",
          9347 => x"1b",
          9348 => x"b3",
          9349 => x"95",
          9350 => x"52",
          9351 => x"ff",
          9352 => x"81",
          9353 => x"1b",
          9354 => x"fd",
          9355 => x"9c",
          9356 => x"8f",
          9357 => x"83",
          9358 => x"06",
          9359 => x"82",
          9360 => x"52",
          9361 => x"51",
          9362 => x"3f",
          9363 => x"1b",
          9364 => x"f3",
          9365 => x"ac",
          9366 => x"8e",
          9367 => x"52",
          9368 => x"ff",
          9369 => x"86",
          9370 => x"51",
          9371 => x"3f",
          9372 => x"80",
          9373 => x"a9",
          9374 => x"1c",
          9375 => x"82",
          9376 => x"80",
          9377 => x"ae",
          9378 => x"b2",
          9379 => x"1b",
          9380 => x"b3",
          9381 => x"ff",
          9382 => x"96",
          9383 => x"8e",
          9384 => x"80",
          9385 => x"34",
          9386 => x"1c",
          9387 => x"82",
          9388 => x"ab",
          9389 => x"8e",
          9390 => x"d4",
          9391 => x"fe",
          9392 => x"59",
          9393 => x"3f",
          9394 => x"53",
          9395 => x"51",
          9396 => x"3f",
          9397 => x"d8",
          9398 => x"e7",
          9399 => x"2e",
          9400 => x"80",
          9401 => x"54",
          9402 => x"53",
          9403 => x"51",
          9404 => x"3f",
          9405 => x"80",
          9406 => x"ff",
          9407 => x"84",
          9408 => x"d2",
          9409 => x"ff",
          9410 => x"86",
          9411 => x"f2",
          9412 => x"1b",
          9413 => x"af",
          9414 => x"52",
          9415 => x"51",
          9416 => x"3f",
          9417 => x"ec",
          9418 => x"8d",
          9419 => x"d4",
          9420 => x"51",
          9421 => x"3f",
          9422 => x"87",
          9423 => x"52",
          9424 => x"89",
          9425 => x"54",
          9426 => x"7a",
          9427 => x"ff",
          9428 => x"65",
          9429 => x"7a",
          9430 => x"bd",
          9431 => x"80",
          9432 => x"2e",
          9433 => x"9a",
          9434 => x"7a",
          9435 => x"d7",
          9436 => x"84",
          9437 => x"8c",
          9438 => x"0a",
          9439 => x"51",
          9440 => x"ff",
          9441 => x"7d",
          9442 => x"38",
          9443 => x"52",
          9444 => x"8c",
          9445 => x"55",
          9446 => x"62",
          9447 => x"74",
          9448 => x"75",
          9449 => x"7e",
          9450 => x"ac",
          9451 => x"c8",
          9452 => x"38",
          9453 => x"82",
          9454 => x"52",
          9455 => x"8c",
          9456 => x"16",
          9457 => x"56",
          9458 => x"38",
          9459 => x"77",
          9460 => x"8d",
          9461 => x"7d",
          9462 => x"38",
          9463 => x"57",
          9464 => x"83",
          9465 => x"76",
          9466 => x"7a",
          9467 => x"ff",
          9468 => x"82",
          9469 => x"81",
          9470 => x"16",
          9471 => x"56",
          9472 => x"38",
          9473 => x"83",
          9474 => x"86",
          9475 => x"ff",
          9476 => x"38",
          9477 => x"82",
          9478 => x"81",
          9479 => x"06",
          9480 => x"fe",
          9481 => x"53",
          9482 => x"51",
          9483 => x"3f",
          9484 => x"52",
          9485 => x"8a",
          9486 => x"be",
          9487 => x"75",
          9488 => x"81",
          9489 => x"0b",
          9490 => x"77",
          9491 => x"75",
          9492 => x"60",
          9493 => x"80",
          9494 => x"75",
          9495 => x"a3",
          9496 => x"85",
          9497 => x"d8",
          9498 => x"2a",
          9499 => x"75",
          9500 => x"82",
          9501 => x"87",
          9502 => x"52",
          9503 => x"51",
          9504 => x"3f",
          9505 => x"ca",
          9506 => x"8a",
          9507 => x"54",
          9508 => x"52",
          9509 => x"86",
          9510 => x"56",
          9511 => x"08",
          9512 => x"53",
          9513 => x"51",
          9514 => x"3f",
          9515 => x"d8",
          9516 => x"38",
          9517 => x"56",
          9518 => x"56",
          9519 => x"d8",
          9520 => x"75",
          9521 => x"0c",
          9522 => x"04",
          9523 => x"7d",
          9524 => x"80",
          9525 => x"05",
          9526 => x"76",
          9527 => x"38",
          9528 => x"11",
          9529 => x"53",
          9530 => x"79",
          9531 => x"3f",
          9532 => x"09",
          9533 => x"38",
          9534 => x"55",
          9535 => x"db",
          9536 => x"70",
          9537 => x"34",
          9538 => x"74",
          9539 => x"81",
          9540 => x"80",
          9541 => x"55",
          9542 => x"76",
          9543 => x"d8",
          9544 => x"3d",
          9545 => x"3d",
          9546 => x"84",
          9547 => x"33",
          9548 => x"8a",
          9549 => x"06",
          9550 => x"52",
          9551 => x"3f",
          9552 => x"56",
          9553 => x"be",
          9554 => x"08",
          9555 => x"05",
          9556 => x"75",
          9557 => x"56",
          9558 => x"a1",
          9559 => x"fc",
          9560 => x"53",
          9561 => x"76",
          9562 => x"c0",
          9563 => x"32",
          9564 => x"72",
          9565 => x"70",
          9566 => x"56",
          9567 => x"18",
          9568 => x"88",
          9569 => x"3d",
          9570 => x"3d",
          9571 => x"11",
          9572 => x"80",
          9573 => x"38",
          9574 => x"05",
          9575 => x"8c",
          9576 => x"08",
          9577 => x"3f",
          9578 => x"08",
          9579 => x"16",
          9580 => x"09",
          9581 => x"38",
          9582 => x"55",
          9583 => x"55",
          9584 => x"c8",
          9585 => x"0d",
          9586 => x"0d",
          9587 => x"cc",
          9588 => x"73",
          9589 => x"c1",
          9590 => x"0c",
          9591 => x"04",
          9592 => x"02",
          9593 => x"33",
          9594 => x"3d",
          9595 => x"54",
          9596 => x"52",
          9597 => x"ae",
          9598 => x"ff",
          9599 => x"3d",
          9600 => x"3d",
          9601 => x"84",
          9602 => x"22",
          9603 => x"52",
          9604 => x"26",
          9605 => x"83",
          9606 => x"52",
          9607 => x"83",
          9608 => x"27",
          9609 => x"b5",
          9610 => x"06",
          9611 => x"80",
          9612 => x"82",
          9613 => x"51",
          9614 => x"9c",
          9615 => x"70",
          9616 => x"06",
          9617 => x"80",
          9618 => x"38",
          9619 => x"cc",
          9620 => x"22",
          9621 => x"39",
          9622 => x"70",
          9623 => x"53",
          9624 => x"d8",
          9625 => x"3d",
          9626 => x"3d",
          9627 => x"05",
          9628 => x"05",
          9629 => x"53",
          9630 => x"70",
          9631 => x"85",
          9632 => x"9a",
          9633 => x"b5",
          9634 => x"06",
          9635 => x"81",
          9636 => x"38",
          9637 => x"ca",
          9638 => x"22",
          9639 => x"82",
          9640 => x"84",
          9641 => x"fb",
          9642 => x"51",
          9643 => x"ff",
          9644 => x"38",
          9645 => x"ff",
          9646 => x"94",
          9647 => x"ff",
          9648 => x"38",
          9649 => x"56",
          9650 => x"05",
          9651 => x"30",
          9652 => x"72",
          9653 => x"51",
          9654 => x"80",
          9655 => x"70",
          9656 => x"22",
          9657 => x"71",
          9658 => x"70",
          9659 => x"55",
          9660 => x"25",
          9661 => x"73",
          9662 => x"dc",
          9663 => x"29",
          9664 => x"05",
          9665 => x"04",
          9666 => x"10",
          9667 => x"22",
          9668 => x"80",
          9669 => x"75",
          9670 => x"72",
          9671 => x"51",
          9672 => x"12",
          9673 => x"e0",
          9674 => x"39",
          9675 => x"95",
          9676 => x"51",
          9677 => x"12",
          9678 => x"ff",
          9679 => x"85",
          9680 => x"12",
          9681 => x"ff",
          9682 => x"8c",
          9683 => x"f8",
          9684 => x"16",
          9685 => x"39",
          9686 => x"82",
          9687 => x"87",
          9688 => x"00",
          9689 => x"ff",
          9690 => x"ff",
          9691 => x"ff",
          9692 => x"00",
          9693 => x"aa",
          9694 => x"2e",
          9695 => x"35",
          9696 => x"3c",
          9697 => x"43",
          9698 => x"4a",
          9699 => x"51",
          9700 => x"58",
          9701 => x"5f",
          9702 => x"66",
          9703 => x"6d",
          9704 => x"74",
          9705 => x"7a",
          9706 => x"80",
          9707 => x"86",
          9708 => x"8c",
          9709 => x"92",
          9710 => x"98",
          9711 => x"9e",
          9712 => x"a4",
          9713 => x"a6",
          9714 => x"ac",
          9715 => x"b2",
          9716 => x"b8",
          9717 => x"be",
          9718 => x"dd",
          9719 => x"dd",
          9720 => x"ee",
          9721 => x"46",
          9722 => x"c5",
          9723 => x"b2",
          9724 => x"b6",
          9725 => x"17",
          9726 => x"f9",
          9727 => x"8f",
          9728 => x"15",
          9729 => x"98",
          9730 => x"b2",
          9731 => x"ee",
          9732 => x"17",
          9733 => x"b6",
          9734 => x"b2",
          9735 => x"b2",
          9736 => x"15",
          9737 => x"8f",
          9738 => x"17",
          9739 => x"46",
          9740 => x"08",
          9741 => x"16",
          9742 => x"22",
          9743 => x"27",
          9744 => x"2c",
          9745 => x"31",
          9746 => x"36",
          9747 => x"3b",
          9748 => x"41",
          9749 => x"31",
          9750 => x"1a",
          9751 => x"1a",
          9752 => x"60",
          9753 => x"1a",
          9754 => x"1a",
          9755 => x"1a",
          9756 => x"1a",
          9757 => x"1a",
          9758 => x"1a",
          9759 => x"1a",
          9760 => x"1d",
          9761 => x"1a",
          9762 => x"48",
          9763 => x"78",
          9764 => x"1a",
          9765 => x"1a",
          9766 => x"1a",
          9767 => x"1a",
          9768 => x"1a",
          9769 => x"1a",
          9770 => x"1a",
          9771 => x"1a",
          9772 => x"1a",
          9773 => x"1a",
          9774 => x"1a",
          9775 => x"1a",
          9776 => x"1a",
          9777 => x"1a",
          9778 => x"1a",
          9779 => x"1a",
          9780 => x"1a",
          9781 => x"1a",
          9782 => x"1a",
          9783 => x"1a",
          9784 => x"1a",
          9785 => x"1a",
          9786 => x"1a",
          9787 => x"1a",
          9788 => x"1a",
          9789 => x"1a",
          9790 => x"1a",
          9791 => x"1a",
          9792 => x"1a",
          9793 => x"1a",
          9794 => x"1a",
          9795 => x"1a",
          9796 => x"1a",
          9797 => x"1a",
          9798 => x"1a",
          9799 => x"1a",
          9800 => x"a8",
          9801 => x"1a",
          9802 => x"1a",
          9803 => x"1a",
          9804 => x"1a",
          9805 => x"16",
          9806 => x"1a",
          9807 => x"1a",
          9808 => x"1a",
          9809 => x"1a",
          9810 => x"1a",
          9811 => x"1a",
          9812 => x"1a",
          9813 => x"1a",
          9814 => x"1a",
          9815 => x"1a",
          9816 => x"d8",
          9817 => x"3f",
          9818 => x"af",
          9819 => x"af",
          9820 => x"af",
          9821 => x"1a",
          9822 => x"3f",
          9823 => x"1a",
          9824 => x"1a",
          9825 => x"98",
          9826 => x"1a",
          9827 => x"1a",
          9828 => x"ec",
          9829 => x"f7",
          9830 => x"1a",
          9831 => x"1a",
          9832 => x"11",
          9833 => x"1a",
          9834 => x"1f",
          9835 => x"1a",
          9836 => x"1a",
          9837 => x"16",
          9838 => x"69",
          9839 => x"00",
          9840 => x"63",
          9841 => x"00",
          9842 => x"69",
          9843 => x"00",
          9844 => x"61",
          9845 => x"00",
          9846 => x"65",
          9847 => x"00",
          9848 => x"65",
          9849 => x"00",
          9850 => x"70",
          9851 => x"00",
          9852 => x"66",
          9853 => x"00",
          9854 => x"6d",
          9855 => x"00",
          9856 => x"00",
          9857 => x"00",
          9858 => x"00",
          9859 => x"00",
          9860 => x"00",
          9861 => x"00",
          9862 => x"00",
          9863 => x"6c",
          9864 => x"00",
          9865 => x"00",
          9866 => x"74",
          9867 => x"00",
          9868 => x"65",
          9869 => x"00",
          9870 => x"6f",
          9871 => x"00",
          9872 => x"74",
          9873 => x"00",
          9874 => x"73",
          9875 => x"00",
          9876 => x"73",
          9877 => x"00",
          9878 => x"6f",
          9879 => x"00",
          9880 => x"00",
          9881 => x"6b",
          9882 => x"72",
          9883 => x"00",
          9884 => x"65",
          9885 => x"6c",
          9886 => x"72",
          9887 => x"00",
          9888 => x"6b",
          9889 => x"74",
          9890 => x"61",
          9891 => x"00",
          9892 => x"66",
          9893 => x"20",
          9894 => x"6e",
          9895 => x"00",
          9896 => x"70",
          9897 => x"20",
          9898 => x"6e",
          9899 => x"00",
          9900 => x"61",
          9901 => x"20",
          9902 => x"65",
          9903 => x"65",
          9904 => x"00",
          9905 => x"65",
          9906 => x"64",
          9907 => x"65",
          9908 => x"00",
          9909 => x"65",
          9910 => x"72",
          9911 => x"79",
          9912 => x"69",
          9913 => x"2e",
          9914 => x"00",
          9915 => x"65",
          9916 => x"6e",
          9917 => x"20",
          9918 => x"61",
          9919 => x"2e",
          9920 => x"00",
          9921 => x"69",
          9922 => x"72",
          9923 => x"20",
          9924 => x"74",
          9925 => x"65",
          9926 => x"00",
          9927 => x"76",
          9928 => x"75",
          9929 => x"72",
          9930 => x"20",
          9931 => x"61",
          9932 => x"2e",
          9933 => x"00",
          9934 => x"6b",
          9935 => x"74",
          9936 => x"61",
          9937 => x"64",
          9938 => x"00",
          9939 => x"63",
          9940 => x"61",
          9941 => x"6c",
          9942 => x"69",
          9943 => x"79",
          9944 => x"6d",
          9945 => x"75",
          9946 => x"6f",
          9947 => x"69",
          9948 => x"00",
          9949 => x"6d",
          9950 => x"61",
          9951 => x"74",
          9952 => x"00",
          9953 => x"65",
          9954 => x"2c",
          9955 => x"65",
          9956 => x"69",
          9957 => x"63",
          9958 => x"65",
          9959 => x"64",
          9960 => x"00",
          9961 => x"65",
          9962 => x"20",
          9963 => x"6b",
          9964 => x"00",
          9965 => x"75",
          9966 => x"63",
          9967 => x"74",
          9968 => x"6d",
          9969 => x"2e",
          9970 => x"00",
          9971 => x"20",
          9972 => x"79",
          9973 => x"65",
          9974 => x"69",
          9975 => x"2e",
          9976 => x"00",
          9977 => x"61",
          9978 => x"65",
          9979 => x"69",
          9980 => x"72",
          9981 => x"74",
          9982 => x"00",
          9983 => x"63",
          9984 => x"2e",
          9985 => x"00",
          9986 => x"6e",
          9987 => x"20",
          9988 => x"6f",
          9989 => x"00",
          9990 => x"75",
          9991 => x"74",
          9992 => x"25",
          9993 => x"74",
          9994 => x"75",
          9995 => x"74",
          9996 => x"73",
          9997 => x"0a",
          9998 => x"00",
          9999 => x"64",
         10000 => x"00",
         10001 => x"30",
         10002 => x"2c",
         10003 => x"25",
         10004 => x"78",
         10005 => x"3d",
         10006 => x"6c",
         10007 => x"5f",
         10008 => x"3d",
         10009 => x"6c",
         10010 => x"30",
         10011 => x"20",
         10012 => x"6c",
         10013 => x"00",
         10014 => x"6c",
         10015 => x"00",
         10016 => x"00",
         10017 => x"58",
         10018 => x"00",
         10019 => x"20",
         10020 => x"20",
         10021 => x"00",
         10022 => x"58",
         10023 => x"00",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"54",
         10028 => x"00",
         10029 => x"20",
         10030 => x"28",
         10031 => x"00",
         10032 => x"30",
         10033 => x"30",
         10034 => x"00",
         10035 => x"35",
         10036 => x"00",
         10037 => x"55",
         10038 => x"65",
         10039 => x"30",
         10040 => x"20",
         10041 => x"25",
         10042 => x"2a",
         10043 => x"00",
         10044 => x"54",
         10045 => x"6e",
         10046 => x"72",
         10047 => x"20",
         10048 => x"64",
         10049 => x"00",
         10050 => x"65",
         10051 => x"6e",
         10052 => x"72",
         10053 => x"00",
         10054 => x"20",
         10055 => x"65",
         10056 => x"70",
         10057 => x"00",
         10058 => x"54",
         10059 => x"44",
         10060 => x"74",
         10061 => x"75",
         10062 => x"00",
         10063 => x"54",
         10064 => x"52",
         10065 => x"74",
         10066 => x"75",
         10067 => x"00",
         10068 => x"54",
         10069 => x"58",
         10070 => x"74",
         10071 => x"75",
         10072 => x"00",
         10073 => x"54",
         10074 => x"58",
         10075 => x"74",
         10076 => x"75",
         10077 => x"00",
         10078 => x"54",
         10079 => x"58",
         10080 => x"74",
         10081 => x"75",
         10082 => x"00",
         10083 => x"54",
         10084 => x"58",
         10085 => x"74",
         10086 => x"75",
         10087 => x"00",
         10088 => x"74",
         10089 => x"20",
         10090 => x"74",
         10091 => x"72",
         10092 => x"00",
         10093 => x"62",
         10094 => x"67",
         10095 => x"6d",
         10096 => x"2e",
         10097 => x"00",
         10098 => x"6f",
         10099 => x"63",
         10100 => x"74",
         10101 => x"00",
         10102 => x"74",
         10103 => x"73",
         10104 => x"00",
         10105 => x"00",
         10106 => x"6c",
         10107 => x"74",
         10108 => x"6e",
         10109 => x"61",
         10110 => x"65",
         10111 => x"20",
         10112 => x"64",
         10113 => x"20",
         10114 => x"61",
         10115 => x"69",
         10116 => x"20",
         10117 => x"75",
         10118 => x"79",
         10119 => x"00",
         10120 => x"00",
         10121 => x"20",
         10122 => x"6b",
         10123 => x"21",
         10124 => x"00",
         10125 => x"74",
         10126 => x"69",
         10127 => x"2e",
         10128 => x"00",
         10129 => x"6c",
         10130 => x"74",
         10131 => x"6e",
         10132 => x"61",
         10133 => x"65",
         10134 => x"00",
         10135 => x"25",
         10136 => x"00",
         10137 => x"00",
         10138 => x"61",
         10139 => x"67",
         10140 => x"2e",
         10141 => x"00",
         10142 => x"79",
         10143 => x"2e",
         10144 => x"00",
         10145 => x"70",
         10146 => x"6e",
         10147 => x"2e",
         10148 => x"00",
         10149 => x"6c",
         10150 => x"30",
         10151 => x"2d",
         10152 => x"38",
         10153 => x"25",
         10154 => x"29",
         10155 => x"00",
         10156 => x"70",
         10157 => x"6d",
         10158 => x"00",
         10159 => x"6d",
         10160 => x"74",
         10161 => x"00",
         10162 => x"6c",
         10163 => x"30",
         10164 => x"00",
         10165 => x"00",
         10166 => x"6c",
         10167 => x"30",
         10168 => x"00",
         10169 => x"6c",
         10170 => x"30",
         10171 => x"2d",
         10172 => x"00",
         10173 => x"61",
         10174 => x"6e",
         10175 => x"6e",
         10176 => x"72",
         10177 => x"73",
         10178 => x"00",
         10179 => x"62",
         10180 => x"67",
         10181 => x"74",
         10182 => x"75",
         10183 => x"00",
         10184 => x"61",
         10185 => x"64",
         10186 => x"72",
         10187 => x"69",
         10188 => x"00",
         10189 => x"62",
         10190 => x"67",
         10191 => x"72",
         10192 => x"69",
         10193 => x"00",
         10194 => x"63",
         10195 => x"6e",
         10196 => x"6f",
         10197 => x"40",
         10198 => x"38",
         10199 => x"2e",
         10200 => x"00",
         10201 => x"6c",
         10202 => x"20",
         10203 => x"65",
         10204 => x"25",
         10205 => x"78",
         10206 => x"2e",
         10207 => x"00",
         10208 => x"6c",
         10209 => x"74",
         10210 => x"65",
         10211 => x"6f",
         10212 => x"28",
         10213 => x"2e",
         10214 => x"00",
         10215 => x"74",
         10216 => x"69",
         10217 => x"61",
         10218 => x"69",
         10219 => x"69",
         10220 => x"2e",
         10221 => x"00",
         10222 => x"64",
         10223 => x"62",
         10224 => x"69",
         10225 => x"2e",
         10226 => x"00",
         10227 => x"00",
         10228 => x"00",
         10229 => x"5c",
         10230 => x"25",
         10231 => x"73",
         10232 => x"00",
         10233 => x"5c",
         10234 => x"25",
         10235 => x"00",
         10236 => x"5c",
         10237 => x"00",
         10238 => x"20",
         10239 => x"6d",
         10240 => x"2e",
         10241 => x"00",
         10242 => x"6e",
         10243 => x"2e",
         10244 => x"00",
         10245 => x"62",
         10246 => x"67",
         10247 => x"74",
         10248 => x"75",
         10249 => x"2e",
         10250 => x"00",
         10251 => x"25",
         10252 => x"64",
         10253 => x"3a",
         10254 => x"25",
         10255 => x"64",
         10256 => x"00",
         10257 => x"20",
         10258 => x"66",
         10259 => x"72",
         10260 => x"6f",
         10261 => x"00",
         10262 => x"72",
         10263 => x"53",
         10264 => x"63",
         10265 => x"69",
         10266 => x"00",
         10267 => x"65",
         10268 => x"65",
         10269 => x"6d",
         10270 => x"6d",
         10271 => x"65",
         10272 => x"00",
         10273 => x"20",
         10274 => x"53",
         10275 => x"4d",
         10276 => x"25",
         10277 => x"3a",
         10278 => x"58",
         10279 => x"00",
         10280 => x"20",
         10281 => x"41",
         10282 => x"20",
         10283 => x"25",
         10284 => x"3a",
         10285 => x"58",
         10286 => x"00",
         10287 => x"20",
         10288 => x"4e",
         10289 => x"41",
         10290 => x"25",
         10291 => x"3a",
         10292 => x"58",
         10293 => x"00",
         10294 => x"20",
         10295 => x"4d",
         10296 => x"20",
         10297 => x"25",
         10298 => x"3a",
         10299 => x"58",
         10300 => x"00",
         10301 => x"20",
         10302 => x"20",
         10303 => x"20",
         10304 => x"25",
         10305 => x"3a",
         10306 => x"58",
         10307 => x"00",
         10308 => x"20",
         10309 => x"43",
         10310 => x"20",
         10311 => x"44",
         10312 => x"63",
         10313 => x"3d",
         10314 => x"64",
         10315 => x"00",
         10316 => x"20",
         10317 => x"45",
         10318 => x"20",
         10319 => x"54",
         10320 => x"72",
         10321 => x"3d",
         10322 => x"64",
         10323 => x"00",
         10324 => x"20",
         10325 => x"52",
         10326 => x"52",
         10327 => x"43",
         10328 => x"6e",
         10329 => x"3d",
         10330 => x"64",
         10331 => x"00",
         10332 => x"20",
         10333 => x"48",
         10334 => x"45",
         10335 => x"53",
         10336 => x"00",
         10337 => x"20",
         10338 => x"49",
         10339 => x"00",
         10340 => x"20",
         10341 => x"54",
         10342 => x"00",
         10343 => x"20",
         10344 => x"00",
         10345 => x"20",
         10346 => x"00",
         10347 => x"72",
         10348 => x"65",
         10349 => x"00",
         10350 => x"20",
         10351 => x"20",
         10352 => x"65",
         10353 => x"65",
         10354 => x"72",
         10355 => x"64",
         10356 => x"73",
         10357 => x"25",
         10358 => x"0a",
         10359 => x"00",
         10360 => x"20",
         10361 => x"20",
         10362 => x"6f",
         10363 => x"53",
         10364 => x"74",
         10365 => x"64",
         10366 => x"73",
         10367 => x"25",
         10368 => x"0a",
         10369 => x"00",
         10370 => x"20",
         10371 => x"63",
         10372 => x"74",
         10373 => x"20",
         10374 => x"72",
         10375 => x"20",
         10376 => x"20",
         10377 => x"25",
         10378 => x"0a",
         10379 => x"00",
         10380 => x"63",
         10381 => x"00",
         10382 => x"20",
         10383 => x"20",
         10384 => x"20",
         10385 => x"20",
         10386 => x"20",
         10387 => x"20",
         10388 => x"20",
         10389 => x"25",
         10390 => x"0a",
         10391 => x"00",
         10392 => x"20",
         10393 => x"74",
         10394 => x"43",
         10395 => x"6b",
         10396 => x"65",
         10397 => x"20",
         10398 => x"20",
         10399 => x"25",
         10400 => x"30",
         10401 => x"48",
         10402 => x"00",
         10403 => x"20",
         10404 => x"41",
         10405 => x"6c",
         10406 => x"20",
         10407 => x"71",
         10408 => x"20",
         10409 => x"20",
         10410 => x"25",
         10411 => x"30",
         10412 => x"48",
         10413 => x"00",
         10414 => x"20",
         10415 => x"68",
         10416 => x"65",
         10417 => x"52",
         10418 => x"43",
         10419 => x"6b",
         10420 => x"65",
         10421 => x"25",
         10422 => x"30",
         10423 => x"48",
         10424 => x"00",
         10425 => x"6c",
         10426 => x"00",
         10427 => x"69",
         10428 => x"00",
         10429 => x"78",
         10430 => x"00",
         10431 => x"00",
         10432 => x"6d",
         10433 => x"00",
         10434 => x"6e",
         10435 => x"00",
         10436 => x"6c",
         10437 => x"00",
         10438 => x"02",
         10439 => x"68",
         10440 => x"00",
         10441 => x"03",
         10442 => x"64",
         10443 => x"00",
         10444 => x"04",
         10445 => x"60",
         10446 => x"00",
         10447 => x"05",
         10448 => x"5c",
         10449 => x"00",
         10450 => x"06",
         10451 => x"58",
         10452 => x"00",
         10453 => x"07",
         10454 => x"54",
         10455 => x"00",
         10456 => x"01",
         10457 => x"50",
         10458 => x"00",
         10459 => x"08",
         10460 => x"4c",
         10461 => x"00",
         10462 => x"0b",
         10463 => x"48",
         10464 => x"00",
         10465 => x"09",
         10466 => x"44",
         10467 => x"00",
         10468 => x"0a",
         10469 => x"40",
         10470 => x"00",
         10471 => x"0d",
         10472 => x"3c",
         10473 => x"00",
         10474 => x"0c",
         10475 => x"38",
         10476 => x"00",
         10477 => x"0e",
         10478 => x"34",
         10479 => x"00",
         10480 => x"0f",
         10481 => x"30",
         10482 => x"00",
         10483 => x"0f",
         10484 => x"2c",
         10485 => x"00",
         10486 => x"10",
         10487 => x"28",
         10488 => x"00",
         10489 => x"11",
         10490 => x"24",
         10491 => x"00",
         10492 => x"12",
         10493 => x"20",
         10494 => x"00",
         10495 => x"13",
         10496 => x"1c",
         10497 => x"00",
         10498 => x"14",
         10499 => x"18",
         10500 => x"00",
         10501 => x"15",
         10502 => x"00",
         10503 => x"00",
         10504 => x"00",
         10505 => x"00",
         10506 => x"7e",
         10507 => x"7e",
         10508 => x"7e",
         10509 => x"00",
         10510 => x"7e",
         10511 => x"7e",
         10512 => x"7e",
         10513 => x"00",
         10514 => x"00",
         10515 => x"00",
         10516 => x"00",
         10517 => x"00",
         10518 => x"00",
         10519 => x"00",
         10520 => x"00",
         10521 => x"00",
         10522 => x"00",
         10523 => x"00",
         10524 => x"74",
         10525 => x"00",
         10526 => x"74",
         10527 => x"00",
         10528 => x"00",
         10529 => x"6c",
         10530 => x"25",
         10531 => x"00",
         10532 => x"6c",
         10533 => x"74",
         10534 => x"65",
         10535 => x"20",
         10536 => x"20",
         10537 => x"74",
         10538 => x"20",
         10539 => x"65",
         10540 => x"20",
         10541 => x"2e",
         10542 => x"00",
         10543 => x"6e",
         10544 => x"6f",
         10545 => x"2f",
         10546 => x"61",
         10547 => x"68",
         10548 => x"6f",
         10549 => x"66",
         10550 => x"2c",
         10551 => x"73",
         10552 => x"69",
         10553 => x"00",
         10554 => x"00",
         10555 => x"3c",
         10556 => x"7f",
         10557 => x"00",
         10558 => x"3d",
         10559 => x"00",
         10560 => x"00",
         10561 => x"33",
         10562 => x"00",
         10563 => x"4d",
         10564 => x"53",
         10565 => x"00",
         10566 => x"4e",
         10567 => x"20",
         10568 => x"46",
         10569 => x"32",
         10570 => x"00",
         10571 => x"4e",
         10572 => x"20",
         10573 => x"46",
         10574 => x"20",
         10575 => x"00",
         10576 => x"e8",
         10577 => x"00",
         10578 => x"00",
         10579 => x"00",
         10580 => x"07",
         10581 => x"12",
         10582 => x"1c",
         10583 => x"00",
         10584 => x"41",
         10585 => x"80",
         10586 => x"49",
         10587 => x"8f",
         10588 => x"4f",
         10589 => x"55",
         10590 => x"9b",
         10591 => x"9f",
         10592 => x"55",
         10593 => x"a7",
         10594 => x"ab",
         10595 => x"af",
         10596 => x"b3",
         10597 => x"b7",
         10598 => x"bb",
         10599 => x"bf",
         10600 => x"c3",
         10601 => x"c7",
         10602 => x"cb",
         10603 => x"cf",
         10604 => x"d3",
         10605 => x"d7",
         10606 => x"db",
         10607 => x"df",
         10608 => x"e3",
         10609 => x"e7",
         10610 => x"eb",
         10611 => x"ef",
         10612 => x"f3",
         10613 => x"f7",
         10614 => x"fb",
         10615 => x"ff",
         10616 => x"3b",
         10617 => x"2f",
         10618 => x"3a",
         10619 => x"7c",
         10620 => x"00",
         10621 => x"04",
         10622 => x"40",
         10623 => x"00",
         10624 => x"00",
         10625 => x"02",
         10626 => x"08",
         10627 => x"20",
         10628 => x"00",
         10629 => x"fc",
         10630 => x"e2",
         10631 => x"e0",
         10632 => x"e7",
         10633 => x"eb",
         10634 => x"ef",
         10635 => x"ec",
         10636 => x"c5",
         10637 => x"e6",
         10638 => x"f4",
         10639 => x"f2",
         10640 => x"f9",
         10641 => x"d6",
         10642 => x"a2",
         10643 => x"a5",
         10644 => x"92",
         10645 => x"ed",
         10646 => x"fa",
         10647 => x"d1",
         10648 => x"ba",
         10649 => x"10",
         10650 => x"bd",
         10651 => x"a1",
         10652 => x"bb",
         10653 => x"92",
         10654 => x"02",
         10655 => x"61",
         10656 => x"56",
         10657 => x"63",
         10658 => x"57",
         10659 => x"5c",
         10660 => x"10",
         10661 => x"34",
         10662 => x"1c",
         10663 => x"3c",
         10664 => x"5f",
         10665 => x"54",
         10666 => x"66",
         10667 => x"50",
         10668 => x"67",
         10669 => x"64",
         10670 => x"59",
         10671 => x"52",
         10672 => x"6b",
         10673 => x"18",
         10674 => x"88",
         10675 => x"8c",
         10676 => x"80",
         10677 => x"df",
         10678 => x"c0",
         10679 => x"c3",
         10680 => x"c4",
         10681 => x"98",
         10682 => x"b4",
         10683 => x"c6",
         10684 => x"29",
         10685 => x"b1",
         10686 => x"64",
         10687 => x"21",
         10688 => x"48",
         10689 => x"19",
         10690 => x"1a",
         10691 => x"b2",
         10692 => x"a0",
         10693 => x"1a",
         10694 => x"17",
         10695 => x"07",
         10696 => x"01",
         10697 => x"00",
         10698 => x"32",
         10699 => x"39",
         10700 => x"4a",
         10701 => x"79",
         10702 => x"80",
         10703 => x"43",
         10704 => x"82",
         10705 => x"84",
         10706 => x"86",
         10707 => x"87",
         10708 => x"8a",
         10709 => x"8b",
         10710 => x"8e",
         10711 => x"90",
         10712 => x"91",
         10713 => x"94",
         10714 => x"96",
         10715 => x"98",
         10716 => x"3d",
         10717 => x"9c",
         10718 => x"20",
         10719 => x"a0",
         10720 => x"a2",
         10721 => x"a4",
         10722 => x"a6",
         10723 => x"a7",
         10724 => x"aa",
         10725 => x"ac",
         10726 => x"ae",
         10727 => x"af",
         10728 => x"b2",
         10729 => x"b3",
         10730 => x"b5",
         10731 => x"b8",
         10732 => x"ba",
         10733 => x"bc",
         10734 => x"be",
         10735 => x"c0",
         10736 => x"c2",
         10737 => x"c4",
         10738 => x"c4",
         10739 => x"c8",
         10740 => x"ca",
         10741 => x"ca",
         10742 => x"10",
         10743 => x"01",
         10744 => x"de",
         10745 => x"f3",
         10746 => x"f1",
         10747 => x"f4",
         10748 => x"28",
         10749 => x"12",
         10750 => x"09",
         10751 => x"3b",
         10752 => x"3d",
         10753 => x"3f",
         10754 => x"41",
         10755 => x"46",
         10756 => x"53",
         10757 => x"81",
         10758 => x"55",
         10759 => x"8a",
         10760 => x"8f",
         10761 => x"90",
         10762 => x"5d",
         10763 => x"5f",
         10764 => x"61",
         10765 => x"94",
         10766 => x"65",
         10767 => x"67",
         10768 => x"96",
         10769 => x"62",
         10770 => x"6d",
         10771 => x"9c",
         10772 => x"71",
         10773 => x"73",
         10774 => x"9f",
         10775 => x"77",
         10776 => x"79",
         10777 => x"7b",
         10778 => x"64",
         10779 => x"7f",
         10780 => x"81",
         10781 => x"a9",
         10782 => x"85",
         10783 => x"87",
         10784 => x"44",
         10785 => x"b2",
         10786 => x"8d",
         10787 => x"8f",
         10788 => x"91",
         10789 => x"7b",
         10790 => x"fd",
         10791 => x"ff",
         10792 => x"04",
         10793 => x"88",
         10794 => x"8a",
         10795 => x"11",
         10796 => x"02",
         10797 => x"a3",
         10798 => x"08",
         10799 => x"03",
         10800 => x"8e",
         10801 => x"d8",
         10802 => x"f2",
         10803 => x"f9",
         10804 => x"f4",
         10805 => x"f6",
         10806 => x"f7",
         10807 => x"fa",
         10808 => x"30",
         10809 => x"50",
         10810 => x"60",
         10811 => x"8a",
         10812 => x"c1",
         10813 => x"cf",
         10814 => x"c0",
         10815 => x"44",
         10816 => x"26",
         10817 => x"00",
         10818 => x"01",
         10819 => x"00",
         10820 => x"a0",
         10821 => x"00",
         10822 => x"10",
         10823 => x"20",
         10824 => x"30",
         10825 => x"40",
         10826 => x"51",
         10827 => x"59",
         10828 => x"5b",
         10829 => x"5d",
         10830 => x"5f",
         10831 => x"08",
         10832 => x"0e",
         10833 => x"bb",
         10834 => x"c9",
         10835 => x"cb",
         10836 => x"db",
         10837 => x"f9",
         10838 => x"eb",
         10839 => x"fb",
         10840 => x"08",
         10841 => x"08",
         10842 => x"08",
         10843 => x"04",
         10844 => x"b9",
         10845 => x"bc",
         10846 => x"01",
         10847 => x"d0",
         10848 => x"e0",
         10849 => x"e5",
         10850 => x"ec",
         10851 => x"01",
         10852 => x"4e",
         10853 => x"32",
         10854 => x"10",
         10855 => x"01",
         10856 => x"d0",
         10857 => x"30",
         10858 => x"60",
         10859 => x"67",
         10860 => x"75",
         10861 => x"80",
         10862 => x"00",
         10863 => x"41",
         10864 => x"00",
         10865 => x"00",
         10866 => x"b8",
         10867 => x"00",
         10868 => x"00",
         10869 => x"00",
         10870 => x"c0",
         10871 => x"00",
         10872 => x"00",
         10873 => x"00",
         10874 => x"c8",
         10875 => x"00",
         10876 => x"00",
         10877 => x"00",
         10878 => x"d0",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"d8",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"e0",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"e8",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"f0",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"f8",
         10899 => x"00",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"04",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"08",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"0c",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"10",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"14",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"18",
         10927 => x"00",
         10928 => x"00",
         10929 => x"00",
         10930 => x"1c",
         10931 => x"00",
         10932 => x"00",
         10933 => x"00",
         10934 => x"24",
         10935 => x"00",
         10936 => x"00",
         10937 => x"00",
         10938 => x"28",
         10939 => x"00",
         10940 => x"00",
         10941 => x"00",
         10942 => x"30",
         10943 => x"00",
         10944 => x"00",
         10945 => x"00",
         10946 => x"38",
         10947 => x"00",
         10948 => x"00",
         10949 => x"00",
         10950 => x"40",
         10951 => x"00",
         10952 => x"00",
         10953 => x"00",
         10954 => x"48",
         10955 => x"00",
         10956 => x"00",
         10957 => x"00",
         10958 => x"50",
         10959 => x"00",
         10960 => x"00",
         10961 => x"00",
         10962 => x"58",
         10963 => x"00",
         10964 => x"00",
         10965 => x"00",
         10966 => x"60",
         10967 => x"00",
         10968 => x"00",
         10969 => x"00",
         10970 => x"00",
         10971 => x"00",
         10972 => x"ff",
         10973 => x"00",
         10974 => x"ff",
         10975 => x"00",
         10976 => x"ff",
         10977 => x"00",
         10978 => x"00",
         10979 => x"00",
         10980 => x"ff",
         10981 => x"00",
         10982 => x"00",
         10983 => x"00",
         10984 => x"00",
         10985 => x"00",
         10986 => x"00",
         10987 => x"00",
         10988 => x"00",
         10989 => x"01",
         10990 => x"01",
         10991 => x"01",
         10992 => x"00",
         10993 => x"00",
         10994 => x"00",
         10995 => x"00",
         10996 => x"00",
         10997 => x"00",
         10998 => x"00",
         10999 => x"00",
         11000 => x"00",
         11001 => x"00",
         11002 => x"00",
         11003 => x"00",
         11004 => x"00",
         11005 => x"00",
         11006 => x"00",
         11007 => x"00",
         11008 => x"00",
         11009 => x"00",
         11010 => x"00",
         11011 => x"00",
         11012 => x"00",
         11013 => x"00",
         11014 => x"00",
         11015 => x"00",
         11016 => x"00",
         11017 => x"70",
         11018 => x"00",
         11019 => x"78",
         11020 => x"00",
         11021 => x"80",
         11022 => x"00",
         11023 => x"00",
         11024 => x"00",
         11025 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"d8",
           386 => x"f9",
           387 => x"d8",
           388 => x"80",
           389 => x"d8",
           390 => x"b2",
           391 => x"d4",
           392 => x"90",
           393 => x"d4",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"84",
           400 => x"82",
           401 => x"94",
           402 => x"d8",
           403 => x"80",
           404 => x"d8",
           405 => x"c2",
           406 => x"d4",
           407 => x"90",
           408 => x"d4",
           409 => x"cc",
           410 => x"d4",
           411 => x"90",
           412 => x"d4",
           413 => x"fb",
           414 => x"d4",
           415 => x"90",
           416 => x"d4",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"84",
           423 => x"82",
           424 => x"97",
           425 => x"d8",
           426 => x"80",
           427 => x"d8",
           428 => x"fc",
           429 => x"d8",
           430 => x"80",
           431 => x"d8",
           432 => x"fd",
           433 => x"d8",
           434 => x"80",
           435 => x"d8",
           436 => x"f4",
           437 => x"d8",
           438 => x"80",
           439 => x"d8",
           440 => x"f6",
           441 => x"d8",
           442 => x"80",
           443 => x"d8",
           444 => x"f8",
           445 => x"d8",
           446 => x"80",
           447 => x"d8",
           448 => x"ee",
           449 => x"d8",
           450 => x"80",
           451 => x"d8",
           452 => x"fb",
           453 => x"d8",
           454 => x"80",
           455 => x"d8",
           456 => x"f3",
           457 => x"d8",
           458 => x"80",
           459 => x"d8",
           460 => x"f6",
           461 => x"d8",
           462 => x"80",
           463 => x"d8",
           464 => x"81",
           465 => x"d8",
           466 => x"80",
           467 => x"d8",
           468 => x"89",
           469 => x"d8",
           470 => x"80",
           471 => x"d8",
           472 => x"fa",
           473 => x"d8",
           474 => x"80",
           475 => x"d8",
           476 => x"84",
           477 => x"d8",
           478 => x"80",
           479 => x"d8",
           480 => x"85",
           481 => x"d8",
           482 => x"80",
           483 => x"d8",
           484 => x"85",
           485 => x"d8",
           486 => x"80",
           487 => x"d8",
           488 => x"8d",
           489 => x"d8",
           490 => x"80",
           491 => x"d8",
           492 => x"8b",
           493 => x"d8",
           494 => x"80",
           495 => x"d8",
           496 => x"90",
           497 => x"d8",
           498 => x"80",
           499 => x"d8",
           500 => x"86",
           501 => x"d8",
           502 => x"80",
           503 => x"d8",
           504 => x"93",
           505 => x"d8",
           506 => x"80",
           507 => x"d8",
           508 => x"94",
           509 => x"d8",
           510 => x"80",
           511 => x"d8",
           512 => x"fc",
           513 => x"d8",
           514 => x"80",
           515 => x"d8",
           516 => x"fb",
           517 => x"d8",
           518 => x"80",
           519 => x"d8",
           520 => x"fd",
           521 => x"d8",
           522 => x"80",
           523 => x"d8",
           524 => x"87",
           525 => x"d8",
           526 => x"80",
           527 => x"d8",
           528 => x"95",
           529 => x"d8",
           530 => x"80",
           531 => x"d8",
           532 => x"97",
           533 => x"d8",
           534 => x"80",
           535 => x"d8",
           536 => x"9a",
           537 => x"d8",
           538 => x"80",
           539 => x"d8",
           540 => x"ed",
           541 => x"d8",
           542 => x"80",
           543 => x"d8",
           544 => x"9d",
           545 => x"d8",
           546 => x"80",
           547 => x"d8",
           548 => x"ab",
           549 => x"d8",
           550 => x"80",
           551 => x"d8",
           552 => x"a9",
           553 => x"d8",
           554 => x"80",
           555 => x"d8",
           556 => x"ad",
           557 => x"d8",
           558 => x"80",
           559 => x"d8",
           560 => x"af",
           561 => x"d8",
           562 => x"80",
           563 => x"d8",
           564 => x"b1",
           565 => x"d8",
           566 => x"80",
           567 => x"d8",
           568 => x"f5",
           569 => x"d8",
           570 => x"80",
           571 => x"d8",
           572 => x"f6",
           573 => x"d8",
           574 => x"80",
           575 => x"d8",
           576 => x"fa",
           577 => x"d8",
           578 => x"80",
           579 => x"d8",
           580 => x"d6",
           581 => x"d8",
           582 => x"80",
           583 => x"d8",
           584 => x"a8",
           585 => x"d8",
           586 => x"80",
           587 => x"d8",
           588 => x"a8",
           589 => x"d8",
           590 => x"80",
           591 => x"d8",
           592 => x"ac",
           593 => x"d8",
           594 => x"80",
           595 => x"d8",
           596 => x"a4",
           597 => x"d8",
           598 => x"80",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"d8",
           623 => x"f4",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"d4",
           631 => x"d8",
           632 => x"3d",
           633 => x"d4",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"d4",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"d4",
           651 => x"d8",
           652 => x"82",
           653 => x"fb",
           654 => x"d8",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"d4",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"d4",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"d8",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"d8",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"d4",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"d4",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"d4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"d8",
           712 => x"05",
           713 => x"d8",
           714 => x"05",
           715 => x"d8",
           716 => x"05",
           717 => x"c8",
           718 => x"0d",
           719 => x"0c",
           720 => x"d4",
           721 => x"d8",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"d8",
           726 => x"05",
           727 => x"d4",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"d8",
           732 => x"05",
           733 => x"d4",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"c8",
           743 => x"d8",
           744 => x"05",
           745 => x"d4",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"d4",
           751 => x"08",
           752 => x"c8",
           753 => x"3d",
           754 => x"d4",
           755 => x"d8",
           756 => x"82",
           757 => x"fb",
           758 => x"d8",
           759 => x"05",
           760 => x"d4",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"d4",
           778 => x"d8",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"d8",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"d8",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"d8",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"d8",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"d8",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"d4",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"d4",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"d4",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"d8",
           848 => x"05",
           849 => x"d4",
           850 => x"33",
           851 => x"d4",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"d8",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"d8",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"d4",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"d8",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"d8",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"b0",
           901 => x"08",
           902 => x"53",
           903 => x"d8",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"d8",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"d4",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"d4",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"d4",
           927 => x"22",
           928 => x"51",
           929 => x"d8",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"d4",
           935 => x"22",
           936 => x"51",
           937 => x"d8",
           938 => x"05",
           939 => x"39",
           940 => x"d8",
           941 => x"05",
           942 => x"d4",
           943 => x"22",
           944 => x"53",
           945 => x"d4",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"d4",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"d4",
           955 => x"0c",
           956 => x"53",
           957 => x"d4",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"d8",
           965 => x"05",
           966 => x"d4",
           967 => x"08",
           968 => x"d8",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"d8",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"d4",
           987 => x"23",
           988 => x"d8",
           989 => x"05",
           990 => x"8a",
           991 => x"c8",
           992 => x"82",
           993 => x"f4",
           994 => x"d8",
           995 => x"05",
           996 => x"d8",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"d4",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"d4",
          1007 => x"0c",
          1008 => x"d8",
          1009 => x"05",
          1010 => x"d4",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"d8",
          1020 => x"05",
          1021 => x"a1",
          1022 => x"d8",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"d4",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"d8",
          1031 => x"05",
          1032 => x"d4",
          1033 => x"22",
          1034 => x"d4",
          1035 => x"22",
          1036 => x"54",
          1037 => x"d8",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"d4",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"d4",
          1050 => x"0c",
          1051 => x"d8",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"d4",
          1061 => x"0c",
          1062 => x"d4",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"d8",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"d8",
          1074 => x"05",
          1075 => x"d8",
          1076 => x"05",
          1077 => x"d4",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"d8",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"d4",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"d4",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"d4",
          1106 => x"0c",
          1107 => x"d8",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"d4",
          1117 => x"0c",
          1118 => x"d4",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"d8",
          1130 => x"05",
          1131 => x"d4",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"f3",
          1137 => x"c8",
          1138 => x"75",
          1139 => x"d4",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"d8",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"d4",
          1154 => x"34",
          1155 => x"d8",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"d4",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"d4",
          1166 => x"08",
          1167 => x"d8",
          1168 => x"05",
          1169 => x"d4",
          1170 => x"22",
          1171 => x"d8",
          1172 => x"05",
          1173 => x"a2",
          1174 => x"d8",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"d4",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"d8",
          1187 => x"05",
          1188 => x"d4",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"d8",
          1193 => x"05",
          1194 => x"51",
          1195 => x"d8",
          1196 => x"05",
          1197 => x"d4",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"d4",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"d4",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"d4",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"d4",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"d8",
          1227 => x"05",
          1228 => x"d4",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"d4",
          1245 => x"23",
          1246 => x"d8",
          1247 => x"05",
          1248 => x"d8",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"d8",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"d4",
          1266 => x"22",
          1267 => x"51",
          1268 => x"d8",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"d4",
          1278 => x"22",
          1279 => x"51",
          1280 => x"d8",
          1281 => x"05",
          1282 => x"d4",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"d4",
          1287 => x"22",
          1288 => x"54",
          1289 => x"d4",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"d4",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"d4",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"d4",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"d8",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"d4",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"d8",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"d4",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"d4",
          1338 => x"08",
          1339 => x"d4",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"d4",
          1348 => x"22",
          1349 => x"54",
          1350 => x"d4",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"d4",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"d4",
          1365 => x"33",
          1366 => x"54",
          1367 => x"d4",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"d4",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"d8",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"d4",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"d8",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"d4",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"d8",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"d4",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"d8",
          1452 => x"05",
          1453 => x"d8",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"d8",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"d8",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"d8",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"d4",
          1494 => x"23",
          1495 => x"d8",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"d4",
          1501 => x"08",
          1502 => x"d4",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"d8",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"d8",
          1513 => x"3d",
          1514 => x"d4",
          1515 => x"d8",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"f4",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"d8",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"d4",
          1531 => x"0d",
          1532 => x"d8",
          1533 => x"05",
          1534 => x"ac",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"d4",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"d4",
          1547 => x"08",
          1548 => x"d8",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"d4",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"d4",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"c8",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"d4",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"d8",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"d4",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"d4",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"d4",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"d8",
          1612 => x"05",
          1613 => x"d4",
          1614 => x"08",
          1615 => x"d4",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"d4",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"d8",
          1631 => x"3d",
          1632 => x"d4",
          1633 => x"d8",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"f4",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"c8",
          1641 => x"d8",
          1642 => x"84",
          1643 => x"d8",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"d8",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"d8",
          1665 => x"05",
          1666 => x"d4",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"d4",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"d4",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"d8",
          1702 => x"05",
          1703 => x"d8",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"d8",
          1709 => x"05",
          1710 => x"c8",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"d4",
          1714 => x"d8",
          1715 => x"3d",
          1716 => x"d4",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"d8",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"d4",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"d8",
          1756 => x"05",
          1757 => x"70",
          1758 => x"d4",
          1759 => x"0c",
          1760 => x"d8",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"d8",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"d4",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"d8",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"d8",
          1791 => x"05",
          1792 => x"d4",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"d4",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"d4",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"d4",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"d4",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"d8",
          1838 => x"05",
          1839 => x"d4",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"d8",
          1849 => x"05",
          1850 => x"d4",
          1851 => x"08",
          1852 => x"d8",
          1853 => x"05",
          1854 => x"81",
          1855 => x"d8",
          1856 => x"05",
          1857 => x"d4",
          1858 => x"08",
          1859 => x"d4",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"d8",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"d8",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"d8",
          1875 => x"05",
          1876 => x"81",
          1877 => x"d8",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"d8",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"d8",
          1886 => x"05",
          1887 => x"d4",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"d4",
          1892 => x"08",
          1893 => x"d8",
          1894 => x"05",
          1895 => x"d4",
          1896 => x"08",
          1897 => x"d8",
          1898 => x"05",
          1899 => x"d4",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"d8",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"d8",
          1909 => x"05",
          1910 => x"71",
          1911 => x"d8",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"d4",
          1917 => x"08",
          1918 => x"c8",
          1919 => x"3d",
          1920 => x"d4",
          1921 => x"d8",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"d8",
          1925 => x"05",
          1926 => x"d4",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"d8",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"d8",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"d4",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"d8",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"d4",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"d4",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"d4",
          1973 => x"08",
          1974 => x"c8",
          1975 => x"3d",
          1976 => x"d4",
          1977 => x"d8",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"d8",
          1981 => x"05",
          1982 => x"d4",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"d8",
          1988 => x"05",
          1989 => x"80",
          1990 => x"d8",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"d8",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"d8",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"d4",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"d8",
          2016 => x"05",
          2017 => x"d8",
          2018 => x"85",
          2019 => x"d8",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"d4",
          2030 => x"08",
          2031 => x"d8",
          2032 => x"05",
          2033 => x"d4",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"d8",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"d4",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"d4",
          2052 => x"08",
          2053 => x"d8",
          2054 => x"05",
          2055 => x"d4",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"d4",
          2069 => x"08",
          2070 => x"d8",
          2071 => x"05",
          2072 => x"d4",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"d4",
          2077 => x"0c",
          2078 => x"d8",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"d8",
          2092 => x"3d",
          2093 => x"d4",
          2094 => x"d8",
          2095 => x"82",
          2096 => x"fd",
          2097 => x"d8",
          2098 => x"05",
          2099 => x"d4",
          2100 => x"0c",
          2101 => x"08",
          2102 => x"8d",
          2103 => x"82",
          2104 => x"fc",
          2105 => x"ec",
          2106 => x"d4",
          2107 => x"08",
          2108 => x"82",
          2109 => x"f8",
          2110 => x"05",
          2111 => x"08",
          2112 => x"70",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"d8",
          2116 => x"05",
          2117 => x"82",
          2118 => x"8c",
          2119 => x"d8",
          2120 => x"05",
          2121 => x"84",
          2122 => x"39",
          2123 => x"08",
          2124 => x"ff",
          2125 => x"d4",
          2126 => x"0c",
          2127 => x"08",
          2128 => x"82",
          2129 => x"88",
          2130 => x"70",
          2131 => x"08",
          2132 => x"51",
          2133 => x"08",
          2134 => x"82",
          2135 => x"85",
          2136 => x"d8",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"d8",
          2143 => x"05",
          2144 => x"d4",
          2145 => x"08",
          2146 => x"d4",
          2147 => x"d4",
          2148 => x"08",
          2149 => x"d8",
          2150 => x"05",
          2151 => x"d4",
          2152 => x"08",
          2153 => x"d8",
          2154 => x"05",
          2155 => x"d4",
          2156 => x"08",
          2157 => x"38",
          2158 => x"08",
          2159 => x"51",
          2160 => x"d4",
          2161 => x"08",
          2162 => x"71",
          2163 => x"d4",
          2164 => x"08",
          2165 => x"d8",
          2166 => x"05",
          2167 => x"39",
          2168 => x"08",
          2169 => x"70",
          2170 => x"0c",
          2171 => x"0d",
          2172 => x"0c",
          2173 => x"d4",
          2174 => x"d8",
          2175 => x"3d",
          2176 => x"82",
          2177 => x"fc",
          2178 => x"d8",
          2179 => x"05",
          2180 => x"b9",
          2181 => x"d4",
          2182 => x"08",
          2183 => x"d4",
          2184 => x"0c",
          2185 => x"d8",
          2186 => x"05",
          2187 => x"d4",
          2188 => x"08",
          2189 => x"0b",
          2190 => x"08",
          2191 => x"82",
          2192 => x"f4",
          2193 => x"d8",
          2194 => x"05",
          2195 => x"d4",
          2196 => x"08",
          2197 => x"38",
          2198 => x"08",
          2199 => x"30",
          2200 => x"08",
          2201 => x"80",
          2202 => x"d4",
          2203 => x"0c",
          2204 => x"08",
          2205 => x"8a",
          2206 => x"82",
          2207 => x"f0",
          2208 => x"d8",
          2209 => x"05",
          2210 => x"d4",
          2211 => x"0c",
          2212 => x"d8",
          2213 => x"05",
          2214 => x"d8",
          2215 => x"05",
          2216 => x"c5",
          2217 => x"c8",
          2218 => x"d8",
          2219 => x"05",
          2220 => x"d8",
          2221 => x"05",
          2222 => x"90",
          2223 => x"d4",
          2224 => x"08",
          2225 => x"d4",
          2226 => x"0c",
          2227 => x"08",
          2228 => x"70",
          2229 => x"0c",
          2230 => x"0d",
          2231 => x"0c",
          2232 => x"d4",
          2233 => x"d8",
          2234 => x"3d",
          2235 => x"82",
          2236 => x"fc",
          2237 => x"d8",
          2238 => x"05",
          2239 => x"99",
          2240 => x"d4",
          2241 => x"08",
          2242 => x"d4",
          2243 => x"0c",
          2244 => x"d8",
          2245 => x"05",
          2246 => x"d4",
          2247 => x"08",
          2248 => x"38",
          2249 => x"08",
          2250 => x"30",
          2251 => x"08",
          2252 => x"81",
          2253 => x"d4",
          2254 => x"08",
          2255 => x"d4",
          2256 => x"08",
          2257 => x"3f",
          2258 => x"08",
          2259 => x"d4",
          2260 => x"0c",
          2261 => x"d4",
          2262 => x"08",
          2263 => x"38",
          2264 => x"08",
          2265 => x"30",
          2266 => x"08",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"82",
          2270 => x"54",
          2271 => x"82",
          2272 => x"04",
          2273 => x"08",
          2274 => x"d4",
          2275 => x"0d",
          2276 => x"d8",
          2277 => x"05",
          2278 => x"d8",
          2279 => x"05",
          2280 => x"c5",
          2281 => x"c8",
          2282 => x"d8",
          2283 => x"85",
          2284 => x"d8",
          2285 => x"82",
          2286 => x"02",
          2287 => x"0c",
          2288 => x"81",
          2289 => x"d4",
          2290 => x"08",
          2291 => x"d4",
          2292 => x"08",
          2293 => x"82",
          2294 => x"70",
          2295 => x"0c",
          2296 => x"0d",
          2297 => x"0c",
          2298 => x"d4",
          2299 => x"d8",
          2300 => x"3d",
          2301 => x"82",
          2302 => x"fc",
          2303 => x"0b",
          2304 => x"08",
          2305 => x"82",
          2306 => x"8c",
          2307 => x"d8",
          2308 => x"05",
          2309 => x"38",
          2310 => x"08",
          2311 => x"80",
          2312 => x"80",
          2313 => x"d4",
          2314 => x"08",
          2315 => x"82",
          2316 => x"8c",
          2317 => x"82",
          2318 => x"8c",
          2319 => x"d8",
          2320 => x"05",
          2321 => x"d8",
          2322 => x"05",
          2323 => x"39",
          2324 => x"08",
          2325 => x"80",
          2326 => x"38",
          2327 => x"08",
          2328 => x"82",
          2329 => x"88",
          2330 => x"ad",
          2331 => x"d4",
          2332 => x"08",
          2333 => x"08",
          2334 => x"31",
          2335 => x"08",
          2336 => x"82",
          2337 => x"f8",
          2338 => x"d8",
          2339 => x"05",
          2340 => x"d8",
          2341 => x"05",
          2342 => x"d4",
          2343 => x"08",
          2344 => x"d8",
          2345 => x"05",
          2346 => x"d4",
          2347 => x"08",
          2348 => x"d8",
          2349 => x"05",
          2350 => x"39",
          2351 => x"08",
          2352 => x"80",
          2353 => x"82",
          2354 => x"88",
          2355 => x"82",
          2356 => x"f4",
          2357 => x"91",
          2358 => x"d4",
          2359 => x"08",
          2360 => x"d4",
          2361 => x"0c",
          2362 => x"d4",
          2363 => x"08",
          2364 => x"0c",
          2365 => x"82",
          2366 => x"04",
          2367 => x"08",
          2368 => x"d4",
          2369 => x"0d",
          2370 => x"d8",
          2371 => x"05",
          2372 => x"d4",
          2373 => x"08",
          2374 => x"0c",
          2375 => x"08",
          2376 => x"70",
          2377 => x"72",
          2378 => x"82",
          2379 => x"f8",
          2380 => x"81",
          2381 => x"72",
          2382 => x"81",
          2383 => x"82",
          2384 => x"88",
          2385 => x"08",
          2386 => x"0c",
          2387 => x"82",
          2388 => x"f8",
          2389 => x"72",
          2390 => x"81",
          2391 => x"81",
          2392 => x"d4",
          2393 => x"34",
          2394 => x"08",
          2395 => x"70",
          2396 => x"71",
          2397 => x"51",
          2398 => x"82",
          2399 => x"f8",
          2400 => x"d8",
          2401 => x"05",
          2402 => x"b0",
          2403 => x"06",
          2404 => x"82",
          2405 => x"88",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"53",
          2409 => x"d8",
          2410 => x"05",
          2411 => x"d4",
          2412 => x"33",
          2413 => x"08",
          2414 => x"82",
          2415 => x"e8",
          2416 => x"e2",
          2417 => x"82",
          2418 => x"e8",
          2419 => x"f8",
          2420 => x"80",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"88",
          2425 => x"08",
          2426 => x"0c",
          2427 => x"53",
          2428 => x"d8",
          2429 => x"05",
          2430 => x"39",
          2431 => x"d8",
          2432 => x"05",
          2433 => x"d4",
          2434 => x"08",
          2435 => x"05",
          2436 => x"08",
          2437 => x"33",
          2438 => x"08",
          2439 => x"80",
          2440 => x"d8",
          2441 => x"05",
          2442 => x"a0",
          2443 => x"81",
          2444 => x"d4",
          2445 => x"0c",
          2446 => x"82",
          2447 => x"f8",
          2448 => x"af",
          2449 => x"38",
          2450 => x"08",
          2451 => x"53",
          2452 => x"83",
          2453 => x"80",
          2454 => x"d4",
          2455 => x"0c",
          2456 => x"88",
          2457 => x"d4",
          2458 => x"34",
          2459 => x"d8",
          2460 => x"05",
          2461 => x"73",
          2462 => x"82",
          2463 => x"f8",
          2464 => x"72",
          2465 => x"38",
          2466 => x"0b",
          2467 => x"08",
          2468 => x"82",
          2469 => x"0b",
          2470 => x"08",
          2471 => x"80",
          2472 => x"d4",
          2473 => x"0c",
          2474 => x"08",
          2475 => x"53",
          2476 => x"81",
          2477 => x"d8",
          2478 => x"05",
          2479 => x"e0",
          2480 => x"38",
          2481 => x"08",
          2482 => x"e0",
          2483 => x"72",
          2484 => x"08",
          2485 => x"82",
          2486 => x"f8",
          2487 => x"11",
          2488 => x"82",
          2489 => x"f8",
          2490 => x"d8",
          2491 => x"05",
          2492 => x"73",
          2493 => x"82",
          2494 => x"f8",
          2495 => x"11",
          2496 => x"82",
          2497 => x"f8",
          2498 => x"d8",
          2499 => x"05",
          2500 => x"89",
          2501 => x"80",
          2502 => x"d4",
          2503 => x"0c",
          2504 => x"82",
          2505 => x"f8",
          2506 => x"d8",
          2507 => x"05",
          2508 => x"72",
          2509 => x"38",
          2510 => x"d8",
          2511 => x"05",
          2512 => x"39",
          2513 => x"08",
          2514 => x"70",
          2515 => x"08",
          2516 => x"29",
          2517 => x"08",
          2518 => x"70",
          2519 => x"d4",
          2520 => x"0c",
          2521 => x"08",
          2522 => x"70",
          2523 => x"71",
          2524 => x"51",
          2525 => x"53",
          2526 => x"d8",
          2527 => x"05",
          2528 => x"39",
          2529 => x"08",
          2530 => x"53",
          2531 => x"90",
          2532 => x"d4",
          2533 => x"08",
          2534 => x"d4",
          2535 => x"0c",
          2536 => x"08",
          2537 => x"82",
          2538 => x"fc",
          2539 => x"0c",
          2540 => x"82",
          2541 => x"ec",
          2542 => x"d8",
          2543 => x"05",
          2544 => x"c8",
          2545 => x"0d",
          2546 => x"0c",
          2547 => x"d4",
          2548 => x"d8",
          2549 => x"3d",
          2550 => x"82",
          2551 => x"f0",
          2552 => x"d8",
          2553 => x"05",
          2554 => x"73",
          2555 => x"d4",
          2556 => x"08",
          2557 => x"53",
          2558 => x"72",
          2559 => x"08",
          2560 => x"72",
          2561 => x"53",
          2562 => x"09",
          2563 => x"38",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"39",
          2568 => x"08",
          2569 => x"53",
          2570 => x"09",
          2571 => x"38",
          2572 => x"d8",
          2573 => x"05",
          2574 => x"d4",
          2575 => x"08",
          2576 => x"05",
          2577 => x"08",
          2578 => x"33",
          2579 => x"08",
          2580 => x"82",
          2581 => x"f8",
          2582 => x"72",
          2583 => x"81",
          2584 => x"38",
          2585 => x"08",
          2586 => x"70",
          2587 => x"71",
          2588 => x"51",
          2589 => x"82",
          2590 => x"f8",
          2591 => x"d8",
          2592 => x"05",
          2593 => x"d4",
          2594 => x"0c",
          2595 => x"08",
          2596 => x"80",
          2597 => x"38",
          2598 => x"08",
          2599 => x"80",
          2600 => x"38",
          2601 => x"90",
          2602 => x"d4",
          2603 => x"34",
          2604 => x"08",
          2605 => x"70",
          2606 => x"71",
          2607 => x"51",
          2608 => x"82",
          2609 => x"f8",
          2610 => x"a4",
          2611 => x"82",
          2612 => x"f4",
          2613 => x"d8",
          2614 => x"05",
          2615 => x"81",
          2616 => x"70",
          2617 => x"72",
          2618 => x"d4",
          2619 => x"34",
          2620 => x"82",
          2621 => x"f8",
          2622 => x"72",
          2623 => x"38",
          2624 => x"d8",
          2625 => x"05",
          2626 => x"39",
          2627 => x"08",
          2628 => x"53",
          2629 => x"90",
          2630 => x"d4",
          2631 => x"33",
          2632 => x"26",
          2633 => x"39",
          2634 => x"d8",
          2635 => x"05",
          2636 => x"39",
          2637 => x"d8",
          2638 => x"05",
          2639 => x"82",
          2640 => x"f8",
          2641 => x"af",
          2642 => x"38",
          2643 => x"08",
          2644 => x"53",
          2645 => x"83",
          2646 => x"80",
          2647 => x"d4",
          2648 => x"0c",
          2649 => x"8a",
          2650 => x"d4",
          2651 => x"34",
          2652 => x"d8",
          2653 => x"05",
          2654 => x"d4",
          2655 => x"33",
          2656 => x"27",
          2657 => x"82",
          2658 => x"f8",
          2659 => x"80",
          2660 => x"94",
          2661 => x"d4",
          2662 => x"33",
          2663 => x"53",
          2664 => x"d4",
          2665 => x"34",
          2666 => x"08",
          2667 => x"d0",
          2668 => x"72",
          2669 => x"08",
          2670 => x"82",
          2671 => x"f8",
          2672 => x"90",
          2673 => x"38",
          2674 => x"08",
          2675 => x"f9",
          2676 => x"72",
          2677 => x"08",
          2678 => x"82",
          2679 => x"f8",
          2680 => x"72",
          2681 => x"38",
          2682 => x"d8",
          2683 => x"05",
          2684 => x"39",
          2685 => x"08",
          2686 => x"82",
          2687 => x"f4",
          2688 => x"54",
          2689 => x"8d",
          2690 => x"82",
          2691 => x"ec",
          2692 => x"f7",
          2693 => x"d4",
          2694 => x"33",
          2695 => x"d4",
          2696 => x"08",
          2697 => x"d4",
          2698 => x"33",
          2699 => x"d8",
          2700 => x"05",
          2701 => x"d4",
          2702 => x"08",
          2703 => x"05",
          2704 => x"08",
          2705 => x"55",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"a5",
          2709 => x"d4",
          2710 => x"33",
          2711 => x"2e",
          2712 => x"d8",
          2713 => x"05",
          2714 => x"d8",
          2715 => x"05",
          2716 => x"d4",
          2717 => x"08",
          2718 => x"08",
          2719 => x"71",
          2720 => x"0b",
          2721 => x"08",
          2722 => x"82",
          2723 => x"ec",
          2724 => x"d8",
          2725 => x"3d",
          2726 => x"d4",
          2727 => x"3d",
          2728 => x"08",
          2729 => x"58",
          2730 => x"80",
          2731 => x"39",
          2732 => x"e6",
          2733 => x"d8",
          2734 => x"78",
          2735 => x"33",
          2736 => x"39",
          2737 => x"73",
          2738 => x"81",
          2739 => x"81",
          2740 => x"39",
          2741 => x"90",
          2742 => x"c8",
          2743 => x"52",
          2744 => x"3f",
          2745 => x"08",
          2746 => x"75",
          2747 => x"a3",
          2748 => x"c8",
          2749 => x"84",
          2750 => x"73",
          2751 => x"b0",
          2752 => x"70",
          2753 => x"58",
          2754 => x"27",
          2755 => x"54",
          2756 => x"c8",
          2757 => x"0d",
          2758 => x"0d",
          2759 => x"93",
          2760 => x"38",
          2761 => x"82",
          2762 => x"52",
          2763 => x"82",
          2764 => x"81",
          2765 => x"b4",
          2766 => x"f9",
          2767 => x"80",
          2768 => x"39",
          2769 => x"51",
          2770 => x"82",
          2771 => x"80",
          2772 => x"b5",
          2773 => x"dd",
          2774 => x"c4",
          2775 => x"39",
          2776 => x"51",
          2777 => x"82",
          2778 => x"80",
          2779 => x"b6",
          2780 => x"c1",
          2781 => x"9c",
          2782 => x"82",
          2783 => x"b5",
          2784 => x"cc",
          2785 => x"82",
          2786 => x"a9",
          2787 => x"84",
          2788 => x"82",
          2789 => x"9d",
          2790 => x"b4",
          2791 => x"82",
          2792 => x"91",
          2793 => x"e4",
          2794 => x"82",
          2795 => x"85",
          2796 => x"88",
          2797 => x"3f",
          2798 => x"04",
          2799 => x"77",
          2800 => x"74",
          2801 => x"8a",
          2802 => x"75",
          2803 => x"51",
          2804 => x"e8",
          2805 => x"ef",
          2806 => x"d8",
          2807 => x"75",
          2808 => x"3f",
          2809 => x"08",
          2810 => x"75",
          2811 => x"98",
          2812 => x"e5",
          2813 => x"0d",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"33",
          2817 => x"68",
          2818 => x"7a",
          2819 => x"51",
          2820 => x"78",
          2821 => x"ff",
          2822 => x"81",
          2823 => x"07",
          2824 => x"06",
          2825 => x"56",
          2826 => x"38",
          2827 => x"52",
          2828 => x"52",
          2829 => x"90",
          2830 => x"c8",
          2831 => x"d8",
          2832 => x"38",
          2833 => x"08",
          2834 => x"88",
          2835 => x"c8",
          2836 => x"3d",
          2837 => x"84",
          2838 => x"52",
          2839 => x"9a",
          2840 => x"d8",
          2841 => x"82",
          2842 => x"90",
          2843 => x"74",
          2844 => x"38",
          2845 => x"19",
          2846 => x"39",
          2847 => x"05",
          2848 => x"c3",
          2849 => x"70",
          2850 => x"25",
          2851 => x"9f",
          2852 => x"51",
          2853 => x"74",
          2854 => x"38",
          2855 => x"53",
          2856 => x"88",
          2857 => x"51",
          2858 => x"76",
          2859 => x"d8",
          2860 => x"3d",
          2861 => x"3d",
          2862 => x"84",
          2863 => x"33",
          2864 => x"59",
          2865 => x"52",
          2866 => x"ad",
          2867 => x"c8",
          2868 => x"38",
          2869 => x"88",
          2870 => x"2e",
          2871 => x"39",
          2872 => x"57",
          2873 => x"56",
          2874 => x"55",
          2875 => x"08",
          2876 => x"ac",
          2877 => x"f4",
          2878 => x"82",
          2879 => x"ff",
          2880 => x"82",
          2881 => x"62",
          2882 => x"82",
          2883 => x"60",
          2884 => x"79",
          2885 => x"c8",
          2886 => x"39",
          2887 => x"82",
          2888 => x"8b",
          2889 => x"f3",
          2890 => x"61",
          2891 => x"05",
          2892 => x"33",
          2893 => x"68",
          2894 => x"5c",
          2895 => x"7a",
          2896 => x"f8",
          2897 => x"91",
          2898 => x"80",
          2899 => x"89",
          2900 => x"74",
          2901 => x"80",
          2902 => x"2e",
          2903 => x"a0",
          2904 => x"80",
          2905 => x"18",
          2906 => x"27",
          2907 => x"22",
          2908 => x"84",
          2909 => x"e1",
          2910 => x"82",
          2911 => x"ff",
          2912 => x"82",
          2913 => x"c3",
          2914 => x"53",
          2915 => x"8e",
          2916 => x"52",
          2917 => x"51",
          2918 => x"3f",
          2919 => x"b9",
          2920 => x"b8",
          2921 => x"15",
          2922 => x"74",
          2923 => x"7a",
          2924 => x"72",
          2925 => x"b9",
          2926 => x"b8",
          2927 => x"39",
          2928 => x"51",
          2929 => x"3f",
          2930 => x"82",
          2931 => x"52",
          2932 => x"df",
          2933 => x"39",
          2934 => x"51",
          2935 => x"3f",
          2936 => x"79",
          2937 => x"38",
          2938 => x"33",
          2939 => x"56",
          2940 => x"83",
          2941 => x"80",
          2942 => x"27",
          2943 => x"53",
          2944 => x"70",
          2945 => x"51",
          2946 => x"2e",
          2947 => x"80",
          2948 => x"38",
          2949 => x"08",
          2950 => x"88",
          2951 => x"ac",
          2952 => x"51",
          2953 => x"81",
          2954 => x"b6",
          2955 => x"a8",
          2956 => x"3f",
          2957 => x"1c",
          2958 => x"80",
          2959 => x"c8",
          2960 => x"70",
          2961 => x"57",
          2962 => x"09",
          2963 => x"38",
          2964 => x"82",
          2965 => x"98",
          2966 => x"2c",
          2967 => x"70",
          2968 => x"32",
          2969 => x"72",
          2970 => x"07",
          2971 => x"58",
          2972 => x"57",
          2973 => x"d8",
          2974 => x"2e",
          2975 => x"85",
          2976 => x"8c",
          2977 => x"53",
          2978 => x"fd",
          2979 => x"53",
          2980 => x"c8",
          2981 => x"0d",
          2982 => x"0d",
          2983 => x"33",
          2984 => x"53",
          2985 => x"52",
          2986 => x"ad",
          2987 => x"a0",
          2988 => x"d9",
          2989 => x"c0",
          2990 => x"cc",
          2991 => x"a1",
          2992 => x"b9",
          2993 => x"b6",
          2994 => x"80",
          2995 => x"a5",
          2996 => x"3d",
          2997 => x"3d",
          2998 => x"96",
          2999 => x"aa",
          3000 => x"51",
          3001 => x"82",
          3002 => x"9d",
          3003 => x"51",
          3004 => x"72",
          3005 => x"81",
          3006 => x"71",
          3007 => x"38",
          3008 => x"a5",
          3009 => x"88",
          3010 => x"3f",
          3011 => x"99",
          3012 => x"2a",
          3013 => x"51",
          3014 => x"2e",
          3015 => x"51",
          3016 => x"82",
          3017 => x"9d",
          3018 => x"51",
          3019 => x"72",
          3020 => x"81",
          3021 => x"71",
          3022 => x"38",
          3023 => x"e9",
          3024 => x"a8",
          3025 => x"3f",
          3026 => x"dd",
          3027 => x"2a",
          3028 => x"51",
          3029 => x"2e",
          3030 => x"51",
          3031 => x"82",
          3032 => x"9c",
          3033 => x"51",
          3034 => x"72",
          3035 => x"81",
          3036 => x"71",
          3037 => x"38",
          3038 => x"ad",
          3039 => x"d0",
          3040 => x"3f",
          3041 => x"a1",
          3042 => x"2a",
          3043 => x"51",
          3044 => x"2e",
          3045 => x"51",
          3046 => x"82",
          3047 => x"9c",
          3048 => x"51",
          3049 => x"72",
          3050 => x"81",
          3051 => x"71",
          3052 => x"38",
          3053 => x"f1",
          3054 => x"f8",
          3055 => x"3f",
          3056 => x"e5",
          3057 => x"2a",
          3058 => x"51",
          3059 => x"2e",
          3060 => x"51",
          3061 => x"82",
          3062 => x"9b",
          3063 => x"51",
          3064 => x"a8",
          3065 => x"3d",
          3066 => x"3d",
          3067 => x"84",
          3068 => x"33",
          3069 => x"56",
          3070 => x"51",
          3071 => x"0b",
          3072 => x"c4",
          3073 => x"a9",
          3074 => x"82",
          3075 => x"82",
          3076 => x"81",
          3077 => x"82",
          3078 => x"30",
          3079 => x"c8",
          3080 => x"25",
          3081 => x"51",
          3082 => x"0b",
          3083 => x"c4",
          3084 => x"82",
          3085 => x"54",
          3086 => x"09",
          3087 => x"38",
          3088 => x"53",
          3089 => x"51",
          3090 => x"3f",
          3091 => x"08",
          3092 => x"38",
          3093 => x"08",
          3094 => x"3f",
          3095 => x"ef",
          3096 => x"9a",
          3097 => x"0b",
          3098 => x"d3",
          3099 => x"0b",
          3100 => x"33",
          3101 => x"2e",
          3102 => x"8c",
          3103 => x"d8",
          3104 => x"75",
          3105 => x"3f",
          3106 => x"d8",
          3107 => x"3d",
          3108 => x"3d",
          3109 => x"71",
          3110 => x"0c",
          3111 => x"52",
          3112 => x"cb",
          3113 => x"d8",
          3114 => x"ff",
          3115 => x"7d",
          3116 => x"06",
          3117 => x"3d",
          3118 => x"82",
          3119 => x"78",
          3120 => x"3f",
          3121 => x"52",
          3122 => x"51",
          3123 => x"3f",
          3124 => x"08",
          3125 => x"38",
          3126 => x"51",
          3127 => x"81",
          3128 => x"82",
          3129 => x"ff",
          3130 => x"96",
          3131 => x"5a",
          3132 => x"79",
          3133 => x"3f",
          3134 => x"84",
          3135 => x"9e",
          3136 => x"c8",
          3137 => x"70",
          3138 => x"59",
          3139 => x"2e",
          3140 => x"78",
          3141 => x"80",
          3142 => x"ab",
          3143 => x"38",
          3144 => x"a4",
          3145 => x"2e",
          3146 => x"78",
          3147 => x"38",
          3148 => x"ff",
          3149 => x"82",
          3150 => x"2e",
          3151 => x"78",
          3152 => x"ad",
          3153 => x"39",
          3154 => x"84",
          3155 => x"bd",
          3156 => x"78",
          3157 => x"a6",
          3158 => x"2e",
          3159 => x"8e",
          3160 => x"bf",
          3161 => x"38",
          3162 => x"2e",
          3163 => x"8e",
          3164 => x"80",
          3165 => x"a2",
          3166 => x"d5",
          3167 => x"78",
          3168 => x"8c",
          3169 => x"80",
          3170 => x"38",
          3171 => x"2e",
          3172 => x"78",
          3173 => x"8b",
          3174 => x"9e",
          3175 => x"d1",
          3176 => x"38",
          3177 => x"2e",
          3178 => x"8e",
          3179 => x"81",
          3180 => x"e4",
          3181 => x"82",
          3182 => x"78",
          3183 => x"8c",
          3184 => x"80",
          3185 => x"93",
          3186 => x"39",
          3187 => x"2e",
          3188 => x"78",
          3189 => x"8d",
          3190 => x"de",
          3191 => x"ff",
          3192 => x"ff",
          3193 => x"eb",
          3194 => x"d8",
          3195 => x"38",
          3196 => x"51",
          3197 => x"b4",
          3198 => x"11",
          3199 => x"05",
          3200 => x"3f",
          3201 => x"08",
          3202 => x"38",
          3203 => x"83",
          3204 => x"02",
          3205 => x"33",
          3206 => x"cf",
          3207 => x"80",
          3208 => x"82",
          3209 => x"81",
          3210 => x"78",
          3211 => x"bc",
          3212 => x"b0",
          3213 => x"fd",
          3214 => x"bc",
          3215 => x"f5",
          3216 => x"ff",
          3217 => x"ff",
          3218 => x"eb",
          3219 => x"d8",
          3220 => x"2e",
          3221 => x"80",
          3222 => x"02",
          3223 => x"33",
          3224 => x"d9",
          3225 => x"c8",
          3226 => x"bc",
          3227 => x"a1",
          3228 => x"ff",
          3229 => x"ff",
          3230 => x"ea",
          3231 => x"d8",
          3232 => x"2e",
          3233 => x"89",
          3234 => x"38",
          3235 => x"fc",
          3236 => x"84",
          3237 => x"b5",
          3238 => x"c8",
          3239 => x"82",
          3240 => x"43",
          3241 => x"bc",
          3242 => x"51",
          3243 => x"3f",
          3244 => x"05",
          3245 => x"52",
          3246 => x"29",
          3247 => x"05",
          3248 => x"a3",
          3249 => x"c8",
          3250 => x"38",
          3251 => x"51",
          3252 => x"81",
          3253 => x"39",
          3254 => x"84",
          3255 => x"c2",
          3256 => x"c8",
          3257 => x"ff",
          3258 => x"5b",
          3259 => x"81",
          3260 => x"c8",
          3261 => x"51",
          3262 => x"80",
          3263 => x"3d",
          3264 => x"51",
          3265 => x"82",
          3266 => x"b5",
          3267 => x"05",
          3268 => x"b2",
          3269 => x"c8",
          3270 => x"ff",
          3271 => x"5a",
          3272 => x"82",
          3273 => x"b5",
          3274 => x"05",
          3275 => x"96",
          3276 => x"ec",
          3277 => x"f8",
          3278 => x"80",
          3279 => x"c8",
          3280 => x"06",
          3281 => x"79",
          3282 => x"f2",
          3283 => x"d8",
          3284 => x"2e",
          3285 => x"82",
          3286 => x"51",
          3287 => x"fb",
          3288 => x"3d",
          3289 => x"53",
          3290 => x"51",
          3291 => x"82",
          3292 => x"80",
          3293 => x"38",
          3294 => x"fc",
          3295 => x"84",
          3296 => x"c9",
          3297 => x"c8",
          3298 => x"fa",
          3299 => x"3d",
          3300 => x"53",
          3301 => x"51",
          3302 => x"82",
          3303 => x"86",
          3304 => x"c8",
          3305 => x"bc",
          3306 => x"ac",
          3307 => x"63",
          3308 => x"7b",
          3309 => x"38",
          3310 => x"7a",
          3311 => x"5c",
          3312 => x"26",
          3313 => x"db",
          3314 => x"ff",
          3315 => x"ff",
          3316 => x"e7",
          3317 => x"d8",
          3318 => x"2e",
          3319 => x"b4",
          3320 => x"11",
          3321 => x"05",
          3322 => x"3f",
          3323 => x"08",
          3324 => x"ef",
          3325 => x"fe",
          3326 => x"ff",
          3327 => x"e7",
          3328 => x"d8",
          3329 => x"2e",
          3330 => x"82",
          3331 => x"ff",
          3332 => x"63",
          3333 => x"27",
          3334 => x"61",
          3335 => x"81",
          3336 => x"79",
          3337 => x"05",
          3338 => x"b4",
          3339 => x"11",
          3340 => x"05",
          3341 => x"3f",
          3342 => x"08",
          3343 => x"a3",
          3344 => x"fe",
          3345 => x"ff",
          3346 => x"e7",
          3347 => x"d8",
          3348 => x"2e",
          3349 => x"b4",
          3350 => x"11",
          3351 => x"05",
          3352 => x"3f",
          3353 => x"08",
          3354 => x"f7",
          3355 => x"84",
          3356 => x"e5",
          3357 => x"79",
          3358 => x"38",
          3359 => x"7b",
          3360 => x"5b",
          3361 => x"92",
          3362 => x"7a",
          3363 => x"53",
          3364 => x"bd",
          3365 => x"aa",
          3366 => x"1a",
          3367 => x"43",
          3368 => x"8a",
          3369 => x"3f",
          3370 => x"b4",
          3371 => x"11",
          3372 => x"05",
          3373 => x"3f",
          3374 => x"08",
          3375 => x"82",
          3376 => x"59",
          3377 => x"89",
          3378 => x"ec",
          3379 => x"cd",
          3380 => x"b5",
          3381 => x"80",
          3382 => x"82",
          3383 => x"44",
          3384 => x"d7",
          3385 => x"78",
          3386 => x"38",
          3387 => x"08",
          3388 => x"82",
          3389 => x"59",
          3390 => x"88",
          3391 => x"84",
          3392 => x"39",
          3393 => x"33",
          3394 => x"2e",
          3395 => x"d7",
          3396 => x"89",
          3397 => x"9c",
          3398 => x"05",
          3399 => x"fe",
          3400 => x"ff",
          3401 => x"e5",
          3402 => x"d8",
          3403 => x"de",
          3404 => x"b4",
          3405 => x"80",
          3406 => x"82",
          3407 => x"43",
          3408 => x"82",
          3409 => x"59",
          3410 => x"88",
          3411 => x"f8",
          3412 => x"39",
          3413 => x"33",
          3414 => x"2e",
          3415 => x"d7",
          3416 => x"aa",
          3417 => x"b7",
          3418 => x"80",
          3419 => x"82",
          3420 => x"43",
          3421 => x"d7",
          3422 => x"78",
          3423 => x"38",
          3424 => x"08",
          3425 => x"82",
          3426 => x"88",
          3427 => x"3d",
          3428 => x"53",
          3429 => x"51",
          3430 => x"82",
          3431 => x"80",
          3432 => x"80",
          3433 => x"7a",
          3434 => x"38",
          3435 => x"90",
          3436 => x"70",
          3437 => x"2a",
          3438 => x"51",
          3439 => x"78",
          3440 => x"38",
          3441 => x"83",
          3442 => x"82",
          3443 => x"c4",
          3444 => x"55",
          3445 => x"53",
          3446 => x"51",
          3447 => x"82",
          3448 => x"87",
          3449 => x"3d",
          3450 => x"53",
          3451 => x"51",
          3452 => x"82",
          3453 => x"80",
          3454 => x"38",
          3455 => x"fc",
          3456 => x"84",
          3457 => x"c5",
          3458 => x"c8",
          3459 => x"a4",
          3460 => x"02",
          3461 => x"33",
          3462 => x"81",
          3463 => x"3d",
          3464 => x"53",
          3465 => x"51",
          3466 => x"82",
          3467 => x"e1",
          3468 => x"39",
          3469 => x"54",
          3470 => x"c8",
          3471 => x"99",
          3472 => x"a8",
          3473 => x"f8",
          3474 => x"ff",
          3475 => x"79",
          3476 => x"59",
          3477 => x"f5",
          3478 => x"79",
          3479 => x"b4",
          3480 => x"11",
          3481 => x"05",
          3482 => x"3f",
          3483 => x"08",
          3484 => x"38",
          3485 => x"80",
          3486 => x"79",
          3487 => x"05",
          3488 => x"39",
          3489 => x"51",
          3490 => x"ff",
          3491 => x"3d",
          3492 => x"53",
          3493 => x"51",
          3494 => x"82",
          3495 => x"80",
          3496 => x"38",
          3497 => x"f0",
          3498 => x"84",
          3499 => x"cc",
          3500 => x"c8",
          3501 => x"a5",
          3502 => x"02",
          3503 => x"79",
          3504 => x"5b",
          3505 => x"b4",
          3506 => x"11",
          3507 => x"05",
          3508 => x"3f",
          3509 => x"08",
          3510 => x"87",
          3511 => x"22",
          3512 => x"bd",
          3513 => x"a5",
          3514 => x"f4",
          3515 => x"80",
          3516 => x"51",
          3517 => x"3f",
          3518 => x"33",
          3519 => x"2e",
          3520 => x"78",
          3521 => x"38",
          3522 => x"41",
          3523 => x"3d",
          3524 => x"53",
          3525 => x"51",
          3526 => x"82",
          3527 => x"80",
          3528 => x"60",
          3529 => x"05",
          3530 => x"82",
          3531 => x"78",
          3532 => x"39",
          3533 => x"51",
          3534 => x"ff",
          3535 => x"3d",
          3536 => x"53",
          3537 => x"51",
          3538 => x"82",
          3539 => x"80",
          3540 => x"38",
          3541 => x"f0",
          3542 => x"84",
          3543 => x"9c",
          3544 => x"c8",
          3545 => x"a0",
          3546 => x"71",
          3547 => x"84",
          3548 => x"3d",
          3549 => x"53",
          3550 => x"51",
          3551 => x"82",
          3552 => x"e5",
          3553 => x"39",
          3554 => x"54",
          3555 => x"e4",
          3556 => x"c5",
          3557 => x"a8",
          3558 => x"f8",
          3559 => x"ff",
          3560 => x"79",
          3561 => x"59",
          3562 => x"f2",
          3563 => x"79",
          3564 => x"b4",
          3565 => x"11",
          3566 => x"05",
          3567 => x"3f",
          3568 => x"08",
          3569 => x"38",
          3570 => x"0c",
          3571 => x"05",
          3572 => x"39",
          3573 => x"51",
          3574 => x"ff",
          3575 => x"bd",
          3576 => x"80",
          3577 => x"98",
          3578 => x"f7",
          3579 => x"8c",
          3580 => x"f0",
          3581 => x"97",
          3582 => x"e7",
          3583 => x"a0",
          3584 => x"e0",
          3585 => x"81",
          3586 => x"94",
          3587 => x"80",
          3588 => x"c0",
          3589 => x"f1",
          3590 => x"be",
          3591 => x"bf",
          3592 => x"80",
          3593 => x"c0",
          3594 => x"8c",
          3595 => x"87",
          3596 => x"0c",
          3597 => x"b4",
          3598 => x"11",
          3599 => x"05",
          3600 => x"3f",
          3601 => x"08",
          3602 => x"97",
          3603 => x"82",
          3604 => x"ff",
          3605 => x"63",
          3606 => x"b4",
          3607 => x"11",
          3608 => x"05",
          3609 => x"3f",
          3610 => x"08",
          3611 => x"f3",
          3612 => x"82",
          3613 => x"ff",
          3614 => x"63",
          3615 => x"82",
          3616 => x"80",
          3617 => x"38",
          3618 => x"08",
          3619 => x"80",
          3620 => x"c5",
          3621 => x"39",
          3622 => x"51",
          3623 => x"3f",
          3624 => x"3f",
          3625 => x"82",
          3626 => x"ff",
          3627 => x"80",
          3628 => x"39",
          3629 => x"f0",
          3630 => x"45",
          3631 => x"78",
          3632 => x"9f",
          3633 => x"06",
          3634 => x"2e",
          3635 => x"b4",
          3636 => x"05",
          3637 => x"3f",
          3638 => x"08",
          3639 => x"7b",
          3640 => x"38",
          3641 => x"89",
          3642 => x"2e",
          3643 => x"ca",
          3644 => x"2e",
          3645 => x"c2",
          3646 => x"cc",
          3647 => x"82",
          3648 => x"80",
          3649 => x"d4",
          3650 => x"ff",
          3651 => x"ff",
          3652 => x"b8",
          3653 => x"b4",
          3654 => x"05",
          3655 => x"3f",
          3656 => x"55",
          3657 => x"54",
          3658 => x"bf",
          3659 => x"3d",
          3660 => x"51",
          3661 => x"3f",
          3662 => x"54",
          3663 => x"bf",
          3664 => x"3d",
          3665 => x"51",
          3666 => x"3f",
          3667 => x"58",
          3668 => x"57",
          3669 => x"55",
          3670 => x"80",
          3671 => x"80",
          3672 => x"3d",
          3673 => x"51",
          3674 => x"82",
          3675 => x"82",
          3676 => x"09",
          3677 => x"72",
          3678 => x"51",
          3679 => x"80",
          3680 => x"26",
          3681 => x"5a",
          3682 => x"59",
          3683 => x"8d",
          3684 => x"70",
          3685 => x"5d",
          3686 => x"c3",
          3687 => x"32",
          3688 => x"07",
          3689 => x"38",
          3690 => x"09",
          3691 => x"b3",
          3692 => x"f8",
          3693 => x"ac",
          3694 => x"39",
          3695 => x"80",
          3696 => x"f8",
          3697 => x"94",
          3698 => x"54",
          3699 => x"80",
          3700 => x"d3",
          3701 => x"d8",
          3702 => x"2b",
          3703 => x"53",
          3704 => x"52",
          3705 => x"9c",
          3706 => x"d8",
          3707 => x"75",
          3708 => x"94",
          3709 => x"54",
          3710 => x"80",
          3711 => x"d3",
          3712 => x"d8",
          3713 => x"2b",
          3714 => x"53",
          3715 => x"52",
          3716 => x"f0",
          3717 => x"d8",
          3718 => x"75",
          3719 => x"83",
          3720 => x"94",
          3721 => x"80",
          3722 => x"c0",
          3723 => x"80",
          3724 => x"80",
          3725 => x"83",
          3726 => x"99",
          3727 => x"5c",
          3728 => x"0b",
          3729 => x"88",
          3730 => x"72",
          3731 => x"ac",
          3732 => x"be",
          3733 => x"3f",
          3734 => x"51",
          3735 => x"3f",
          3736 => x"51",
          3737 => x"3f",
          3738 => x"51",
          3739 => x"81",
          3740 => x"3f",
          3741 => x"80",
          3742 => x"0d",
          3743 => x"53",
          3744 => x"52",
          3745 => x"82",
          3746 => x"81",
          3747 => x"07",
          3748 => x"52",
          3749 => x"e8",
          3750 => x"d8",
          3751 => x"3d",
          3752 => x"3d",
          3753 => x"08",
          3754 => x"73",
          3755 => x"74",
          3756 => x"38",
          3757 => x"70",
          3758 => x"81",
          3759 => x"81",
          3760 => x"39",
          3761 => x"70",
          3762 => x"81",
          3763 => x"81",
          3764 => x"54",
          3765 => x"81",
          3766 => x"06",
          3767 => x"39",
          3768 => x"80",
          3769 => x"54",
          3770 => x"83",
          3771 => x"70",
          3772 => x"38",
          3773 => x"98",
          3774 => x"52",
          3775 => x"52",
          3776 => x"2e",
          3777 => x"54",
          3778 => x"84",
          3779 => x"38",
          3780 => x"52",
          3781 => x"2e",
          3782 => x"83",
          3783 => x"70",
          3784 => x"30",
          3785 => x"76",
          3786 => x"51",
          3787 => x"88",
          3788 => x"70",
          3789 => x"34",
          3790 => x"72",
          3791 => x"d8",
          3792 => x"3d",
          3793 => x"3d",
          3794 => x"72",
          3795 => x"91",
          3796 => x"fc",
          3797 => x"51",
          3798 => x"82",
          3799 => x"85",
          3800 => x"83",
          3801 => x"72",
          3802 => x"0c",
          3803 => x"04",
          3804 => x"76",
          3805 => x"ff",
          3806 => x"81",
          3807 => x"26",
          3808 => x"83",
          3809 => x"05",
          3810 => x"70",
          3811 => x"8a",
          3812 => x"33",
          3813 => x"70",
          3814 => x"fe",
          3815 => x"33",
          3816 => x"70",
          3817 => x"f2",
          3818 => x"33",
          3819 => x"70",
          3820 => x"e6",
          3821 => x"22",
          3822 => x"74",
          3823 => x"80",
          3824 => x"13",
          3825 => x"52",
          3826 => x"26",
          3827 => x"81",
          3828 => x"98",
          3829 => x"22",
          3830 => x"bc",
          3831 => x"33",
          3832 => x"b8",
          3833 => x"33",
          3834 => x"b4",
          3835 => x"33",
          3836 => x"b0",
          3837 => x"33",
          3838 => x"ac",
          3839 => x"33",
          3840 => x"a8",
          3841 => x"c0",
          3842 => x"73",
          3843 => x"a0",
          3844 => x"87",
          3845 => x"0c",
          3846 => x"82",
          3847 => x"86",
          3848 => x"f3",
          3849 => x"5b",
          3850 => x"9c",
          3851 => x"0c",
          3852 => x"bc",
          3853 => x"7b",
          3854 => x"98",
          3855 => x"79",
          3856 => x"87",
          3857 => x"08",
          3858 => x"1c",
          3859 => x"98",
          3860 => x"79",
          3861 => x"87",
          3862 => x"08",
          3863 => x"1c",
          3864 => x"98",
          3865 => x"79",
          3866 => x"87",
          3867 => x"08",
          3868 => x"1c",
          3869 => x"98",
          3870 => x"79",
          3871 => x"80",
          3872 => x"83",
          3873 => x"59",
          3874 => x"ff",
          3875 => x"1b",
          3876 => x"1b",
          3877 => x"1b",
          3878 => x"1b",
          3879 => x"1b",
          3880 => x"83",
          3881 => x"52",
          3882 => x"51",
          3883 => x"3f",
          3884 => x"04",
          3885 => x"02",
          3886 => x"82",
          3887 => x"70",
          3888 => x"58",
          3889 => x"c0",
          3890 => x"75",
          3891 => x"38",
          3892 => x"94",
          3893 => x"70",
          3894 => x"81",
          3895 => x"52",
          3896 => x"8c",
          3897 => x"2a",
          3898 => x"51",
          3899 => x"38",
          3900 => x"70",
          3901 => x"51",
          3902 => x"8d",
          3903 => x"2a",
          3904 => x"51",
          3905 => x"be",
          3906 => x"ff",
          3907 => x"c0",
          3908 => x"70",
          3909 => x"38",
          3910 => x"90",
          3911 => x"0c",
          3912 => x"c8",
          3913 => x"0d",
          3914 => x"0d",
          3915 => x"33",
          3916 => x"9f",
          3917 => x"52",
          3918 => x"e8",
          3919 => x"0d",
          3920 => x"0d",
          3921 => x"33",
          3922 => x"2e",
          3923 => x"87",
          3924 => x"8d",
          3925 => x"82",
          3926 => x"70",
          3927 => x"58",
          3928 => x"94",
          3929 => x"80",
          3930 => x"87",
          3931 => x"53",
          3932 => x"96",
          3933 => x"06",
          3934 => x"72",
          3935 => x"38",
          3936 => x"70",
          3937 => x"53",
          3938 => x"74",
          3939 => x"81",
          3940 => x"72",
          3941 => x"38",
          3942 => x"70",
          3943 => x"53",
          3944 => x"38",
          3945 => x"06",
          3946 => x"94",
          3947 => x"80",
          3948 => x"87",
          3949 => x"54",
          3950 => x"80",
          3951 => x"c8",
          3952 => x"0d",
          3953 => x"0d",
          3954 => x"74",
          3955 => x"ff",
          3956 => x"57",
          3957 => x"80",
          3958 => x"81",
          3959 => x"15",
          3960 => x"33",
          3961 => x"06",
          3962 => x"58",
          3963 => x"84",
          3964 => x"2e",
          3965 => x"c0",
          3966 => x"70",
          3967 => x"2a",
          3968 => x"53",
          3969 => x"80",
          3970 => x"71",
          3971 => x"81",
          3972 => x"70",
          3973 => x"81",
          3974 => x"06",
          3975 => x"80",
          3976 => x"71",
          3977 => x"81",
          3978 => x"70",
          3979 => x"74",
          3980 => x"51",
          3981 => x"80",
          3982 => x"2e",
          3983 => x"c0",
          3984 => x"77",
          3985 => x"17",
          3986 => x"81",
          3987 => x"53",
          3988 => x"86",
          3989 => x"d8",
          3990 => x"3d",
          3991 => x"3d",
          3992 => x"e8",
          3993 => x"ff",
          3994 => x"87",
          3995 => x"51",
          3996 => x"86",
          3997 => x"94",
          3998 => x"08",
          3999 => x"70",
          4000 => x"51",
          4001 => x"2e",
          4002 => x"81",
          4003 => x"87",
          4004 => x"52",
          4005 => x"86",
          4006 => x"94",
          4007 => x"08",
          4008 => x"06",
          4009 => x"0c",
          4010 => x"0d",
          4011 => x"3f",
          4012 => x"08",
          4013 => x"82",
          4014 => x"04",
          4015 => x"82",
          4016 => x"70",
          4017 => x"52",
          4018 => x"94",
          4019 => x"80",
          4020 => x"87",
          4021 => x"52",
          4022 => x"82",
          4023 => x"06",
          4024 => x"ff",
          4025 => x"2e",
          4026 => x"81",
          4027 => x"87",
          4028 => x"52",
          4029 => x"86",
          4030 => x"94",
          4031 => x"08",
          4032 => x"70",
          4033 => x"53",
          4034 => x"d8",
          4035 => x"3d",
          4036 => x"3d",
          4037 => x"9e",
          4038 => x"9c",
          4039 => x"51",
          4040 => x"2e",
          4041 => x"87",
          4042 => x"08",
          4043 => x"0c",
          4044 => x"a8",
          4045 => x"f0",
          4046 => x"9e",
          4047 => x"d6",
          4048 => x"c0",
          4049 => x"82",
          4050 => x"87",
          4051 => x"08",
          4052 => x"0c",
          4053 => x"a0",
          4054 => x"80",
          4055 => x"9e",
          4056 => x"d7",
          4057 => x"c0",
          4058 => x"82",
          4059 => x"87",
          4060 => x"08",
          4061 => x"0c",
          4062 => x"b8",
          4063 => x"90",
          4064 => x"9e",
          4065 => x"d7",
          4066 => x"c0",
          4067 => x"82",
          4068 => x"87",
          4069 => x"08",
          4070 => x"0c",
          4071 => x"80",
          4072 => x"82",
          4073 => x"87",
          4074 => x"08",
          4075 => x"0c",
          4076 => x"88",
          4077 => x"a8",
          4078 => x"9e",
          4079 => x"d7",
          4080 => x"0b",
          4081 => x"34",
          4082 => x"c0",
          4083 => x"70",
          4084 => x"06",
          4085 => x"70",
          4086 => x"38",
          4087 => x"82",
          4088 => x"80",
          4089 => x"9e",
          4090 => x"88",
          4091 => x"51",
          4092 => x"80",
          4093 => x"81",
          4094 => x"d7",
          4095 => x"0b",
          4096 => x"90",
          4097 => x"80",
          4098 => x"52",
          4099 => x"2e",
          4100 => x"52",
          4101 => x"b3",
          4102 => x"87",
          4103 => x"08",
          4104 => x"80",
          4105 => x"52",
          4106 => x"83",
          4107 => x"71",
          4108 => x"34",
          4109 => x"c0",
          4110 => x"70",
          4111 => x"06",
          4112 => x"70",
          4113 => x"38",
          4114 => x"82",
          4115 => x"80",
          4116 => x"9e",
          4117 => x"90",
          4118 => x"51",
          4119 => x"80",
          4120 => x"81",
          4121 => x"d7",
          4122 => x"0b",
          4123 => x"90",
          4124 => x"80",
          4125 => x"52",
          4126 => x"2e",
          4127 => x"52",
          4128 => x"b7",
          4129 => x"87",
          4130 => x"08",
          4131 => x"80",
          4132 => x"52",
          4133 => x"83",
          4134 => x"71",
          4135 => x"34",
          4136 => x"c0",
          4137 => x"70",
          4138 => x"06",
          4139 => x"70",
          4140 => x"38",
          4141 => x"82",
          4142 => x"80",
          4143 => x"9e",
          4144 => x"80",
          4145 => x"51",
          4146 => x"80",
          4147 => x"81",
          4148 => x"d7",
          4149 => x"0b",
          4150 => x"90",
          4151 => x"80",
          4152 => x"52",
          4153 => x"83",
          4154 => x"71",
          4155 => x"34",
          4156 => x"90",
          4157 => x"80",
          4158 => x"2a",
          4159 => x"70",
          4160 => x"34",
          4161 => x"c0",
          4162 => x"70",
          4163 => x"51",
          4164 => x"80",
          4165 => x"81",
          4166 => x"d7",
          4167 => x"c0",
          4168 => x"70",
          4169 => x"70",
          4170 => x"51",
          4171 => x"d7",
          4172 => x"0b",
          4173 => x"90",
          4174 => x"06",
          4175 => x"70",
          4176 => x"38",
          4177 => x"82",
          4178 => x"87",
          4179 => x"08",
          4180 => x"51",
          4181 => x"d7",
          4182 => x"3d",
          4183 => x"3d",
          4184 => x"c4",
          4185 => x"f1",
          4186 => x"b0",
          4187 => x"80",
          4188 => x"82",
          4189 => x"ff",
          4190 => x"82",
          4191 => x"ff",
          4192 => x"82",
          4193 => x"54",
          4194 => x"94",
          4195 => x"8c",
          4196 => x"90",
          4197 => x"52",
          4198 => x"51",
          4199 => x"3f",
          4200 => x"33",
          4201 => x"2e",
          4202 => x"d7",
          4203 => x"d7",
          4204 => x"54",
          4205 => x"a0",
          4206 => x"9d",
          4207 => x"b4",
          4208 => x"80",
          4209 => x"82",
          4210 => x"82",
          4211 => x"11",
          4212 => x"c1",
          4213 => x"90",
          4214 => x"d7",
          4215 => x"73",
          4216 => x"38",
          4217 => x"08",
          4218 => x"08",
          4219 => x"82",
          4220 => x"ff",
          4221 => x"82",
          4222 => x"54",
          4223 => x"94",
          4224 => x"fc",
          4225 => x"80",
          4226 => x"52",
          4227 => x"51",
          4228 => x"3f",
          4229 => x"33",
          4230 => x"2e",
          4231 => x"d7",
          4232 => x"82",
          4233 => x"ff",
          4234 => x"82",
          4235 => x"54",
          4236 => x"8e",
          4237 => x"c0",
          4238 => x"c2",
          4239 => x"8f",
          4240 => x"d7",
          4241 => x"73",
          4242 => x"38",
          4243 => x"33",
          4244 => x"d0",
          4245 => x"81",
          4246 => x"b1",
          4247 => x"80",
          4248 => x"82",
          4249 => x"ff",
          4250 => x"82",
          4251 => x"54",
          4252 => x"89",
          4253 => x"84",
          4254 => x"e8",
          4255 => x"b8",
          4256 => x"80",
          4257 => x"82",
          4258 => x"ff",
          4259 => x"82",
          4260 => x"54",
          4261 => x"89",
          4262 => x"9c",
          4263 => x"c4",
          4264 => x"ba",
          4265 => x"80",
          4266 => x"82",
          4267 => x"ff",
          4268 => x"82",
          4269 => x"ff",
          4270 => x"82",
          4271 => x"52",
          4272 => x"51",
          4273 => x"3f",
          4274 => x"08",
          4275 => x"e0",
          4276 => x"85",
          4277 => x"9c",
          4278 => x"c4",
          4279 => x"8d",
          4280 => x"c4",
          4281 => x"a9",
          4282 => x"d7",
          4283 => x"82",
          4284 => x"ff",
          4285 => x"82",
          4286 => x"56",
          4287 => x"52",
          4288 => x"80",
          4289 => x"c8",
          4290 => x"c0",
          4291 => x"31",
          4292 => x"d8",
          4293 => x"82",
          4294 => x"ff",
          4295 => x"82",
          4296 => x"54",
          4297 => x"a9",
          4298 => x"a8",
          4299 => x"84",
          4300 => x"51",
          4301 => x"82",
          4302 => x"bd",
          4303 => x"76",
          4304 => x"54",
          4305 => x"08",
          4306 => x"8c",
          4307 => x"89",
          4308 => x"b2",
          4309 => x"80",
          4310 => x"82",
          4311 => x"56",
          4312 => x"52",
          4313 => x"9c",
          4314 => x"c8",
          4315 => x"c0",
          4316 => x"31",
          4317 => x"d8",
          4318 => x"82",
          4319 => x"ff",
          4320 => x"8a",
          4321 => x"fe",
          4322 => x"0d",
          4323 => x"0d",
          4324 => x"33",
          4325 => x"71",
          4326 => x"38",
          4327 => x"82",
          4328 => x"52",
          4329 => x"82",
          4330 => x"9d",
          4331 => x"ec",
          4332 => x"82",
          4333 => x"91",
          4334 => x"fc",
          4335 => x"82",
          4336 => x"85",
          4337 => x"88",
          4338 => x"8d",
          4339 => x"0d",
          4340 => x"80",
          4341 => x"3d",
          4342 => x"96",
          4343 => x"52",
          4344 => x"0c",
          4345 => x"70",
          4346 => x"0c",
          4347 => x"3d",
          4348 => x"3d",
          4349 => x"96",
          4350 => x"82",
          4351 => x"52",
          4352 => x"73",
          4353 => x"d7",
          4354 => x"70",
          4355 => x"0c",
          4356 => x"83",
          4357 => x"80",
          4358 => x"96",
          4359 => x"82",
          4360 => x"87",
          4361 => x"0c",
          4362 => x"0d",
          4363 => x"70",
          4364 => x"98",
          4365 => x"2c",
          4366 => x"70",
          4367 => x"53",
          4368 => x"51",
          4369 => x"c6",
          4370 => x"55",
          4371 => x"25",
          4372 => x"c6",
          4373 => x"12",
          4374 => x"97",
          4375 => x"33",
          4376 => x"70",
          4377 => x"81",
          4378 => x"81",
          4379 => x"d8",
          4380 => x"3d",
          4381 => x"3d",
          4382 => x"84",
          4383 => x"33",
          4384 => x"56",
          4385 => x"2e",
          4386 => x"f4",
          4387 => x"88",
          4388 => x"9f",
          4389 => x"ac",
          4390 => x"51",
          4391 => x"3f",
          4392 => x"08",
          4393 => x"ff",
          4394 => x"73",
          4395 => x"53",
          4396 => x"72",
          4397 => x"53",
          4398 => x"51",
          4399 => x"3f",
          4400 => x"87",
          4401 => x"f6",
          4402 => x"02",
          4403 => x"05",
          4404 => x"05",
          4405 => x"82",
          4406 => x"70",
          4407 => x"d7",
          4408 => x"08",
          4409 => x"5a",
          4410 => x"80",
          4411 => x"74",
          4412 => x"3f",
          4413 => x"33",
          4414 => x"82",
          4415 => x"81",
          4416 => x"58",
          4417 => x"fb",
          4418 => x"c8",
          4419 => x"82",
          4420 => x"70",
          4421 => x"d7",
          4422 => x"08",
          4423 => x"74",
          4424 => x"38",
          4425 => x"52",
          4426 => x"b3",
          4427 => x"d8",
          4428 => x"05",
          4429 => x"d8",
          4430 => x"81",
          4431 => x"93",
          4432 => x"38",
          4433 => x"d8",
          4434 => x"80",
          4435 => x"82",
          4436 => x"56",
          4437 => x"ac",
          4438 => x"98",
          4439 => x"a4",
          4440 => x"fc",
          4441 => x"53",
          4442 => x"51",
          4443 => x"3f",
          4444 => x"08",
          4445 => x"81",
          4446 => x"82",
          4447 => x"51",
          4448 => x"3f",
          4449 => x"04",
          4450 => x"82",
          4451 => x"93",
          4452 => x"52",
          4453 => x"89",
          4454 => x"99",
          4455 => x"73",
          4456 => x"84",
          4457 => x"73",
          4458 => x"38",
          4459 => x"d8",
          4460 => x"d8",
          4461 => x"71",
          4462 => x"38",
          4463 => x"f0",
          4464 => x"d8",
          4465 => x"99",
          4466 => x"0b",
          4467 => x"0c",
          4468 => x"04",
          4469 => x"81",
          4470 => x"82",
          4471 => x"51",
          4472 => x"3f",
          4473 => x"08",
          4474 => x"82",
          4475 => x"53",
          4476 => x"88",
          4477 => x"56",
          4478 => x"3f",
          4479 => x"08",
          4480 => x"38",
          4481 => x"af",
          4482 => x"d8",
          4483 => x"80",
          4484 => x"c8",
          4485 => x"38",
          4486 => x"08",
          4487 => x"17",
          4488 => x"74",
          4489 => x"76",
          4490 => x"82",
          4491 => x"57",
          4492 => x"3f",
          4493 => x"09",
          4494 => x"af",
          4495 => x"0d",
          4496 => x"0d",
          4497 => x"ad",
          4498 => x"5a",
          4499 => x"58",
          4500 => x"d8",
          4501 => x"80",
          4502 => x"82",
          4503 => x"81",
          4504 => x"0b",
          4505 => x"08",
          4506 => x"f8",
          4507 => x"70",
          4508 => x"9c",
          4509 => x"d8",
          4510 => x"2e",
          4511 => x"51",
          4512 => x"3f",
          4513 => x"08",
          4514 => x"55",
          4515 => x"d8",
          4516 => x"8e",
          4517 => x"c8",
          4518 => x"70",
          4519 => x"80",
          4520 => x"09",
          4521 => x"72",
          4522 => x"51",
          4523 => x"77",
          4524 => x"73",
          4525 => x"82",
          4526 => x"8c",
          4527 => x"51",
          4528 => x"3f",
          4529 => x"08",
          4530 => x"38",
          4531 => x"51",
          4532 => x"3f",
          4533 => x"09",
          4534 => x"38",
          4535 => x"51",
          4536 => x"3f",
          4537 => x"ae",
          4538 => x"3d",
          4539 => x"d8",
          4540 => x"34",
          4541 => x"82",
          4542 => x"a9",
          4543 => x"f6",
          4544 => x"7e",
          4545 => x"72",
          4546 => x"5a",
          4547 => x"2e",
          4548 => x"a2",
          4549 => x"78",
          4550 => x"76",
          4551 => x"81",
          4552 => x"70",
          4553 => x"58",
          4554 => x"2e",
          4555 => x"86",
          4556 => x"26",
          4557 => x"54",
          4558 => x"82",
          4559 => x"70",
          4560 => x"ff",
          4561 => x"82",
          4562 => x"53",
          4563 => x"08",
          4564 => x"bf",
          4565 => x"c8",
          4566 => x"38",
          4567 => x"55",
          4568 => x"88",
          4569 => x"2e",
          4570 => x"39",
          4571 => x"ac",
          4572 => x"5a",
          4573 => x"11",
          4574 => x"51",
          4575 => x"82",
          4576 => x"80",
          4577 => x"ff",
          4578 => x"52",
          4579 => x"b1",
          4580 => x"c8",
          4581 => x"06",
          4582 => x"38",
          4583 => x"39",
          4584 => x"81",
          4585 => x"54",
          4586 => x"ff",
          4587 => x"54",
          4588 => x"c8",
          4589 => x"0d",
          4590 => x"0d",
          4591 => x"b2",
          4592 => x"3d",
          4593 => x"5a",
          4594 => x"3d",
          4595 => x"a0",
          4596 => x"9c",
          4597 => x"73",
          4598 => x"73",
          4599 => x"33",
          4600 => x"83",
          4601 => x"76",
          4602 => x"bc",
          4603 => x"76",
          4604 => x"73",
          4605 => x"ad",
          4606 => x"98",
          4607 => x"d8",
          4608 => x"d8",
          4609 => x"d8",
          4610 => x"2e",
          4611 => x"93",
          4612 => x"82",
          4613 => x"51",
          4614 => x"3f",
          4615 => x"08",
          4616 => x"38",
          4617 => x"51",
          4618 => x"3f",
          4619 => x"82",
          4620 => x"5b",
          4621 => x"08",
          4622 => x"52",
          4623 => x"52",
          4624 => x"89",
          4625 => x"c8",
          4626 => x"d8",
          4627 => x"2e",
          4628 => x"80",
          4629 => x"d8",
          4630 => x"ff",
          4631 => x"82",
          4632 => x"55",
          4633 => x"d8",
          4634 => x"a9",
          4635 => x"c8",
          4636 => x"70",
          4637 => x"80",
          4638 => x"53",
          4639 => x"06",
          4640 => x"f8",
          4641 => x"1b",
          4642 => x"06",
          4643 => x"7b",
          4644 => x"80",
          4645 => x"2e",
          4646 => x"ff",
          4647 => x"39",
          4648 => x"98",
          4649 => x"38",
          4650 => x"08",
          4651 => x"38",
          4652 => x"8f",
          4653 => x"84",
          4654 => x"c8",
          4655 => x"70",
          4656 => x"59",
          4657 => x"ee",
          4658 => x"ff",
          4659 => x"84",
          4660 => x"2b",
          4661 => x"82",
          4662 => x"70",
          4663 => x"97",
          4664 => x"2c",
          4665 => x"29",
          4666 => x"05",
          4667 => x"70",
          4668 => x"51",
          4669 => x"51",
          4670 => x"81",
          4671 => x"2e",
          4672 => x"77",
          4673 => x"38",
          4674 => x"0a",
          4675 => x"0a",
          4676 => x"2c",
          4677 => x"75",
          4678 => x"38",
          4679 => x"52",
          4680 => x"85",
          4681 => x"c8",
          4682 => x"06",
          4683 => x"2e",
          4684 => x"82",
          4685 => x"81",
          4686 => x"74",
          4687 => x"29",
          4688 => x"05",
          4689 => x"70",
          4690 => x"56",
          4691 => x"95",
          4692 => x"76",
          4693 => x"77",
          4694 => x"3f",
          4695 => x"08",
          4696 => x"54",
          4697 => x"d3",
          4698 => x"75",
          4699 => x"ca",
          4700 => x"55",
          4701 => x"84",
          4702 => x"2b",
          4703 => x"82",
          4704 => x"70",
          4705 => x"98",
          4706 => x"11",
          4707 => x"82",
          4708 => x"33",
          4709 => x"51",
          4710 => x"55",
          4711 => x"09",
          4712 => x"92",
          4713 => x"98",
          4714 => x"0c",
          4715 => x"f0",
          4716 => x"0b",
          4717 => x"34",
          4718 => x"82",
          4719 => x"75",
          4720 => x"34",
          4721 => x"34",
          4722 => x"7e",
          4723 => x"26",
          4724 => x"73",
          4725 => x"af",
          4726 => x"73",
          4727 => x"f0",
          4728 => x"73",
          4729 => x"cb",
          4730 => x"88",
          4731 => x"75",
          4732 => x"74",
          4733 => x"98",
          4734 => x"73",
          4735 => x"38",
          4736 => x"73",
          4737 => x"34",
          4738 => x"0a",
          4739 => x"0a",
          4740 => x"2c",
          4741 => x"33",
          4742 => x"df",
          4743 => x"8c",
          4744 => x"56",
          4745 => x"f0",
          4746 => x"1a",
          4747 => x"33",
          4748 => x"f0",
          4749 => x"73",
          4750 => x"38",
          4751 => x"73",
          4752 => x"34",
          4753 => x"33",
          4754 => x"0a",
          4755 => x"0a",
          4756 => x"2c",
          4757 => x"33",
          4758 => x"56",
          4759 => x"a8",
          4760 => x"ac",
          4761 => x"1a",
          4762 => x"54",
          4763 => x"3f",
          4764 => x"0a",
          4765 => x"0a",
          4766 => x"2c",
          4767 => x"33",
          4768 => x"73",
          4769 => x"38",
          4770 => x"33",
          4771 => x"70",
          4772 => x"f0",
          4773 => x"51",
          4774 => x"77",
          4775 => x"38",
          4776 => x"08",
          4777 => x"ff",
          4778 => x"74",
          4779 => x"29",
          4780 => x"05",
          4781 => x"82",
          4782 => x"56",
          4783 => x"75",
          4784 => x"fb",
          4785 => x"7a",
          4786 => x"81",
          4787 => x"f0",
          4788 => x"52",
          4789 => x"51",
          4790 => x"81",
          4791 => x"f0",
          4792 => x"81",
          4793 => x"55",
          4794 => x"fb",
          4795 => x"f0",
          4796 => x"05",
          4797 => x"f0",
          4798 => x"15",
          4799 => x"f0",
          4800 => x"f4",
          4801 => x"88",
          4802 => x"a7",
          4803 => x"8c",
          4804 => x"2b",
          4805 => x"82",
          4806 => x"57",
          4807 => x"74",
          4808 => x"38",
          4809 => x"81",
          4810 => x"34",
          4811 => x"08",
          4812 => x"51",
          4813 => x"3f",
          4814 => x"0a",
          4815 => x"0a",
          4816 => x"2c",
          4817 => x"33",
          4818 => x"75",
          4819 => x"38",
          4820 => x"08",
          4821 => x"ff",
          4822 => x"82",
          4823 => x"70",
          4824 => x"98",
          4825 => x"88",
          4826 => x"56",
          4827 => x"24",
          4828 => x"82",
          4829 => x"52",
          4830 => x"9c",
          4831 => x"81",
          4832 => x"81",
          4833 => x"70",
          4834 => x"f0",
          4835 => x"51",
          4836 => x"25",
          4837 => x"9b",
          4838 => x"88",
          4839 => x"54",
          4840 => x"82",
          4841 => x"52",
          4842 => x"9c",
          4843 => x"f0",
          4844 => x"51",
          4845 => x"82",
          4846 => x"81",
          4847 => x"73",
          4848 => x"f0",
          4849 => x"73",
          4850 => x"38",
          4851 => x"52",
          4852 => x"f3",
          4853 => x"80",
          4854 => x"0b",
          4855 => x"34",
          4856 => x"f0",
          4857 => x"82",
          4858 => x"af",
          4859 => x"82",
          4860 => x"54",
          4861 => x"f9",
          4862 => x"f4",
          4863 => x"88",
          4864 => x"af",
          4865 => x"8c",
          4866 => x"54",
          4867 => x"8c",
          4868 => x"ff",
          4869 => x"39",
          4870 => x"33",
          4871 => x"33",
          4872 => x"75",
          4873 => x"38",
          4874 => x"73",
          4875 => x"34",
          4876 => x"70",
          4877 => x"81",
          4878 => x"51",
          4879 => x"25",
          4880 => x"1a",
          4881 => x"33",
          4882 => x"f4",
          4883 => x"73",
          4884 => x"9a",
          4885 => x"81",
          4886 => x"81",
          4887 => x"70",
          4888 => x"f0",
          4889 => x"51",
          4890 => x"24",
          4891 => x"f4",
          4892 => x"a0",
          4893 => x"bb",
          4894 => x"8c",
          4895 => x"2b",
          4896 => x"82",
          4897 => x"57",
          4898 => x"74",
          4899 => x"a3",
          4900 => x"ac",
          4901 => x"51",
          4902 => x"3f",
          4903 => x"0a",
          4904 => x"0a",
          4905 => x"2c",
          4906 => x"33",
          4907 => x"75",
          4908 => x"38",
          4909 => x"82",
          4910 => x"70",
          4911 => x"82",
          4912 => x"59",
          4913 => x"77",
          4914 => x"38",
          4915 => x"08",
          4916 => x"54",
          4917 => x"8c",
          4918 => x"70",
          4919 => x"ff",
          4920 => x"82",
          4921 => x"70",
          4922 => x"82",
          4923 => x"58",
          4924 => x"75",
          4925 => x"f7",
          4926 => x"f0",
          4927 => x"52",
          4928 => x"51",
          4929 => x"80",
          4930 => x"8c",
          4931 => x"82",
          4932 => x"f7",
          4933 => x"b0",
          4934 => x"94",
          4935 => x"80",
          4936 => x"74",
          4937 => x"de",
          4938 => x"c8",
          4939 => x"88",
          4940 => x"c8",
          4941 => x"06",
          4942 => x"74",
          4943 => x"ff",
          4944 => x"93",
          4945 => x"39",
          4946 => x"82",
          4947 => x"fc",
          4948 => x"54",
          4949 => x"a7",
          4950 => x"ff",
          4951 => x"82",
          4952 => x"82",
          4953 => x"82",
          4954 => x"81",
          4955 => x"05",
          4956 => x"79",
          4957 => x"ee",
          4958 => x"54",
          4959 => x"73",
          4960 => x"80",
          4961 => x"38",
          4962 => x"a0",
          4963 => x"39",
          4964 => x"09",
          4965 => x"38",
          4966 => x"08",
          4967 => x"2e",
          4968 => x"51",
          4969 => x"3f",
          4970 => x"08",
          4971 => x"34",
          4972 => x"08",
          4973 => x"81",
          4974 => x"52",
          4975 => x"a2",
          4976 => x"c3",
          4977 => x"29",
          4978 => x"05",
          4979 => x"54",
          4980 => x"ab",
          4981 => x"ff",
          4982 => x"82",
          4983 => x"82",
          4984 => x"82",
          4985 => x"81",
          4986 => x"05",
          4987 => x"79",
          4988 => x"f2",
          4989 => x"54",
          4990 => x"06",
          4991 => x"74",
          4992 => x"34",
          4993 => x"82",
          4994 => x"82",
          4995 => x"52",
          4996 => x"e2",
          4997 => x"39",
          4998 => x"33",
          4999 => x"06",
          5000 => x"33",
          5001 => x"74",
          5002 => x"87",
          5003 => x"ac",
          5004 => x"14",
          5005 => x"f0",
          5006 => x"1a",
          5007 => x"54",
          5008 => x"3f",
          5009 => x"82",
          5010 => x"54",
          5011 => x"f4",
          5012 => x"f4",
          5013 => x"88",
          5014 => x"d7",
          5015 => x"8c",
          5016 => x"54",
          5017 => x"8c",
          5018 => x"39",
          5019 => x"83",
          5020 => x"82",
          5021 => x"84",
          5022 => x"d8",
          5023 => x"80",
          5024 => x"83",
          5025 => x"ff",
          5026 => x"82",
          5027 => x"54",
          5028 => x"74",
          5029 => x"76",
          5030 => x"82",
          5031 => x"54",
          5032 => x"34",
          5033 => x"34",
          5034 => x"08",
          5035 => x"15",
          5036 => x"15",
          5037 => x"c0",
          5038 => x"bc",
          5039 => x"fe",
          5040 => x"70",
          5041 => x"06",
          5042 => x"58",
          5043 => x"74",
          5044 => x"73",
          5045 => x"82",
          5046 => x"70",
          5047 => x"d8",
          5048 => x"f8",
          5049 => x"55",
          5050 => x"34",
          5051 => x"34",
          5052 => x"04",
          5053 => x"73",
          5054 => x"84",
          5055 => x"38",
          5056 => x"2a",
          5057 => x"83",
          5058 => x"51",
          5059 => x"82",
          5060 => x"83",
          5061 => x"f9",
          5062 => x"a6",
          5063 => x"84",
          5064 => x"22",
          5065 => x"d8",
          5066 => x"83",
          5067 => x"74",
          5068 => x"11",
          5069 => x"12",
          5070 => x"2b",
          5071 => x"05",
          5072 => x"71",
          5073 => x"06",
          5074 => x"2a",
          5075 => x"59",
          5076 => x"57",
          5077 => x"71",
          5078 => x"81",
          5079 => x"d8",
          5080 => x"75",
          5081 => x"54",
          5082 => x"34",
          5083 => x"34",
          5084 => x"08",
          5085 => x"33",
          5086 => x"71",
          5087 => x"70",
          5088 => x"ff",
          5089 => x"52",
          5090 => x"05",
          5091 => x"ff",
          5092 => x"2a",
          5093 => x"71",
          5094 => x"72",
          5095 => x"53",
          5096 => x"34",
          5097 => x"08",
          5098 => x"76",
          5099 => x"17",
          5100 => x"0d",
          5101 => x"0d",
          5102 => x"08",
          5103 => x"9e",
          5104 => x"83",
          5105 => x"86",
          5106 => x"12",
          5107 => x"2b",
          5108 => x"07",
          5109 => x"52",
          5110 => x"05",
          5111 => x"85",
          5112 => x"88",
          5113 => x"88",
          5114 => x"56",
          5115 => x"13",
          5116 => x"13",
          5117 => x"c0",
          5118 => x"84",
          5119 => x"12",
          5120 => x"2b",
          5121 => x"07",
          5122 => x"52",
          5123 => x"12",
          5124 => x"33",
          5125 => x"07",
          5126 => x"54",
          5127 => x"70",
          5128 => x"73",
          5129 => x"82",
          5130 => x"13",
          5131 => x"12",
          5132 => x"2b",
          5133 => x"ff",
          5134 => x"88",
          5135 => x"53",
          5136 => x"73",
          5137 => x"14",
          5138 => x"0d",
          5139 => x"0d",
          5140 => x"22",
          5141 => x"08",
          5142 => x"71",
          5143 => x"81",
          5144 => x"88",
          5145 => x"88",
          5146 => x"33",
          5147 => x"71",
          5148 => x"90",
          5149 => x"5f",
          5150 => x"5a",
          5151 => x"54",
          5152 => x"80",
          5153 => x"51",
          5154 => x"82",
          5155 => x"70",
          5156 => x"81",
          5157 => x"8b",
          5158 => x"2b",
          5159 => x"70",
          5160 => x"33",
          5161 => x"07",
          5162 => x"8f",
          5163 => x"51",
          5164 => x"53",
          5165 => x"72",
          5166 => x"2a",
          5167 => x"82",
          5168 => x"83",
          5169 => x"d8",
          5170 => x"16",
          5171 => x"12",
          5172 => x"2b",
          5173 => x"07",
          5174 => x"55",
          5175 => x"33",
          5176 => x"71",
          5177 => x"70",
          5178 => x"06",
          5179 => x"57",
          5180 => x"52",
          5181 => x"71",
          5182 => x"88",
          5183 => x"fb",
          5184 => x"d8",
          5185 => x"84",
          5186 => x"22",
          5187 => x"72",
          5188 => x"33",
          5189 => x"71",
          5190 => x"83",
          5191 => x"5b",
          5192 => x"52",
          5193 => x"33",
          5194 => x"71",
          5195 => x"02",
          5196 => x"05",
          5197 => x"70",
          5198 => x"51",
          5199 => x"71",
          5200 => x"81",
          5201 => x"d8",
          5202 => x"15",
          5203 => x"12",
          5204 => x"2b",
          5205 => x"07",
          5206 => x"52",
          5207 => x"12",
          5208 => x"33",
          5209 => x"07",
          5210 => x"54",
          5211 => x"70",
          5212 => x"72",
          5213 => x"82",
          5214 => x"14",
          5215 => x"83",
          5216 => x"88",
          5217 => x"d8",
          5218 => x"54",
          5219 => x"04",
          5220 => x"7b",
          5221 => x"08",
          5222 => x"70",
          5223 => x"06",
          5224 => x"53",
          5225 => x"82",
          5226 => x"76",
          5227 => x"11",
          5228 => x"83",
          5229 => x"8b",
          5230 => x"2b",
          5231 => x"70",
          5232 => x"33",
          5233 => x"71",
          5234 => x"53",
          5235 => x"53",
          5236 => x"59",
          5237 => x"25",
          5238 => x"80",
          5239 => x"51",
          5240 => x"81",
          5241 => x"14",
          5242 => x"33",
          5243 => x"71",
          5244 => x"76",
          5245 => x"2a",
          5246 => x"58",
          5247 => x"14",
          5248 => x"ff",
          5249 => x"87",
          5250 => x"d8",
          5251 => x"19",
          5252 => x"85",
          5253 => x"88",
          5254 => x"88",
          5255 => x"5b",
          5256 => x"84",
          5257 => x"85",
          5258 => x"d8",
          5259 => x"53",
          5260 => x"14",
          5261 => x"87",
          5262 => x"d8",
          5263 => x"76",
          5264 => x"75",
          5265 => x"82",
          5266 => x"18",
          5267 => x"12",
          5268 => x"2b",
          5269 => x"80",
          5270 => x"88",
          5271 => x"55",
          5272 => x"74",
          5273 => x"15",
          5274 => x"0d",
          5275 => x"0d",
          5276 => x"d8",
          5277 => x"38",
          5278 => x"71",
          5279 => x"38",
          5280 => x"8c",
          5281 => x"0d",
          5282 => x"0d",
          5283 => x"58",
          5284 => x"82",
          5285 => x"83",
          5286 => x"82",
          5287 => x"84",
          5288 => x"12",
          5289 => x"2b",
          5290 => x"59",
          5291 => x"81",
          5292 => x"75",
          5293 => x"cb",
          5294 => x"29",
          5295 => x"81",
          5296 => x"88",
          5297 => x"81",
          5298 => x"79",
          5299 => x"ff",
          5300 => x"7f",
          5301 => x"51",
          5302 => x"77",
          5303 => x"38",
          5304 => x"85",
          5305 => x"5a",
          5306 => x"33",
          5307 => x"71",
          5308 => x"57",
          5309 => x"38",
          5310 => x"ff",
          5311 => x"7a",
          5312 => x"80",
          5313 => x"82",
          5314 => x"11",
          5315 => x"12",
          5316 => x"2b",
          5317 => x"ff",
          5318 => x"52",
          5319 => x"55",
          5320 => x"83",
          5321 => x"80",
          5322 => x"26",
          5323 => x"74",
          5324 => x"2e",
          5325 => x"77",
          5326 => x"81",
          5327 => x"75",
          5328 => x"3f",
          5329 => x"82",
          5330 => x"79",
          5331 => x"f7",
          5332 => x"d8",
          5333 => x"1c",
          5334 => x"87",
          5335 => x"8b",
          5336 => x"2b",
          5337 => x"5e",
          5338 => x"7a",
          5339 => x"ff",
          5340 => x"88",
          5341 => x"56",
          5342 => x"15",
          5343 => x"ff",
          5344 => x"85",
          5345 => x"d8",
          5346 => x"83",
          5347 => x"72",
          5348 => x"33",
          5349 => x"71",
          5350 => x"70",
          5351 => x"5b",
          5352 => x"56",
          5353 => x"19",
          5354 => x"19",
          5355 => x"c0",
          5356 => x"84",
          5357 => x"12",
          5358 => x"2b",
          5359 => x"07",
          5360 => x"55",
          5361 => x"78",
          5362 => x"76",
          5363 => x"82",
          5364 => x"70",
          5365 => x"84",
          5366 => x"12",
          5367 => x"2b",
          5368 => x"2a",
          5369 => x"52",
          5370 => x"84",
          5371 => x"85",
          5372 => x"d8",
          5373 => x"84",
          5374 => x"82",
          5375 => x"8d",
          5376 => x"fe",
          5377 => x"52",
          5378 => x"08",
          5379 => x"dc",
          5380 => x"71",
          5381 => x"38",
          5382 => x"ed",
          5383 => x"c8",
          5384 => x"82",
          5385 => x"84",
          5386 => x"ee",
          5387 => x"66",
          5388 => x"70",
          5389 => x"d8",
          5390 => x"2e",
          5391 => x"84",
          5392 => x"3f",
          5393 => x"7e",
          5394 => x"3f",
          5395 => x"08",
          5396 => x"39",
          5397 => x"7b",
          5398 => x"3f",
          5399 => x"ba",
          5400 => x"f5",
          5401 => x"d8",
          5402 => x"ff",
          5403 => x"d8",
          5404 => x"71",
          5405 => x"70",
          5406 => x"06",
          5407 => x"73",
          5408 => x"81",
          5409 => x"88",
          5410 => x"75",
          5411 => x"ff",
          5412 => x"88",
          5413 => x"73",
          5414 => x"70",
          5415 => x"33",
          5416 => x"07",
          5417 => x"53",
          5418 => x"48",
          5419 => x"54",
          5420 => x"56",
          5421 => x"80",
          5422 => x"76",
          5423 => x"06",
          5424 => x"83",
          5425 => x"42",
          5426 => x"33",
          5427 => x"71",
          5428 => x"70",
          5429 => x"70",
          5430 => x"33",
          5431 => x"71",
          5432 => x"53",
          5433 => x"56",
          5434 => x"25",
          5435 => x"75",
          5436 => x"ff",
          5437 => x"54",
          5438 => x"81",
          5439 => x"18",
          5440 => x"2e",
          5441 => x"8f",
          5442 => x"f6",
          5443 => x"83",
          5444 => x"58",
          5445 => x"7f",
          5446 => x"74",
          5447 => x"78",
          5448 => x"3f",
          5449 => x"7f",
          5450 => x"75",
          5451 => x"38",
          5452 => x"11",
          5453 => x"33",
          5454 => x"07",
          5455 => x"f4",
          5456 => x"52",
          5457 => x"b7",
          5458 => x"c8",
          5459 => x"ff",
          5460 => x"7c",
          5461 => x"2b",
          5462 => x"08",
          5463 => x"53",
          5464 => x"8e",
          5465 => x"d8",
          5466 => x"84",
          5467 => x"ff",
          5468 => x"5c",
          5469 => x"60",
          5470 => x"74",
          5471 => x"38",
          5472 => x"c9",
          5473 => x"c0",
          5474 => x"11",
          5475 => x"33",
          5476 => x"07",
          5477 => x"f4",
          5478 => x"52",
          5479 => x"df",
          5480 => x"c8",
          5481 => x"ff",
          5482 => x"7c",
          5483 => x"2b",
          5484 => x"08",
          5485 => x"53",
          5486 => x"8d",
          5487 => x"d8",
          5488 => x"84",
          5489 => x"05",
          5490 => x"73",
          5491 => x"06",
          5492 => x"7b",
          5493 => x"f9",
          5494 => x"d8",
          5495 => x"82",
          5496 => x"80",
          5497 => x"7d",
          5498 => x"82",
          5499 => x"51",
          5500 => x"3f",
          5501 => x"98",
          5502 => x"7a",
          5503 => x"38",
          5504 => x"52",
          5505 => x"8f",
          5506 => x"83",
          5507 => x"c0",
          5508 => x"05",
          5509 => x"3f",
          5510 => x"82",
          5511 => x"94",
          5512 => x"fc",
          5513 => x"77",
          5514 => x"54",
          5515 => x"82",
          5516 => x"55",
          5517 => x"08",
          5518 => x"38",
          5519 => x"52",
          5520 => x"08",
          5521 => x"9f",
          5522 => x"d8",
          5523 => x"3d",
          5524 => x"3d",
          5525 => x"05",
          5526 => x"52",
          5527 => x"87",
          5528 => x"c4",
          5529 => x"71",
          5530 => x"0c",
          5531 => x"04",
          5532 => x"02",
          5533 => x"02",
          5534 => x"05",
          5535 => x"83",
          5536 => x"26",
          5537 => x"72",
          5538 => x"c0",
          5539 => x"53",
          5540 => x"74",
          5541 => x"38",
          5542 => x"73",
          5543 => x"c0",
          5544 => x"51",
          5545 => x"85",
          5546 => x"98",
          5547 => x"52",
          5548 => x"82",
          5549 => x"70",
          5550 => x"38",
          5551 => x"8c",
          5552 => x"ec",
          5553 => x"fc",
          5554 => x"52",
          5555 => x"87",
          5556 => x"08",
          5557 => x"2e",
          5558 => x"82",
          5559 => x"34",
          5560 => x"13",
          5561 => x"82",
          5562 => x"86",
          5563 => x"f3",
          5564 => x"62",
          5565 => x"05",
          5566 => x"57",
          5567 => x"83",
          5568 => x"fe",
          5569 => x"d8",
          5570 => x"06",
          5571 => x"71",
          5572 => x"71",
          5573 => x"2b",
          5574 => x"80",
          5575 => x"92",
          5576 => x"c0",
          5577 => x"41",
          5578 => x"5a",
          5579 => x"87",
          5580 => x"0c",
          5581 => x"84",
          5582 => x"08",
          5583 => x"70",
          5584 => x"53",
          5585 => x"2e",
          5586 => x"08",
          5587 => x"70",
          5588 => x"34",
          5589 => x"80",
          5590 => x"53",
          5591 => x"2e",
          5592 => x"53",
          5593 => x"26",
          5594 => x"80",
          5595 => x"87",
          5596 => x"08",
          5597 => x"38",
          5598 => x"8c",
          5599 => x"80",
          5600 => x"78",
          5601 => x"99",
          5602 => x"0c",
          5603 => x"8c",
          5604 => x"08",
          5605 => x"51",
          5606 => x"38",
          5607 => x"8d",
          5608 => x"17",
          5609 => x"81",
          5610 => x"53",
          5611 => x"2e",
          5612 => x"fc",
          5613 => x"52",
          5614 => x"7d",
          5615 => x"ed",
          5616 => x"80",
          5617 => x"71",
          5618 => x"38",
          5619 => x"53",
          5620 => x"c8",
          5621 => x"0d",
          5622 => x"0d",
          5623 => x"02",
          5624 => x"05",
          5625 => x"58",
          5626 => x"80",
          5627 => x"fc",
          5628 => x"d8",
          5629 => x"06",
          5630 => x"71",
          5631 => x"81",
          5632 => x"38",
          5633 => x"2b",
          5634 => x"80",
          5635 => x"92",
          5636 => x"c0",
          5637 => x"40",
          5638 => x"5a",
          5639 => x"c0",
          5640 => x"76",
          5641 => x"76",
          5642 => x"75",
          5643 => x"2a",
          5644 => x"51",
          5645 => x"80",
          5646 => x"7a",
          5647 => x"5c",
          5648 => x"81",
          5649 => x"81",
          5650 => x"06",
          5651 => x"80",
          5652 => x"87",
          5653 => x"08",
          5654 => x"38",
          5655 => x"8c",
          5656 => x"80",
          5657 => x"77",
          5658 => x"99",
          5659 => x"0c",
          5660 => x"8c",
          5661 => x"08",
          5662 => x"51",
          5663 => x"38",
          5664 => x"8d",
          5665 => x"70",
          5666 => x"84",
          5667 => x"5b",
          5668 => x"2e",
          5669 => x"fc",
          5670 => x"52",
          5671 => x"7d",
          5672 => x"f8",
          5673 => x"80",
          5674 => x"71",
          5675 => x"38",
          5676 => x"53",
          5677 => x"c8",
          5678 => x"0d",
          5679 => x"0d",
          5680 => x"05",
          5681 => x"02",
          5682 => x"05",
          5683 => x"54",
          5684 => x"fe",
          5685 => x"c8",
          5686 => x"53",
          5687 => x"80",
          5688 => x"0b",
          5689 => x"8c",
          5690 => x"71",
          5691 => x"dc",
          5692 => x"24",
          5693 => x"84",
          5694 => x"92",
          5695 => x"54",
          5696 => x"8d",
          5697 => x"39",
          5698 => x"80",
          5699 => x"cb",
          5700 => x"70",
          5701 => x"81",
          5702 => x"52",
          5703 => x"8a",
          5704 => x"98",
          5705 => x"71",
          5706 => x"c0",
          5707 => x"52",
          5708 => x"81",
          5709 => x"c0",
          5710 => x"53",
          5711 => x"82",
          5712 => x"71",
          5713 => x"39",
          5714 => x"39",
          5715 => x"77",
          5716 => x"81",
          5717 => x"72",
          5718 => x"84",
          5719 => x"73",
          5720 => x"0c",
          5721 => x"04",
          5722 => x"74",
          5723 => x"71",
          5724 => x"2b",
          5725 => x"c8",
          5726 => x"84",
          5727 => x"fd",
          5728 => x"83",
          5729 => x"12",
          5730 => x"2b",
          5731 => x"07",
          5732 => x"70",
          5733 => x"2b",
          5734 => x"07",
          5735 => x"0c",
          5736 => x"56",
          5737 => x"3d",
          5738 => x"3d",
          5739 => x"84",
          5740 => x"22",
          5741 => x"72",
          5742 => x"54",
          5743 => x"2a",
          5744 => x"34",
          5745 => x"04",
          5746 => x"73",
          5747 => x"70",
          5748 => x"05",
          5749 => x"88",
          5750 => x"72",
          5751 => x"54",
          5752 => x"2a",
          5753 => x"70",
          5754 => x"34",
          5755 => x"51",
          5756 => x"83",
          5757 => x"fe",
          5758 => x"75",
          5759 => x"51",
          5760 => x"92",
          5761 => x"81",
          5762 => x"73",
          5763 => x"55",
          5764 => x"51",
          5765 => x"3d",
          5766 => x"3d",
          5767 => x"76",
          5768 => x"72",
          5769 => x"05",
          5770 => x"11",
          5771 => x"38",
          5772 => x"04",
          5773 => x"78",
          5774 => x"56",
          5775 => x"81",
          5776 => x"74",
          5777 => x"56",
          5778 => x"31",
          5779 => x"52",
          5780 => x"80",
          5781 => x"71",
          5782 => x"38",
          5783 => x"c8",
          5784 => x"0d",
          5785 => x"0d",
          5786 => x"51",
          5787 => x"73",
          5788 => x"81",
          5789 => x"33",
          5790 => x"38",
          5791 => x"d8",
          5792 => x"3d",
          5793 => x"0b",
          5794 => x"0c",
          5795 => x"0d",
          5796 => x"70",
          5797 => x"52",
          5798 => x"55",
          5799 => x"3f",
          5800 => x"d8",
          5801 => x"38",
          5802 => x"98",
          5803 => x"52",
          5804 => x"f7",
          5805 => x"d8",
          5806 => x"ff",
          5807 => x"72",
          5808 => x"38",
          5809 => x"72",
          5810 => x"d8",
          5811 => x"3d",
          5812 => x"3d",
          5813 => x"80",
          5814 => x"33",
          5815 => x"7a",
          5816 => x"38",
          5817 => x"16",
          5818 => x"16",
          5819 => x"17",
          5820 => x"f9",
          5821 => x"d8",
          5822 => x"2e",
          5823 => x"b7",
          5824 => x"c8",
          5825 => x"34",
          5826 => x"70",
          5827 => x"31",
          5828 => x"59",
          5829 => x"77",
          5830 => x"82",
          5831 => x"74",
          5832 => x"81",
          5833 => x"81",
          5834 => x"53",
          5835 => x"16",
          5836 => x"a5",
          5837 => x"81",
          5838 => x"d8",
          5839 => x"3d",
          5840 => x"3d",
          5841 => x"56",
          5842 => x"74",
          5843 => x"2e",
          5844 => x"51",
          5845 => x"82",
          5846 => x"57",
          5847 => x"08",
          5848 => x"54",
          5849 => x"16",
          5850 => x"33",
          5851 => x"3f",
          5852 => x"08",
          5853 => x"38",
          5854 => x"57",
          5855 => x"0c",
          5856 => x"c8",
          5857 => x"0d",
          5858 => x"0d",
          5859 => x"57",
          5860 => x"82",
          5861 => x"58",
          5862 => x"08",
          5863 => x"76",
          5864 => x"83",
          5865 => x"06",
          5866 => x"84",
          5867 => x"78",
          5868 => x"81",
          5869 => x"38",
          5870 => x"82",
          5871 => x"52",
          5872 => x"52",
          5873 => x"3f",
          5874 => x"52",
          5875 => x"51",
          5876 => x"84",
          5877 => x"d2",
          5878 => x"fb",
          5879 => x"8a",
          5880 => x"52",
          5881 => x"51",
          5882 => x"94",
          5883 => x"84",
          5884 => x"fb",
          5885 => x"17",
          5886 => x"a4",
          5887 => x"c8",
          5888 => x"08",
          5889 => x"b4",
          5890 => x"55",
          5891 => x"81",
          5892 => x"f7",
          5893 => x"84",
          5894 => x"53",
          5895 => x"17",
          5896 => x"99",
          5897 => x"c8",
          5898 => x"83",
          5899 => x"77",
          5900 => x"0c",
          5901 => x"04",
          5902 => x"77",
          5903 => x"12",
          5904 => x"55",
          5905 => x"56",
          5906 => x"8d",
          5907 => x"22",
          5908 => x"b0",
          5909 => x"57",
          5910 => x"d8",
          5911 => x"3d",
          5912 => x"3d",
          5913 => x"70",
          5914 => x"57",
          5915 => x"81",
          5916 => x"9c",
          5917 => x"81",
          5918 => x"74",
          5919 => x"72",
          5920 => x"f5",
          5921 => x"24",
          5922 => x"81",
          5923 => x"81",
          5924 => x"83",
          5925 => x"38",
          5926 => x"76",
          5927 => x"70",
          5928 => x"16",
          5929 => x"74",
          5930 => x"96",
          5931 => x"c8",
          5932 => x"38",
          5933 => x"06",
          5934 => x"33",
          5935 => x"89",
          5936 => x"08",
          5937 => x"54",
          5938 => x"fc",
          5939 => x"d8",
          5940 => x"fe",
          5941 => x"ff",
          5942 => x"11",
          5943 => x"2b",
          5944 => x"81",
          5945 => x"2a",
          5946 => x"51",
          5947 => x"e2",
          5948 => x"ff",
          5949 => x"da",
          5950 => x"2a",
          5951 => x"05",
          5952 => x"fc",
          5953 => x"d8",
          5954 => x"c6",
          5955 => x"83",
          5956 => x"05",
          5957 => x"f8",
          5958 => x"d8",
          5959 => x"ff",
          5960 => x"ae",
          5961 => x"2a",
          5962 => x"05",
          5963 => x"fc",
          5964 => x"d8",
          5965 => x"38",
          5966 => x"83",
          5967 => x"05",
          5968 => x"f8",
          5969 => x"d8",
          5970 => x"0a",
          5971 => x"39",
          5972 => x"82",
          5973 => x"89",
          5974 => x"f8",
          5975 => x"7c",
          5976 => x"56",
          5977 => x"77",
          5978 => x"38",
          5979 => x"08",
          5980 => x"38",
          5981 => x"72",
          5982 => x"9d",
          5983 => x"24",
          5984 => x"81",
          5985 => x"82",
          5986 => x"83",
          5987 => x"38",
          5988 => x"76",
          5989 => x"70",
          5990 => x"18",
          5991 => x"76",
          5992 => x"9e",
          5993 => x"c8",
          5994 => x"d8",
          5995 => x"d9",
          5996 => x"ff",
          5997 => x"05",
          5998 => x"81",
          5999 => x"54",
          6000 => x"80",
          6001 => x"77",
          6002 => x"f0",
          6003 => x"8f",
          6004 => x"51",
          6005 => x"34",
          6006 => x"17",
          6007 => x"2a",
          6008 => x"05",
          6009 => x"fa",
          6010 => x"d8",
          6011 => x"82",
          6012 => x"81",
          6013 => x"83",
          6014 => x"b8",
          6015 => x"2a",
          6016 => x"8f",
          6017 => x"2a",
          6018 => x"f0",
          6019 => x"06",
          6020 => x"72",
          6021 => x"ec",
          6022 => x"2a",
          6023 => x"05",
          6024 => x"fa",
          6025 => x"d8",
          6026 => x"82",
          6027 => x"80",
          6028 => x"83",
          6029 => x"52",
          6030 => x"fe",
          6031 => x"b8",
          6032 => x"e6",
          6033 => x"76",
          6034 => x"17",
          6035 => x"75",
          6036 => x"3f",
          6037 => x"08",
          6038 => x"c8",
          6039 => x"77",
          6040 => x"77",
          6041 => x"fc",
          6042 => x"b8",
          6043 => x"51",
          6044 => x"8b",
          6045 => x"c8",
          6046 => x"06",
          6047 => x"72",
          6048 => x"3f",
          6049 => x"17",
          6050 => x"d8",
          6051 => x"3d",
          6052 => x"3d",
          6053 => x"7e",
          6054 => x"56",
          6055 => x"75",
          6056 => x"74",
          6057 => x"27",
          6058 => x"80",
          6059 => x"ff",
          6060 => x"75",
          6061 => x"3f",
          6062 => x"08",
          6063 => x"c8",
          6064 => x"38",
          6065 => x"54",
          6066 => x"81",
          6067 => x"39",
          6068 => x"08",
          6069 => x"39",
          6070 => x"51",
          6071 => x"82",
          6072 => x"58",
          6073 => x"08",
          6074 => x"c7",
          6075 => x"c8",
          6076 => x"d2",
          6077 => x"c8",
          6078 => x"cf",
          6079 => x"74",
          6080 => x"fc",
          6081 => x"d8",
          6082 => x"38",
          6083 => x"fe",
          6084 => x"08",
          6085 => x"74",
          6086 => x"38",
          6087 => x"17",
          6088 => x"33",
          6089 => x"73",
          6090 => x"77",
          6091 => x"26",
          6092 => x"80",
          6093 => x"d8",
          6094 => x"3d",
          6095 => x"3d",
          6096 => x"71",
          6097 => x"5b",
          6098 => x"90",
          6099 => x"77",
          6100 => x"38",
          6101 => x"78",
          6102 => x"81",
          6103 => x"79",
          6104 => x"f9",
          6105 => x"55",
          6106 => x"c8",
          6107 => x"e0",
          6108 => x"c8",
          6109 => x"d8",
          6110 => x"2e",
          6111 => x"9c",
          6112 => x"d8",
          6113 => x"82",
          6114 => x"58",
          6115 => x"70",
          6116 => x"80",
          6117 => x"38",
          6118 => x"09",
          6119 => x"e2",
          6120 => x"56",
          6121 => x"76",
          6122 => x"82",
          6123 => x"7a",
          6124 => x"3f",
          6125 => x"d8",
          6126 => x"2e",
          6127 => x"86",
          6128 => x"c8",
          6129 => x"d8",
          6130 => x"70",
          6131 => x"07",
          6132 => x"7c",
          6133 => x"c8",
          6134 => x"51",
          6135 => x"81",
          6136 => x"d8",
          6137 => x"2e",
          6138 => x"17",
          6139 => x"74",
          6140 => x"73",
          6141 => x"27",
          6142 => x"58",
          6143 => x"80",
          6144 => x"56",
          6145 => x"9c",
          6146 => x"26",
          6147 => x"56",
          6148 => x"81",
          6149 => x"52",
          6150 => x"c6",
          6151 => x"c8",
          6152 => x"b8",
          6153 => x"82",
          6154 => x"81",
          6155 => x"06",
          6156 => x"d8",
          6157 => x"82",
          6158 => x"09",
          6159 => x"72",
          6160 => x"70",
          6161 => x"51",
          6162 => x"80",
          6163 => x"78",
          6164 => x"06",
          6165 => x"73",
          6166 => x"39",
          6167 => x"52",
          6168 => x"f7",
          6169 => x"c8",
          6170 => x"c8",
          6171 => x"82",
          6172 => x"07",
          6173 => x"55",
          6174 => x"2e",
          6175 => x"80",
          6176 => x"75",
          6177 => x"76",
          6178 => x"3f",
          6179 => x"08",
          6180 => x"38",
          6181 => x"0c",
          6182 => x"fe",
          6183 => x"08",
          6184 => x"74",
          6185 => x"ff",
          6186 => x"0c",
          6187 => x"81",
          6188 => x"84",
          6189 => x"39",
          6190 => x"81",
          6191 => x"8c",
          6192 => x"8c",
          6193 => x"c8",
          6194 => x"39",
          6195 => x"55",
          6196 => x"c8",
          6197 => x"0d",
          6198 => x"0d",
          6199 => x"55",
          6200 => x"82",
          6201 => x"58",
          6202 => x"d8",
          6203 => x"d8",
          6204 => x"74",
          6205 => x"3f",
          6206 => x"08",
          6207 => x"08",
          6208 => x"59",
          6209 => x"77",
          6210 => x"70",
          6211 => x"8a",
          6212 => x"84",
          6213 => x"56",
          6214 => x"58",
          6215 => x"97",
          6216 => x"75",
          6217 => x"52",
          6218 => x"51",
          6219 => x"82",
          6220 => x"80",
          6221 => x"8a",
          6222 => x"32",
          6223 => x"72",
          6224 => x"2a",
          6225 => x"56",
          6226 => x"c8",
          6227 => x"0d",
          6228 => x"0d",
          6229 => x"08",
          6230 => x"74",
          6231 => x"26",
          6232 => x"74",
          6233 => x"72",
          6234 => x"74",
          6235 => x"88",
          6236 => x"73",
          6237 => x"33",
          6238 => x"27",
          6239 => x"16",
          6240 => x"9b",
          6241 => x"2a",
          6242 => x"88",
          6243 => x"58",
          6244 => x"80",
          6245 => x"16",
          6246 => x"0c",
          6247 => x"8a",
          6248 => x"89",
          6249 => x"72",
          6250 => x"38",
          6251 => x"51",
          6252 => x"82",
          6253 => x"54",
          6254 => x"08",
          6255 => x"38",
          6256 => x"d8",
          6257 => x"8b",
          6258 => x"08",
          6259 => x"08",
          6260 => x"82",
          6261 => x"74",
          6262 => x"cb",
          6263 => x"75",
          6264 => x"3f",
          6265 => x"08",
          6266 => x"73",
          6267 => x"98",
          6268 => x"82",
          6269 => x"2e",
          6270 => x"39",
          6271 => x"39",
          6272 => x"13",
          6273 => x"74",
          6274 => x"16",
          6275 => x"18",
          6276 => x"77",
          6277 => x"0c",
          6278 => x"04",
          6279 => x"7a",
          6280 => x"12",
          6281 => x"59",
          6282 => x"80",
          6283 => x"86",
          6284 => x"98",
          6285 => x"14",
          6286 => x"55",
          6287 => x"81",
          6288 => x"83",
          6289 => x"77",
          6290 => x"81",
          6291 => x"0c",
          6292 => x"55",
          6293 => x"76",
          6294 => x"17",
          6295 => x"74",
          6296 => x"9b",
          6297 => x"39",
          6298 => x"ff",
          6299 => x"2a",
          6300 => x"81",
          6301 => x"52",
          6302 => x"e6",
          6303 => x"c8",
          6304 => x"55",
          6305 => x"d8",
          6306 => x"80",
          6307 => x"55",
          6308 => x"08",
          6309 => x"f4",
          6310 => x"08",
          6311 => x"08",
          6312 => x"38",
          6313 => x"77",
          6314 => x"84",
          6315 => x"39",
          6316 => x"52",
          6317 => x"86",
          6318 => x"c8",
          6319 => x"55",
          6320 => x"08",
          6321 => x"c4",
          6322 => x"82",
          6323 => x"81",
          6324 => x"81",
          6325 => x"c8",
          6326 => x"b0",
          6327 => x"c8",
          6328 => x"51",
          6329 => x"82",
          6330 => x"a0",
          6331 => x"15",
          6332 => x"75",
          6333 => x"3f",
          6334 => x"08",
          6335 => x"76",
          6336 => x"77",
          6337 => x"9c",
          6338 => x"55",
          6339 => x"c8",
          6340 => x"0d",
          6341 => x"0d",
          6342 => x"08",
          6343 => x"80",
          6344 => x"fc",
          6345 => x"d8",
          6346 => x"82",
          6347 => x"80",
          6348 => x"d8",
          6349 => x"98",
          6350 => x"78",
          6351 => x"3f",
          6352 => x"08",
          6353 => x"c8",
          6354 => x"38",
          6355 => x"08",
          6356 => x"70",
          6357 => x"58",
          6358 => x"2e",
          6359 => x"83",
          6360 => x"82",
          6361 => x"55",
          6362 => x"81",
          6363 => x"07",
          6364 => x"2e",
          6365 => x"16",
          6366 => x"2e",
          6367 => x"88",
          6368 => x"82",
          6369 => x"56",
          6370 => x"51",
          6371 => x"82",
          6372 => x"54",
          6373 => x"08",
          6374 => x"9b",
          6375 => x"2e",
          6376 => x"83",
          6377 => x"73",
          6378 => x"0c",
          6379 => x"04",
          6380 => x"76",
          6381 => x"54",
          6382 => x"82",
          6383 => x"83",
          6384 => x"76",
          6385 => x"53",
          6386 => x"2e",
          6387 => x"90",
          6388 => x"51",
          6389 => x"82",
          6390 => x"90",
          6391 => x"53",
          6392 => x"c8",
          6393 => x"0d",
          6394 => x"0d",
          6395 => x"83",
          6396 => x"54",
          6397 => x"55",
          6398 => x"3f",
          6399 => x"51",
          6400 => x"2e",
          6401 => x"8b",
          6402 => x"2a",
          6403 => x"51",
          6404 => x"86",
          6405 => x"fd",
          6406 => x"54",
          6407 => x"53",
          6408 => x"71",
          6409 => x"05",
          6410 => x"05",
          6411 => x"05",
          6412 => x"06",
          6413 => x"51",
          6414 => x"e4",
          6415 => x"d8",
          6416 => x"3d",
          6417 => x"3d",
          6418 => x"40",
          6419 => x"08",
          6420 => x"ff",
          6421 => x"98",
          6422 => x"2e",
          6423 => x"98",
          6424 => x"7d",
          6425 => x"3f",
          6426 => x"08",
          6427 => x"c8",
          6428 => x"38",
          6429 => x"70",
          6430 => x"73",
          6431 => x"5b",
          6432 => x"8b",
          6433 => x"06",
          6434 => x"06",
          6435 => x"86",
          6436 => x"d8",
          6437 => x"73",
          6438 => x"09",
          6439 => x"38",
          6440 => x"d8",
          6441 => x"73",
          6442 => x"81",
          6443 => x"81",
          6444 => x"07",
          6445 => x"38",
          6446 => x"08",
          6447 => x"54",
          6448 => x"2e",
          6449 => x"83",
          6450 => x"75",
          6451 => x"38",
          6452 => x"81",
          6453 => x"8f",
          6454 => x"06",
          6455 => x"73",
          6456 => x"81",
          6457 => x"72",
          6458 => x"38",
          6459 => x"74",
          6460 => x"70",
          6461 => x"ac",
          6462 => x"5d",
          6463 => x"2e",
          6464 => x"81",
          6465 => x"15",
          6466 => x"73",
          6467 => x"06",
          6468 => x"8c",
          6469 => x"16",
          6470 => x"cc",
          6471 => x"c8",
          6472 => x"ff",
          6473 => x"80",
          6474 => x"33",
          6475 => x"06",
          6476 => x"05",
          6477 => x"7b",
          6478 => x"ca",
          6479 => x"75",
          6480 => x"a4",
          6481 => x"c8",
          6482 => x"ff",
          6483 => x"80",
          6484 => x"73",
          6485 => x"80",
          6486 => x"10",
          6487 => x"53",
          6488 => x"81",
          6489 => x"39",
          6490 => x"ff",
          6491 => x"06",
          6492 => x"17",
          6493 => x"27",
          6494 => x"33",
          6495 => x"70",
          6496 => x"54",
          6497 => x"2e",
          6498 => x"81",
          6499 => x"38",
          6500 => x"53",
          6501 => x"ff",
          6502 => x"ff",
          6503 => x"84",
          6504 => x"53",
          6505 => x"39",
          6506 => x"74",
          6507 => x"3f",
          6508 => x"08",
          6509 => x"53",
          6510 => x"a7",
          6511 => x"ac",
          6512 => x"39",
          6513 => x"51",
          6514 => x"82",
          6515 => x"5b",
          6516 => x"08",
          6517 => x"19",
          6518 => x"38",
          6519 => x"0b",
          6520 => x"7a",
          6521 => x"0c",
          6522 => x"04",
          6523 => x"60",
          6524 => x"59",
          6525 => x"51",
          6526 => x"82",
          6527 => x"58",
          6528 => x"08",
          6529 => x"81",
          6530 => x"5c",
          6531 => x"1a",
          6532 => x"08",
          6533 => x"ea",
          6534 => x"d8",
          6535 => x"82",
          6536 => x"83",
          6537 => x"19",
          6538 => x"57",
          6539 => x"38",
          6540 => x"f6",
          6541 => x"33",
          6542 => x"81",
          6543 => x"54",
          6544 => x"34",
          6545 => x"2e",
          6546 => x"74",
          6547 => x"81",
          6548 => x"74",
          6549 => x"38",
          6550 => x"38",
          6551 => x"09",
          6552 => x"f7",
          6553 => x"33",
          6554 => x"70",
          6555 => x"55",
          6556 => x"a1",
          6557 => x"2a",
          6558 => x"51",
          6559 => x"2e",
          6560 => x"17",
          6561 => x"bf",
          6562 => x"1c",
          6563 => x"0c",
          6564 => x"75",
          6565 => x"81",
          6566 => x"38",
          6567 => x"56",
          6568 => x"09",
          6569 => x"ac",
          6570 => x"08",
          6571 => x"5d",
          6572 => x"82",
          6573 => x"83",
          6574 => x"55",
          6575 => x"38",
          6576 => x"bf",
          6577 => x"f3",
          6578 => x"81",
          6579 => x"82",
          6580 => x"33",
          6581 => x"e5",
          6582 => x"d8",
          6583 => x"ff",
          6584 => x"79",
          6585 => x"38",
          6586 => x"26",
          6587 => x"75",
          6588 => x"b4",
          6589 => x"c8",
          6590 => x"1e",
          6591 => x"55",
          6592 => x"55",
          6593 => x"3f",
          6594 => x"c8",
          6595 => x"81",
          6596 => x"38",
          6597 => x"39",
          6598 => x"ff",
          6599 => x"06",
          6600 => x"1b",
          6601 => x"27",
          6602 => x"76",
          6603 => x"2a",
          6604 => x"51",
          6605 => x"80",
          6606 => x"73",
          6607 => x"38",
          6608 => x"70",
          6609 => x"73",
          6610 => x"1c",
          6611 => x"06",
          6612 => x"39",
          6613 => x"73",
          6614 => x"7b",
          6615 => x"51",
          6616 => x"82",
          6617 => x"81",
          6618 => x"73",
          6619 => x"38",
          6620 => x"81",
          6621 => x"95",
          6622 => x"a0",
          6623 => x"19",
          6624 => x"b0",
          6625 => x"c8",
          6626 => x"9e",
          6627 => x"5c",
          6628 => x"1a",
          6629 => x"78",
          6630 => x"3f",
          6631 => x"08",
          6632 => x"c8",
          6633 => x"fc",
          6634 => x"82",
          6635 => x"90",
          6636 => x"ee",
          6637 => x"70",
          6638 => x"33",
          6639 => x"56",
          6640 => x"55",
          6641 => x"38",
          6642 => x"08",
          6643 => x"56",
          6644 => x"2e",
          6645 => x"1d",
          6646 => x"70",
          6647 => x"5d",
          6648 => x"53",
          6649 => x"53",
          6650 => x"53",
          6651 => x"87",
          6652 => x"cb",
          6653 => x"06",
          6654 => x"2e",
          6655 => x"80",
          6656 => x"1b",
          6657 => x"8c",
          6658 => x"56",
          6659 => x"7d",
          6660 => x"e3",
          6661 => x"7b",
          6662 => x"38",
          6663 => x"22",
          6664 => x"ff",
          6665 => x"73",
          6666 => x"38",
          6667 => x"ff",
          6668 => x"59",
          6669 => x"74",
          6670 => x"10",
          6671 => x"2a",
          6672 => x"70",
          6673 => x"56",
          6674 => x"80",
          6675 => x"75",
          6676 => x"32",
          6677 => x"57",
          6678 => x"db",
          6679 => x"75",
          6680 => x"84",
          6681 => x"57",
          6682 => x"07",
          6683 => x"b9",
          6684 => x"38",
          6685 => x"73",
          6686 => x"16",
          6687 => x"84",
          6688 => x"56",
          6689 => x"94",
          6690 => x"17",
          6691 => x"74",
          6692 => x"27",
          6693 => x"33",
          6694 => x"2e",
          6695 => x"19",
          6696 => x"54",
          6697 => x"82",
          6698 => x"80",
          6699 => x"ff",
          6700 => x"74",
          6701 => x"81",
          6702 => x"15",
          6703 => x"27",
          6704 => x"19",
          6705 => x"54",
          6706 => x"3d",
          6707 => x"05",
          6708 => x"81",
          6709 => x"a0",
          6710 => x"26",
          6711 => x"17",
          6712 => x"33",
          6713 => x"75",
          6714 => x"75",
          6715 => x"79",
          6716 => x"3f",
          6717 => x"08",
          6718 => x"1b",
          6719 => x"7b",
          6720 => x"38",
          6721 => x"80",
          6722 => x"f0",
          6723 => x"c8",
          6724 => x"d8",
          6725 => x"2e",
          6726 => x"82",
          6727 => x"80",
          6728 => x"ab",
          6729 => x"80",
          6730 => x"70",
          6731 => x"81",
          6732 => x"5e",
          6733 => x"80",
          6734 => x"8d",
          6735 => x"51",
          6736 => x"3f",
          6737 => x"08",
          6738 => x"52",
          6739 => x"c5",
          6740 => x"c8",
          6741 => x"d8",
          6742 => x"9e",
          6743 => x"59",
          6744 => x"81",
          6745 => x"85",
          6746 => x"08",
          6747 => x"54",
          6748 => x"dd",
          6749 => x"c8",
          6750 => x"d8",
          6751 => x"fa",
          6752 => x"51",
          6753 => x"82",
          6754 => x"81",
          6755 => x"98",
          6756 => x"7b",
          6757 => x"3f",
          6758 => x"08",
          6759 => x"c8",
          6760 => x"38",
          6761 => x"9c",
          6762 => x"81",
          6763 => x"57",
          6764 => x"17",
          6765 => x"8b",
          6766 => x"d8",
          6767 => x"17",
          6768 => x"c8",
          6769 => x"16",
          6770 => x"3f",
          6771 => x"f3",
          6772 => x"55",
          6773 => x"ff",
          6774 => x"74",
          6775 => x"22",
          6776 => x"51",
          6777 => x"82",
          6778 => x"33",
          6779 => x"df",
          6780 => x"85",
          6781 => x"ff",
          6782 => x"57",
          6783 => x"d4",
          6784 => x"ff",
          6785 => x"38",
          6786 => x"70",
          6787 => x"73",
          6788 => x"80",
          6789 => x"77",
          6790 => x"0b",
          6791 => x"80",
          6792 => x"ef",
          6793 => x"d8",
          6794 => x"82",
          6795 => x"80",
          6796 => x"19",
          6797 => x"d7",
          6798 => x"08",
          6799 => x"e2",
          6800 => x"d8",
          6801 => x"82",
          6802 => x"ae",
          6803 => x"82",
          6804 => x"52",
          6805 => x"51",
          6806 => x"8b",
          6807 => x"52",
          6808 => x"51",
          6809 => x"9c",
          6810 => x"1b",
          6811 => x"55",
          6812 => x"16",
          6813 => x"83",
          6814 => x"55",
          6815 => x"c8",
          6816 => x"0d",
          6817 => x"0d",
          6818 => x"90",
          6819 => x"13",
          6820 => x"57",
          6821 => x"2e",
          6822 => x"52",
          6823 => x"b1",
          6824 => x"c8",
          6825 => x"d8",
          6826 => x"c9",
          6827 => x"08",
          6828 => x"e1",
          6829 => x"d8",
          6830 => x"82",
          6831 => x"ab",
          6832 => x"08",
          6833 => x"34",
          6834 => x"17",
          6835 => x"08",
          6836 => x"38",
          6837 => x"08",
          6838 => x"ee",
          6839 => x"d8",
          6840 => x"82",
          6841 => x"80",
          6842 => x"73",
          6843 => x"81",
          6844 => x"82",
          6845 => x"d8",
          6846 => x"3d",
          6847 => x"3d",
          6848 => x"71",
          6849 => x"5c",
          6850 => x"19",
          6851 => x"08",
          6852 => x"e2",
          6853 => x"08",
          6854 => x"bb",
          6855 => x"71",
          6856 => x"08",
          6857 => x"57",
          6858 => x"72",
          6859 => x"9d",
          6860 => x"14",
          6861 => x"1b",
          6862 => x"7a",
          6863 => x"d0",
          6864 => x"83",
          6865 => x"51",
          6866 => x"ff",
          6867 => x"74",
          6868 => x"39",
          6869 => x"11",
          6870 => x"31",
          6871 => x"83",
          6872 => x"90",
          6873 => x"51",
          6874 => x"3f",
          6875 => x"08",
          6876 => x"06",
          6877 => x"75",
          6878 => x"81",
          6879 => x"38",
          6880 => x"53",
          6881 => x"74",
          6882 => x"82",
          6883 => x"74",
          6884 => x"70",
          6885 => x"25",
          6886 => x"07",
          6887 => x"73",
          6888 => x"38",
          6889 => x"39",
          6890 => x"81",
          6891 => x"57",
          6892 => x"1d",
          6893 => x"11",
          6894 => x"54",
          6895 => x"f1",
          6896 => x"70",
          6897 => x"30",
          6898 => x"51",
          6899 => x"94",
          6900 => x"0b",
          6901 => x"80",
          6902 => x"58",
          6903 => x"1c",
          6904 => x"33",
          6905 => x"56",
          6906 => x"2e",
          6907 => x"85",
          6908 => x"06",
          6909 => x"e5",
          6910 => x"32",
          6911 => x"72",
          6912 => x"51",
          6913 => x"8b",
          6914 => x"72",
          6915 => x"38",
          6916 => x"81",
          6917 => x"81",
          6918 => x"76",
          6919 => x"58",
          6920 => x"57",
          6921 => x"ff",
          6922 => x"17",
          6923 => x"80",
          6924 => x"34",
          6925 => x"53",
          6926 => x"38",
          6927 => x"bf",
          6928 => x"34",
          6929 => x"e1",
          6930 => x"89",
          6931 => x"5a",
          6932 => x"2e",
          6933 => x"96",
          6934 => x"55",
          6935 => x"ff",
          6936 => x"55",
          6937 => x"aa",
          6938 => x"08",
          6939 => x"51",
          6940 => x"27",
          6941 => x"84",
          6942 => x"39",
          6943 => x"53",
          6944 => x"53",
          6945 => x"8a",
          6946 => x"70",
          6947 => x"06",
          6948 => x"76",
          6949 => x"58",
          6950 => x"81",
          6951 => x"71",
          6952 => x"55",
          6953 => x"b5",
          6954 => x"94",
          6955 => x"0b",
          6956 => x"9c",
          6957 => x"11",
          6958 => x"72",
          6959 => x"89",
          6960 => x"1c",
          6961 => x"13",
          6962 => x"34",
          6963 => x"9c",
          6964 => x"d9",
          6965 => x"d8",
          6966 => x"0c",
          6967 => x"d9",
          6968 => x"d8",
          6969 => x"19",
          6970 => x"51",
          6971 => x"82",
          6972 => x"84",
          6973 => x"3d",
          6974 => x"3d",
          6975 => x"08",
          6976 => x"64",
          6977 => x"55",
          6978 => x"2e",
          6979 => x"55",
          6980 => x"2e",
          6981 => x"80",
          6982 => x"7f",
          6983 => x"88",
          6984 => x"39",
          6985 => x"80",
          6986 => x"56",
          6987 => x"af",
          6988 => x"06",
          6989 => x"56",
          6990 => x"32",
          6991 => x"80",
          6992 => x"51",
          6993 => x"dc",
          6994 => x"1f",
          6995 => x"33",
          6996 => x"9f",
          6997 => x"ff",
          6998 => x"1f",
          6999 => x"7d",
          7000 => x"3f",
          7001 => x"08",
          7002 => x"39",
          7003 => x"08",
          7004 => x"5b",
          7005 => x"92",
          7006 => x"51",
          7007 => x"82",
          7008 => x"ff",
          7009 => x"38",
          7010 => x"0b",
          7011 => x"08",
          7012 => x"78",
          7013 => x"d8",
          7014 => x"2a",
          7015 => x"75",
          7016 => x"59",
          7017 => x"08",
          7018 => x"06",
          7019 => x"70",
          7020 => x"27",
          7021 => x"07",
          7022 => x"56",
          7023 => x"75",
          7024 => x"ae",
          7025 => x"ff",
          7026 => x"75",
          7027 => x"ec",
          7028 => x"3f",
          7029 => x"08",
          7030 => x"78",
          7031 => x"81",
          7032 => x"10",
          7033 => x"74",
          7034 => x"59",
          7035 => x"81",
          7036 => x"61",
          7037 => x"56",
          7038 => x"2e",
          7039 => x"83",
          7040 => x"73",
          7041 => x"70",
          7042 => x"25",
          7043 => x"51",
          7044 => x"38",
          7045 => x"76",
          7046 => x"57",
          7047 => x"09",
          7048 => x"38",
          7049 => x"73",
          7050 => x"38",
          7051 => x"78",
          7052 => x"81",
          7053 => x"38",
          7054 => x"54",
          7055 => x"09",
          7056 => x"c1",
          7057 => x"54",
          7058 => x"09",
          7059 => x"38",
          7060 => x"54",
          7061 => x"80",
          7062 => x"56",
          7063 => x"78",
          7064 => x"38",
          7065 => x"75",
          7066 => x"57",
          7067 => x"58",
          7068 => x"e9",
          7069 => x"07",
          7070 => x"1f",
          7071 => x"39",
          7072 => x"a8",
          7073 => x"1a",
          7074 => x"74",
          7075 => x"71",
          7076 => x"70",
          7077 => x"2a",
          7078 => x"58",
          7079 => x"ae",
          7080 => x"73",
          7081 => x"19",
          7082 => x"38",
          7083 => x"11",
          7084 => x"74",
          7085 => x"38",
          7086 => x"90",
          7087 => x"07",
          7088 => x"39",
          7089 => x"70",
          7090 => x"06",
          7091 => x"73",
          7092 => x"81",
          7093 => x"81",
          7094 => x"1b",
          7095 => x"55",
          7096 => x"2e",
          7097 => x"8f",
          7098 => x"ff",
          7099 => x"73",
          7100 => x"81",
          7101 => x"76",
          7102 => x"78",
          7103 => x"38",
          7104 => x"05",
          7105 => x"54",
          7106 => x"9d",
          7107 => x"1a",
          7108 => x"ff",
          7109 => x"80",
          7110 => x"fe",
          7111 => x"55",
          7112 => x"2e",
          7113 => x"eb",
          7114 => x"a0",
          7115 => x"51",
          7116 => x"80",
          7117 => x"88",
          7118 => x"1a",
          7119 => x"1f",
          7120 => x"75",
          7121 => x"94",
          7122 => x"2e",
          7123 => x"ae",
          7124 => x"70",
          7125 => x"51",
          7126 => x"2e",
          7127 => x"80",
          7128 => x"76",
          7129 => x"d1",
          7130 => x"73",
          7131 => x"26",
          7132 => x"5b",
          7133 => x"70",
          7134 => x"07",
          7135 => x"7e",
          7136 => x"55",
          7137 => x"2e",
          7138 => x"8b",
          7139 => x"38",
          7140 => x"8b",
          7141 => x"07",
          7142 => x"26",
          7143 => x"78",
          7144 => x"8b",
          7145 => x"81",
          7146 => x"5f",
          7147 => x"80",
          7148 => x"af",
          7149 => x"07",
          7150 => x"52",
          7151 => x"cc",
          7152 => x"d8",
          7153 => x"ff",
          7154 => x"87",
          7155 => x"06",
          7156 => x"73",
          7157 => x"38",
          7158 => x"06",
          7159 => x"11",
          7160 => x"81",
          7161 => x"a4",
          7162 => x"54",
          7163 => x"8a",
          7164 => x"07",
          7165 => x"fe",
          7166 => x"18",
          7167 => x"88",
          7168 => x"73",
          7169 => x"18",
          7170 => x"39",
          7171 => x"92",
          7172 => x"82",
          7173 => x"d4",
          7174 => x"d8",
          7175 => x"2e",
          7176 => x"df",
          7177 => x"58",
          7178 => x"ff",
          7179 => x"73",
          7180 => x"38",
          7181 => x"5c",
          7182 => x"54",
          7183 => x"8e",
          7184 => x"07",
          7185 => x"83",
          7186 => x"58",
          7187 => x"18",
          7188 => x"75",
          7189 => x"18",
          7190 => x"39",
          7191 => x"54",
          7192 => x"2e",
          7193 => x"86",
          7194 => x"a0",
          7195 => x"88",
          7196 => x"06",
          7197 => x"82",
          7198 => x"06",
          7199 => x"06",
          7200 => x"2e",
          7201 => x"83",
          7202 => x"83",
          7203 => x"06",
          7204 => x"82",
          7205 => x"81",
          7206 => x"06",
          7207 => x"9f",
          7208 => x"06",
          7209 => x"2e",
          7210 => x"90",
          7211 => x"82",
          7212 => x"06",
          7213 => x"80",
          7214 => x"76",
          7215 => x"76",
          7216 => x"7d",
          7217 => x"3f",
          7218 => x"08",
          7219 => x"56",
          7220 => x"c8",
          7221 => x"be",
          7222 => x"c8",
          7223 => x"09",
          7224 => x"e8",
          7225 => x"2a",
          7226 => x"76",
          7227 => x"51",
          7228 => x"2e",
          7229 => x"81",
          7230 => x"80",
          7231 => x"38",
          7232 => x"ab",
          7233 => x"56",
          7234 => x"74",
          7235 => x"73",
          7236 => x"56",
          7237 => x"82",
          7238 => x"06",
          7239 => x"ac",
          7240 => x"33",
          7241 => x"70",
          7242 => x"55",
          7243 => x"2e",
          7244 => x"1e",
          7245 => x"06",
          7246 => x"05",
          7247 => x"e4",
          7248 => x"d8",
          7249 => x"1f",
          7250 => x"39",
          7251 => x"c8",
          7252 => x"0d",
          7253 => x"0d",
          7254 => x"7b",
          7255 => x"73",
          7256 => x"55",
          7257 => x"2e",
          7258 => x"75",
          7259 => x"57",
          7260 => x"26",
          7261 => x"ba",
          7262 => x"70",
          7263 => x"ba",
          7264 => x"06",
          7265 => x"73",
          7266 => x"70",
          7267 => x"51",
          7268 => x"89",
          7269 => x"82",
          7270 => x"ff",
          7271 => x"56",
          7272 => x"2e",
          7273 => x"80",
          7274 => x"c0",
          7275 => x"08",
          7276 => x"76",
          7277 => x"58",
          7278 => x"81",
          7279 => x"ff",
          7280 => x"53",
          7281 => x"26",
          7282 => x"13",
          7283 => x"06",
          7284 => x"9f",
          7285 => x"99",
          7286 => x"e0",
          7287 => x"ff",
          7288 => x"72",
          7289 => x"2a",
          7290 => x"72",
          7291 => x"06",
          7292 => x"ff",
          7293 => x"30",
          7294 => x"70",
          7295 => x"07",
          7296 => x"9f",
          7297 => x"54",
          7298 => x"80",
          7299 => x"81",
          7300 => x"59",
          7301 => x"25",
          7302 => x"8b",
          7303 => x"24",
          7304 => x"76",
          7305 => x"78",
          7306 => x"82",
          7307 => x"51",
          7308 => x"c8",
          7309 => x"0d",
          7310 => x"0d",
          7311 => x"0b",
          7312 => x"ff",
          7313 => x"0c",
          7314 => x"51",
          7315 => x"84",
          7316 => x"c8",
          7317 => x"38",
          7318 => x"51",
          7319 => x"82",
          7320 => x"83",
          7321 => x"54",
          7322 => x"82",
          7323 => x"09",
          7324 => x"e3",
          7325 => x"b8",
          7326 => x"57",
          7327 => x"2e",
          7328 => x"83",
          7329 => x"74",
          7330 => x"70",
          7331 => x"25",
          7332 => x"51",
          7333 => x"38",
          7334 => x"2e",
          7335 => x"b5",
          7336 => x"82",
          7337 => x"80",
          7338 => x"cf",
          7339 => x"d8",
          7340 => x"82",
          7341 => x"80",
          7342 => x"85",
          7343 => x"84",
          7344 => x"16",
          7345 => x"3f",
          7346 => x"08",
          7347 => x"c8",
          7348 => x"83",
          7349 => x"74",
          7350 => x"0c",
          7351 => x"04",
          7352 => x"61",
          7353 => x"80",
          7354 => x"58",
          7355 => x"0c",
          7356 => x"e1",
          7357 => x"c8",
          7358 => x"56",
          7359 => x"d8",
          7360 => x"87",
          7361 => x"d8",
          7362 => x"29",
          7363 => x"05",
          7364 => x"53",
          7365 => x"80",
          7366 => x"38",
          7367 => x"76",
          7368 => x"74",
          7369 => x"72",
          7370 => x"38",
          7371 => x"51",
          7372 => x"82",
          7373 => x"81",
          7374 => x"81",
          7375 => x"72",
          7376 => x"80",
          7377 => x"38",
          7378 => x"70",
          7379 => x"53",
          7380 => x"86",
          7381 => x"af",
          7382 => x"34",
          7383 => x"34",
          7384 => x"14",
          7385 => x"88",
          7386 => x"c8",
          7387 => x"06",
          7388 => x"54",
          7389 => x"72",
          7390 => x"76",
          7391 => x"38",
          7392 => x"70",
          7393 => x"53",
          7394 => x"85",
          7395 => x"70",
          7396 => x"5b",
          7397 => x"82",
          7398 => x"81",
          7399 => x"76",
          7400 => x"81",
          7401 => x"38",
          7402 => x"56",
          7403 => x"83",
          7404 => x"70",
          7405 => x"80",
          7406 => x"83",
          7407 => x"cb",
          7408 => x"d8",
          7409 => x"76",
          7410 => x"05",
          7411 => x"16",
          7412 => x"56",
          7413 => x"d7",
          7414 => x"8d",
          7415 => x"72",
          7416 => x"54",
          7417 => x"57",
          7418 => x"95",
          7419 => x"73",
          7420 => x"3f",
          7421 => x"08",
          7422 => x"57",
          7423 => x"89",
          7424 => x"56",
          7425 => x"d7",
          7426 => x"76",
          7427 => x"f9",
          7428 => x"76",
          7429 => x"f1",
          7430 => x"14",
          7431 => x"3f",
          7432 => x"08",
          7433 => x"06",
          7434 => x"80",
          7435 => x"06",
          7436 => x"80",
          7437 => x"ca",
          7438 => x"d8",
          7439 => x"ff",
          7440 => x"77",
          7441 => x"dc",
          7442 => x"b3",
          7443 => x"c8",
          7444 => x"a0",
          7445 => x"c8",
          7446 => x"15",
          7447 => x"14",
          7448 => x"70",
          7449 => x"51",
          7450 => x"56",
          7451 => x"84",
          7452 => x"81",
          7453 => x"71",
          7454 => x"16",
          7455 => x"53",
          7456 => x"23",
          7457 => x"8b",
          7458 => x"73",
          7459 => x"80",
          7460 => x"8d",
          7461 => x"39",
          7462 => x"51",
          7463 => x"82",
          7464 => x"53",
          7465 => x"08",
          7466 => x"72",
          7467 => x"8d",
          7468 => x"d5",
          7469 => x"14",
          7470 => x"3f",
          7471 => x"08",
          7472 => x"06",
          7473 => x"38",
          7474 => x"51",
          7475 => x"82",
          7476 => x"55",
          7477 => x"51",
          7478 => x"82",
          7479 => x"83",
          7480 => x"53",
          7481 => x"80",
          7482 => x"38",
          7483 => x"78",
          7484 => x"2a",
          7485 => x"78",
          7486 => x"8d",
          7487 => x"22",
          7488 => x"31",
          7489 => x"fc",
          7490 => x"c8",
          7491 => x"d8",
          7492 => x"2e",
          7493 => x"82",
          7494 => x"80",
          7495 => x"f5",
          7496 => x"83",
          7497 => x"ff",
          7498 => x"38",
          7499 => x"9f",
          7500 => x"38",
          7501 => x"39",
          7502 => x"80",
          7503 => x"38",
          7504 => x"9c",
          7505 => x"a4",
          7506 => x"1c",
          7507 => x"0c",
          7508 => x"17",
          7509 => x"76",
          7510 => x"81",
          7511 => x"80",
          7512 => x"c8",
          7513 => x"d8",
          7514 => x"ff",
          7515 => x"8d",
          7516 => x"95",
          7517 => x"91",
          7518 => x"14",
          7519 => x"3f",
          7520 => x"08",
          7521 => x"74",
          7522 => x"a2",
          7523 => x"79",
          7524 => x"f5",
          7525 => x"ac",
          7526 => x"15",
          7527 => x"2e",
          7528 => x"10",
          7529 => x"2a",
          7530 => x"05",
          7531 => x"ff",
          7532 => x"53",
          7533 => x"a0",
          7534 => x"81",
          7535 => x"0b",
          7536 => x"ff",
          7537 => x"0c",
          7538 => x"84",
          7539 => x"83",
          7540 => x"06",
          7541 => x"80",
          7542 => x"c7",
          7543 => x"d8",
          7544 => x"ff",
          7545 => x"72",
          7546 => x"81",
          7547 => x"38",
          7548 => x"73",
          7549 => x"3f",
          7550 => x"08",
          7551 => x"82",
          7552 => x"84",
          7553 => x"b6",
          7554 => x"dc",
          7555 => x"c8",
          7556 => x"ff",
          7557 => x"82",
          7558 => x"09",
          7559 => x"c8",
          7560 => x"51",
          7561 => x"82",
          7562 => x"84",
          7563 => x"d2",
          7564 => x"06",
          7565 => x"9c",
          7566 => x"c3",
          7567 => x"c8",
          7568 => x"85",
          7569 => x"09",
          7570 => x"38",
          7571 => x"51",
          7572 => x"82",
          7573 => x"94",
          7574 => x"a4",
          7575 => x"9f",
          7576 => x"c8",
          7577 => x"0c",
          7578 => x"82",
          7579 => x"81",
          7580 => x"82",
          7581 => x"72",
          7582 => x"82",
          7583 => x"8c",
          7584 => x"0b",
          7585 => x"80",
          7586 => x"d8",
          7587 => x"3d",
          7588 => x"3d",
          7589 => x"89",
          7590 => x"2e",
          7591 => x"08",
          7592 => x"2e",
          7593 => x"33",
          7594 => x"2e",
          7595 => x"13",
          7596 => x"22",
          7597 => x"76",
          7598 => x"06",
          7599 => x"13",
          7600 => x"bf",
          7601 => x"d8",
          7602 => x"06",
          7603 => x"38",
          7604 => x"54",
          7605 => x"80",
          7606 => x"71",
          7607 => x"82",
          7608 => x"87",
          7609 => x"fa",
          7610 => x"ab",
          7611 => x"58",
          7612 => x"05",
          7613 => x"dd",
          7614 => x"80",
          7615 => x"c8",
          7616 => x"38",
          7617 => x"08",
          7618 => x"f0",
          7619 => x"08",
          7620 => x"80",
          7621 => x"80",
          7622 => x"54",
          7623 => x"84",
          7624 => x"34",
          7625 => x"75",
          7626 => x"2e",
          7627 => x"53",
          7628 => x"53",
          7629 => x"f7",
          7630 => x"d8",
          7631 => x"73",
          7632 => x"0c",
          7633 => x"04",
          7634 => x"68",
          7635 => x"80",
          7636 => x"59",
          7637 => x"78",
          7638 => x"c8",
          7639 => x"06",
          7640 => x"3d",
          7641 => x"9a",
          7642 => x"52",
          7643 => x"3f",
          7644 => x"08",
          7645 => x"c8",
          7646 => x"38",
          7647 => x"52",
          7648 => x"52",
          7649 => x"3f",
          7650 => x"08",
          7651 => x"c8",
          7652 => x"02",
          7653 => x"33",
          7654 => x"55",
          7655 => x"25",
          7656 => x"55",
          7657 => x"54",
          7658 => x"81",
          7659 => x"80",
          7660 => x"74",
          7661 => x"81",
          7662 => x"75",
          7663 => x"3f",
          7664 => x"08",
          7665 => x"02",
          7666 => x"91",
          7667 => x"81",
          7668 => x"82",
          7669 => x"06",
          7670 => x"80",
          7671 => x"88",
          7672 => x"39",
          7673 => x"58",
          7674 => x"38",
          7675 => x"70",
          7676 => x"54",
          7677 => x"81",
          7678 => x"52",
          7679 => x"b0",
          7680 => x"c8",
          7681 => x"88",
          7682 => x"62",
          7683 => x"c3",
          7684 => x"54",
          7685 => x"15",
          7686 => x"62",
          7687 => x"d7",
          7688 => x"52",
          7689 => x"51",
          7690 => x"7a",
          7691 => x"83",
          7692 => x"80",
          7693 => x"38",
          7694 => x"08",
          7695 => x"53",
          7696 => x"3d",
          7697 => x"cc",
          7698 => x"d8",
          7699 => x"82",
          7700 => x"82",
          7701 => x"39",
          7702 => x"38",
          7703 => x"33",
          7704 => x"70",
          7705 => x"55",
          7706 => x"2e",
          7707 => x"55",
          7708 => x"77",
          7709 => x"81",
          7710 => x"73",
          7711 => x"38",
          7712 => x"54",
          7713 => x"a0",
          7714 => x"82",
          7715 => x"52",
          7716 => x"ae",
          7717 => x"c8",
          7718 => x"18",
          7719 => x"55",
          7720 => x"c8",
          7721 => x"38",
          7722 => x"70",
          7723 => x"54",
          7724 => x"86",
          7725 => x"c0",
          7726 => x"b4",
          7727 => x"1b",
          7728 => x"1b",
          7729 => x"70",
          7730 => x"e4",
          7731 => x"c8",
          7732 => x"c8",
          7733 => x"0c",
          7734 => x"52",
          7735 => x"3f",
          7736 => x"08",
          7737 => x"08",
          7738 => x"77",
          7739 => x"86",
          7740 => x"1a",
          7741 => x"1a",
          7742 => x"91",
          7743 => x"0b",
          7744 => x"80",
          7745 => x"0c",
          7746 => x"70",
          7747 => x"54",
          7748 => x"81",
          7749 => x"d8",
          7750 => x"2e",
          7751 => x"82",
          7752 => x"94",
          7753 => x"17",
          7754 => x"2b",
          7755 => x"57",
          7756 => x"52",
          7757 => x"aa",
          7758 => x"c8",
          7759 => x"d8",
          7760 => x"26",
          7761 => x"55",
          7762 => x"08",
          7763 => x"81",
          7764 => x"79",
          7765 => x"31",
          7766 => x"70",
          7767 => x"25",
          7768 => x"76",
          7769 => x"81",
          7770 => x"55",
          7771 => x"38",
          7772 => x"0c",
          7773 => x"75",
          7774 => x"54",
          7775 => x"a2",
          7776 => x"7a",
          7777 => x"3f",
          7778 => x"08",
          7779 => x"55",
          7780 => x"89",
          7781 => x"c8",
          7782 => x"1a",
          7783 => x"80",
          7784 => x"54",
          7785 => x"c8",
          7786 => x"0d",
          7787 => x"0d",
          7788 => x"64",
          7789 => x"59",
          7790 => x"90",
          7791 => x"52",
          7792 => x"ce",
          7793 => x"c8",
          7794 => x"d8",
          7795 => x"38",
          7796 => x"55",
          7797 => x"86",
          7798 => x"82",
          7799 => x"19",
          7800 => x"55",
          7801 => x"80",
          7802 => x"38",
          7803 => x"0b",
          7804 => x"82",
          7805 => x"39",
          7806 => x"1a",
          7807 => x"82",
          7808 => x"19",
          7809 => x"08",
          7810 => x"7c",
          7811 => x"74",
          7812 => x"2e",
          7813 => x"94",
          7814 => x"83",
          7815 => x"56",
          7816 => x"38",
          7817 => x"22",
          7818 => x"89",
          7819 => x"55",
          7820 => x"75",
          7821 => x"19",
          7822 => x"39",
          7823 => x"52",
          7824 => x"9e",
          7825 => x"c8",
          7826 => x"75",
          7827 => x"38",
          7828 => x"ff",
          7829 => x"98",
          7830 => x"19",
          7831 => x"51",
          7832 => x"82",
          7833 => x"80",
          7834 => x"38",
          7835 => x"08",
          7836 => x"2a",
          7837 => x"80",
          7838 => x"38",
          7839 => x"8a",
          7840 => x"5c",
          7841 => x"27",
          7842 => x"7a",
          7843 => x"54",
          7844 => x"52",
          7845 => x"51",
          7846 => x"3f",
          7847 => x"08",
          7848 => x"7e",
          7849 => x"56",
          7850 => x"2e",
          7851 => x"16",
          7852 => x"55",
          7853 => x"95",
          7854 => x"53",
          7855 => x"b4",
          7856 => x"31",
          7857 => x"05",
          7858 => x"ab",
          7859 => x"2b",
          7860 => x"76",
          7861 => x"94",
          7862 => x"ff",
          7863 => x"71",
          7864 => x"7b",
          7865 => x"38",
          7866 => x"19",
          7867 => x"51",
          7868 => x"82",
          7869 => x"fd",
          7870 => x"53",
          7871 => x"83",
          7872 => x"b8",
          7873 => x"51",
          7874 => x"3f",
          7875 => x"7e",
          7876 => x"0c",
          7877 => x"1b",
          7878 => x"1c",
          7879 => x"fd",
          7880 => x"56",
          7881 => x"c8",
          7882 => x"0d",
          7883 => x"0d",
          7884 => x"64",
          7885 => x"58",
          7886 => x"90",
          7887 => x"52",
          7888 => x"ce",
          7889 => x"c8",
          7890 => x"d8",
          7891 => x"38",
          7892 => x"55",
          7893 => x"86",
          7894 => x"83",
          7895 => x"18",
          7896 => x"2a",
          7897 => x"51",
          7898 => x"56",
          7899 => x"83",
          7900 => x"39",
          7901 => x"19",
          7902 => x"83",
          7903 => x"0b",
          7904 => x"81",
          7905 => x"39",
          7906 => x"7c",
          7907 => x"74",
          7908 => x"38",
          7909 => x"7b",
          7910 => x"f2",
          7911 => x"08",
          7912 => x"06",
          7913 => x"82",
          7914 => x"8a",
          7915 => x"05",
          7916 => x"06",
          7917 => x"bf",
          7918 => x"38",
          7919 => x"55",
          7920 => x"7a",
          7921 => x"98",
          7922 => x"77",
          7923 => x"3f",
          7924 => x"08",
          7925 => x"c8",
          7926 => x"82",
          7927 => x"81",
          7928 => x"38",
          7929 => x"ff",
          7930 => x"98",
          7931 => x"18",
          7932 => x"74",
          7933 => x"7e",
          7934 => x"08",
          7935 => x"2e",
          7936 => x"8e",
          7937 => x"ff",
          7938 => x"82",
          7939 => x"fe",
          7940 => x"18",
          7941 => x"51",
          7942 => x"82",
          7943 => x"80",
          7944 => x"38",
          7945 => x"08",
          7946 => x"2a",
          7947 => x"80",
          7948 => x"38",
          7949 => x"8a",
          7950 => x"5b",
          7951 => x"27",
          7952 => x"7b",
          7953 => x"54",
          7954 => x"52",
          7955 => x"51",
          7956 => x"3f",
          7957 => x"08",
          7958 => x"7e",
          7959 => x"78",
          7960 => x"74",
          7961 => x"38",
          7962 => x"b4",
          7963 => x"31",
          7964 => x"05",
          7965 => x"51",
          7966 => x"3f",
          7967 => x"0b",
          7968 => x"78",
          7969 => x"80",
          7970 => x"18",
          7971 => x"08",
          7972 => x"7e",
          7973 => x"ba",
          7974 => x"c8",
          7975 => x"38",
          7976 => x"12",
          7977 => x"9c",
          7978 => x"18",
          7979 => x"06",
          7980 => x"31",
          7981 => x"76",
          7982 => x"7b",
          7983 => x"08",
          7984 => x"ff",
          7985 => x"82",
          7986 => x"fd",
          7987 => x"53",
          7988 => x"18",
          7989 => x"06",
          7990 => x"51",
          7991 => x"3f",
          7992 => x"0b",
          7993 => x"7b",
          7994 => x"08",
          7995 => x"76",
          7996 => x"08",
          7997 => x"1c",
          7998 => x"08",
          7999 => x"5c",
          8000 => x"83",
          8001 => x"74",
          8002 => x"fd",
          8003 => x"18",
          8004 => x"07",
          8005 => x"19",
          8006 => x"75",
          8007 => x"0c",
          8008 => x"04",
          8009 => x"7a",
          8010 => x"05",
          8011 => x"56",
          8012 => x"82",
          8013 => x"57",
          8014 => x"08",
          8015 => x"90",
          8016 => x"86",
          8017 => x"06",
          8018 => x"73",
          8019 => x"ee",
          8020 => x"08",
          8021 => x"ff",
          8022 => x"82",
          8023 => x"57",
          8024 => x"08",
          8025 => x"a4",
          8026 => x"11",
          8027 => x"55",
          8028 => x"16",
          8029 => x"08",
          8030 => x"75",
          8031 => x"e9",
          8032 => x"08",
          8033 => x"51",
          8034 => x"3f",
          8035 => x"0a",
          8036 => x"51",
          8037 => x"3f",
          8038 => x"15",
          8039 => x"8a",
          8040 => x"81",
          8041 => x"34",
          8042 => x"bb",
          8043 => x"d8",
          8044 => x"17",
          8045 => x"06",
          8046 => x"90",
          8047 => x"82",
          8048 => x"8a",
          8049 => x"fc",
          8050 => x"70",
          8051 => x"d4",
          8052 => x"c8",
          8053 => x"d8",
          8054 => x"38",
          8055 => x"05",
          8056 => x"f1",
          8057 => x"d8",
          8058 => x"82",
          8059 => x"87",
          8060 => x"c8",
          8061 => x"72",
          8062 => x"0c",
          8063 => x"04",
          8064 => x"84",
          8065 => x"cd",
          8066 => x"80",
          8067 => x"c8",
          8068 => x"38",
          8069 => x"08",
          8070 => x"34",
          8071 => x"82",
          8072 => x"83",
          8073 => x"ee",
          8074 => x"53",
          8075 => x"05",
          8076 => x"51",
          8077 => x"82",
          8078 => x"55",
          8079 => x"08",
          8080 => x"76",
          8081 => x"94",
          8082 => x"51",
          8083 => x"82",
          8084 => x"55",
          8085 => x"08",
          8086 => x"80",
          8087 => x"70",
          8088 => x"56",
          8089 => x"89",
          8090 => x"98",
          8091 => x"b2",
          8092 => x"05",
          8093 => x"2a",
          8094 => x"51",
          8095 => x"80",
          8096 => x"76",
          8097 => x"52",
          8098 => x"3f",
          8099 => x"08",
          8100 => x"8e",
          8101 => x"c8",
          8102 => x"09",
          8103 => x"38",
          8104 => x"82",
          8105 => x"94",
          8106 => x"ff",
          8107 => x"80",
          8108 => x"80",
          8109 => x"5b",
          8110 => x"34",
          8111 => x"df",
          8112 => x"05",
          8113 => x"3d",
          8114 => x"3f",
          8115 => x"08",
          8116 => x"c8",
          8117 => x"38",
          8118 => x"3d",
          8119 => x"98",
          8120 => x"d8",
          8121 => x"58",
          8122 => x"08",
          8123 => x"2e",
          8124 => x"a0",
          8125 => x"3d",
          8126 => x"c4",
          8127 => x"d8",
          8128 => x"82",
          8129 => x"82",
          8130 => x"d9",
          8131 => x"7b",
          8132 => x"ae",
          8133 => x"c8",
          8134 => x"d8",
          8135 => x"d8",
          8136 => x"3d",
          8137 => x"51",
          8138 => x"82",
          8139 => x"80",
          8140 => x"76",
          8141 => x"c4",
          8142 => x"d8",
          8143 => x"82",
          8144 => x"82",
          8145 => x"52",
          8146 => x"fa",
          8147 => x"c8",
          8148 => x"d8",
          8149 => x"38",
          8150 => x"08",
          8151 => x"c8",
          8152 => x"82",
          8153 => x"2e",
          8154 => x"52",
          8155 => x"ac",
          8156 => x"c8",
          8157 => x"d8",
          8158 => x"2e",
          8159 => x"84",
          8160 => x"06",
          8161 => x"57",
          8162 => x"76",
          8163 => x"80",
          8164 => x"b8",
          8165 => x"51",
          8166 => x"76",
          8167 => x"11",
          8168 => x"51",
          8169 => x"73",
          8170 => x"38",
          8171 => x"05",
          8172 => x"81",
          8173 => x"56",
          8174 => x"f5",
          8175 => x"54",
          8176 => x"81",
          8177 => x"80",
          8178 => x"78",
          8179 => x"55",
          8180 => x"e1",
          8181 => x"ff",
          8182 => x"58",
          8183 => x"74",
          8184 => x"75",
          8185 => x"18",
          8186 => x"08",
          8187 => x"af",
          8188 => x"f4",
          8189 => x"2e",
          8190 => x"8d",
          8191 => x"80",
          8192 => x"11",
          8193 => x"74",
          8194 => x"82",
          8195 => x"70",
          8196 => x"ca",
          8197 => x"08",
          8198 => x"5c",
          8199 => x"73",
          8200 => x"38",
          8201 => x"1a",
          8202 => x"55",
          8203 => x"38",
          8204 => x"73",
          8205 => x"38",
          8206 => x"76",
          8207 => x"74",
          8208 => x"33",
          8209 => x"05",
          8210 => x"15",
          8211 => x"ba",
          8212 => x"05",
          8213 => x"ff",
          8214 => x"06",
          8215 => x"57",
          8216 => x"e0",
          8217 => x"81",
          8218 => x"73",
          8219 => x"81",
          8220 => x"7a",
          8221 => x"38",
          8222 => x"76",
          8223 => x"0c",
          8224 => x"0d",
          8225 => x"0d",
          8226 => x"3d",
          8227 => x"71",
          8228 => x"eb",
          8229 => x"d8",
          8230 => x"82",
          8231 => x"82",
          8232 => x"15",
          8233 => x"82",
          8234 => x"15",
          8235 => x"76",
          8236 => x"90",
          8237 => x"81",
          8238 => x"06",
          8239 => x"72",
          8240 => x"56",
          8241 => x"54",
          8242 => x"17",
          8243 => x"78",
          8244 => x"38",
          8245 => x"22",
          8246 => x"59",
          8247 => x"78",
          8248 => x"76",
          8249 => x"51",
          8250 => x"3f",
          8251 => x"08",
          8252 => x"54",
          8253 => x"53",
          8254 => x"3f",
          8255 => x"08",
          8256 => x"38",
          8257 => x"75",
          8258 => x"18",
          8259 => x"31",
          8260 => x"57",
          8261 => x"b2",
          8262 => x"08",
          8263 => x"38",
          8264 => x"51",
          8265 => x"3f",
          8266 => x"08",
          8267 => x"c8",
          8268 => x"81",
          8269 => x"d8",
          8270 => x"2e",
          8271 => x"82",
          8272 => x"88",
          8273 => x"98",
          8274 => x"80",
          8275 => x"38",
          8276 => x"80",
          8277 => x"77",
          8278 => x"08",
          8279 => x"0c",
          8280 => x"70",
          8281 => x"81",
          8282 => x"5a",
          8283 => x"2e",
          8284 => x"52",
          8285 => x"bb",
          8286 => x"d8",
          8287 => x"82",
          8288 => x"95",
          8289 => x"c8",
          8290 => x"39",
          8291 => x"51",
          8292 => x"3f",
          8293 => x"08",
          8294 => x"2e",
          8295 => x"74",
          8296 => x"79",
          8297 => x"14",
          8298 => x"38",
          8299 => x"0c",
          8300 => x"94",
          8301 => x"94",
          8302 => x"83",
          8303 => x"72",
          8304 => x"38",
          8305 => x"51",
          8306 => x"3f",
          8307 => x"08",
          8308 => x"0b",
          8309 => x"82",
          8310 => x"39",
          8311 => x"16",
          8312 => x"bb",
          8313 => x"2a",
          8314 => x"08",
          8315 => x"15",
          8316 => x"15",
          8317 => x"90",
          8318 => x"16",
          8319 => x"33",
          8320 => x"53",
          8321 => x"34",
          8322 => x"06",
          8323 => x"2e",
          8324 => x"9c",
          8325 => x"85",
          8326 => x"16",
          8327 => x"72",
          8328 => x"0c",
          8329 => x"04",
          8330 => x"79",
          8331 => x"75",
          8332 => x"8b",
          8333 => x"89",
          8334 => x"52",
          8335 => x"05",
          8336 => x"3f",
          8337 => x"08",
          8338 => x"c8",
          8339 => x"38",
          8340 => x"7a",
          8341 => x"d5",
          8342 => x"d8",
          8343 => x"82",
          8344 => x"80",
          8345 => x"16",
          8346 => x"2b",
          8347 => x"74",
          8348 => x"86",
          8349 => x"84",
          8350 => x"06",
          8351 => x"73",
          8352 => x"38",
          8353 => x"52",
          8354 => x"a4",
          8355 => x"c8",
          8356 => x"0c",
          8357 => x"14",
          8358 => x"23",
          8359 => x"51",
          8360 => x"3f",
          8361 => x"08",
          8362 => x"2e",
          8363 => x"85",
          8364 => x"86",
          8365 => x"2e",
          8366 => x"76",
          8367 => x"73",
          8368 => x"0c",
          8369 => x"04",
          8370 => x"76",
          8371 => x"05",
          8372 => x"53",
          8373 => x"82",
          8374 => x"87",
          8375 => x"c8",
          8376 => x"86",
          8377 => x"fb",
          8378 => x"79",
          8379 => x"05",
          8380 => x"56",
          8381 => x"3f",
          8382 => x"08",
          8383 => x"c8",
          8384 => x"38",
          8385 => x"82",
          8386 => x"52",
          8387 => x"bc",
          8388 => x"d8",
          8389 => x"80",
          8390 => x"d8",
          8391 => x"73",
          8392 => x"3f",
          8393 => x"08",
          8394 => x"c8",
          8395 => x"09",
          8396 => x"38",
          8397 => x"39",
          8398 => x"08",
          8399 => x"52",
          8400 => x"ba",
          8401 => x"73",
          8402 => x"d0",
          8403 => x"c8",
          8404 => x"70",
          8405 => x"07",
          8406 => x"82",
          8407 => x"06",
          8408 => x"54",
          8409 => x"c8",
          8410 => x"0d",
          8411 => x"0d",
          8412 => x"53",
          8413 => x"53",
          8414 => x"56",
          8415 => x"82",
          8416 => x"55",
          8417 => x"08",
          8418 => x"52",
          8419 => x"ea",
          8420 => x"c8",
          8421 => x"d8",
          8422 => x"38",
          8423 => x"05",
          8424 => x"2b",
          8425 => x"80",
          8426 => x"86",
          8427 => x"76",
          8428 => x"38",
          8429 => x"51",
          8430 => x"74",
          8431 => x"0c",
          8432 => x"04",
          8433 => x"63",
          8434 => x"80",
          8435 => x"ec",
          8436 => x"3d",
          8437 => x"3f",
          8438 => x"08",
          8439 => x"c8",
          8440 => x"38",
          8441 => x"73",
          8442 => x"08",
          8443 => x"13",
          8444 => x"58",
          8445 => x"26",
          8446 => x"7c",
          8447 => x"39",
          8448 => x"ce",
          8449 => x"81",
          8450 => x"d8",
          8451 => x"33",
          8452 => x"81",
          8453 => x"06",
          8454 => x"82",
          8455 => x"76",
          8456 => x"f0",
          8457 => x"b0",
          8458 => x"d8",
          8459 => x"2e",
          8460 => x"d8",
          8461 => x"2e",
          8462 => x"d8",
          8463 => x"70",
          8464 => x"08",
          8465 => x"7a",
          8466 => x"7f",
          8467 => x"54",
          8468 => x"77",
          8469 => x"80",
          8470 => x"15",
          8471 => x"c8",
          8472 => x"75",
          8473 => x"52",
          8474 => x"52",
          8475 => x"d2",
          8476 => x"c8",
          8477 => x"d8",
          8478 => x"d6",
          8479 => x"33",
          8480 => x"1a",
          8481 => x"54",
          8482 => x"09",
          8483 => x"38",
          8484 => x"ff",
          8485 => x"82",
          8486 => x"83",
          8487 => x"70",
          8488 => x"25",
          8489 => x"59",
          8490 => x"9b",
          8491 => x"51",
          8492 => x"3f",
          8493 => x"08",
          8494 => x"70",
          8495 => x"25",
          8496 => x"59",
          8497 => x"75",
          8498 => x"7a",
          8499 => x"ff",
          8500 => x"7c",
          8501 => x"94",
          8502 => x"11",
          8503 => x"56",
          8504 => x"15",
          8505 => x"d8",
          8506 => x"3d",
          8507 => x"3d",
          8508 => x"3d",
          8509 => x"70",
          8510 => x"96",
          8511 => x"c8",
          8512 => x"d8",
          8513 => x"aa",
          8514 => x"33",
          8515 => x"a2",
          8516 => x"33",
          8517 => x"70",
          8518 => x"55",
          8519 => x"73",
          8520 => x"90",
          8521 => x"08",
          8522 => x"18",
          8523 => x"82",
          8524 => x"38",
          8525 => x"08",
          8526 => x"08",
          8527 => x"ff",
          8528 => x"82",
          8529 => x"74",
          8530 => x"56",
          8531 => x"98",
          8532 => x"76",
          8533 => x"8a",
          8534 => x"c8",
          8535 => x"09",
          8536 => x"38",
          8537 => x"d8",
          8538 => x"2e",
          8539 => x"85",
          8540 => x"a4",
          8541 => x"38",
          8542 => x"d8",
          8543 => x"15",
          8544 => x"38",
          8545 => x"53",
          8546 => x"08",
          8547 => x"ff",
          8548 => x"82",
          8549 => x"56",
          8550 => x"8c",
          8551 => x"17",
          8552 => x"07",
          8553 => x"18",
          8554 => x"2e",
          8555 => x"91",
          8556 => x"55",
          8557 => x"c8",
          8558 => x"0d",
          8559 => x"0d",
          8560 => x"3d",
          8561 => x"52",
          8562 => x"da",
          8563 => x"d8",
          8564 => x"82",
          8565 => x"81",
          8566 => x"46",
          8567 => x"52",
          8568 => x"52",
          8569 => x"3f",
          8570 => x"08",
          8571 => x"c8",
          8572 => x"38",
          8573 => x"05",
          8574 => x"2a",
          8575 => x"51",
          8576 => x"55",
          8577 => x"38",
          8578 => x"54",
          8579 => x"81",
          8580 => x"80",
          8581 => x"70",
          8582 => x"54",
          8583 => x"81",
          8584 => x"52",
          8585 => x"bb",
          8586 => x"d8",
          8587 => x"84",
          8588 => x"06",
          8589 => x"73",
          8590 => x"d6",
          8591 => x"82",
          8592 => x"98",
          8593 => x"81",
          8594 => x"5a",
          8595 => x"08",
          8596 => x"8a",
          8597 => x"54",
          8598 => x"3f",
          8599 => x"08",
          8600 => x"c8",
          8601 => x"38",
          8602 => x"08",
          8603 => x"ff",
          8604 => x"82",
          8605 => x"55",
          8606 => x"08",
          8607 => x"55",
          8608 => x"82",
          8609 => x"84",
          8610 => x"82",
          8611 => x"80",
          8612 => x"51",
          8613 => x"82",
          8614 => x"82",
          8615 => x"30",
          8616 => x"c8",
          8617 => x"25",
          8618 => x"75",
          8619 => x"38",
          8620 => x"90",
          8621 => x"75",
          8622 => x"ff",
          8623 => x"82",
          8624 => x"55",
          8625 => x"78",
          8626 => x"bd",
          8627 => x"c8",
          8628 => x"82",
          8629 => x"a2",
          8630 => x"e8",
          8631 => x"53",
          8632 => x"bc",
          8633 => x"3d",
          8634 => x"3f",
          8635 => x"08",
          8636 => x"c8",
          8637 => x"38",
          8638 => x"52",
          8639 => x"52",
          8640 => x"3f",
          8641 => x"08",
          8642 => x"c8",
          8643 => x"88",
          8644 => x"39",
          8645 => x"08",
          8646 => x"81",
          8647 => x"38",
          8648 => x"05",
          8649 => x"2a",
          8650 => x"55",
          8651 => x"81",
          8652 => x"5a",
          8653 => x"3d",
          8654 => x"ff",
          8655 => x"82",
          8656 => x"75",
          8657 => x"d8",
          8658 => x"38",
          8659 => x"d8",
          8660 => x"2e",
          8661 => x"83",
          8662 => x"82",
          8663 => x"ff",
          8664 => x"06",
          8665 => x"54",
          8666 => x"73",
          8667 => x"82",
          8668 => x"52",
          8669 => x"b2",
          8670 => x"d8",
          8671 => x"82",
          8672 => x"81",
          8673 => x"53",
          8674 => x"19",
          8675 => x"8a",
          8676 => x"ae",
          8677 => x"34",
          8678 => x"0b",
          8679 => x"34",
          8680 => x"0a",
          8681 => x"19",
          8682 => x"9c",
          8683 => x"78",
          8684 => x"51",
          8685 => x"3f",
          8686 => x"b8",
          8687 => x"d8",
          8688 => x"a4",
          8689 => x"54",
          8690 => x"d9",
          8691 => x"53",
          8692 => x"11",
          8693 => x"b8",
          8694 => x"54",
          8695 => x"15",
          8696 => x"ff",
          8697 => x"82",
          8698 => x"54",
          8699 => x"08",
          8700 => x"88",
          8701 => x"64",
          8702 => x"ff",
          8703 => x"75",
          8704 => x"78",
          8705 => x"e1",
          8706 => x"90",
          8707 => x"34",
          8708 => x"0b",
          8709 => x"78",
          8710 => x"ed",
          8711 => x"c8",
          8712 => x"39",
          8713 => x"52",
          8714 => x"ac",
          8715 => x"82",
          8716 => x"9a",
          8717 => x"d8",
          8718 => x"3d",
          8719 => x"d2",
          8720 => x"53",
          8721 => x"fc",
          8722 => x"3d",
          8723 => x"3f",
          8724 => x"08",
          8725 => x"c8",
          8726 => x"38",
          8727 => x"3d",
          8728 => x"3d",
          8729 => x"c9",
          8730 => x"d8",
          8731 => x"82",
          8732 => x"82",
          8733 => x"81",
          8734 => x"81",
          8735 => x"86",
          8736 => x"af",
          8737 => x"a5",
          8738 => x"aa",
          8739 => x"05",
          8740 => x"e3",
          8741 => x"77",
          8742 => x"70",
          8743 => x"a2",
          8744 => x"3d",
          8745 => x"51",
          8746 => x"82",
          8747 => x"55",
          8748 => x"08",
          8749 => x"a1",
          8750 => x"09",
          8751 => x"38",
          8752 => x"08",
          8753 => x"88",
          8754 => x"39",
          8755 => x"08",
          8756 => x"81",
          8757 => x"38",
          8758 => x"bd",
          8759 => x"d8",
          8760 => x"82",
          8761 => x"81",
          8762 => x"56",
          8763 => x"3d",
          8764 => x"52",
          8765 => x"ff",
          8766 => x"02",
          8767 => x"8b",
          8768 => x"16",
          8769 => x"2a",
          8770 => x"51",
          8771 => x"89",
          8772 => x"07",
          8773 => x"17",
          8774 => x"81",
          8775 => x"34",
          8776 => x"70",
          8777 => x"81",
          8778 => x"55",
          8779 => x"80",
          8780 => x"64",
          8781 => x"38",
          8782 => x"51",
          8783 => x"3f",
          8784 => x"08",
          8785 => x"ff",
          8786 => x"82",
          8787 => x"c8",
          8788 => x"80",
          8789 => x"d8",
          8790 => x"78",
          8791 => x"e2",
          8792 => x"c8",
          8793 => x"d8",
          8794 => x"55",
          8795 => x"08",
          8796 => x"81",
          8797 => x"73",
          8798 => x"81",
          8799 => x"63",
          8800 => x"76",
          8801 => x"e1",
          8802 => x"81",
          8803 => x"34",
          8804 => x"d8",
          8805 => x"38",
          8806 => x"e9",
          8807 => x"c8",
          8808 => x"d8",
          8809 => x"38",
          8810 => x"a3",
          8811 => x"d8",
          8812 => x"74",
          8813 => x"0c",
          8814 => x"04",
          8815 => x"02",
          8816 => x"33",
          8817 => x"80",
          8818 => x"57",
          8819 => x"96",
          8820 => x"52",
          8821 => x"d2",
          8822 => x"d8",
          8823 => x"82",
          8824 => x"80",
          8825 => x"5a",
          8826 => x"3d",
          8827 => x"c6",
          8828 => x"d8",
          8829 => x"82",
          8830 => x"b8",
          8831 => x"cf",
          8832 => x"a0",
          8833 => x"55",
          8834 => x"75",
          8835 => x"71",
          8836 => x"33",
          8837 => x"74",
          8838 => x"57",
          8839 => x"8b",
          8840 => x"54",
          8841 => x"15",
          8842 => x"ff",
          8843 => x"82",
          8844 => x"55",
          8845 => x"c8",
          8846 => x"0d",
          8847 => x"0d",
          8848 => x"53",
          8849 => x"05",
          8850 => x"51",
          8851 => x"82",
          8852 => x"55",
          8853 => x"08",
          8854 => x"76",
          8855 => x"94",
          8856 => x"51",
          8857 => x"82",
          8858 => x"55",
          8859 => x"08",
          8860 => x"80",
          8861 => x"81",
          8862 => x"86",
          8863 => x"38",
          8864 => x"86",
          8865 => x"90",
          8866 => x"54",
          8867 => x"ff",
          8868 => x"76",
          8869 => x"83",
          8870 => x"51",
          8871 => x"3f",
          8872 => x"08",
          8873 => x"d8",
          8874 => x"3d",
          8875 => x"3d",
          8876 => x"5c",
          8877 => x"99",
          8878 => x"52",
          8879 => x"d0",
          8880 => x"d8",
          8881 => x"d8",
          8882 => x"70",
          8883 => x"08",
          8884 => x"51",
          8885 => x"80",
          8886 => x"38",
          8887 => x"06",
          8888 => x"80",
          8889 => x"38",
          8890 => x"5f",
          8891 => x"3d",
          8892 => x"ff",
          8893 => x"82",
          8894 => x"57",
          8895 => x"08",
          8896 => x"74",
          8897 => x"ff",
          8898 => x"82",
          8899 => x"57",
          8900 => x"08",
          8901 => x"d8",
          8902 => x"d8",
          8903 => x"5b",
          8904 => x"18",
          8905 => x"18",
          8906 => x"74",
          8907 => x"81",
          8908 => x"78",
          8909 => x"8b",
          8910 => x"54",
          8911 => x"75",
          8912 => x"38",
          8913 => x"1b",
          8914 => x"55",
          8915 => x"2e",
          8916 => x"39",
          8917 => x"09",
          8918 => x"38",
          8919 => x"80",
          8920 => x"70",
          8921 => x"25",
          8922 => x"80",
          8923 => x"38",
          8924 => x"bc",
          8925 => x"11",
          8926 => x"ff",
          8927 => x"82",
          8928 => x"57",
          8929 => x"08",
          8930 => x"70",
          8931 => x"80",
          8932 => x"83",
          8933 => x"80",
          8934 => x"84",
          8935 => x"a7",
          8936 => x"b8",
          8937 => x"9b",
          8938 => x"d8",
          8939 => x"0c",
          8940 => x"c8",
          8941 => x"0d",
          8942 => x"0d",
          8943 => x"3d",
          8944 => x"52",
          8945 => x"ce",
          8946 => x"d8",
          8947 => x"d8",
          8948 => x"54",
          8949 => x"08",
          8950 => x"8b",
          8951 => x"8a",
          8952 => x"58",
          8953 => x"3f",
          8954 => x"33",
          8955 => x"9f",
          8956 => x"86",
          8957 => x"9d",
          8958 => x"9d",
          8959 => x"d8",
          8960 => x"ff",
          8961 => x"c4",
          8962 => x"c8",
          8963 => x"98",
          8964 => x"52",
          8965 => x"08",
          8966 => x"3f",
          8967 => x"08",
          8968 => x"06",
          8969 => x"2e",
          8970 => x"52",
          8971 => x"51",
          8972 => x"3f",
          8973 => x"08",
          8974 => x"ff",
          8975 => x"38",
          8976 => x"88",
          8977 => x"8a",
          8978 => x"38",
          8979 => x"e7",
          8980 => x"75",
          8981 => x"74",
          8982 => x"73",
          8983 => x"05",
          8984 => x"16",
          8985 => x"70",
          8986 => x"34",
          8987 => x"70",
          8988 => x"56",
          8989 => x"fe",
          8990 => x"3d",
          8991 => x"55",
          8992 => x"2e",
          8993 => x"75",
          8994 => x"38",
          8995 => x"55",
          8996 => x"33",
          8997 => x"a0",
          8998 => x"06",
          8999 => x"16",
          9000 => x"38",
          9001 => x"42",
          9002 => x"3d",
          9003 => x"ff",
          9004 => x"82",
          9005 => x"54",
          9006 => x"08",
          9007 => x"81",
          9008 => x"ff",
          9009 => x"82",
          9010 => x"54",
          9011 => x"08",
          9012 => x"80",
          9013 => x"54",
          9014 => x"80",
          9015 => x"d8",
          9016 => x"2e",
          9017 => x"80",
          9018 => x"54",
          9019 => x"80",
          9020 => x"52",
          9021 => x"ac",
          9022 => x"d8",
          9023 => x"82",
          9024 => x"b1",
          9025 => x"82",
          9026 => x"52",
          9027 => x"9a",
          9028 => x"54",
          9029 => x"15",
          9030 => x"77",
          9031 => x"ff",
          9032 => x"78",
          9033 => x"83",
          9034 => x"51",
          9035 => x"3f",
          9036 => x"08",
          9037 => x"74",
          9038 => x"0c",
          9039 => x"04",
          9040 => x"60",
          9041 => x"05",
          9042 => x"33",
          9043 => x"05",
          9044 => x"40",
          9045 => x"ba",
          9046 => x"c8",
          9047 => x"d8",
          9048 => x"bd",
          9049 => x"33",
          9050 => x"b5",
          9051 => x"2e",
          9052 => x"1a",
          9053 => x"90",
          9054 => x"33",
          9055 => x"70",
          9056 => x"55",
          9057 => x"38",
          9058 => x"97",
          9059 => x"82",
          9060 => x"58",
          9061 => x"7e",
          9062 => x"70",
          9063 => x"55",
          9064 => x"56",
          9065 => x"dc",
          9066 => x"7d",
          9067 => x"70",
          9068 => x"2a",
          9069 => x"08",
          9070 => x"08",
          9071 => x"5d",
          9072 => x"77",
          9073 => x"9c",
          9074 => x"26",
          9075 => x"57",
          9076 => x"59",
          9077 => x"52",
          9078 => x"9d",
          9079 => x"15",
          9080 => x"9c",
          9081 => x"26",
          9082 => x"55",
          9083 => x"08",
          9084 => x"99",
          9085 => x"c8",
          9086 => x"ff",
          9087 => x"d8",
          9088 => x"38",
          9089 => x"75",
          9090 => x"81",
          9091 => x"93",
          9092 => x"80",
          9093 => x"2e",
          9094 => x"ff",
          9095 => x"58",
          9096 => x"7d",
          9097 => x"38",
          9098 => x"55",
          9099 => x"b4",
          9100 => x"56",
          9101 => x"09",
          9102 => x"38",
          9103 => x"53",
          9104 => x"51",
          9105 => x"3f",
          9106 => x"08",
          9107 => x"c8",
          9108 => x"38",
          9109 => x"ff",
          9110 => x"5c",
          9111 => x"84",
          9112 => x"5c",
          9113 => x"12",
          9114 => x"80",
          9115 => x"78",
          9116 => x"7c",
          9117 => x"90",
          9118 => x"c0",
          9119 => x"90",
          9120 => x"15",
          9121 => x"94",
          9122 => x"54",
          9123 => x"91",
          9124 => x"31",
          9125 => x"84",
          9126 => x"07",
          9127 => x"16",
          9128 => x"73",
          9129 => x"0c",
          9130 => x"04",
          9131 => x"6b",
          9132 => x"05",
          9133 => x"33",
          9134 => x"5a",
          9135 => x"95",
          9136 => x"80",
          9137 => x"c8",
          9138 => x"f8",
          9139 => x"c8",
          9140 => x"82",
          9141 => x"70",
          9142 => x"74",
          9143 => x"38",
          9144 => x"82",
          9145 => x"81",
          9146 => x"81",
          9147 => x"ff",
          9148 => x"82",
          9149 => x"81",
          9150 => x"81",
          9151 => x"83",
          9152 => x"c0",
          9153 => x"2a",
          9154 => x"51",
          9155 => x"74",
          9156 => x"99",
          9157 => x"53",
          9158 => x"51",
          9159 => x"3f",
          9160 => x"08",
          9161 => x"55",
          9162 => x"92",
          9163 => x"80",
          9164 => x"38",
          9165 => x"06",
          9166 => x"2e",
          9167 => x"48",
          9168 => x"87",
          9169 => x"79",
          9170 => x"78",
          9171 => x"26",
          9172 => x"19",
          9173 => x"74",
          9174 => x"38",
          9175 => x"e4",
          9176 => x"2a",
          9177 => x"70",
          9178 => x"59",
          9179 => x"7a",
          9180 => x"56",
          9181 => x"80",
          9182 => x"51",
          9183 => x"74",
          9184 => x"99",
          9185 => x"53",
          9186 => x"51",
          9187 => x"3f",
          9188 => x"d8",
          9189 => x"ac",
          9190 => x"2a",
          9191 => x"82",
          9192 => x"43",
          9193 => x"83",
          9194 => x"66",
          9195 => x"60",
          9196 => x"90",
          9197 => x"31",
          9198 => x"80",
          9199 => x"8a",
          9200 => x"56",
          9201 => x"26",
          9202 => x"77",
          9203 => x"81",
          9204 => x"74",
          9205 => x"38",
          9206 => x"55",
          9207 => x"83",
          9208 => x"81",
          9209 => x"80",
          9210 => x"38",
          9211 => x"55",
          9212 => x"5e",
          9213 => x"89",
          9214 => x"5a",
          9215 => x"09",
          9216 => x"e1",
          9217 => x"38",
          9218 => x"57",
          9219 => x"cc",
          9220 => x"5a",
          9221 => x"9d",
          9222 => x"26",
          9223 => x"cc",
          9224 => x"10",
          9225 => x"22",
          9226 => x"74",
          9227 => x"38",
          9228 => x"ee",
          9229 => x"66",
          9230 => x"c8",
          9231 => x"c8",
          9232 => x"84",
          9233 => x"89",
          9234 => x"a0",
          9235 => x"82",
          9236 => x"fc",
          9237 => x"56",
          9238 => x"f0",
          9239 => x"80",
          9240 => x"d3",
          9241 => x"38",
          9242 => x"57",
          9243 => x"cb",
          9244 => x"5a",
          9245 => x"9d",
          9246 => x"26",
          9247 => x"cb",
          9248 => x"10",
          9249 => x"22",
          9250 => x"74",
          9251 => x"38",
          9252 => x"ee",
          9253 => x"66",
          9254 => x"e8",
          9255 => x"c8",
          9256 => x"05",
          9257 => x"c8",
          9258 => x"26",
          9259 => x"0b",
          9260 => x"08",
          9261 => x"c8",
          9262 => x"11",
          9263 => x"05",
          9264 => x"83",
          9265 => x"2a",
          9266 => x"a0",
          9267 => x"7d",
          9268 => x"69",
          9269 => x"05",
          9270 => x"72",
          9271 => x"5c",
          9272 => x"59",
          9273 => x"2e",
          9274 => x"89",
          9275 => x"60",
          9276 => x"84",
          9277 => x"5d",
          9278 => x"18",
          9279 => x"68",
          9280 => x"74",
          9281 => x"af",
          9282 => x"31",
          9283 => x"53",
          9284 => x"52",
          9285 => x"ec",
          9286 => x"c8",
          9287 => x"83",
          9288 => x"06",
          9289 => x"d8",
          9290 => x"ff",
          9291 => x"dd",
          9292 => x"83",
          9293 => x"2a",
          9294 => x"be",
          9295 => x"39",
          9296 => x"09",
          9297 => x"c5",
          9298 => x"f5",
          9299 => x"c8",
          9300 => x"38",
          9301 => x"79",
          9302 => x"80",
          9303 => x"38",
          9304 => x"96",
          9305 => x"06",
          9306 => x"2e",
          9307 => x"5e",
          9308 => x"82",
          9309 => x"9f",
          9310 => x"38",
          9311 => x"38",
          9312 => x"81",
          9313 => x"fc",
          9314 => x"ab",
          9315 => x"7d",
          9316 => x"81",
          9317 => x"7d",
          9318 => x"78",
          9319 => x"74",
          9320 => x"8e",
          9321 => x"9c",
          9322 => x"53",
          9323 => x"51",
          9324 => x"3f",
          9325 => x"ca",
          9326 => x"51",
          9327 => x"3f",
          9328 => x"8b",
          9329 => x"8f",
          9330 => x"8d",
          9331 => x"83",
          9332 => x"52",
          9333 => x"ff",
          9334 => x"81",
          9335 => x"34",
          9336 => x"70",
          9337 => x"2a",
          9338 => x"54",
          9339 => x"1b",
          9340 => x"b6",
          9341 => x"74",
          9342 => x"26",
          9343 => x"83",
          9344 => x"52",
          9345 => x"ff",
          9346 => x"8a",
          9347 => x"a0",
          9348 => x"8f",
          9349 => x"0b",
          9350 => x"bf",
          9351 => x"51",
          9352 => x"3f",
          9353 => x"9a",
          9354 => x"8e",
          9355 => x"52",
          9356 => x"ff",
          9357 => x"7d",
          9358 => x"81",
          9359 => x"38",
          9360 => x"0a",
          9361 => x"1b",
          9362 => x"fc",
          9363 => x"a4",
          9364 => x"8e",
          9365 => x"52",
          9366 => x"ff",
          9367 => x"81",
          9368 => x"51",
          9369 => x"3f",
          9370 => x"1b",
          9371 => x"ba",
          9372 => x"0b",
          9373 => x"34",
          9374 => x"c2",
          9375 => x"53",
          9376 => x"52",
          9377 => x"51",
          9378 => x"88",
          9379 => x"a7",
          9380 => x"8e",
          9381 => x"83",
          9382 => x"52",
          9383 => x"ff",
          9384 => x"ff",
          9385 => x"1c",
          9386 => x"a6",
          9387 => x"53",
          9388 => x"52",
          9389 => x"ff",
          9390 => x"82",
          9391 => x"83",
          9392 => x"52",
          9393 => x"e2",
          9394 => x"60",
          9395 => x"7e",
          9396 => x"85",
          9397 => x"82",
          9398 => x"83",
          9399 => x"83",
          9400 => x"06",
          9401 => x"75",
          9402 => x"05",
          9403 => x"7e",
          9404 => x"e5",
          9405 => x"53",
          9406 => x"51",
          9407 => x"3f",
          9408 => x"a4",
          9409 => x"51",
          9410 => x"3f",
          9411 => x"e4",
          9412 => x"e4",
          9413 => x"8d",
          9414 => x"18",
          9415 => x"1b",
          9416 => x"a4",
          9417 => x"83",
          9418 => x"ff",
          9419 => x"82",
          9420 => x"78",
          9421 => x"f2",
          9422 => x"60",
          9423 => x"7a",
          9424 => x"ff",
          9425 => x"75",
          9426 => x"53",
          9427 => x"51",
          9428 => x"3f",
          9429 => x"52",
          9430 => x"8d",
          9431 => x"56",
          9432 => x"83",
          9433 => x"06",
          9434 => x"52",
          9435 => x"8c",
          9436 => x"52",
          9437 => x"ff",
          9438 => x"f0",
          9439 => x"1b",
          9440 => x"87",
          9441 => x"55",
          9442 => x"83",
          9443 => x"74",
          9444 => x"ff",
          9445 => x"7c",
          9446 => x"74",
          9447 => x"38",
          9448 => x"54",
          9449 => x"52",
          9450 => x"88",
          9451 => x"d8",
          9452 => x"87",
          9453 => x"53",
          9454 => x"08",
          9455 => x"ff",
          9456 => x"76",
          9457 => x"31",
          9458 => x"cd",
          9459 => x"58",
          9460 => x"ff",
          9461 => x"55",
          9462 => x"83",
          9463 => x"61",
          9464 => x"26",
          9465 => x"57",
          9466 => x"53",
          9467 => x"51",
          9468 => x"3f",
          9469 => x"08",
          9470 => x"76",
          9471 => x"31",
          9472 => x"db",
          9473 => x"7d",
          9474 => x"38",
          9475 => x"83",
          9476 => x"8a",
          9477 => x"7d",
          9478 => x"38",
          9479 => x"81",
          9480 => x"80",
          9481 => x"80",
          9482 => x"7a",
          9483 => x"ea",
          9484 => x"d5",
          9485 => x"ff",
          9486 => x"83",
          9487 => x"77",
          9488 => x"0b",
          9489 => x"81",
          9490 => x"34",
          9491 => x"34",
          9492 => x"34",
          9493 => x"56",
          9494 => x"52",
          9495 => x"9e",
          9496 => x"0b",
          9497 => x"82",
          9498 => x"82",
          9499 => x"56",
          9500 => x"34",
          9501 => x"08",
          9502 => x"60",
          9503 => x"1b",
          9504 => x"c4",
          9505 => x"83",
          9506 => x"ff",
          9507 => x"81",
          9508 => x"7a",
          9509 => x"ff",
          9510 => x"81",
          9511 => x"c8",
          9512 => x"80",
          9513 => x"7e",
          9514 => x"91",
          9515 => x"82",
          9516 => x"90",
          9517 => x"8e",
          9518 => x"81",
          9519 => x"82",
          9520 => x"56",
          9521 => x"c8",
          9522 => x"0d",
          9523 => x"0d",
          9524 => x"59",
          9525 => x"ff",
          9526 => x"57",
          9527 => x"b4",
          9528 => x"f8",
          9529 => x"81",
          9530 => x"52",
          9531 => x"bd",
          9532 => x"2e",
          9533 => x"9c",
          9534 => x"33",
          9535 => x"2e",
          9536 => x"76",
          9537 => x"58",
          9538 => x"57",
          9539 => x"09",
          9540 => x"38",
          9541 => x"78",
          9542 => x"38",
          9543 => x"82",
          9544 => x"8d",
          9545 => x"f7",
          9546 => x"02",
          9547 => x"05",
          9548 => x"77",
          9549 => x"81",
          9550 => x"8d",
          9551 => x"e7",
          9552 => x"08",
          9553 => x"24",
          9554 => x"17",
          9555 => x"8c",
          9556 => x"77",
          9557 => x"16",
          9558 => x"25",
          9559 => x"3d",
          9560 => x"75",
          9561 => x"52",
          9562 => x"cb",
          9563 => x"76",
          9564 => x"70",
          9565 => x"2a",
          9566 => x"51",
          9567 => x"84",
          9568 => x"19",
          9569 => x"8b",
          9570 => x"f9",
          9571 => x"84",
          9572 => x"56",
          9573 => x"a7",
          9574 => x"fc",
          9575 => x"53",
          9576 => x"75",
          9577 => x"85",
          9578 => x"c8",
          9579 => x"84",
          9580 => x"2e",
          9581 => x"87",
          9582 => x"08",
          9583 => x"ff",
          9584 => x"d8",
          9585 => x"3d",
          9586 => x"3d",
          9587 => x"80",
          9588 => x"52",
          9589 => x"88",
          9590 => x"74",
          9591 => x"0d",
          9592 => x"0d",
          9593 => x"05",
          9594 => x"86",
          9595 => x"54",
          9596 => x"73",
          9597 => x"fe",
          9598 => x"51",
          9599 => x"98",
          9600 => x"fd",
          9601 => x"02",
          9602 => x"05",
          9603 => x"80",
          9604 => x"ff",
          9605 => x"72",
          9606 => x"06",
          9607 => x"39",
          9608 => x"73",
          9609 => x"83",
          9610 => x"81",
          9611 => x"70",
          9612 => x"38",
          9613 => x"22",
          9614 => x"2e",
          9615 => x"12",
          9616 => x"ff",
          9617 => x"71",
          9618 => x"8d",
          9619 => x"82",
          9620 => x"70",
          9621 => x"e1",
          9622 => x"12",
          9623 => x"06",
          9624 => x"82",
          9625 => x"85",
          9626 => x"fe",
          9627 => x"92",
          9628 => x"84",
          9629 => x"22",
          9630 => x"53",
          9631 => x"26",
          9632 => x"53",
          9633 => x"83",
          9634 => x"81",
          9635 => x"70",
          9636 => x"8b",
          9637 => x"82",
          9638 => x"70",
          9639 => x"72",
          9640 => x"0c",
          9641 => x"04",
          9642 => x"77",
          9643 => x"ff",
          9644 => x"a7",
          9645 => x"ff",
          9646 => x"ce",
          9647 => x"9f",
          9648 => x"85",
          9649 => x"88",
          9650 => x"82",
          9651 => x"70",
          9652 => x"25",
          9653 => x"07",
          9654 => x"70",
          9655 => x"75",
          9656 => x"57",
          9657 => x"2a",
          9658 => x"06",
          9659 => x"52",
          9660 => x"71",
          9661 => x"38",
          9662 => x"80",
          9663 => x"84",
          9664 => x"b0",
          9665 => x"08",
          9666 => x"31",
          9667 => x"70",
          9668 => x"51",
          9669 => x"71",
          9670 => x"06",
          9671 => x"51",
          9672 => x"f0",
          9673 => x"39",
          9674 => x"9a",
          9675 => x"51",
          9676 => x"12",
          9677 => x"88",
          9678 => x"39",
          9679 => x"51",
          9680 => x"a0",
          9681 => x"83",
          9682 => x"52",
          9683 => x"fe",
          9684 => x"10",
          9685 => x"f1",
          9686 => x"70",
          9687 => x"0c",
          9688 => x"04",
          9689 => x"ff",
          9690 => x"ff",
          9691 => x"00",
          9692 => x"ff",
          9693 => x"2b",
          9694 => x"2b",
          9695 => x"2b",
          9696 => x"2b",
          9697 => x"2b",
          9698 => x"2b",
          9699 => x"2b",
          9700 => x"2b",
          9701 => x"2b",
          9702 => x"2b",
          9703 => x"2b",
          9704 => x"2b",
          9705 => x"2b",
          9706 => x"2b",
          9707 => x"2b",
          9708 => x"2b",
          9709 => x"2b",
          9710 => x"2b",
          9711 => x"2b",
          9712 => x"2b",
          9713 => x"43",
          9714 => x"43",
          9715 => x"43",
          9716 => x"43",
          9717 => x"43",
          9718 => x"49",
          9719 => x"4a",
          9720 => x"4b",
          9721 => x"4e",
          9722 => x"4a",
          9723 => x"48",
          9724 => x"4c",
          9725 => x"4e",
          9726 => x"4c",
          9727 => x"4d",
          9728 => x"4d",
          9729 => x"4b",
          9730 => x"48",
          9731 => x"4b",
          9732 => x"4c",
          9733 => x"4c",
          9734 => x"48",
          9735 => x"48",
          9736 => x"4d",
          9737 => x"4d",
          9738 => x"4e",
          9739 => x"4e",
          9740 => x"97",
          9741 => x"97",
          9742 => x"97",
          9743 => x"97",
          9744 => x"97",
          9745 => x"97",
          9746 => x"97",
          9747 => x"97",
          9748 => x"97",
          9749 => x"0e",
          9750 => x"17",
          9751 => x"17",
          9752 => x"0e",
          9753 => x"17",
          9754 => x"17",
          9755 => x"17",
          9756 => x"17",
          9757 => x"17",
          9758 => x"17",
          9759 => x"17",
          9760 => x"0e",
          9761 => x"17",
          9762 => x"0e",
          9763 => x"0e",
          9764 => x"17",
          9765 => x"17",
          9766 => x"17",
          9767 => x"17",
          9768 => x"17",
          9769 => x"17",
          9770 => x"17",
          9771 => x"17",
          9772 => x"17",
          9773 => x"17",
          9774 => x"17",
          9775 => x"17",
          9776 => x"17",
          9777 => x"17",
          9778 => x"17",
          9779 => x"17",
          9780 => x"17",
          9781 => x"17",
          9782 => x"17",
          9783 => x"17",
          9784 => x"17",
          9785 => x"17",
          9786 => x"17",
          9787 => x"17",
          9788 => x"17",
          9789 => x"17",
          9790 => x"17",
          9791 => x"17",
          9792 => x"17",
          9793 => x"17",
          9794 => x"17",
          9795 => x"17",
          9796 => x"17",
          9797 => x"17",
          9798 => x"17",
          9799 => x"17",
          9800 => x"0f",
          9801 => x"17",
          9802 => x"17",
          9803 => x"17",
          9804 => x"17",
          9805 => x"11",
          9806 => x"17",
          9807 => x"17",
          9808 => x"17",
          9809 => x"17",
          9810 => x"17",
          9811 => x"17",
          9812 => x"17",
          9813 => x"17",
          9814 => x"17",
          9815 => x"17",
          9816 => x"0e",
          9817 => x"10",
          9818 => x"0e",
          9819 => x"0e",
          9820 => x"0e",
          9821 => x"17",
          9822 => x"10",
          9823 => x"17",
          9824 => x"17",
          9825 => x"0e",
          9826 => x"17",
          9827 => x"17",
          9828 => x"10",
          9829 => x"10",
          9830 => x"17",
          9831 => x"17",
          9832 => x"0f",
          9833 => x"17",
          9834 => x"11",
          9835 => x"17",
          9836 => x"17",
          9837 => x"11",
          9838 => x"6e",
          9839 => x"00",
          9840 => x"6f",
          9841 => x"00",
          9842 => x"6e",
          9843 => x"00",
          9844 => x"6f",
          9845 => x"00",
          9846 => x"78",
          9847 => x"00",
          9848 => x"6c",
          9849 => x"00",
          9850 => x"6f",
          9851 => x"00",
          9852 => x"69",
          9853 => x"00",
          9854 => x"75",
          9855 => x"00",
          9856 => x"62",
          9857 => x"68",
          9858 => x"77",
          9859 => x"64",
          9860 => x"65",
          9861 => x"64",
          9862 => x"65",
          9863 => x"6c",
          9864 => x"00",
          9865 => x"70",
          9866 => x"73",
          9867 => x"74",
          9868 => x"73",
          9869 => x"00",
          9870 => x"66",
          9871 => x"00",
          9872 => x"73",
          9873 => x"00",
          9874 => x"61",
          9875 => x"00",
          9876 => x"61",
          9877 => x"00",
          9878 => x"6c",
          9879 => x"00",
          9880 => x"00",
          9881 => x"73",
          9882 => x"72",
          9883 => x"00",
          9884 => x"74",
          9885 => x"61",
          9886 => x"72",
          9887 => x"2e",
          9888 => x"73",
          9889 => x"6f",
          9890 => x"65",
          9891 => x"2e",
          9892 => x"20",
          9893 => x"65",
          9894 => x"75",
          9895 => x"00",
          9896 => x"20",
          9897 => x"68",
          9898 => x"75",
          9899 => x"00",
          9900 => x"76",
          9901 => x"64",
          9902 => x"6c",
          9903 => x"6d",
          9904 => x"00",
          9905 => x"63",
          9906 => x"20",
          9907 => x"69",
          9908 => x"00",
          9909 => x"6c",
          9910 => x"6c",
          9911 => x"64",
          9912 => x"78",
          9913 => x"73",
          9914 => x"00",
          9915 => x"6c",
          9916 => x"61",
          9917 => x"65",
          9918 => x"76",
          9919 => x"64",
          9920 => x"00",
          9921 => x"20",
          9922 => x"77",
          9923 => x"65",
          9924 => x"6f",
          9925 => x"74",
          9926 => x"00",
          9927 => x"69",
          9928 => x"6e",
          9929 => x"65",
          9930 => x"73",
          9931 => x"76",
          9932 => x"64",
          9933 => x"00",
          9934 => x"73",
          9935 => x"6f",
          9936 => x"6e",
          9937 => x"65",
          9938 => x"00",
          9939 => x"20",
          9940 => x"70",
          9941 => x"62",
          9942 => x"66",
          9943 => x"73",
          9944 => x"65",
          9945 => x"6f",
          9946 => x"20",
          9947 => x"64",
          9948 => x"2e",
          9949 => x"72",
          9950 => x"20",
          9951 => x"72",
          9952 => x"2e",
          9953 => x"6d",
          9954 => x"74",
          9955 => x"70",
          9956 => x"74",
          9957 => x"20",
          9958 => x"63",
          9959 => x"65",
          9960 => x"00",
          9961 => x"6c",
          9962 => x"73",
          9963 => x"63",
          9964 => x"2e",
          9965 => x"73",
          9966 => x"69",
          9967 => x"6e",
          9968 => x"65",
          9969 => x"79",
          9970 => x"00",
          9971 => x"6f",
          9972 => x"6e",
          9973 => x"70",
          9974 => x"66",
          9975 => x"73",
          9976 => x"00",
          9977 => x"72",
          9978 => x"74",
          9979 => x"20",
          9980 => x"6f",
          9981 => x"63",
          9982 => x"00",
          9983 => x"63",
          9984 => x"73",
          9985 => x"00",
          9986 => x"6b",
          9987 => x"6e",
          9988 => x"72",
          9989 => x"00",
          9990 => x"6c",
          9991 => x"79",
          9992 => x"20",
          9993 => x"61",
          9994 => x"6c",
          9995 => x"79",
          9996 => x"2f",
          9997 => x"2e",
          9998 => x"00",
          9999 => x"61",
         10000 => x"00",
         10001 => x"25",
         10002 => x"78",
         10003 => x"3d",
         10004 => x"6c",
         10005 => x"32",
         10006 => x"38",
         10007 => x"20",
         10008 => x"42",
         10009 => x"38",
         10010 => x"25",
         10011 => x"78",
         10012 => x"38",
         10013 => x"00",
         10014 => x"38",
         10015 => x"00",
         10016 => x"20",
         10017 => x"34",
         10018 => x"00",
         10019 => x"20",
         10020 => x"20",
         10021 => x"00",
         10022 => x"32",
         10023 => x"00",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"55",
         10028 => x"00",
         10029 => x"2a",
         10030 => x"20",
         10031 => x"00",
         10032 => x"2f",
         10033 => x"32",
         10034 => x"00",
         10035 => x"2e",
         10036 => x"00",
         10037 => x"50",
         10038 => x"72",
         10039 => x"25",
         10040 => x"29",
         10041 => x"20",
         10042 => x"2a",
         10043 => x"00",
         10044 => x"55",
         10045 => x"49",
         10046 => x"72",
         10047 => x"74",
         10048 => x"6e",
         10049 => x"72",
         10050 => x"6d",
         10051 => x"69",
         10052 => x"72",
         10053 => x"74",
         10054 => x"32",
         10055 => x"74",
         10056 => x"75",
         10057 => x"00",
         10058 => x"43",
         10059 => x"52",
         10060 => x"6e",
         10061 => x"72",
         10062 => x"00",
         10063 => x"43",
         10064 => x"57",
         10065 => x"6e",
         10066 => x"72",
         10067 => x"00",
         10068 => x"52",
         10069 => x"52",
         10070 => x"6e",
         10071 => x"72",
         10072 => x"00",
         10073 => x"52",
         10074 => x"54",
         10075 => x"6e",
         10076 => x"72",
         10077 => x"00",
         10078 => x"52",
         10079 => x"52",
         10080 => x"6e",
         10081 => x"72",
         10082 => x"00",
         10083 => x"52",
         10084 => x"54",
         10085 => x"6e",
         10086 => x"72",
         10087 => x"00",
         10088 => x"74",
         10089 => x"67",
         10090 => x"20",
         10091 => x"65",
         10092 => x"2e",
         10093 => x"61",
         10094 => x"6e",
         10095 => x"69",
         10096 => x"2e",
         10097 => x"00",
         10098 => x"74",
         10099 => x"65",
         10100 => x"61",
         10101 => x"00",
         10102 => x"75",
         10103 => x"68",
         10104 => x"00",
         10105 => x"00",
         10106 => x"69",
         10107 => x"20",
         10108 => x"69",
         10109 => x"69",
         10110 => x"73",
         10111 => x"64",
         10112 => x"72",
         10113 => x"2c",
         10114 => x"65",
         10115 => x"20",
         10116 => x"74",
         10117 => x"6e",
         10118 => x"6c",
         10119 => x"00",
         10120 => x"00",
         10121 => x"64",
         10122 => x"73",
         10123 => x"64",
         10124 => x"00",
         10125 => x"69",
         10126 => x"6c",
         10127 => x"64",
         10128 => x"00",
         10129 => x"69",
         10130 => x"20",
         10131 => x"69",
         10132 => x"69",
         10133 => x"73",
         10134 => x"00",
         10135 => x"3d",
         10136 => x"00",
         10137 => x"3a",
         10138 => x"65",
         10139 => x"6e",
         10140 => x"2e",
         10141 => x"00",
         10142 => x"70",
         10143 => x"67",
         10144 => x"00",
         10145 => x"6d",
         10146 => x"69",
         10147 => x"2e",
         10148 => x"00",
         10149 => x"38",
         10150 => x"25",
         10151 => x"29",
         10152 => x"30",
         10153 => x"28",
         10154 => x"78",
         10155 => x"00",
         10156 => x"6d",
         10157 => x"65",
         10158 => x"79",
         10159 => x"6f",
         10160 => x"65",
         10161 => x"00",
         10162 => x"38",
         10163 => x"25",
         10164 => x"2d",
         10165 => x"3f",
         10166 => x"38",
         10167 => x"25",
         10168 => x"2d",
         10169 => x"38",
         10170 => x"25",
         10171 => x"58",
         10172 => x"00",
         10173 => x"73",
         10174 => x"69",
         10175 => x"69",
         10176 => x"72",
         10177 => x"74",
         10178 => x"00",
         10179 => x"61",
         10180 => x"6e",
         10181 => x"6e",
         10182 => x"72",
         10183 => x"73",
         10184 => x"73",
         10185 => x"65",
         10186 => x"61",
         10187 => x"66",
         10188 => x"00",
         10189 => x"61",
         10190 => x"6e",
         10191 => x"61",
         10192 => x"66",
         10193 => x"00",
         10194 => x"65",
         10195 => x"69",
         10196 => x"63",
         10197 => x"20",
         10198 => x"30",
         10199 => x"20",
         10200 => x"0a",
         10201 => x"6c",
         10202 => x"67",
         10203 => x"64",
         10204 => x"20",
         10205 => x"6c",
         10206 => x"2e",
         10207 => x"00",
         10208 => x"6c",
         10209 => x"65",
         10210 => x"6e",
         10211 => x"63",
         10212 => x"20",
         10213 => x"29",
         10214 => x"00",
         10215 => x"73",
         10216 => x"74",
         10217 => x"20",
         10218 => x"6c",
         10219 => x"74",
         10220 => x"2e",
         10221 => x"00",
         10222 => x"6c",
         10223 => x"65",
         10224 => x"74",
         10225 => x"2e",
         10226 => x"00",
         10227 => x"55",
         10228 => x"6e",
         10229 => x"3a",
         10230 => x"5c",
         10231 => x"25",
         10232 => x"00",
         10233 => x"3a",
         10234 => x"5c",
         10235 => x"00",
         10236 => x"3a",
         10237 => x"00",
         10238 => x"64",
         10239 => x"6d",
         10240 => x"64",
         10241 => x"00",
         10242 => x"6e",
         10243 => x"67",
         10244 => x"00",
         10245 => x"61",
         10246 => x"6e",
         10247 => x"6e",
         10248 => x"72",
         10249 => x"73",
         10250 => x"00",
         10251 => x"2f",
         10252 => x"25",
         10253 => x"64",
         10254 => x"3a",
         10255 => x"25",
         10256 => x"0a",
         10257 => x"43",
         10258 => x"6e",
         10259 => x"75",
         10260 => x"69",
         10261 => x"00",
         10262 => x"66",
         10263 => x"20",
         10264 => x"20",
         10265 => x"66",
         10266 => x"00",
         10267 => x"44",
         10268 => x"63",
         10269 => x"69",
         10270 => x"65",
         10271 => x"74",
         10272 => x"00",
         10273 => x"20",
         10274 => x"20",
         10275 => x"41",
         10276 => x"28",
         10277 => x"58",
         10278 => x"38",
         10279 => x"0a",
         10280 => x"20",
         10281 => x"52",
         10282 => x"20",
         10283 => x"28",
         10284 => x"58",
         10285 => x"38",
         10286 => x"0a",
         10287 => x"20",
         10288 => x"53",
         10289 => x"52",
         10290 => x"28",
         10291 => x"58",
         10292 => x"38",
         10293 => x"0a",
         10294 => x"20",
         10295 => x"41",
         10296 => x"20",
         10297 => x"28",
         10298 => x"58",
         10299 => x"38",
         10300 => x"0a",
         10301 => x"20",
         10302 => x"4d",
         10303 => x"20",
         10304 => x"28",
         10305 => x"58",
         10306 => x"38",
         10307 => x"0a",
         10308 => x"20",
         10309 => x"20",
         10310 => x"44",
         10311 => x"28",
         10312 => x"69",
         10313 => x"20",
         10314 => x"32",
         10315 => x"0a",
         10316 => x"20",
         10317 => x"4d",
         10318 => x"20",
         10319 => x"28",
         10320 => x"65",
         10321 => x"20",
         10322 => x"32",
         10323 => x"0a",
         10324 => x"20",
         10325 => x"54",
         10326 => x"54",
         10327 => x"28",
         10328 => x"6e",
         10329 => x"73",
         10330 => x"32",
         10331 => x"0a",
         10332 => x"20",
         10333 => x"53",
         10334 => x"4e",
         10335 => x"55",
         10336 => x"00",
         10337 => x"20",
         10338 => x"20",
         10339 => x"00",
         10340 => x"20",
         10341 => x"43",
         10342 => x"00",
         10343 => x"20",
         10344 => x"32",
         10345 => x"20",
         10346 => x"49",
         10347 => x"64",
         10348 => x"73",
         10349 => x"00",
         10350 => x"20",
         10351 => x"55",
         10352 => x"73",
         10353 => x"56",
         10354 => x"6f",
         10355 => x"64",
         10356 => x"73",
         10357 => x"20",
         10358 => x"58",
         10359 => x"00",
         10360 => x"20",
         10361 => x"55",
         10362 => x"6d",
         10363 => x"20",
         10364 => x"72",
         10365 => x"64",
         10366 => x"73",
         10367 => x"20",
         10368 => x"58",
         10369 => x"00",
         10370 => x"20",
         10371 => x"61",
         10372 => x"53",
         10373 => x"74",
         10374 => x"64",
         10375 => x"73",
         10376 => x"20",
         10377 => x"20",
         10378 => x"58",
         10379 => x"00",
         10380 => x"73",
         10381 => x"00",
         10382 => x"20",
         10383 => x"55",
         10384 => x"20",
         10385 => x"20",
         10386 => x"20",
         10387 => x"20",
         10388 => x"20",
         10389 => x"20",
         10390 => x"58",
         10391 => x"00",
         10392 => x"20",
         10393 => x"73",
         10394 => x"20",
         10395 => x"63",
         10396 => x"72",
         10397 => x"20",
         10398 => x"20",
         10399 => x"20",
         10400 => x"25",
         10401 => x"4d",
         10402 => x"00",
         10403 => x"20",
         10404 => x"52",
         10405 => x"43",
         10406 => x"6b",
         10407 => x"65",
         10408 => x"20",
         10409 => x"20",
         10410 => x"20",
         10411 => x"25",
         10412 => x"4d",
         10413 => x"00",
         10414 => x"20",
         10415 => x"73",
         10416 => x"6e",
         10417 => x"44",
         10418 => x"20",
         10419 => x"63",
         10420 => x"72",
         10421 => x"20",
         10422 => x"25",
         10423 => x"4d",
         10424 => x"00",
         10425 => x"61",
         10426 => x"00",
         10427 => x"64",
         10428 => x"00",
         10429 => x"65",
         10430 => x"00",
         10431 => x"4f",
         10432 => x"4f",
         10433 => x"00",
         10434 => x"6b",
         10435 => x"6e",
         10436 => x"a4",
         10437 => x"00",
         10438 => x"00",
         10439 => x"a4",
         10440 => x"00",
         10441 => x"00",
         10442 => x"a4",
         10443 => x"00",
         10444 => x"00",
         10445 => x"a4",
         10446 => x"00",
         10447 => x"00",
         10448 => x"a4",
         10449 => x"00",
         10450 => x"00",
         10451 => x"a4",
         10452 => x"00",
         10453 => x"00",
         10454 => x"a4",
         10455 => x"00",
         10456 => x"00",
         10457 => x"a4",
         10458 => x"00",
         10459 => x"00",
         10460 => x"a4",
         10461 => x"00",
         10462 => x"00",
         10463 => x"a4",
         10464 => x"00",
         10465 => x"00",
         10466 => x"a4",
         10467 => x"00",
         10468 => x"00",
         10469 => x"a4",
         10470 => x"00",
         10471 => x"00",
         10472 => x"a4",
         10473 => x"00",
         10474 => x"00",
         10475 => x"a4",
         10476 => x"00",
         10477 => x"00",
         10478 => x"a4",
         10479 => x"00",
         10480 => x"00",
         10481 => x"a4",
         10482 => x"00",
         10483 => x"00",
         10484 => x"a4",
         10485 => x"00",
         10486 => x"00",
         10487 => x"a4",
         10488 => x"00",
         10489 => x"00",
         10490 => x"a4",
         10491 => x"00",
         10492 => x"00",
         10493 => x"a4",
         10494 => x"00",
         10495 => x"00",
         10496 => x"a4",
         10497 => x"00",
         10498 => x"00",
         10499 => x"a4",
         10500 => x"00",
         10501 => x"00",
         10502 => x"44",
         10503 => x"43",
         10504 => x"42",
         10505 => x"41",
         10506 => x"36",
         10507 => x"35",
         10508 => x"34",
         10509 => x"46",
         10510 => x"33",
         10511 => x"32",
         10512 => x"31",
         10513 => x"00",
         10514 => x"00",
         10515 => x"00",
         10516 => x"00",
         10517 => x"00",
         10518 => x"00",
         10519 => x"00",
         10520 => x"00",
         10521 => x"00",
         10522 => x"00",
         10523 => x"00",
         10524 => x"73",
         10525 => x"79",
         10526 => x"73",
         10527 => x"00",
         10528 => x"00",
         10529 => x"34",
         10530 => x"20",
         10531 => x"00",
         10532 => x"69",
         10533 => x"20",
         10534 => x"72",
         10535 => x"74",
         10536 => x"65",
         10537 => x"73",
         10538 => x"79",
         10539 => x"6c",
         10540 => x"6f",
         10541 => x"46",
         10542 => x"00",
         10543 => x"6e",
         10544 => x"20",
         10545 => x"6e",
         10546 => x"65",
         10547 => x"20",
         10548 => x"74",
         10549 => x"20",
         10550 => x"65",
         10551 => x"69",
         10552 => x"6c",
         10553 => x"2e",
         10554 => x"00",
         10555 => x"3a",
         10556 => x"7c",
         10557 => x"00",
         10558 => x"3b",
         10559 => x"00",
         10560 => x"54",
         10561 => x"54",
         10562 => x"00",
         10563 => x"90",
         10564 => x"4f",
         10565 => x"30",
         10566 => x"20",
         10567 => x"45",
         10568 => x"20",
         10569 => x"33",
         10570 => x"20",
         10571 => x"20",
         10572 => x"45",
         10573 => x"20",
         10574 => x"20",
         10575 => x"20",
         10576 => x"a4",
         10577 => x"00",
         10578 => x"00",
         10579 => x"00",
         10580 => x"05",
         10581 => x"10",
         10582 => x"18",
         10583 => x"00",
         10584 => x"45",
         10585 => x"8f",
         10586 => x"45",
         10587 => x"8e",
         10588 => x"92",
         10589 => x"55",
         10590 => x"9a",
         10591 => x"9e",
         10592 => x"4f",
         10593 => x"a6",
         10594 => x"aa",
         10595 => x"ae",
         10596 => x"b2",
         10597 => x"b6",
         10598 => x"ba",
         10599 => x"be",
         10600 => x"c2",
         10601 => x"c6",
         10602 => x"ca",
         10603 => x"ce",
         10604 => x"d2",
         10605 => x"d6",
         10606 => x"da",
         10607 => x"de",
         10608 => x"e2",
         10609 => x"e6",
         10610 => x"ea",
         10611 => x"ee",
         10612 => x"f2",
         10613 => x"f6",
         10614 => x"fa",
         10615 => x"fe",
         10616 => x"2c",
         10617 => x"5d",
         10618 => x"2a",
         10619 => x"3f",
         10620 => x"00",
         10621 => x"00",
         10622 => x"00",
         10623 => x"02",
         10624 => x"00",
         10625 => x"00",
         10626 => x"00",
         10627 => x"00",
         10628 => x"00",
         10629 => x"00",
         10630 => x"00",
         10631 => x"00",
         10632 => x"00",
         10633 => x"00",
         10634 => x"00",
         10635 => x"00",
         10636 => x"00",
         10637 => x"00",
         10638 => x"00",
         10639 => x"00",
         10640 => x"00",
         10641 => x"00",
         10642 => x"00",
         10643 => x"00",
         10644 => x"01",
         10645 => x"00",
         10646 => x"00",
         10647 => x"00",
         10648 => x"00",
         10649 => x"23",
         10650 => x"00",
         10651 => x"00",
         10652 => x"00",
         10653 => x"25",
         10654 => x"25",
         10655 => x"25",
         10656 => x"25",
         10657 => x"25",
         10658 => x"25",
         10659 => x"25",
         10660 => x"25",
         10661 => x"25",
         10662 => x"25",
         10663 => x"25",
         10664 => x"25",
         10665 => x"25",
         10666 => x"25",
         10667 => x"25",
         10668 => x"25",
         10669 => x"25",
         10670 => x"25",
         10671 => x"25",
         10672 => x"25",
         10673 => x"25",
         10674 => x"25",
         10675 => x"25",
         10676 => x"25",
         10677 => x"00",
         10678 => x"03",
         10679 => x"03",
         10680 => x"03",
         10681 => x"03",
         10682 => x"03",
         10683 => x"03",
         10684 => x"22",
         10685 => x"00",
         10686 => x"22",
         10687 => x"23",
         10688 => x"22",
         10689 => x"22",
         10690 => x"22",
         10691 => x"00",
         10692 => x"00",
         10693 => x"03",
         10694 => x"03",
         10695 => x"03",
         10696 => x"00",
         10697 => x"01",
         10698 => x"01",
         10699 => x"01",
         10700 => x"01",
         10701 => x"01",
         10702 => x"01",
         10703 => x"02",
         10704 => x"01",
         10705 => x"01",
         10706 => x"01",
         10707 => x"01",
         10708 => x"01",
         10709 => x"01",
         10710 => x"01",
         10711 => x"01",
         10712 => x"01",
         10713 => x"01",
         10714 => x"01",
         10715 => x"01",
         10716 => x"02",
         10717 => x"01",
         10718 => x"02",
         10719 => x"01",
         10720 => x"01",
         10721 => x"01",
         10722 => x"01",
         10723 => x"01",
         10724 => x"01",
         10725 => x"01",
         10726 => x"01",
         10727 => x"01",
         10728 => x"01",
         10729 => x"01",
         10730 => x"01",
         10731 => x"01",
         10732 => x"01",
         10733 => x"01",
         10734 => x"01",
         10735 => x"01",
         10736 => x"01",
         10737 => x"01",
         10738 => x"01",
         10739 => x"01",
         10740 => x"01",
         10741 => x"01",
         10742 => x"01",
         10743 => x"00",
         10744 => x"01",
         10745 => x"01",
         10746 => x"01",
         10747 => x"01",
         10748 => x"01",
         10749 => x"01",
         10750 => x"00",
         10751 => x"02",
         10752 => x"02",
         10753 => x"02",
         10754 => x"02",
         10755 => x"02",
         10756 => x"02",
         10757 => x"01",
         10758 => x"02",
         10759 => x"01",
         10760 => x"01",
         10761 => x"01",
         10762 => x"02",
         10763 => x"02",
         10764 => x"02",
         10765 => x"01",
         10766 => x"02",
         10767 => x"02",
         10768 => x"01",
         10769 => x"2c",
         10770 => x"02",
         10771 => x"01",
         10772 => x"02",
         10773 => x"02",
         10774 => x"01",
         10775 => x"02",
         10776 => x"02",
         10777 => x"02",
         10778 => x"2c",
         10779 => x"02",
         10780 => x"02",
         10781 => x"01",
         10782 => x"02",
         10783 => x"02",
         10784 => x"02",
         10785 => x"01",
         10786 => x"02",
         10787 => x"02",
         10788 => x"02",
         10789 => x"03",
         10790 => x"03",
         10791 => x"03",
         10792 => x"00",
         10793 => x"03",
         10794 => x"03",
         10795 => x"03",
         10796 => x"00",
         10797 => x"03",
         10798 => x"03",
         10799 => x"00",
         10800 => x"03",
         10801 => x"03",
         10802 => x"03",
         10803 => x"03",
         10804 => x"03",
         10805 => x"03",
         10806 => x"03",
         10807 => x"03",
         10808 => x"04",
         10809 => x"04",
         10810 => x"04",
         10811 => x"04",
         10812 => x"04",
         10813 => x"04",
         10814 => x"04",
         10815 => x"01",
         10816 => x"04",
         10817 => x"00",
         10818 => x"00",
         10819 => x"1e",
         10820 => x"1e",
         10821 => x"1f",
         10822 => x"1f",
         10823 => x"1f",
         10824 => x"1f",
         10825 => x"1f",
         10826 => x"1f",
         10827 => x"1f",
         10828 => x"1f",
         10829 => x"1f",
         10830 => x"1f",
         10831 => x"06",
         10832 => x"00",
         10833 => x"1f",
         10834 => x"1f",
         10835 => x"1f",
         10836 => x"1f",
         10837 => x"1f",
         10838 => x"1f",
         10839 => x"1f",
         10840 => x"06",
         10841 => x"06",
         10842 => x"06",
         10843 => x"00",
         10844 => x"1f",
         10845 => x"1f",
         10846 => x"00",
         10847 => x"1f",
         10848 => x"1f",
         10849 => x"1f",
         10850 => x"1f",
         10851 => x"00",
         10852 => x"21",
         10853 => x"21",
         10854 => x"02",
         10855 => x"00",
         10856 => x"24",
         10857 => x"2c",
         10858 => x"2c",
         10859 => x"2c",
         10860 => x"2c",
         10861 => x"2c",
         10862 => x"2d",
         10863 => x"ff",
         10864 => x"00",
         10865 => x"00",
         10866 => x"99",
         10867 => x"01",
         10868 => x"00",
         10869 => x"00",
         10870 => x"99",
         10871 => x"01",
         10872 => x"00",
         10873 => x"00",
         10874 => x"99",
         10875 => x"03",
         10876 => x"00",
         10877 => x"00",
         10878 => x"99",
         10879 => x"03",
         10880 => x"00",
         10881 => x"00",
         10882 => x"99",
         10883 => x"03",
         10884 => x"00",
         10885 => x"00",
         10886 => x"99",
         10887 => x"04",
         10888 => x"00",
         10889 => x"00",
         10890 => x"99",
         10891 => x"04",
         10892 => x"00",
         10893 => x"00",
         10894 => x"99",
         10895 => x"04",
         10896 => x"00",
         10897 => x"00",
         10898 => x"99",
         10899 => x"04",
         10900 => x"00",
         10901 => x"00",
         10902 => x"9a",
         10903 => x"04",
         10904 => x"00",
         10905 => x"00",
         10906 => x"9a",
         10907 => x"04",
         10908 => x"00",
         10909 => x"00",
         10910 => x"9a",
         10911 => x"04",
         10912 => x"00",
         10913 => x"00",
         10914 => x"9a",
         10915 => x"05",
         10916 => x"00",
         10917 => x"00",
         10918 => x"9a",
         10919 => x"05",
         10920 => x"00",
         10921 => x"00",
         10922 => x"9a",
         10923 => x"05",
         10924 => x"00",
         10925 => x"00",
         10926 => x"9a",
         10927 => x"05",
         10928 => x"00",
         10929 => x"00",
         10930 => x"9a",
         10931 => x"07",
         10932 => x"00",
         10933 => x"00",
         10934 => x"9a",
         10935 => x"07",
         10936 => x"00",
         10937 => x"00",
         10938 => x"9a",
         10939 => x"08",
         10940 => x"00",
         10941 => x"00",
         10942 => x"9a",
         10943 => x"08",
         10944 => x"00",
         10945 => x"00",
         10946 => x"9a",
         10947 => x"08",
         10948 => x"00",
         10949 => x"00",
         10950 => x"9a",
         10951 => x"08",
         10952 => x"00",
         10953 => x"00",
         10954 => x"9a",
         10955 => x"09",
         10956 => x"00",
         10957 => x"00",
         10958 => x"9a",
         10959 => x"09",
         10960 => x"00",
         10961 => x"00",
         10962 => x"9a",
         10963 => x"09",
         10964 => x"00",
         10965 => x"00",
         10966 => x"9a",
         10967 => x"09",
         10968 => x"00",
         10969 => x"00",
         10970 => x"00",
         10971 => x"00",
         10972 => x"7f",
         10973 => x"00",
         10974 => x"7f",
         10975 => x"00",
         10976 => x"7f",
         10977 => x"00",
         10978 => x"00",
         10979 => x"00",
         10980 => x"ff",
         10981 => x"00",
         10982 => x"00",
         10983 => x"78",
         10984 => x"00",
         10985 => x"e1",
         10986 => x"e1",
         10987 => x"e1",
         10988 => x"00",
         10989 => x"01",
         10990 => x"01",
         10991 => x"10",
         10992 => x"00",
         10993 => x"00",
         10994 => x"00",
         10995 => x"00",
         10996 => x"00",
         10997 => x"00",
         10998 => x"00",
         10999 => x"00",
         11000 => x"00",
         11001 => x"00",
         11002 => x"00",
         11003 => x"00",
         11004 => x"00",
         11005 => x"00",
         11006 => x"00",
         11007 => x"00",
         11008 => x"00",
         11009 => x"00",
         11010 => x"00",
         11011 => x"00",
         11012 => x"00",
         11013 => x"00",
         11014 => x"00",
         11015 => x"00",
         11016 => x"00",
         11017 => x"a4",
         11018 => x"00",
         11019 => x"a4",
         11020 => x"00",
         11021 => x"a4",
         11022 => x"00",
         11023 => x"00",
         11024 => x"00",
         11025 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"84",
           389 => x"82",
           390 => x"b3",
           391 => x"d8",
           392 => x"80",
           393 => x"d8",
           394 => x"e3",
           395 => x"d4",
           396 => x"90",
           397 => x"d4",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"84",
           404 => x"82",
           405 => x"b1",
           406 => x"d8",
           407 => x"80",
           408 => x"d8",
           409 => x"cf",
           410 => x"d8",
           411 => x"80",
           412 => x"d8",
           413 => x"c9",
           414 => x"d8",
           415 => x"80",
           416 => x"d8",
           417 => x"d8",
           418 => x"d4",
           419 => x"90",
           420 => x"d4",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"84",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"84",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"84",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"84",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"84",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"84",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"84",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"84",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"84",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"84",
           463 => x"82",
           464 => x"82",
           465 => x"82",
           466 => x"84",
           467 => x"82",
           468 => x"82",
           469 => x"82",
           470 => x"84",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"84",
           475 => x"82",
           476 => x"82",
           477 => x"82",
           478 => x"84",
           479 => x"82",
           480 => x"82",
           481 => x"82",
           482 => x"84",
           483 => x"82",
           484 => x"82",
           485 => x"82",
           486 => x"84",
           487 => x"82",
           488 => x"82",
           489 => x"82",
           490 => x"84",
           491 => x"82",
           492 => x"82",
           493 => x"82",
           494 => x"84",
           495 => x"82",
           496 => x"82",
           497 => x"82",
           498 => x"84",
           499 => x"82",
           500 => x"82",
           501 => x"82",
           502 => x"84",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"84",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"84",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"84",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"84",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"84",
           523 => x"82",
           524 => x"82",
           525 => x"82",
           526 => x"84",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"84",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"84",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"84",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"84",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"84",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"84",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"84",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"84",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"84",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"84",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"84",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"84",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"84",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"84",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"84",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"84",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"84",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"84",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"bb",
           630 => x"d8",
           631 => x"82",
           632 => x"fb",
           633 => x"d8",
           634 => x"05",
           635 => x"d4",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"c8",
           644 => x"d8",
           645 => x"05",
           646 => x"d4",
           647 => x"08",
           648 => x"c8",
           649 => x"87",
           650 => x"d8",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"d8",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"d4",
           670 => x"0c",
           671 => x"d8",
           672 => x"05",
           673 => x"d4",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"d4",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"d8",
           696 => x"05",
           697 => x"d4",
           698 => x"08",
           699 => x"73",
           700 => x"d4",
           701 => x"08",
           702 => x"d8",
           703 => x"05",
           704 => x"d4",
           705 => x"08",
           706 => x"d8",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"d8",
           718 => x"3d",
           719 => x"d4",
           720 => x"d8",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"d8",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"d8",
           734 => x"05",
           735 => x"d4",
           736 => x"08",
           737 => x"d4",
           738 => x"08",
           739 => x"d4",
           740 => x"70",
           741 => x"81",
           742 => x"d8",
           743 => x"82",
           744 => x"dc",
           745 => x"d8",
           746 => x"05",
           747 => x"d4",
           748 => x"08",
           749 => x"80",
           750 => x"d8",
           751 => x"05",
           752 => x"d8",
           753 => x"8e",
           754 => x"d8",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"d8",
           761 => x"05",
           762 => x"d4",
           763 => x"08",
           764 => x"d4",
           765 => x"08",
           766 => x"d4",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"d4",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"d4",
           777 => x"d8",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"d4",
           797 => x"08",
           798 => x"53",
           799 => x"d4",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"d4",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"d4",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"d8",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"d4",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"d8",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"d8",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"d8",
           850 => x"05",
           851 => x"d8",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"d4",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"d8",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"d4",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"d8",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"d8",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"d8",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"d8",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"d8",
           943 => x"05",
           944 => x"51",
           945 => x"d8",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"d8",
           951 => x"05",
           952 => x"d4",
           953 => x"08",
           954 => x"d8",
           955 => x"05",
           956 => x"51",
           957 => x"d8",
           958 => x"05",
           959 => x"d4",
           960 => x"22",
           961 => x"53",
           962 => x"d4",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"d8",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"d4",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"d8",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"d8",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"d8",
          1003 => x"05",
          1004 => x"d4",
          1005 => x"08",
          1006 => x"d8",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"d8",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"d4",
          1025 => x"23",
          1026 => x"d8",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"c8",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"d8",
          1033 => x"05",
          1034 => x"d8",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"d4",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"d8",
          1046 => x"05",
          1047 => x"d4",
          1048 => x"08",
          1049 => x"d8",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"d4",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"d4",
          1059 => x"0c",
          1060 => x"d8",
          1061 => x"05",
          1062 => x"d8",
          1063 => x"05",
          1064 => x"d4",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"d8",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"d4",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"d4",
          1093 => x"34",
          1094 => x"d8",
          1095 => x"05",
          1096 => x"d4",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"d8",
          1102 => x"05",
          1103 => x"d4",
          1104 => x"08",
          1105 => x"d8",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"d4",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"d4",
          1115 => x"0c",
          1116 => x"d8",
          1117 => x"05",
          1118 => x"d8",
          1119 => x"05",
          1120 => x"d4",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"d4",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"d8",
          1132 => x"05",
          1133 => x"d4",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a3",
          1137 => x"d8",
          1138 => x"72",
          1139 => x"d8",
          1140 => x"05",
          1141 => x"d4",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"d8",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"d8",
          1160 => x"05",
          1161 => x"d4",
          1162 => x"08",
          1163 => x"d4",
          1164 => x"33",
          1165 => x"d8",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"d8",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"d8",
          1182 => x"05",
          1183 => x"d8",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"d8",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"d8",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"d8",
          1206 => x"05",
          1207 => x"d4",
          1208 => x"08",
          1209 => x"d8",
          1210 => x"05",
          1211 => x"d4",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"d8",
          1216 => x"05",
          1217 => x"53",
          1218 => x"d4",
          1219 => x"23",
          1220 => x"d8",
          1221 => x"05",
          1222 => x"53",
          1223 => x"d4",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"d8",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"d4",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"d4",
          1242 => x"22",
          1243 => x"51",
          1244 => x"d8",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"d8",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"d8",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"d8",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"d8",
          1287 => x"05",
          1288 => x"54",
          1289 => x"d8",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"d8",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"d4",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"d8",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"d8",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"d8",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"d4",
          1331 => x"08",
          1332 => x"89",
          1333 => x"d8",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"d8",
          1338 => x"05",
          1339 => x"d8",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"d4",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"d8",
          1348 => x"05",
          1349 => x"54",
          1350 => x"d8",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"d8",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"d4",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"d8",
          1365 => x"05",
          1366 => x"54",
          1367 => x"d8",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"d8",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"d4",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"d8",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"d4",
          1416 => x"08",
          1417 => x"d4",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"d8",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"d4",
          1439 => x"08",
          1440 => x"d4",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"d8",
          1449 => x"05",
          1450 => x"d8",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"d4",
          1468 => x"22",
          1469 => x"54",
          1470 => x"d4",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"d4",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"d4",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"d4",
          1492 => x"23",
          1493 => x"d8",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"d8",
          1501 => x"05",
          1502 => x"d8",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"d8",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"d4",
          1530 => x"d8",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"f4",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"d8",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"d8",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"ac",
          1556 => x"ac",
          1557 => x"d8",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"c8",
          1562 => x"80",
          1563 => x"38",
          1564 => x"d8",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"d8",
          1572 => x"72",
          1573 => x"38",
          1574 => x"d8",
          1575 => x"05",
          1576 => x"d4",
          1577 => x"08",
          1578 => x"d4",
          1579 => x"0c",
          1580 => x"d4",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"d4",
          1587 => x"0d",
          1588 => x"d8",
          1589 => x"05",
          1590 => x"d4",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"d8",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"d4",
          1606 => x"0c",
          1607 => x"d8",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"d8",
          1614 => x"05",
          1615 => x"d8",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"c8",
          1620 => x"80",
          1621 => x"38",
          1622 => x"d8",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"d8",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"d8",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"d4",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"d4",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"d8",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"d8",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"d8",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"d4",
          1683 => x"08",
          1684 => x"d4",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"d4",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"d8",
          1711 => x"3d",
          1712 => x"d4",
          1713 => x"d8",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"d8",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"d4",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"d4",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"d8",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"d4",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"d4",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"d8",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"d8",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"d4",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"d8",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"d8",
          1801 => x"05",
          1802 => x"52",
          1803 => x"d4",
          1804 => x"34",
          1805 => x"d8",
          1806 => x"05",
          1807 => x"52",
          1808 => x"d4",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"d4",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"d8",
          1827 => x"05",
          1828 => x"c8",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"d4",
          1832 => x"d8",
          1833 => x"3d",
          1834 => x"d4",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"d8",
          1840 => x"05",
          1841 => x"d4",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"d4",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"d8",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"d8",
          1858 => x"05",
          1859 => x"d8",
          1860 => x"05",
          1861 => x"d4",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"d8",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"d8",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"d8",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"d8",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"d4",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"d8",
          1917 => x"05",
          1918 => x"d8",
          1919 => x"85",
          1920 => x"d8",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"d8",
          1927 => x"05",
          1928 => x"d4",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"d4",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"d4",
          1950 => x"d8",
          1951 => x"3d",
          1952 => x"d4",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"d4",
          1959 => x"08",
          1960 => x"d8",
          1961 => x"05",
          1962 => x"d4",
          1963 => x"08",
          1964 => x"72",
          1965 => x"d4",
          1966 => x"08",
          1967 => x"d8",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"d8",
          1973 => x"05",
          1974 => x"d8",
          1975 => x"84",
          1976 => x"d8",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"d8",
          1983 => x"05",
          1984 => x"d4",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"d8",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"d4",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"d4",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"d4",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"d8",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"d8",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"d4",
          2043 => x"08",
          2044 => x"d8",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"d8",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"d8",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"d8",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"d8",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"d8",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"d4",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"d4",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"d8",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"88",
          2099 => x"d8",
          2100 => x"05",
          2101 => x"d4",
          2102 => x"08",
          2103 => x"0b",
          2104 => x"08",
          2105 => x"80",
          2106 => x"d8",
          2107 => x"05",
          2108 => x"33",
          2109 => x"08",
          2110 => x"81",
          2111 => x"d4",
          2112 => x"0c",
          2113 => x"06",
          2114 => x"80",
          2115 => x"82",
          2116 => x"8c",
          2117 => x"05",
          2118 => x"08",
          2119 => x"82",
          2120 => x"8c",
          2121 => x"2e",
          2122 => x"be",
          2123 => x"d4",
          2124 => x"08",
          2125 => x"d8",
          2126 => x"05",
          2127 => x"d4",
          2128 => x"08",
          2129 => x"08",
          2130 => x"31",
          2131 => x"d4",
          2132 => x"0c",
          2133 => x"d4",
          2134 => x"08",
          2135 => x"0c",
          2136 => x"82",
          2137 => x"04",
          2138 => x"08",
          2139 => x"d4",
          2140 => x"0d",
          2141 => x"08",
          2142 => x"82",
          2143 => x"fc",
          2144 => x"d8",
          2145 => x"05",
          2146 => x"80",
          2147 => x"d8",
          2148 => x"05",
          2149 => x"82",
          2150 => x"90",
          2151 => x"d8",
          2152 => x"05",
          2153 => x"82",
          2154 => x"90",
          2155 => x"d8",
          2156 => x"05",
          2157 => x"a9",
          2158 => x"d4",
          2159 => x"08",
          2160 => x"d8",
          2161 => x"05",
          2162 => x"71",
          2163 => x"d8",
          2164 => x"05",
          2165 => x"82",
          2166 => x"fc",
          2167 => x"be",
          2168 => x"d4",
          2169 => x"08",
          2170 => x"c8",
          2171 => x"3d",
          2172 => x"d4",
          2173 => x"d8",
          2174 => x"82",
          2175 => x"f9",
          2176 => x"0b",
          2177 => x"08",
          2178 => x"82",
          2179 => x"88",
          2180 => x"25",
          2181 => x"d8",
          2182 => x"05",
          2183 => x"d8",
          2184 => x"05",
          2185 => x"82",
          2186 => x"f4",
          2187 => x"d8",
          2188 => x"05",
          2189 => x"81",
          2190 => x"d4",
          2191 => x"0c",
          2192 => x"08",
          2193 => x"82",
          2194 => x"fc",
          2195 => x"d8",
          2196 => x"05",
          2197 => x"b9",
          2198 => x"d4",
          2199 => x"08",
          2200 => x"d4",
          2201 => x"0c",
          2202 => x"d8",
          2203 => x"05",
          2204 => x"d4",
          2205 => x"08",
          2206 => x"0b",
          2207 => x"08",
          2208 => x"82",
          2209 => x"f0",
          2210 => x"d8",
          2211 => x"05",
          2212 => x"82",
          2213 => x"8c",
          2214 => x"82",
          2215 => x"88",
          2216 => x"82",
          2217 => x"d8",
          2218 => x"82",
          2219 => x"f8",
          2220 => x"82",
          2221 => x"fc",
          2222 => x"2e",
          2223 => x"d8",
          2224 => x"05",
          2225 => x"d8",
          2226 => x"05",
          2227 => x"d4",
          2228 => x"08",
          2229 => x"c8",
          2230 => x"3d",
          2231 => x"d4",
          2232 => x"d8",
          2233 => x"82",
          2234 => x"fb",
          2235 => x"0b",
          2236 => x"08",
          2237 => x"82",
          2238 => x"88",
          2239 => x"25",
          2240 => x"d8",
          2241 => x"05",
          2242 => x"d8",
          2243 => x"05",
          2244 => x"82",
          2245 => x"fc",
          2246 => x"d8",
          2247 => x"05",
          2248 => x"90",
          2249 => x"d4",
          2250 => x"08",
          2251 => x"d4",
          2252 => x"0c",
          2253 => x"d8",
          2254 => x"05",
          2255 => x"d8",
          2256 => x"05",
          2257 => x"a2",
          2258 => x"c8",
          2259 => x"d8",
          2260 => x"05",
          2261 => x"d8",
          2262 => x"05",
          2263 => x"90",
          2264 => x"d4",
          2265 => x"08",
          2266 => x"d4",
          2267 => x"0c",
          2268 => x"08",
          2269 => x"70",
          2270 => x"0c",
          2271 => x"0d",
          2272 => x"0c",
          2273 => x"d4",
          2274 => x"d8",
          2275 => x"3d",
          2276 => x"82",
          2277 => x"8c",
          2278 => x"82",
          2279 => x"88",
          2280 => x"80",
          2281 => x"d8",
          2282 => x"82",
          2283 => x"54",
          2284 => x"82",
          2285 => x"04",
          2286 => x"08",
          2287 => x"d4",
          2288 => x"0d",
          2289 => x"d8",
          2290 => x"05",
          2291 => x"d8",
          2292 => x"05",
          2293 => x"3f",
          2294 => x"08",
          2295 => x"c8",
          2296 => x"3d",
          2297 => x"d4",
          2298 => x"d8",
          2299 => x"82",
          2300 => x"fd",
          2301 => x"0b",
          2302 => x"08",
          2303 => x"80",
          2304 => x"d4",
          2305 => x"0c",
          2306 => x"08",
          2307 => x"82",
          2308 => x"88",
          2309 => x"b9",
          2310 => x"d4",
          2311 => x"08",
          2312 => x"38",
          2313 => x"d8",
          2314 => x"05",
          2315 => x"38",
          2316 => x"08",
          2317 => x"10",
          2318 => x"08",
          2319 => x"82",
          2320 => x"fc",
          2321 => x"82",
          2322 => x"fc",
          2323 => x"b8",
          2324 => x"d4",
          2325 => x"08",
          2326 => x"e1",
          2327 => x"d4",
          2328 => x"08",
          2329 => x"08",
          2330 => x"26",
          2331 => x"d8",
          2332 => x"05",
          2333 => x"d4",
          2334 => x"08",
          2335 => x"d4",
          2336 => x"0c",
          2337 => x"08",
          2338 => x"82",
          2339 => x"fc",
          2340 => x"82",
          2341 => x"f8",
          2342 => x"d8",
          2343 => x"05",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"d8",
          2347 => x"05",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"95",
          2351 => x"d4",
          2352 => x"08",
          2353 => x"38",
          2354 => x"08",
          2355 => x"70",
          2356 => x"08",
          2357 => x"51",
          2358 => x"d8",
          2359 => x"05",
          2360 => x"d8",
          2361 => x"05",
          2362 => x"d8",
          2363 => x"05",
          2364 => x"c8",
          2365 => x"0d",
          2366 => x"0c",
          2367 => x"d4",
          2368 => x"d8",
          2369 => x"3d",
          2370 => x"82",
          2371 => x"f0",
          2372 => x"d8",
          2373 => x"05",
          2374 => x"73",
          2375 => x"d4",
          2376 => x"08",
          2377 => x"53",
          2378 => x"72",
          2379 => x"08",
          2380 => x"72",
          2381 => x"53",
          2382 => x"09",
          2383 => x"38",
          2384 => x"08",
          2385 => x"70",
          2386 => x"71",
          2387 => x"39",
          2388 => x"08",
          2389 => x"53",
          2390 => x"09",
          2391 => x"38",
          2392 => x"d8",
          2393 => x"05",
          2394 => x"d4",
          2395 => x"08",
          2396 => x"05",
          2397 => x"08",
          2398 => x"33",
          2399 => x"08",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"72",
          2403 => x"81",
          2404 => x"38",
          2405 => x"08",
          2406 => x"70",
          2407 => x"71",
          2408 => x"51",
          2409 => x"82",
          2410 => x"f8",
          2411 => x"d8",
          2412 => x"05",
          2413 => x"d4",
          2414 => x"0c",
          2415 => x"08",
          2416 => x"80",
          2417 => x"38",
          2418 => x"08",
          2419 => x"80",
          2420 => x"38",
          2421 => x"90",
          2422 => x"d4",
          2423 => x"34",
          2424 => x"08",
          2425 => x"70",
          2426 => x"71",
          2427 => x"51",
          2428 => x"82",
          2429 => x"f8",
          2430 => x"a4",
          2431 => x"82",
          2432 => x"f4",
          2433 => x"d8",
          2434 => x"05",
          2435 => x"81",
          2436 => x"70",
          2437 => x"72",
          2438 => x"d4",
          2439 => x"34",
          2440 => x"82",
          2441 => x"f8",
          2442 => x"72",
          2443 => x"38",
          2444 => x"d8",
          2445 => x"05",
          2446 => x"39",
          2447 => x"08",
          2448 => x"53",
          2449 => x"90",
          2450 => x"d4",
          2451 => x"33",
          2452 => x"26",
          2453 => x"39",
          2454 => x"d8",
          2455 => x"05",
          2456 => x"39",
          2457 => x"d8",
          2458 => x"05",
          2459 => x"82",
          2460 => x"f8",
          2461 => x"af",
          2462 => x"38",
          2463 => x"08",
          2464 => x"53",
          2465 => x"83",
          2466 => x"80",
          2467 => x"d4",
          2468 => x"0c",
          2469 => x"8a",
          2470 => x"d4",
          2471 => x"34",
          2472 => x"d8",
          2473 => x"05",
          2474 => x"d4",
          2475 => x"33",
          2476 => x"27",
          2477 => x"82",
          2478 => x"f8",
          2479 => x"80",
          2480 => x"94",
          2481 => x"d4",
          2482 => x"33",
          2483 => x"53",
          2484 => x"d4",
          2485 => x"34",
          2486 => x"08",
          2487 => x"d0",
          2488 => x"72",
          2489 => x"08",
          2490 => x"82",
          2491 => x"f8",
          2492 => x"90",
          2493 => x"38",
          2494 => x"08",
          2495 => x"f9",
          2496 => x"72",
          2497 => x"08",
          2498 => x"82",
          2499 => x"f8",
          2500 => x"72",
          2501 => x"38",
          2502 => x"d8",
          2503 => x"05",
          2504 => x"39",
          2505 => x"08",
          2506 => x"82",
          2507 => x"f4",
          2508 => x"54",
          2509 => x"8d",
          2510 => x"82",
          2511 => x"ec",
          2512 => x"f7",
          2513 => x"d4",
          2514 => x"33",
          2515 => x"d4",
          2516 => x"08",
          2517 => x"d4",
          2518 => x"33",
          2519 => x"d8",
          2520 => x"05",
          2521 => x"d4",
          2522 => x"08",
          2523 => x"05",
          2524 => x"08",
          2525 => x"55",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"a5",
          2529 => x"d4",
          2530 => x"33",
          2531 => x"2e",
          2532 => x"d8",
          2533 => x"05",
          2534 => x"d8",
          2535 => x"05",
          2536 => x"d4",
          2537 => x"08",
          2538 => x"08",
          2539 => x"71",
          2540 => x"0b",
          2541 => x"08",
          2542 => x"82",
          2543 => x"ec",
          2544 => x"d8",
          2545 => x"3d",
          2546 => x"d4",
          2547 => x"d8",
          2548 => x"82",
          2549 => x"f7",
          2550 => x"0b",
          2551 => x"08",
          2552 => x"82",
          2553 => x"8c",
          2554 => x"80",
          2555 => x"d8",
          2556 => x"05",
          2557 => x"51",
          2558 => x"53",
          2559 => x"d4",
          2560 => x"34",
          2561 => x"06",
          2562 => x"2e",
          2563 => x"91",
          2564 => x"d4",
          2565 => x"08",
          2566 => x"05",
          2567 => x"ce",
          2568 => x"d4",
          2569 => x"33",
          2570 => x"2e",
          2571 => x"a4",
          2572 => x"82",
          2573 => x"f0",
          2574 => x"d8",
          2575 => x"05",
          2576 => x"81",
          2577 => x"70",
          2578 => x"72",
          2579 => x"d4",
          2580 => x"34",
          2581 => x"08",
          2582 => x"53",
          2583 => x"09",
          2584 => x"dc",
          2585 => x"d4",
          2586 => x"08",
          2587 => x"05",
          2588 => x"08",
          2589 => x"33",
          2590 => x"08",
          2591 => x"82",
          2592 => x"f8",
          2593 => x"d8",
          2594 => x"05",
          2595 => x"d4",
          2596 => x"08",
          2597 => x"b6",
          2598 => x"d4",
          2599 => x"08",
          2600 => x"84",
          2601 => x"39",
          2602 => x"d8",
          2603 => x"05",
          2604 => x"d4",
          2605 => x"08",
          2606 => x"05",
          2607 => x"08",
          2608 => x"33",
          2609 => x"08",
          2610 => x"81",
          2611 => x"0b",
          2612 => x"08",
          2613 => x"82",
          2614 => x"88",
          2615 => x"08",
          2616 => x"0c",
          2617 => x"53",
          2618 => x"d8",
          2619 => x"05",
          2620 => x"39",
          2621 => x"08",
          2622 => x"53",
          2623 => x"8d",
          2624 => x"82",
          2625 => x"ec",
          2626 => x"80",
          2627 => x"d4",
          2628 => x"33",
          2629 => x"27",
          2630 => x"d8",
          2631 => x"05",
          2632 => x"b9",
          2633 => x"8d",
          2634 => x"82",
          2635 => x"ec",
          2636 => x"d8",
          2637 => x"82",
          2638 => x"f4",
          2639 => x"39",
          2640 => x"08",
          2641 => x"53",
          2642 => x"90",
          2643 => x"d4",
          2644 => x"33",
          2645 => x"26",
          2646 => x"39",
          2647 => x"d8",
          2648 => x"05",
          2649 => x"39",
          2650 => x"d8",
          2651 => x"05",
          2652 => x"82",
          2653 => x"fc",
          2654 => x"d8",
          2655 => x"05",
          2656 => x"73",
          2657 => x"38",
          2658 => x"08",
          2659 => x"53",
          2660 => x"27",
          2661 => x"d8",
          2662 => x"05",
          2663 => x"51",
          2664 => x"d8",
          2665 => x"05",
          2666 => x"d4",
          2667 => x"33",
          2668 => x"53",
          2669 => x"d4",
          2670 => x"34",
          2671 => x"08",
          2672 => x"53",
          2673 => x"ad",
          2674 => x"d4",
          2675 => x"33",
          2676 => x"53",
          2677 => x"d4",
          2678 => x"34",
          2679 => x"08",
          2680 => x"53",
          2681 => x"8d",
          2682 => x"82",
          2683 => x"ec",
          2684 => x"98",
          2685 => x"d4",
          2686 => x"33",
          2687 => x"08",
          2688 => x"54",
          2689 => x"26",
          2690 => x"0b",
          2691 => x"08",
          2692 => x"80",
          2693 => x"d8",
          2694 => x"05",
          2695 => x"d8",
          2696 => x"05",
          2697 => x"d8",
          2698 => x"05",
          2699 => x"82",
          2700 => x"fc",
          2701 => x"d8",
          2702 => x"05",
          2703 => x"81",
          2704 => x"70",
          2705 => x"52",
          2706 => x"33",
          2707 => x"08",
          2708 => x"fe",
          2709 => x"d8",
          2710 => x"05",
          2711 => x"80",
          2712 => x"82",
          2713 => x"fc",
          2714 => x"82",
          2715 => x"fc",
          2716 => x"d8",
          2717 => x"05",
          2718 => x"d4",
          2719 => x"08",
          2720 => x"81",
          2721 => x"d4",
          2722 => x"0c",
          2723 => x"08",
          2724 => x"82",
          2725 => x"8b",
          2726 => x"d8",
          2727 => x"f9",
          2728 => x"70",
          2729 => x"56",
          2730 => x"2e",
          2731 => x"95",
          2732 => x"51",
          2733 => x"82",
          2734 => x"15",
          2735 => x"16",
          2736 => x"cd",
          2737 => x"54",
          2738 => x"09",
          2739 => x"38",
          2740 => x"f1",
          2741 => x"76",
          2742 => x"d3",
          2743 => x"08",
          2744 => x"a3",
          2745 => x"c8",
          2746 => x"52",
          2747 => x"e9",
          2748 => x"d8",
          2749 => x"38",
          2750 => x"54",
          2751 => x"ff",
          2752 => x"17",
          2753 => x"06",
          2754 => x"77",
          2755 => x"ff",
          2756 => x"d8",
          2757 => x"3d",
          2758 => x"3d",
          2759 => x"71",
          2760 => x"8e",
          2761 => x"29",
          2762 => x"05",
          2763 => x"04",
          2764 => x"51",
          2765 => x"82",
          2766 => x"80",
          2767 => x"b5",
          2768 => x"f2",
          2769 => x"90",
          2770 => x"39",
          2771 => x"51",
          2772 => x"82",
          2773 => x"80",
          2774 => x"b5",
          2775 => x"d6",
          2776 => x"d4",
          2777 => x"39",
          2778 => x"51",
          2779 => x"82",
          2780 => x"80",
          2781 => x"b6",
          2782 => x"39",
          2783 => x"51",
          2784 => x"b6",
          2785 => x"39",
          2786 => x"51",
          2787 => x"b7",
          2788 => x"39",
          2789 => x"51",
          2790 => x"b7",
          2791 => x"39",
          2792 => x"51",
          2793 => x"b7",
          2794 => x"39",
          2795 => x"51",
          2796 => x"b8",
          2797 => x"ad",
          2798 => x"0d",
          2799 => x"0d",
          2800 => x"56",
          2801 => x"26",
          2802 => x"52",
          2803 => x"29",
          2804 => x"87",
          2805 => x"51",
          2806 => x"82",
          2807 => x"52",
          2808 => x"a1",
          2809 => x"c8",
          2810 => x"53",
          2811 => x"b8",
          2812 => x"bb",
          2813 => x"3d",
          2814 => x"3d",
          2815 => x"84",
          2816 => x"05",
          2817 => x"80",
          2818 => x"70",
          2819 => x"25",
          2820 => x"59",
          2821 => x"87",
          2822 => x"38",
          2823 => x"76",
          2824 => x"ff",
          2825 => x"93",
          2826 => x"82",
          2827 => x"76",
          2828 => x"70",
          2829 => x"96",
          2830 => x"d8",
          2831 => x"82",
          2832 => x"b9",
          2833 => x"c8",
          2834 => x"98",
          2835 => x"d8",
          2836 => x"96",
          2837 => x"54",
          2838 => x"77",
          2839 => x"81",
          2840 => x"82",
          2841 => x"57",
          2842 => x"08",
          2843 => x"55",
          2844 => x"89",
          2845 => x"75",
          2846 => x"d7",
          2847 => x"d8",
          2848 => x"a2",
          2849 => x"30",
          2850 => x"80",
          2851 => x"70",
          2852 => x"06",
          2853 => x"56",
          2854 => x"90",
          2855 => x"bc",
          2856 => x"98",
          2857 => x"78",
          2858 => x"3f",
          2859 => x"82",
          2860 => x"96",
          2861 => x"f7",
          2862 => x"02",
          2863 => x"05",
          2864 => x"ff",
          2865 => x"7c",
          2866 => x"fe",
          2867 => x"d8",
          2868 => x"cb",
          2869 => x"2e",
          2870 => x"81",
          2871 => x"bf",
          2872 => x"a8",
          2873 => x"a8",
          2874 => x"a8",
          2875 => x"b0",
          2876 => x"f4",
          2877 => x"82",
          2878 => x"52",
          2879 => x"51",
          2880 => x"3f",
          2881 => x"56",
          2882 => x"54",
          2883 => x"53",
          2884 => x"51",
          2885 => x"d8",
          2886 => x"83",
          2887 => x"78",
          2888 => x"0c",
          2889 => x"04",
          2890 => x"7f",
          2891 => x"8c",
          2892 => x"05",
          2893 => x"15",
          2894 => x"5c",
          2895 => x"5e",
          2896 => x"b8",
          2897 => x"b9",
          2898 => x"b9",
          2899 => x"b9",
          2900 => x"55",
          2901 => x"81",
          2902 => x"90",
          2903 => x"7b",
          2904 => x"38",
          2905 => x"74",
          2906 => x"7a",
          2907 => x"72",
          2908 => x"b9",
          2909 => x"b8",
          2910 => x"39",
          2911 => x"51",
          2912 => x"3f",
          2913 => x"80",
          2914 => x"18",
          2915 => x"27",
          2916 => x"08",
          2917 => x"f8",
          2918 => x"be",
          2919 => x"82",
          2920 => x"ff",
          2921 => x"84",
          2922 => x"39",
          2923 => x"72",
          2924 => x"38",
          2925 => x"82",
          2926 => x"ff",
          2927 => x"89",
          2928 => x"a0",
          2929 => x"92",
          2930 => x"55",
          2931 => x"08",
          2932 => x"d7",
          2933 => x"fc",
          2934 => x"a4",
          2935 => x"fa",
          2936 => x"74",
          2937 => x"c6",
          2938 => x"70",
          2939 => x"80",
          2940 => x"27",
          2941 => x"56",
          2942 => x"74",
          2943 => x"81",
          2944 => x"06",
          2945 => x"06",
          2946 => x"80",
          2947 => x"73",
          2948 => x"8a",
          2949 => x"ac",
          2950 => x"51",
          2951 => x"f4",
          2952 => x"a0",
          2953 => x"3f",
          2954 => x"ff",
          2955 => x"b9",
          2956 => x"b1",
          2957 => x"79",
          2958 => x"a1",
          2959 => x"d8",
          2960 => x"2b",
          2961 => x"51",
          2962 => x"2e",
          2963 => x"aa",
          2964 => x"3f",
          2965 => x"08",
          2966 => x"98",
          2967 => x"32",
          2968 => x"9b",
          2969 => x"70",
          2970 => x"75",
          2971 => x"58",
          2972 => x"51",
          2973 => x"24",
          2974 => x"9b",
          2975 => x"06",
          2976 => x"53",
          2977 => x"1e",
          2978 => x"26",
          2979 => x"ff",
          2980 => x"d8",
          2981 => x"3d",
          2982 => x"3d",
          2983 => x"05",
          2984 => x"ac",
          2985 => x"b4",
          2986 => x"b6",
          2987 => x"d7",
          2988 => x"a9",
          2989 => x"b9",
          2990 => x"b9",
          2991 => x"d7",
          2992 => x"82",
          2993 => x"ff",
          2994 => x"74",
          2995 => x"38",
          2996 => x"86",
          2997 => x"fe",
          2998 => x"c0",
          2999 => x"53",
          3000 => x"81",
          3001 => x"3f",
          3002 => x"51",
          3003 => x"80",
          3004 => x"3f",
          3005 => x"70",
          3006 => x"52",
          3007 => x"92",
          3008 => x"9c",
          3009 => x"ba",
          3010 => x"ba",
          3011 => x"9c",
          3012 => x"82",
          3013 => x"06",
          3014 => x"80",
          3015 => x"81",
          3016 => x"3f",
          3017 => x"51",
          3018 => x"80",
          3019 => x"3f",
          3020 => x"70",
          3021 => x"52",
          3022 => x"92",
          3023 => x"9b",
          3024 => x"ba",
          3025 => x"fe",
          3026 => x"9b",
          3027 => x"84",
          3028 => x"06",
          3029 => x"80",
          3030 => x"81",
          3031 => x"3f",
          3032 => x"51",
          3033 => x"80",
          3034 => x"3f",
          3035 => x"70",
          3036 => x"52",
          3037 => x"92",
          3038 => x"9b",
          3039 => x"ba",
          3040 => x"c2",
          3041 => x"9b",
          3042 => x"86",
          3043 => x"06",
          3044 => x"80",
          3045 => x"81",
          3046 => x"3f",
          3047 => x"51",
          3048 => x"80",
          3049 => x"3f",
          3050 => x"70",
          3051 => x"52",
          3052 => x"92",
          3053 => x"9a",
          3054 => x"ba",
          3055 => x"86",
          3056 => x"9a",
          3057 => x"88",
          3058 => x"06",
          3059 => x"80",
          3060 => x"81",
          3061 => x"3f",
          3062 => x"51",
          3063 => x"80",
          3064 => x"3f",
          3065 => x"84",
          3066 => x"fb",
          3067 => x"02",
          3068 => x"05",
          3069 => x"56",
          3070 => x"75",
          3071 => x"3f",
          3072 => x"d3",
          3073 => x"73",
          3074 => x"53",
          3075 => x"52",
          3076 => x"51",
          3077 => x"3f",
          3078 => x"08",
          3079 => x"d8",
          3080 => x"80",
          3081 => x"31",
          3082 => x"73",
          3083 => x"d3",
          3084 => x"0b",
          3085 => x"33",
          3086 => x"2e",
          3087 => x"af",
          3088 => x"d8",
          3089 => x"75",
          3090 => x"82",
          3091 => x"c8",
          3092 => x"8b",
          3093 => x"c8",
          3094 => x"89",
          3095 => x"82",
          3096 => x"81",
          3097 => x"82",
          3098 => x"82",
          3099 => x"0b",
          3100 => x"c4",
          3101 => x"82",
          3102 => x"06",
          3103 => x"bb",
          3104 => x"52",
          3105 => x"b2",
          3106 => x"82",
          3107 => x"87",
          3108 => x"ce",
          3109 => x"70",
          3110 => x"d4",
          3111 => x"81",
          3112 => x"80",
          3113 => x"82",
          3114 => x"81",
          3115 => x"78",
          3116 => x"81",
          3117 => x"96",
          3118 => x"53",
          3119 => x"52",
          3120 => x"a3",
          3121 => x"78",
          3122 => x"f4",
          3123 => x"98",
          3124 => x"c8",
          3125 => x"88",
          3126 => x"e8",
          3127 => x"39",
          3128 => x"5d",
          3129 => x"51",
          3130 => x"3f",
          3131 => x"46",
          3132 => x"52",
          3133 => x"f3",
          3134 => x"ff",
          3135 => x"f3",
          3136 => x"d8",
          3137 => x"2b",
          3138 => x"51",
          3139 => x"c1",
          3140 => x"38",
          3141 => x"24",
          3142 => x"78",
          3143 => x"b9",
          3144 => x"24",
          3145 => x"82",
          3146 => x"38",
          3147 => x"8a",
          3148 => x"2e",
          3149 => x"8f",
          3150 => x"84",
          3151 => x"38",
          3152 => x"82",
          3153 => x"f3",
          3154 => x"2e",
          3155 => x"78",
          3156 => x"38",
          3157 => x"83",
          3158 => x"bc",
          3159 => x"38",
          3160 => x"78",
          3161 => x"c4",
          3162 => x"c0",
          3163 => x"38",
          3164 => x"78",
          3165 => x"8d",
          3166 => x"80",
          3167 => x"38",
          3168 => x"2e",
          3169 => x"78",
          3170 => x"92",
          3171 => x"c2",
          3172 => x"38",
          3173 => x"2e",
          3174 => x"8e",
          3175 => x"80",
          3176 => x"ca",
          3177 => x"d4",
          3178 => x"38",
          3179 => x"78",
          3180 => x"8d",
          3181 => x"81",
          3182 => x"38",
          3183 => x"2e",
          3184 => x"78",
          3185 => x"8d",
          3186 => x"ef",
          3187 => x"83",
          3188 => x"38",
          3189 => x"2e",
          3190 => x"8d",
          3191 => x"3d",
          3192 => x"53",
          3193 => x"51",
          3194 => x"82",
          3195 => x"88",
          3196 => x"a4",
          3197 => x"39",
          3198 => x"fc",
          3199 => x"84",
          3200 => x"ca",
          3201 => x"c8",
          3202 => x"88",
          3203 => x"25",
          3204 => x"43",
          3205 => x"05",
          3206 => x"80",
          3207 => x"51",
          3208 => x"3f",
          3209 => x"08",
          3210 => x"59",
          3211 => x"82",
          3212 => x"cb",
          3213 => x"5e",
          3214 => x"82",
          3215 => x"8e",
          3216 => x"3d",
          3217 => x"53",
          3218 => x"51",
          3219 => x"82",
          3220 => x"80",
          3221 => x"38",
          3222 => x"52",
          3223 => x"05",
          3224 => x"cc",
          3225 => x"d8",
          3226 => x"82",
          3227 => x"8c",
          3228 => x"3d",
          3229 => x"53",
          3230 => x"51",
          3231 => x"82",
          3232 => x"80",
          3233 => x"63",
          3234 => x"d8",
          3235 => x"fe",
          3236 => x"ff",
          3237 => x"ea",
          3238 => x"d8",
          3239 => x"38",
          3240 => x"08",
          3241 => x"82",
          3242 => x"79",
          3243 => x"92",
          3244 => x"cb",
          3245 => x"79",
          3246 => x"b8",
          3247 => x"f4",
          3248 => x"88",
          3249 => x"d8",
          3250 => x"8c",
          3251 => x"b4",
          3252 => x"3f",
          3253 => x"8c",
          3254 => x"ff",
          3255 => x"8f",
          3256 => x"d8",
          3257 => x"3d",
          3258 => x"52",
          3259 => x"3f",
          3260 => x"d8",
          3261 => x"7a",
          3262 => x"3f",
          3263 => x"b4",
          3264 => x"05",
          3265 => x"3f",
          3266 => x"08",
          3267 => x"84",
          3268 => x"90",
          3269 => x"d8",
          3270 => x"3d",
          3271 => x"52",
          3272 => x"3f",
          3273 => x"08",
          3274 => x"84",
          3275 => x"90",
          3276 => x"d6",
          3277 => x"d8",
          3278 => x"56",
          3279 => x"d8",
          3280 => x"ff",
          3281 => x"53",
          3282 => x"51",
          3283 => x"82",
          3284 => x"80",
          3285 => x"38",
          3286 => x"08",
          3287 => x"3f",
          3288 => x"b4",
          3289 => x"11",
          3290 => x"05",
          3291 => x"3f",
          3292 => x"08",
          3293 => x"ec",
          3294 => x"fe",
          3295 => x"ff",
          3296 => x"e8",
          3297 => x"d8",
          3298 => x"2e",
          3299 => x"b4",
          3300 => x"11",
          3301 => x"05",
          3302 => x"3f",
          3303 => x"08",
          3304 => x"d8",
          3305 => x"82",
          3306 => x"ff",
          3307 => x"63",
          3308 => x"79",
          3309 => x"ec",
          3310 => x"78",
          3311 => x"05",
          3312 => x"7a",
          3313 => x"81",
          3314 => x"3d",
          3315 => x"53",
          3316 => x"51",
          3317 => x"82",
          3318 => x"80",
          3319 => x"38",
          3320 => x"fc",
          3321 => x"84",
          3322 => x"e2",
          3323 => x"c8",
          3324 => x"f9",
          3325 => x"3d",
          3326 => x"53",
          3327 => x"51",
          3328 => x"82",
          3329 => x"80",
          3330 => x"38",
          3331 => x"51",
          3332 => x"3f",
          3333 => x"63",
          3334 => x"38",
          3335 => x"70",
          3336 => x"33",
          3337 => x"81",
          3338 => x"39",
          3339 => x"80",
          3340 => x"84",
          3341 => x"96",
          3342 => x"c8",
          3343 => x"f9",
          3344 => x"3d",
          3345 => x"53",
          3346 => x"51",
          3347 => x"82",
          3348 => x"80",
          3349 => x"38",
          3350 => x"f8",
          3351 => x"84",
          3352 => x"ea",
          3353 => x"c8",
          3354 => x"f8",
          3355 => x"bd",
          3356 => x"aa",
          3357 => x"5a",
          3358 => x"a8",
          3359 => x"33",
          3360 => x"5a",
          3361 => x"2e",
          3362 => x"55",
          3363 => x"33",
          3364 => x"82",
          3365 => x"ff",
          3366 => x"81",
          3367 => x"05",
          3368 => x"39",
          3369 => x"df",
          3370 => x"39",
          3371 => x"80",
          3372 => x"84",
          3373 => x"96",
          3374 => x"c8",
          3375 => x"38",
          3376 => x"33",
          3377 => x"2e",
          3378 => x"d6",
          3379 => x"80",
          3380 => x"d7",
          3381 => x"78",
          3382 => x"38",
          3383 => x"08",
          3384 => x"82",
          3385 => x"59",
          3386 => x"88",
          3387 => x"fc",
          3388 => x"39",
          3389 => x"33",
          3390 => x"2e",
          3391 => x"d7",
          3392 => x"9a",
          3393 => x"b2",
          3394 => x"80",
          3395 => x"82",
          3396 => x"44",
          3397 => x"d7",
          3398 => x"80",
          3399 => x"3d",
          3400 => x"53",
          3401 => x"51",
          3402 => x"82",
          3403 => x"80",
          3404 => x"d7",
          3405 => x"78",
          3406 => x"38",
          3407 => x"08",
          3408 => x"39",
          3409 => x"33",
          3410 => x"2e",
          3411 => x"d6",
          3412 => x"bb",
          3413 => x"b6",
          3414 => x"80",
          3415 => x"82",
          3416 => x"43",
          3417 => x"d7",
          3418 => x"78",
          3419 => x"38",
          3420 => x"08",
          3421 => x"82",
          3422 => x"59",
          3423 => x"88",
          3424 => x"90",
          3425 => x"39",
          3426 => x"08",
          3427 => x"b4",
          3428 => x"11",
          3429 => x"05",
          3430 => x"3f",
          3431 => x"08",
          3432 => x"38",
          3433 => x"5c",
          3434 => x"83",
          3435 => x"7a",
          3436 => x"30",
          3437 => x"9f",
          3438 => x"06",
          3439 => x"5a",
          3440 => x"88",
          3441 => x"2e",
          3442 => x"42",
          3443 => x"51",
          3444 => x"a0",
          3445 => x"61",
          3446 => x"63",
          3447 => x"3f",
          3448 => x"51",
          3449 => x"b4",
          3450 => x"11",
          3451 => x"05",
          3452 => x"3f",
          3453 => x"08",
          3454 => x"e8",
          3455 => x"fe",
          3456 => x"ff",
          3457 => x"e3",
          3458 => x"d8",
          3459 => x"2e",
          3460 => x"59",
          3461 => x"05",
          3462 => x"63",
          3463 => x"b4",
          3464 => x"11",
          3465 => x"05",
          3466 => x"3f",
          3467 => x"08",
          3468 => x"b0",
          3469 => x"33",
          3470 => x"bd",
          3471 => x"a7",
          3472 => x"f4",
          3473 => x"80",
          3474 => x"51",
          3475 => x"3f",
          3476 => x"33",
          3477 => x"2e",
          3478 => x"9f",
          3479 => x"38",
          3480 => x"fc",
          3481 => x"84",
          3482 => x"e2",
          3483 => x"c8",
          3484 => x"91",
          3485 => x"02",
          3486 => x"33",
          3487 => x"81",
          3488 => x"b1",
          3489 => x"d4",
          3490 => x"3f",
          3491 => x"b4",
          3492 => x"11",
          3493 => x"05",
          3494 => x"3f",
          3495 => x"08",
          3496 => x"c0",
          3497 => x"fe",
          3498 => x"ff",
          3499 => x"dc",
          3500 => x"d8",
          3501 => x"2e",
          3502 => x"59",
          3503 => x"22",
          3504 => x"05",
          3505 => x"41",
          3506 => x"f0",
          3507 => x"84",
          3508 => x"a9",
          3509 => x"c8",
          3510 => x"f4",
          3511 => x"70",
          3512 => x"82",
          3513 => x"ff",
          3514 => x"82",
          3515 => x"53",
          3516 => x"79",
          3517 => x"b7",
          3518 => x"79",
          3519 => x"ae",
          3520 => x"38",
          3521 => x"87",
          3522 => x"05",
          3523 => x"b4",
          3524 => x"11",
          3525 => x"05",
          3526 => x"3f",
          3527 => x"08",
          3528 => x"38",
          3529 => x"be",
          3530 => x"70",
          3531 => x"23",
          3532 => x"aa",
          3533 => x"d4",
          3534 => x"3f",
          3535 => x"b4",
          3536 => x"11",
          3537 => x"05",
          3538 => x"3f",
          3539 => x"08",
          3540 => x"90",
          3541 => x"fe",
          3542 => x"ff",
          3543 => x"db",
          3544 => x"d8",
          3545 => x"2e",
          3546 => x"60",
          3547 => x"60",
          3548 => x"b4",
          3549 => x"11",
          3550 => x"05",
          3551 => x"3f",
          3552 => x"08",
          3553 => x"dc",
          3554 => x"08",
          3555 => x"bd",
          3556 => x"a4",
          3557 => x"f4",
          3558 => x"80",
          3559 => x"51",
          3560 => x"3f",
          3561 => x"33",
          3562 => x"2e",
          3563 => x"9f",
          3564 => x"38",
          3565 => x"f0",
          3566 => x"84",
          3567 => x"bd",
          3568 => x"c8",
          3569 => x"8d",
          3570 => x"71",
          3571 => x"84",
          3572 => x"b5",
          3573 => x"d4",
          3574 => x"3f",
          3575 => x"82",
          3576 => x"c0",
          3577 => x"51",
          3578 => x"f1",
          3579 => x"be",
          3580 => x"bf",
          3581 => x"51",
          3582 => x"f1",
          3583 => x"be",
          3584 => x"bf",
          3585 => x"80",
          3586 => x"c0",
          3587 => x"84",
          3588 => x"87",
          3589 => x"0c",
          3590 => x"82",
          3591 => x"ff",
          3592 => x"8c",
          3593 => x"87",
          3594 => x"0c",
          3595 => x"0b",
          3596 => x"94",
          3597 => x"39",
          3598 => x"80",
          3599 => x"84",
          3600 => x"8a",
          3601 => x"c8",
          3602 => x"f1",
          3603 => x"52",
          3604 => x"51",
          3605 => x"3f",
          3606 => x"04",
          3607 => x"80",
          3608 => x"84",
          3609 => x"e6",
          3610 => x"c8",
          3611 => x"f0",
          3612 => x"52",
          3613 => x"51",
          3614 => x"3f",
          3615 => x"2d",
          3616 => x"08",
          3617 => x"dc",
          3618 => x"c8",
          3619 => x"bf",
          3620 => x"a2",
          3621 => x"cc",
          3622 => x"9c",
          3623 => x"c5",
          3624 => x"97",
          3625 => x"39",
          3626 => x"51",
          3627 => x"3f",
          3628 => x"a6",
          3629 => x"3f",
          3630 => x"79",
          3631 => x"59",
          3632 => x"f0",
          3633 => x"7d",
          3634 => x"80",
          3635 => x"38",
          3636 => x"84",
          3637 => x"cb",
          3638 => x"c8",
          3639 => x"5c",
          3640 => x"b2",
          3641 => x"24",
          3642 => x"81",
          3643 => x"80",
          3644 => x"83",
          3645 => x"80",
          3646 => x"bf",
          3647 => x"55",
          3648 => x"54",
          3649 => x"bf",
          3650 => x"3d",
          3651 => x"51",
          3652 => x"3f",
          3653 => x"52",
          3654 => x"b0",
          3655 => x"d5",
          3656 => x"7a",
          3657 => x"d0",
          3658 => x"82",
          3659 => x"b4",
          3660 => x"05",
          3661 => x"8a",
          3662 => x"7a",
          3663 => x"82",
          3664 => x"b4",
          3665 => x"05",
          3666 => x"f6",
          3667 => x"ec",
          3668 => x"f8",
          3669 => x"64",
          3670 => x"84",
          3671 => x"84",
          3672 => x"b4",
          3673 => x"05",
          3674 => x"3f",
          3675 => x"08",
          3676 => x"08",
          3677 => x"70",
          3678 => x"25",
          3679 => x"5f",
          3680 => x"83",
          3681 => x"81",
          3682 => x"06",
          3683 => x"2e",
          3684 => x"1c",
          3685 => x"06",
          3686 => x"fe",
          3687 => x"81",
          3688 => x"32",
          3689 => x"8a",
          3690 => x"2e",
          3691 => x"ee",
          3692 => x"bf",
          3693 => x"bc",
          3694 => x"a8",
          3695 => x"0d",
          3696 => x"d8",
          3697 => x"c0",
          3698 => x"08",
          3699 => x"84",
          3700 => x"51",
          3701 => x"82",
          3702 => x"90",
          3703 => x"55",
          3704 => x"80",
          3705 => x"d3",
          3706 => x"82",
          3707 => x"07",
          3708 => x"c0",
          3709 => x"08",
          3710 => x"84",
          3711 => x"51",
          3712 => x"82",
          3713 => x"90",
          3714 => x"55",
          3715 => x"80",
          3716 => x"d2",
          3717 => x"82",
          3718 => x"07",
          3719 => x"80",
          3720 => x"c0",
          3721 => x"8c",
          3722 => x"87",
          3723 => x"0c",
          3724 => x"5a",
          3725 => x"5b",
          3726 => x"05",
          3727 => x"80",
          3728 => x"a8",
          3729 => x"70",
          3730 => x"70",
          3731 => x"f4",
          3732 => x"89",
          3733 => x"c0",
          3734 => x"88",
          3735 => x"85",
          3736 => x"94",
          3737 => x"fd",
          3738 => x"d5",
          3739 => x"3f",
          3740 => x"a6",
          3741 => x"3f",
          3742 => x"3d",
          3743 => x"83",
          3744 => x"2b",
          3745 => x"3f",
          3746 => x"08",
          3747 => x"72",
          3748 => x"54",
          3749 => x"25",
          3750 => x"82",
          3751 => x"84",
          3752 => x"fc",
          3753 => x"70",
          3754 => x"80",
          3755 => x"72",
          3756 => x"8a",
          3757 => x"51",
          3758 => x"09",
          3759 => x"38",
          3760 => x"f1",
          3761 => x"51",
          3762 => x"09",
          3763 => x"38",
          3764 => x"81",
          3765 => x"73",
          3766 => x"81",
          3767 => x"84",
          3768 => x"52",
          3769 => x"52",
          3770 => x"2e",
          3771 => x"54",
          3772 => x"9d",
          3773 => x"38",
          3774 => x"12",
          3775 => x"33",
          3776 => x"a0",
          3777 => x"81",
          3778 => x"2e",
          3779 => x"ea",
          3780 => x"33",
          3781 => x"a0",
          3782 => x"06",
          3783 => x"54",
          3784 => x"70",
          3785 => x"25",
          3786 => x"51",
          3787 => x"2e",
          3788 => x"72",
          3789 => x"54",
          3790 => x"0c",
          3791 => x"82",
          3792 => x"86",
          3793 => x"fc",
          3794 => x"53",
          3795 => x"2e",
          3796 => x"3d",
          3797 => x"72",
          3798 => x"3f",
          3799 => x"08",
          3800 => x"53",
          3801 => x"53",
          3802 => x"c8",
          3803 => x"0d",
          3804 => x"0d",
          3805 => x"33",
          3806 => x"53",
          3807 => x"8b",
          3808 => x"38",
          3809 => x"ff",
          3810 => x"52",
          3811 => x"81",
          3812 => x"13",
          3813 => x"52",
          3814 => x"80",
          3815 => x"13",
          3816 => x"52",
          3817 => x"80",
          3818 => x"13",
          3819 => x"52",
          3820 => x"80",
          3821 => x"13",
          3822 => x"52",
          3823 => x"26",
          3824 => x"8a",
          3825 => x"87",
          3826 => x"e7",
          3827 => x"38",
          3828 => x"c0",
          3829 => x"72",
          3830 => x"98",
          3831 => x"13",
          3832 => x"98",
          3833 => x"13",
          3834 => x"98",
          3835 => x"13",
          3836 => x"98",
          3837 => x"13",
          3838 => x"98",
          3839 => x"13",
          3840 => x"98",
          3841 => x"87",
          3842 => x"0c",
          3843 => x"98",
          3844 => x"0b",
          3845 => x"9c",
          3846 => x"71",
          3847 => x"0c",
          3848 => x"04",
          3849 => x"7f",
          3850 => x"98",
          3851 => x"7d",
          3852 => x"98",
          3853 => x"7d",
          3854 => x"c0",
          3855 => x"5a",
          3856 => x"34",
          3857 => x"b4",
          3858 => x"83",
          3859 => x"c0",
          3860 => x"5a",
          3861 => x"34",
          3862 => x"ac",
          3863 => x"85",
          3864 => x"c0",
          3865 => x"5a",
          3866 => x"34",
          3867 => x"a4",
          3868 => x"88",
          3869 => x"c0",
          3870 => x"5a",
          3871 => x"23",
          3872 => x"79",
          3873 => x"06",
          3874 => x"ff",
          3875 => x"86",
          3876 => x"85",
          3877 => x"84",
          3878 => x"83",
          3879 => x"82",
          3880 => x"7d",
          3881 => x"06",
          3882 => x"ac",
          3883 => x"aa",
          3884 => x"0d",
          3885 => x"0d",
          3886 => x"33",
          3887 => x"33",
          3888 => x"06",
          3889 => x"87",
          3890 => x"51",
          3891 => x"86",
          3892 => x"94",
          3893 => x"08",
          3894 => x"70",
          3895 => x"54",
          3896 => x"2e",
          3897 => x"91",
          3898 => x"06",
          3899 => x"d7",
          3900 => x"32",
          3901 => x"51",
          3902 => x"2e",
          3903 => x"93",
          3904 => x"06",
          3905 => x"ff",
          3906 => x"81",
          3907 => x"87",
          3908 => x"52",
          3909 => x"86",
          3910 => x"94",
          3911 => x"72",
          3912 => x"d8",
          3913 => x"3d",
          3914 => x"3d",
          3915 => x"05",
          3916 => x"70",
          3917 => x"52",
          3918 => x"d6",
          3919 => x"3d",
          3920 => x"3d",
          3921 => x"05",
          3922 => x"8a",
          3923 => x"06",
          3924 => x"52",
          3925 => x"3f",
          3926 => x"33",
          3927 => x"06",
          3928 => x"c0",
          3929 => x"76",
          3930 => x"38",
          3931 => x"94",
          3932 => x"70",
          3933 => x"81",
          3934 => x"54",
          3935 => x"8c",
          3936 => x"2a",
          3937 => x"51",
          3938 => x"38",
          3939 => x"70",
          3940 => x"53",
          3941 => x"8d",
          3942 => x"2a",
          3943 => x"51",
          3944 => x"be",
          3945 => x"ff",
          3946 => x"c0",
          3947 => x"72",
          3948 => x"38",
          3949 => x"90",
          3950 => x"0c",
          3951 => x"d8",
          3952 => x"3d",
          3953 => x"3d",
          3954 => x"80",
          3955 => x"81",
          3956 => x"53",
          3957 => x"2e",
          3958 => x"71",
          3959 => x"81",
          3960 => x"e8",
          3961 => x"ff",
          3962 => x"55",
          3963 => x"94",
          3964 => x"80",
          3965 => x"87",
          3966 => x"51",
          3967 => x"96",
          3968 => x"06",
          3969 => x"70",
          3970 => x"38",
          3971 => x"70",
          3972 => x"51",
          3973 => x"72",
          3974 => x"81",
          3975 => x"70",
          3976 => x"38",
          3977 => x"70",
          3978 => x"51",
          3979 => x"38",
          3980 => x"06",
          3981 => x"94",
          3982 => x"80",
          3983 => x"87",
          3984 => x"52",
          3985 => x"81",
          3986 => x"70",
          3987 => x"53",
          3988 => x"ff",
          3989 => x"82",
          3990 => x"89",
          3991 => x"fe",
          3992 => x"d6",
          3993 => x"81",
          3994 => x"52",
          3995 => x"84",
          3996 => x"2e",
          3997 => x"c0",
          3998 => x"70",
          3999 => x"2a",
          4000 => x"51",
          4001 => x"80",
          4002 => x"71",
          4003 => x"51",
          4004 => x"80",
          4005 => x"2e",
          4006 => x"c0",
          4007 => x"71",
          4008 => x"ff",
          4009 => x"c8",
          4010 => x"3d",
          4011 => x"af",
          4012 => x"c8",
          4013 => x"06",
          4014 => x"0c",
          4015 => x"0d",
          4016 => x"33",
          4017 => x"06",
          4018 => x"c0",
          4019 => x"70",
          4020 => x"38",
          4021 => x"94",
          4022 => x"70",
          4023 => x"81",
          4024 => x"51",
          4025 => x"80",
          4026 => x"72",
          4027 => x"51",
          4028 => x"80",
          4029 => x"2e",
          4030 => x"c0",
          4031 => x"71",
          4032 => x"2b",
          4033 => x"51",
          4034 => x"82",
          4035 => x"84",
          4036 => x"ff",
          4037 => x"c0",
          4038 => x"70",
          4039 => x"06",
          4040 => x"80",
          4041 => x"38",
          4042 => x"a4",
          4043 => x"ec",
          4044 => x"9e",
          4045 => x"d6",
          4046 => x"c0",
          4047 => x"82",
          4048 => x"87",
          4049 => x"08",
          4050 => x"0c",
          4051 => x"9c",
          4052 => x"fc",
          4053 => x"9e",
          4054 => x"d7",
          4055 => x"c0",
          4056 => x"82",
          4057 => x"87",
          4058 => x"08",
          4059 => x"0c",
          4060 => x"b4",
          4061 => x"8c",
          4062 => x"9e",
          4063 => x"d7",
          4064 => x"c0",
          4065 => x"82",
          4066 => x"87",
          4067 => x"08",
          4068 => x"0c",
          4069 => x"c4",
          4070 => x"9c",
          4071 => x"9e",
          4072 => x"70",
          4073 => x"23",
          4074 => x"84",
          4075 => x"a4",
          4076 => x"9e",
          4077 => x"d7",
          4078 => x"c0",
          4079 => x"82",
          4080 => x"81",
          4081 => x"b0",
          4082 => x"87",
          4083 => x"08",
          4084 => x"0a",
          4085 => x"52",
          4086 => x"83",
          4087 => x"71",
          4088 => x"34",
          4089 => x"c0",
          4090 => x"70",
          4091 => x"06",
          4092 => x"70",
          4093 => x"38",
          4094 => x"82",
          4095 => x"80",
          4096 => x"9e",
          4097 => x"90",
          4098 => x"51",
          4099 => x"80",
          4100 => x"81",
          4101 => x"d7",
          4102 => x"0b",
          4103 => x"90",
          4104 => x"80",
          4105 => x"52",
          4106 => x"2e",
          4107 => x"52",
          4108 => x"b4",
          4109 => x"87",
          4110 => x"08",
          4111 => x"80",
          4112 => x"52",
          4113 => x"83",
          4114 => x"71",
          4115 => x"34",
          4116 => x"c0",
          4117 => x"70",
          4118 => x"06",
          4119 => x"70",
          4120 => x"38",
          4121 => x"82",
          4122 => x"80",
          4123 => x"9e",
          4124 => x"84",
          4125 => x"51",
          4126 => x"80",
          4127 => x"81",
          4128 => x"d7",
          4129 => x"0b",
          4130 => x"90",
          4131 => x"80",
          4132 => x"52",
          4133 => x"2e",
          4134 => x"52",
          4135 => x"b8",
          4136 => x"87",
          4137 => x"08",
          4138 => x"80",
          4139 => x"52",
          4140 => x"83",
          4141 => x"71",
          4142 => x"34",
          4143 => x"c0",
          4144 => x"70",
          4145 => x"06",
          4146 => x"70",
          4147 => x"38",
          4148 => x"82",
          4149 => x"80",
          4150 => x"9e",
          4151 => x"a0",
          4152 => x"52",
          4153 => x"2e",
          4154 => x"52",
          4155 => x"bb",
          4156 => x"9e",
          4157 => x"98",
          4158 => x"8a",
          4159 => x"51",
          4160 => x"bc",
          4161 => x"87",
          4162 => x"08",
          4163 => x"06",
          4164 => x"70",
          4165 => x"38",
          4166 => x"82",
          4167 => x"87",
          4168 => x"08",
          4169 => x"06",
          4170 => x"51",
          4171 => x"82",
          4172 => x"80",
          4173 => x"9e",
          4174 => x"88",
          4175 => x"52",
          4176 => x"83",
          4177 => x"71",
          4178 => x"34",
          4179 => x"90",
          4180 => x"06",
          4181 => x"82",
          4182 => x"83",
          4183 => x"fb",
          4184 => x"c0",
          4185 => x"90",
          4186 => x"d7",
          4187 => x"73",
          4188 => x"38",
          4189 => x"51",
          4190 => x"3f",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"33",
          4194 => x"2e",
          4195 => x"d7",
          4196 => x"d7",
          4197 => x"54",
          4198 => x"84",
          4199 => x"ba",
          4200 => x"b7",
          4201 => x"80",
          4202 => x"82",
          4203 => x"82",
          4204 => x"11",
          4205 => x"c1",
          4206 => x"90",
          4207 => x"d7",
          4208 => x"73",
          4209 => x"38",
          4210 => x"08",
          4211 => x"08",
          4212 => x"82",
          4213 => x"ff",
          4214 => x"82",
          4215 => x"54",
          4216 => x"94",
          4217 => x"f4",
          4218 => x"f8",
          4219 => x"52",
          4220 => x"51",
          4221 => x"3f",
          4222 => x"33",
          4223 => x"2e",
          4224 => x"d6",
          4225 => x"d7",
          4226 => x"54",
          4227 => x"f4",
          4228 => x"c6",
          4229 => x"bb",
          4230 => x"80",
          4231 => x"82",
          4232 => x"52",
          4233 => x"51",
          4234 => x"3f",
          4235 => x"33",
          4236 => x"2e",
          4237 => x"d7",
          4238 => x"82",
          4239 => x"ff",
          4240 => x"82",
          4241 => x"54",
          4242 => x"8e",
          4243 => x"be",
          4244 => x"c2",
          4245 => x"8f",
          4246 => x"d7",
          4247 => x"73",
          4248 => x"38",
          4249 => x"51",
          4250 => x"3f",
          4251 => x"33",
          4252 => x"2e",
          4253 => x"c3",
          4254 => x"aa",
          4255 => x"d7",
          4256 => x"73",
          4257 => x"38",
          4258 => x"51",
          4259 => x"3f",
          4260 => x"33",
          4261 => x"2e",
          4262 => x"c3",
          4263 => x"aa",
          4264 => x"d7",
          4265 => x"73",
          4266 => x"38",
          4267 => x"51",
          4268 => x"3f",
          4269 => x"51",
          4270 => x"3f",
          4271 => x"08",
          4272 => x"b8",
          4273 => x"92",
          4274 => x"98",
          4275 => x"c3",
          4276 => x"8e",
          4277 => x"d7",
          4278 => x"82",
          4279 => x"ff",
          4280 => x"82",
          4281 => x"ff",
          4282 => x"82",
          4283 => x"52",
          4284 => x"51",
          4285 => x"3f",
          4286 => x"08",
          4287 => x"c0",
          4288 => x"c1",
          4289 => x"d8",
          4290 => x"84",
          4291 => x"71",
          4292 => x"82",
          4293 => x"52",
          4294 => x"51",
          4295 => x"3f",
          4296 => x"33",
          4297 => x"2e",
          4298 => x"d7",
          4299 => x"bd",
          4300 => x"75",
          4301 => x"3f",
          4302 => x"08",
          4303 => x"29",
          4304 => x"54",
          4305 => x"c8",
          4306 => x"c5",
          4307 => x"8d",
          4308 => x"d7",
          4309 => x"73",
          4310 => x"38",
          4311 => x"08",
          4312 => x"c0",
          4313 => x"c0",
          4314 => x"d8",
          4315 => x"84",
          4316 => x"71",
          4317 => x"82",
          4318 => x"52",
          4319 => x"51",
          4320 => x"3f",
          4321 => x"ab",
          4322 => x"3d",
          4323 => x"3d",
          4324 => x"05",
          4325 => x"52",
          4326 => x"aa",
          4327 => x"29",
          4328 => x"05",
          4329 => x"04",
          4330 => x"51",
          4331 => x"c5",
          4332 => x"39",
          4333 => x"51",
          4334 => x"c5",
          4335 => x"39",
          4336 => x"51",
          4337 => x"c6",
          4338 => x"8c",
          4339 => x"3d",
          4340 => x"88",
          4341 => x"ff",
          4342 => x"c0",
          4343 => x"08",
          4344 => x"72",
          4345 => x"07",
          4346 => x"c4",
          4347 => x"83",
          4348 => x"ff",
          4349 => x"c0",
          4350 => x"08",
          4351 => x"0c",
          4352 => x"0c",
          4353 => x"82",
          4354 => x"06",
          4355 => x"c4",
          4356 => x"51",
          4357 => x"04",
          4358 => x"c0",
          4359 => x"04",
          4360 => x"08",
          4361 => x"84",
          4362 => x"3d",
          4363 => x"2b",
          4364 => x"79",
          4365 => x"98",
          4366 => x"13",
          4367 => x"51",
          4368 => x"51",
          4369 => x"82",
          4370 => x"33",
          4371 => x"74",
          4372 => x"82",
          4373 => x"08",
          4374 => x"05",
          4375 => x"71",
          4376 => x"52",
          4377 => x"09",
          4378 => x"38",
          4379 => x"82",
          4380 => x"85",
          4381 => x"fb",
          4382 => x"02",
          4383 => x"05",
          4384 => x"55",
          4385 => x"80",
          4386 => x"82",
          4387 => x"52",
          4388 => x"aa",
          4389 => x"f4",
          4390 => x"a0",
          4391 => x"94",
          4392 => x"ac",
          4393 => x"51",
          4394 => x"3f",
          4395 => x"05",
          4396 => x"34",
          4397 => x"06",
          4398 => x"77",
          4399 => x"9a",
          4400 => x"34",
          4401 => x"04",
          4402 => x"7c",
          4403 => x"b7",
          4404 => x"88",
          4405 => x"33",
          4406 => x"33",
          4407 => x"82",
          4408 => x"70",
          4409 => x"59",
          4410 => x"74",
          4411 => x"38",
          4412 => x"fa",
          4413 => x"a0",
          4414 => x"29",
          4415 => x"05",
          4416 => x"54",
          4417 => x"9d",
          4418 => x"d8",
          4419 => x"0c",
          4420 => x"33",
          4421 => x"82",
          4422 => x"70",
          4423 => x"5a",
          4424 => x"a7",
          4425 => x"78",
          4426 => x"ff",
          4427 => x"82",
          4428 => x"81",
          4429 => x"82",
          4430 => x"74",
          4431 => x"55",
          4432 => x"87",
          4433 => x"82",
          4434 => x"77",
          4435 => x"38",
          4436 => x"08",
          4437 => x"2e",
          4438 => x"d8",
          4439 => x"74",
          4440 => x"3d",
          4441 => x"76",
          4442 => x"75",
          4443 => x"be",
          4444 => x"9c",
          4445 => x"51",
          4446 => x"3f",
          4447 => x"08",
          4448 => x"a1",
          4449 => x"0d",
          4450 => x"0d",
          4451 => x"53",
          4452 => x"08",
          4453 => x"2e",
          4454 => x"51",
          4455 => x"80",
          4456 => x"14",
          4457 => x"54",
          4458 => x"e6",
          4459 => x"82",
          4460 => x"82",
          4461 => x"52",
          4462 => x"95",
          4463 => x"80",
          4464 => x"82",
          4465 => x"51",
          4466 => x"80",
          4467 => x"9c",
          4468 => x"0d",
          4469 => x"0d",
          4470 => x"52",
          4471 => x"08",
          4472 => x"a2",
          4473 => x"c8",
          4474 => x"38",
          4475 => x"08",
          4476 => x"52",
          4477 => x"52",
          4478 => x"d2",
          4479 => x"c8",
          4480 => x"ba",
          4481 => x"ff",
          4482 => x"82",
          4483 => x"55",
          4484 => x"d8",
          4485 => x"9d",
          4486 => x"c8",
          4487 => x"70",
          4488 => x"80",
          4489 => x"53",
          4490 => x"17",
          4491 => x"52",
          4492 => x"a6",
          4493 => x"2e",
          4494 => x"ff",
          4495 => x"3d",
          4496 => x"3d",
          4497 => x"08",
          4498 => x"5a",
          4499 => x"58",
          4500 => x"82",
          4501 => x"51",
          4502 => x"3f",
          4503 => x"08",
          4504 => x"ff",
          4505 => x"9c",
          4506 => x"80",
          4507 => x"3d",
          4508 => x"81",
          4509 => x"82",
          4510 => x"80",
          4511 => x"75",
          4512 => x"83",
          4513 => x"c8",
          4514 => x"58",
          4515 => x"82",
          4516 => x"25",
          4517 => x"d8",
          4518 => x"05",
          4519 => x"55",
          4520 => x"74",
          4521 => x"70",
          4522 => x"2a",
          4523 => x"78",
          4524 => x"38",
          4525 => x"38",
          4526 => x"08",
          4527 => x"53",
          4528 => x"c2",
          4529 => x"c8",
          4530 => x"89",
          4531 => x"90",
          4532 => x"86",
          4533 => x"2e",
          4534 => x"9b",
          4535 => x"79",
          4536 => x"91",
          4537 => x"ff",
          4538 => x"ab",
          4539 => x"82",
          4540 => x"74",
          4541 => x"77",
          4542 => x"0c",
          4543 => x"04",
          4544 => x"7c",
          4545 => x"71",
          4546 => x"59",
          4547 => x"a0",
          4548 => x"06",
          4549 => x"33",
          4550 => x"77",
          4551 => x"38",
          4552 => x"5b",
          4553 => x"56",
          4554 => x"a0",
          4555 => x"06",
          4556 => x"75",
          4557 => x"80",
          4558 => x"29",
          4559 => x"05",
          4560 => x"55",
          4561 => x"3f",
          4562 => x"08",
          4563 => x"74",
          4564 => x"b0",
          4565 => x"d8",
          4566 => x"c5",
          4567 => x"33",
          4568 => x"2e",
          4569 => x"82",
          4570 => x"b5",
          4571 => x"3f",
          4572 => x"1a",
          4573 => x"fc",
          4574 => x"05",
          4575 => x"3f",
          4576 => x"08",
          4577 => x"38",
          4578 => x"78",
          4579 => x"fd",
          4580 => x"d8",
          4581 => x"ff",
          4582 => x"85",
          4583 => x"91",
          4584 => x"70",
          4585 => x"51",
          4586 => x"27",
          4587 => x"80",
          4588 => x"d8",
          4589 => x"3d",
          4590 => x"3d",
          4591 => x"08",
          4592 => x"b4",
          4593 => x"5f",
          4594 => x"af",
          4595 => x"d8",
          4596 => x"d8",
          4597 => x"5b",
          4598 => x"38",
          4599 => x"98",
          4600 => x"73",
          4601 => x"55",
          4602 => x"81",
          4603 => x"70",
          4604 => x"56",
          4605 => x"81",
          4606 => x"51",
          4607 => x"82",
          4608 => x"82",
          4609 => x"82",
          4610 => x"80",
          4611 => x"38",
          4612 => x"52",
          4613 => x"08",
          4614 => x"ad",
          4615 => x"c8",
          4616 => x"8c",
          4617 => x"bc",
          4618 => x"b9",
          4619 => x"39",
          4620 => x"08",
          4621 => x"9c",
          4622 => x"f8",
          4623 => x"70",
          4624 => x"99",
          4625 => x"d8",
          4626 => x"82",
          4627 => x"74",
          4628 => x"06",
          4629 => x"82",
          4630 => x"51",
          4631 => x"3f",
          4632 => x"08",
          4633 => x"82",
          4634 => x"25",
          4635 => x"d8",
          4636 => x"05",
          4637 => x"55",
          4638 => x"80",
          4639 => x"ff",
          4640 => x"51",
          4641 => x"81",
          4642 => x"ff",
          4643 => x"93",
          4644 => x"38",
          4645 => x"ff",
          4646 => x"06",
          4647 => x"86",
          4648 => x"d8",
          4649 => x"8c",
          4650 => x"9c",
          4651 => x"84",
          4652 => x"3f",
          4653 => x"ec",
          4654 => x"d8",
          4655 => x"2b",
          4656 => x"51",
          4657 => x"2e",
          4658 => x"81",
          4659 => x"f0",
          4660 => x"98",
          4661 => x"2c",
          4662 => x"33",
          4663 => x"70",
          4664 => x"98",
          4665 => x"84",
          4666 => x"90",
          4667 => x"15",
          4668 => x"51",
          4669 => x"59",
          4670 => x"58",
          4671 => x"78",
          4672 => x"38",
          4673 => x"b4",
          4674 => x"80",
          4675 => x"ff",
          4676 => x"98",
          4677 => x"80",
          4678 => x"ce",
          4679 => x"74",
          4680 => x"f6",
          4681 => x"d8",
          4682 => x"ff",
          4683 => x"80",
          4684 => x"74",
          4685 => x"34",
          4686 => x"39",
          4687 => x"0a",
          4688 => x"0a",
          4689 => x"2c",
          4690 => x"06",
          4691 => x"73",
          4692 => x"38",
          4693 => x"52",
          4694 => x"ce",
          4695 => x"c8",
          4696 => x"06",
          4697 => x"38",
          4698 => x"56",
          4699 => x"80",
          4700 => x"1c",
          4701 => x"f0",
          4702 => x"98",
          4703 => x"2c",
          4704 => x"33",
          4705 => x"70",
          4706 => x"10",
          4707 => x"2b",
          4708 => x"11",
          4709 => x"51",
          4710 => x"51",
          4711 => x"2e",
          4712 => x"fe",
          4713 => x"c6",
          4714 => x"7d",
          4715 => x"82",
          4716 => x"80",
          4717 => x"80",
          4718 => x"75",
          4719 => x"34",
          4720 => x"80",
          4721 => x"3d",
          4722 => x"0c",
          4723 => x"95",
          4724 => x"38",
          4725 => x"82",
          4726 => x"54",
          4727 => x"82",
          4728 => x"54",
          4729 => x"fd",
          4730 => x"f0",
          4731 => x"73",
          4732 => x"38",
          4733 => x"70",
          4734 => x"55",
          4735 => x"9e",
          4736 => x"54",
          4737 => x"15",
          4738 => x"80",
          4739 => x"ff",
          4740 => x"98",
          4741 => x"8c",
          4742 => x"55",
          4743 => x"f0",
          4744 => x"11",
          4745 => x"82",
          4746 => x"73",
          4747 => x"3d",
          4748 => x"82",
          4749 => x"54",
          4750 => x"89",
          4751 => x"54",
          4752 => x"88",
          4753 => x"8c",
          4754 => x"80",
          4755 => x"ff",
          4756 => x"98",
          4757 => x"88",
          4758 => x"56",
          4759 => x"25",
          4760 => x"f4",
          4761 => x"74",
          4762 => x"52",
          4763 => x"c4",
          4764 => x"80",
          4765 => x"80",
          4766 => x"98",
          4767 => x"88",
          4768 => x"55",
          4769 => x"da",
          4770 => x"8c",
          4771 => x"2b",
          4772 => x"82",
          4773 => x"5a",
          4774 => x"74",
          4775 => x"94",
          4776 => x"ac",
          4777 => x"51",
          4778 => x"3f",
          4779 => x"0a",
          4780 => x"0a",
          4781 => x"2c",
          4782 => x"33",
          4783 => x"73",
          4784 => x"38",
          4785 => x"83",
          4786 => x"0b",
          4787 => x"82",
          4788 => x"80",
          4789 => x"b8",
          4790 => x"3f",
          4791 => x"82",
          4792 => x"70",
          4793 => x"55",
          4794 => x"2e",
          4795 => x"82",
          4796 => x"ff",
          4797 => x"82",
          4798 => x"ff",
          4799 => x"82",
          4800 => x"82",
          4801 => x"52",
          4802 => x"9d",
          4803 => x"f0",
          4804 => x"98",
          4805 => x"2c",
          4806 => x"33",
          4807 => x"57",
          4808 => x"ad",
          4809 => x"54",
          4810 => x"74",
          4811 => x"ac",
          4812 => x"33",
          4813 => x"fc",
          4814 => x"80",
          4815 => x"80",
          4816 => x"98",
          4817 => x"88",
          4818 => x"55",
          4819 => x"d5",
          4820 => x"ac",
          4821 => x"51",
          4822 => x"3f",
          4823 => x"33",
          4824 => x"70",
          4825 => x"f0",
          4826 => x"51",
          4827 => x"74",
          4828 => x"38",
          4829 => x"08",
          4830 => x"ff",
          4831 => x"74",
          4832 => x"29",
          4833 => x"05",
          4834 => x"82",
          4835 => x"58",
          4836 => x"75",
          4837 => x"fa",
          4838 => x"f0",
          4839 => x"05",
          4840 => x"34",
          4841 => x"08",
          4842 => x"ff",
          4843 => x"82",
          4844 => x"79",
          4845 => x"3f",
          4846 => x"08",
          4847 => x"54",
          4848 => x"82",
          4849 => x"54",
          4850 => x"8f",
          4851 => x"73",
          4852 => x"f1",
          4853 => x"39",
          4854 => x"80",
          4855 => x"8c",
          4856 => x"82",
          4857 => x"79",
          4858 => x"0c",
          4859 => x"04",
          4860 => x"33",
          4861 => x"2e",
          4862 => x"82",
          4863 => x"52",
          4864 => x"9b",
          4865 => x"f0",
          4866 => x"05",
          4867 => x"f0",
          4868 => x"81",
          4869 => x"dd",
          4870 => x"8c",
          4871 => x"88",
          4872 => x"73",
          4873 => x"8c",
          4874 => x"54",
          4875 => x"88",
          4876 => x"2b",
          4877 => x"75",
          4878 => x"56",
          4879 => x"74",
          4880 => x"74",
          4881 => x"14",
          4882 => x"82",
          4883 => x"52",
          4884 => x"ff",
          4885 => x"74",
          4886 => x"29",
          4887 => x"05",
          4888 => x"82",
          4889 => x"58",
          4890 => x"75",
          4891 => x"82",
          4892 => x"52",
          4893 => x"9a",
          4894 => x"f0",
          4895 => x"98",
          4896 => x"2c",
          4897 => x"33",
          4898 => x"57",
          4899 => x"f8",
          4900 => x"f4",
          4901 => x"88",
          4902 => x"98",
          4903 => x"80",
          4904 => x"80",
          4905 => x"98",
          4906 => x"88",
          4907 => x"55",
          4908 => x"de",
          4909 => x"39",
          4910 => x"33",
          4911 => x"06",
          4912 => x"33",
          4913 => x"74",
          4914 => x"e8",
          4915 => x"ac",
          4916 => x"14",
          4917 => x"f0",
          4918 => x"1a",
          4919 => x"54",
          4920 => x"3f",
          4921 => x"33",
          4922 => x"06",
          4923 => x"33",
          4924 => x"75",
          4925 => x"38",
          4926 => x"82",
          4927 => x"80",
          4928 => x"b8",
          4929 => x"3f",
          4930 => x"f0",
          4931 => x"0b",
          4932 => x"34",
          4933 => x"7a",
          4934 => x"d8",
          4935 => x"74",
          4936 => x"38",
          4937 => x"a1",
          4938 => x"d8",
          4939 => x"f0",
          4940 => x"d8",
          4941 => x"ff",
          4942 => x"53",
          4943 => x"51",
          4944 => x"3f",
          4945 => x"c0",
          4946 => x"29",
          4947 => x"05",
          4948 => x"56",
          4949 => x"2e",
          4950 => x"51",
          4951 => x"3f",
          4952 => x"08",
          4953 => x"34",
          4954 => x"08",
          4955 => x"81",
          4956 => x"52",
          4957 => x"a2",
          4958 => x"1b",
          4959 => x"39",
          4960 => x"74",
          4961 => x"ac",
          4962 => x"ff",
          4963 => x"99",
          4964 => x"2e",
          4965 => x"ae",
          4966 => x"c8",
          4967 => x"80",
          4968 => x"74",
          4969 => x"df",
          4970 => x"c8",
          4971 => x"88",
          4972 => x"c8",
          4973 => x"06",
          4974 => x"74",
          4975 => x"ff",
          4976 => x"80",
          4977 => x"84",
          4978 => x"cc",
          4979 => x"56",
          4980 => x"2e",
          4981 => x"51",
          4982 => x"3f",
          4983 => x"08",
          4984 => x"34",
          4985 => x"08",
          4986 => x"81",
          4987 => x"52",
          4988 => x"a1",
          4989 => x"1b",
          4990 => x"ff",
          4991 => x"39",
          4992 => x"88",
          4993 => x"34",
          4994 => x"53",
          4995 => x"33",
          4996 => x"ec",
          4997 => x"9c",
          4998 => x"8c",
          4999 => x"ff",
          5000 => x"88",
          5001 => x"54",
          5002 => x"f5",
          5003 => x"f4",
          5004 => x"81",
          5005 => x"82",
          5006 => x"74",
          5007 => x"52",
          5008 => x"f0",
          5009 => x"39",
          5010 => x"33",
          5011 => x"2e",
          5012 => x"82",
          5013 => x"52",
          5014 => x"96",
          5015 => x"f0",
          5016 => x"05",
          5017 => x"f0",
          5018 => x"c8",
          5019 => x"0d",
          5020 => x"0b",
          5021 => x"0c",
          5022 => x"82",
          5023 => x"a0",
          5024 => x"52",
          5025 => x"51",
          5026 => x"3f",
          5027 => x"08",
          5028 => x"77",
          5029 => x"57",
          5030 => x"34",
          5031 => x"08",
          5032 => x"15",
          5033 => x"15",
          5034 => x"c0",
          5035 => x"86",
          5036 => x"87",
          5037 => x"d8",
          5038 => x"d8",
          5039 => x"05",
          5040 => x"07",
          5041 => x"ff",
          5042 => x"2a",
          5043 => x"56",
          5044 => x"34",
          5045 => x"34",
          5046 => x"22",
          5047 => x"82",
          5048 => x"05",
          5049 => x"55",
          5050 => x"15",
          5051 => x"15",
          5052 => x"0d",
          5053 => x"0d",
          5054 => x"51",
          5055 => x"8f",
          5056 => x"83",
          5057 => x"70",
          5058 => x"06",
          5059 => x"70",
          5060 => x"0c",
          5061 => x"04",
          5062 => x"02",
          5063 => x"02",
          5064 => x"05",
          5065 => x"82",
          5066 => x"71",
          5067 => x"11",
          5068 => x"73",
          5069 => x"81",
          5070 => x"88",
          5071 => x"a4",
          5072 => x"22",
          5073 => x"ff",
          5074 => x"88",
          5075 => x"52",
          5076 => x"5b",
          5077 => x"55",
          5078 => x"70",
          5079 => x"82",
          5080 => x"14",
          5081 => x"52",
          5082 => x"15",
          5083 => x"15",
          5084 => x"c0",
          5085 => x"70",
          5086 => x"33",
          5087 => x"07",
          5088 => x"8f",
          5089 => x"51",
          5090 => x"71",
          5091 => x"ff",
          5092 => x"88",
          5093 => x"51",
          5094 => x"34",
          5095 => x"06",
          5096 => x"12",
          5097 => x"c0",
          5098 => x"71",
          5099 => x"81",
          5100 => x"3d",
          5101 => x"3d",
          5102 => x"c0",
          5103 => x"05",
          5104 => x"70",
          5105 => x"11",
          5106 => x"87",
          5107 => x"8b",
          5108 => x"2b",
          5109 => x"59",
          5110 => x"72",
          5111 => x"33",
          5112 => x"71",
          5113 => x"70",
          5114 => x"56",
          5115 => x"84",
          5116 => x"85",
          5117 => x"d8",
          5118 => x"14",
          5119 => x"85",
          5120 => x"8b",
          5121 => x"2b",
          5122 => x"57",
          5123 => x"86",
          5124 => x"13",
          5125 => x"2b",
          5126 => x"2a",
          5127 => x"52",
          5128 => x"34",
          5129 => x"34",
          5130 => x"08",
          5131 => x"81",
          5132 => x"88",
          5133 => x"81",
          5134 => x"70",
          5135 => x"51",
          5136 => x"71",
          5137 => x"81",
          5138 => x"3d",
          5139 => x"3d",
          5140 => x"05",
          5141 => x"c0",
          5142 => x"2b",
          5143 => x"33",
          5144 => x"71",
          5145 => x"70",
          5146 => x"70",
          5147 => x"33",
          5148 => x"71",
          5149 => x"53",
          5150 => x"52",
          5151 => x"53",
          5152 => x"25",
          5153 => x"72",
          5154 => x"3f",
          5155 => x"08",
          5156 => x"33",
          5157 => x"71",
          5158 => x"83",
          5159 => x"11",
          5160 => x"12",
          5161 => x"2b",
          5162 => x"2b",
          5163 => x"06",
          5164 => x"51",
          5165 => x"53",
          5166 => x"88",
          5167 => x"72",
          5168 => x"73",
          5169 => x"82",
          5170 => x"70",
          5171 => x"81",
          5172 => x"8b",
          5173 => x"2b",
          5174 => x"57",
          5175 => x"70",
          5176 => x"33",
          5177 => x"07",
          5178 => x"ff",
          5179 => x"2a",
          5180 => x"58",
          5181 => x"34",
          5182 => x"34",
          5183 => x"04",
          5184 => x"82",
          5185 => x"02",
          5186 => x"05",
          5187 => x"2b",
          5188 => x"11",
          5189 => x"33",
          5190 => x"71",
          5191 => x"59",
          5192 => x"56",
          5193 => x"71",
          5194 => x"33",
          5195 => x"07",
          5196 => x"a2",
          5197 => x"07",
          5198 => x"53",
          5199 => x"53",
          5200 => x"70",
          5201 => x"82",
          5202 => x"70",
          5203 => x"81",
          5204 => x"8b",
          5205 => x"2b",
          5206 => x"57",
          5207 => x"82",
          5208 => x"13",
          5209 => x"2b",
          5210 => x"2a",
          5211 => x"52",
          5212 => x"34",
          5213 => x"34",
          5214 => x"08",
          5215 => x"33",
          5216 => x"71",
          5217 => x"82",
          5218 => x"52",
          5219 => x"0d",
          5220 => x"0d",
          5221 => x"c0",
          5222 => x"2a",
          5223 => x"ff",
          5224 => x"57",
          5225 => x"3f",
          5226 => x"08",
          5227 => x"71",
          5228 => x"33",
          5229 => x"71",
          5230 => x"83",
          5231 => x"11",
          5232 => x"12",
          5233 => x"2b",
          5234 => x"07",
          5235 => x"51",
          5236 => x"55",
          5237 => x"80",
          5238 => x"82",
          5239 => x"75",
          5240 => x"3f",
          5241 => x"84",
          5242 => x"15",
          5243 => x"2b",
          5244 => x"07",
          5245 => x"88",
          5246 => x"55",
          5247 => x"86",
          5248 => x"81",
          5249 => x"75",
          5250 => x"82",
          5251 => x"70",
          5252 => x"33",
          5253 => x"71",
          5254 => x"70",
          5255 => x"57",
          5256 => x"72",
          5257 => x"73",
          5258 => x"82",
          5259 => x"18",
          5260 => x"86",
          5261 => x"0b",
          5262 => x"82",
          5263 => x"53",
          5264 => x"34",
          5265 => x"34",
          5266 => x"08",
          5267 => x"81",
          5268 => x"88",
          5269 => x"82",
          5270 => x"70",
          5271 => x"51",
          5272 => x"74",
          5273 => x"81",
          5274 => x"3d",
          5275 => x"3d",
          5276 => x"82",
          5277 => x"84",
          5278 => x"3f",
          5279 => x"86",
          5280 => x"fe",
          5281 => x"3d",
          5282 => x"3d",
          5283 => x"52",
          5284 => x"3f",
          5285 => x"08",
          5286 => x"06",
          5287 => x"08",
          5288 => x"85",
          5289 => x"88",
          5290 => x"5f",
          5291 => x"5a",
          5292 => x"59",
          5293 => x"80",
          5294 => x"88",
          5295 => x"33",
          5296 => x"71",
          5297 => x"70",
          5298 => x"06",
          5299 => x"83",
          5300 => x"70",
          5301 => x"53",
          5302 => x"55",
          5303 => x"8a",
          5304 => x"2e",
          5305 => x"78",
          5306 => x"15",
          5307 => x"33",
          5308 => x"07",
          5309 => x"c2",
          5310 => x"ff",
          5311 => x"38",
          5312 => x"56",
          5313 => x"2b",
          5314 => x"08",
          5315 => x"81",
          5316 => x"88",
          5317 => x"81",
          5318 => x"51",
          5319 => x"5c",
          5320 => x"2e",
          5321 => x"55",
          5322 => x"78",
          5323 => x"38",
          5324 => x"80",
          5325 => x"38",
          5326 => x"09",
          5327 => x"38",
          5328 => x"f2",
          5329 => x"39",
          5330 => x"53",
          5331 => x"51",
          5332 => x"82",
          5333 => x"70",
          5334 => x"33",
          5335 => x"71",
          5336 => x"83",
          5337 => x"5a",
          5338 => x"05",
          5339 => x"83",
          5340 => x"70",
          5341 => x"59",
          5342 => x"84",
          5343 => x"81",
          5344 => x"76",
          5345 => x"82",
          5346 => x"75",
          5347 => x"11",
          5348 => x"11",
          5349 => x"33",
          5350 => x"07",
          5351 => x"53",
          5352 => x"5a",
          5353 => x"86",
          5354 => x"87",
          5355 => x"d8",
          5356 => x"1c",
          5357 => x"85",
          5358 => x"8b",
          5359 => x"2b",
          5360 => x"5a",
          5361 => x"54",
          5362 => x"34",
          5363 => x"34",
          5364 => x"08",
          5365 => x"1d",
          5366 => x"85",
          5367 => x"88",
          5368 => x"88",
          5369 => x"5f",
          5370 => x"73",
          5371 => x"75",
          5372 => x"82",
          5373 => x"1b",
          5374 => x"73",
          5375 => x"0c",
          5376 => x"04",
          5377 => x"74",
          5378 => x"c0",
          5379 => x"f4",
          5380 => x"53",
          5381 => x"8b",
          5382 => x"fc",
          5383 => x"d8",
          5384 => x"72",
          5385 => x"0c",
          5386 => x"04",
          5387 => x"64",
          5388 => x"80",
          5389 => x"82",
          5390 => x"60",
          5391 => x"06",
          5392 => x"a9",
          5393 => x"38",
          5394 => x"b8",
          5395 => x"c8",
          5396 => x"c7",
          5397 => x"38",
          5398 => x"92",
          5399 => x"83",
          5400 => x"51",
          5401 => x"82",
          5402 => x"83",
          5403 => x"82",
          5404 => x"7d",
          5405 => x"2a",
          5406 => x"ff",
          5407 => x"2b",
          5408 => x"33",
          5409 => x"71",
          5410 => x"70",
          5411 => x"83",
          5412 => x"70",
          5413 => x"05",
          5414 => x"1a",
          5415 => x"12",
          5416 => x"2b",
          5417 => x"2b",
          5418 => x"53",
          5419 => x"5c",
          5420 => x"5c",
          5421 => x"73",
          5422 => x"38",
          5423 => x"ff",
          5424 => x"70",
          5425 => x"06",
          5426 => x"16",
          5427 => x"33",
          5428 => x"07",
          5429 => x"1c",
          5430 => x"12",
          5431 => x"2b",
          5432 => x"07",
          5433 => x"52",
          5434 => x"80",
          5435 => x"78",
          5436 => x"83",
          5437 => x"41",
          5438 => x"27",
          5439 => x"60",
          5440 => x"7b",
          5441 => x"06",
          5442 => x"51",
          5443 => x"7a",
          5444 => x"06",
          5445 => x"39",
          5446 => x"7a",
          5447 => x"38",
          5448 => x"aa",
          5449 => x"39",
          5450 => x"7a",
          5451 => x"c8",
          5452 => x"82",
          5453 => x"12",
          5454 => x"2b",
          5455 => x"54",
          5456 => x"80",
          5457 => x"f7",
          5458 => x"d8",
          5459 => x"ff",
          5460 => x"54",
          5461 => x"83",
          5462 => x"c0",
          5463 => x"05",
          5464 => x"ff",
          5465 => x"82",
          5466 => x"14",
          5467 => x"83",
          5468 => x"59",
          5469 => x"39",
          5470 => x"7a",
          5471 => x"d4",
          5472 => x"f5",
          5473 => x"d8",
          5474 => x"82",
          5475 => x"12",
          5476 => x"2b",
          5477 => x"54",
          5478 => x"80",
          5479 => x"f6",
          5480 => x"d8",
          5481 => x"ff",
          5482 => x"54",
          5483 => x"83",
          5484 => x"c0",
          5485 => x"05",
          5486 => x"ff",
          5487 => x"82",
          5488 => x"14",
          5489 => x"62",
          5490 => x"5c",
          5491 => x"ff",
          5492 => x"39",
          5493 => x"54",
          5494 => x"82",
          5495 => x"5c",
          5496 => x"08",
          5497 => x"38",
          5498 => x"52",
          5499 => x"08",
          5500 => x"f3",
          5501 => x"f7",
          5502 => x"58",
          5503 => x"99",
          5504 => x"7a",
          5505 => x"f2",
          5506 => x"19",
          5507 => x"d8",
          5508 => x"84",
          5509 => x"f9",
          5510 => x"73",
          5511 => x"0c",
          5512 => x"04",
          5513 => x"77",
          5514 => x"52",
          5515 => x"3f",
          5516 => x"08",
          5517 => x"c8",
          5518 => x"8e",
          5519 => x"80",
          5520 => x"c8",
          5521 => x"96",
          5522 => x"82",
          5523 => x"86",
          5524 => x"ff",
          5525 => x"8f",
          5526 => x"81",
          5527 => x"26",
          5528 => x"d8",
          5529 => x"52",
          5530 => x"c8",
          5531 => x"0d",
          5532 => x"0d",
          5533 => x"33",
          5534 => x"9f",
          5535 => x"53",
          5536 => x"81",
          5537 => x"38",
          5538 => x"87",
          5539 => x"11",
          5540 => x"54",
          5541 => x"84",
          5542 => x"54",
          5543 => x"87",
          5544 => x"11",
          5545 => x"0c",
          5546 => x"c0",
          5547 => x"70",
          5548 => x"70",
          5549 => x"51",
          5550 => x"8a",
          5551 => x"98",
          5552 => x"70",
          5553 => x"08",
          5554 => x"06",
          5555 => x"38",
          5556 => x"8c",
          5557 => x"80",
          5558 => x"71",
          5559 => x"14",
          5560 => x"c4",
          5561 => x"70",
          5562 => x"0c",
          5563 => x"04",
          5564 => x"60",
          5565 => x"8c",
          5566 => x"33",
          5567 => x"5b",
          5568 => x"5a",
          5569 => x"82",
          5570 => x"81",
          5571 => x"52",
          5572 => x"38",
          5573 => x"84",
          5574 => x"92",
          5575 => x"c0",
          5576 => x"87",
          5577 => x"13",
          5578 => x"57",
          5579 => x"0b",
          5580 => x"8c",
          5581 => x"0c",
          5582 => x"75",
          5583 => x"2a",
          5584 => x"51",
          5585 => x"80",
          5586 => x"7b",
          5587 => x"7b",
          5588 => x"5d",
          5589 => x"59",
          5590 => x"06",
          5591 => x"73",
          5592 => x"81",
          5593 => x"ff",
          5594 => x"72",
          5595 => x"38",
          5596 => x"8c",
          5597 => x"c3",
          5598 => x"98",
          5599 => x"71",
          5600 => x"38",
          5601 => x"2e",
          5602 => x"76",
          5603 => x"92",
          5604 => x"72",
          5605 => x"06",
          5606 => x"f7",
          5607 => x"5a",
          5608 => x"80",
          5609 => x"70",
          5610 => x"5a",
          5611 => x"80",
          5612 => x"73",
          5613 => x"06",
          5614 => x"38",
          5615 => x"fe",
          5616 => x"fc",
          5617 => x"52",
          5618 => x"83",
          5619 => x"71",
          5620 => x"d8",
          5621 => x"3d",
          5622 => x"3d",
          5623 => x"64",
          5624 => x"bf",
          5625 => x"40",
          5626 => x"59",
          5627 => x"58",
          5628 => x"82",
          5629 => x"81",
          5630 => x"52",
          5631 => x"09",
          5632 => x"b1",
          5633 => x"84",
          5634 => x"92",
          5635 => x"c0",
          5636 => x"87",
          5637 => x"13",
          5638 => x"56",
          5639 => x"87",
          5640 => x"0c",
          5641 => x"82",
          5642 => x"58",
          5643 => x"84",
          5644 => x"06",
          5645 => x"71",
          5646 => x"38",
          5647 => x"05",
          5648 => x"0c",
          5649 => x"73",
          5650 => x"81",
          5651 => x"71",
          5652 => x"38",
          5653 => x"8c",
          5654 => x"d0",
          5655 => x"98",
          5656 => x"71",
          5657 => x"38",
          5658 => x"2e",
          5659 => x"76",
          5660 => x"92",
          5661 => x"72",
          5662 => x"06",
          5663 => x"f7",
          5664 => x"59",
          5665 => x"1a",
          5666 => x"06",
          5667 => x"59",
          5668 => x"80",
          5669 => x"73",
          5670 => x"06",
          5671 => x"38",
          5672 => x"fe",
          5673 => x"fc",
          5674 => x"52",
          5675 => x"83",
          5676 => x"71",
          5677 => x"d8",
          5678 => x"3d",
          5679 => x"3d",
          5680 => x"84",
          5681 => x"33",
          5682 => x"a7",
          5683 => x"54",
          5684 => x"fa",
          5685 => x"d8",
          5686 => x"06",
          5687 => x"72",
          5688 => x"85",
          5689 => x"98",
          5690 => x"56",
          5691 => x"80",
          5692 => x"76",
          5693 => x"74",
          5694 => x"c0",
          5695 => x"54",
          5696 => x"2e",
          5697 => x"d4",
          5698 => x"2e",
          5699 => x"80",
          5700 => x"08",
          5701 => x"70",
          5702 => x"51",
          5703 => x"2e",
          5704 => x"c0",
          5705 => x"52",
          5706 => x"87",
          5707 => x"08",
          5708 => x"38",
          5709 => x"87",
          5710 => x"14",
          5711 => x"70",
          5712 => x"52",
          5713 => x"96",
          5714 => x"92",
          5715 => x"0a",
          5716 => x"39",
          5717 => x"0c",
          5718 => x"39",
          5719 => x"54",
          5720 => x"c8",
          5721 => x"0d",
          5722 => x"0d",
          5723 => x"33",
          5724 => x"88",
          5725 => x"d8",
          5726 => x"51",
          5727 => x"04",
          5728 => x"75",
          5729 => x"82",
          5730 => x"90",
          5731 => x"2b",
          5732 => x"33",
          5733 => x"88",
          5734 => x"71",
          5735 => x"c8",
          5736 => x"54",
          5737 => x"85",
          5738 => x"ff",
          5739 => x"02",
          5740 => x"05",
          5741 => x"70",
          5742 => x"05",
          5743 => x"88",
          5744 => x"72",
          5745 => x"0d",
          5746 => x"0d",
          5747 => x"52",
          5748 => x"81",
          5749 => x"70",
          5750 => x"70",
          5751 => x"05",
          5752 => x"88",
          5753 => x"72",
          5754 => x"54",
          5755 => x"2a",
          5756 => x"34",
          5757 => x"04",
          5758 => x"76",
          5759 => x"54",
          5760 => x"2e",
          5761 => x"70",
          5762 => x"33",
          5763 => x"05",
          5764 => x"11",
          5765 => x"84",
          5766 => x"fe",
          5767 => x"77",
          5768 => x"53",
          5769 => x"81",
          5770 => x"ff",
          5771 => x"f4",
          5772 => x"0d",
          5773 => x"0d",
          5774 => x"56",
          5775 => x"70",
          5776 => x"33",
          5777 => x"05",
          5778 => x"71",
          5779 => x"56",
          5780 => x"72",
          5781 => x"38",
          5782 => x"e2",
          5783 => x"d8",
          5784 => x"3d",
          5785 => x"3d",
          5786 => x"54",
          5787 => x"71",
          5788 => x"38",
          5789 => x"70",
          5790 => x"f3",
          5791 => x"82",
          5792 => x"84",
          5793 => x"80",
          5794 => x"c8",
          5795 => x"3d",
          5796 => x"08",
          5797 => x"05",
          5798 => x"54",
          5799 => x"e7",
          5800 => x"82",
          5801 => x"a2",
          5802 => x"2e",
          5803 => x"b5",
          5804 => x"80",
          5805 => x"82",
          5806 => x"83",
          5807 => x"53",
          5808 => x"86",
          5809 => x"0c",
          5810 => x"82",
          5811 => x"87",
          5812 => x"f7",
          5813 => x"56",
          5814 => x"17",
          5815 => x"74",
          5816 => x"d6",
          5817 => x"b4",
          5818 => x"b8",
          5819 => x"81",
          5820 => x"59",
          5821 => x"82",
          5822 => x"7a",
          5823 => x"06",
          5824 => x"d8",
          5825 => x"17",
          5826 => x"08",
          5827 => x"08",
          5828 => x"08",
          5829 => x"74",
          5830 => x"38",
          5831 => x"55",
          5832 => x"09",
          5833 => x"38",
          5834 => x"18",
          5835 => x"81",
          5836 => x"f9",
          5837 => x"39",
          5838 => x"82",
          5839 => x"8b",
          5840 => x"fa",
          5841 => x"7a",
          5842 => x"57",
          5843 => x"08",
          5844 => x"75",
          5845 => x"3f",
          5846 => x"08",
          5847 => x"c8",
          5848 => x"81",
          5849 => x"b8",
          5850 => x"16",
          5851 => x"80",
          5852 => x"c8",
          5853 => x"85",
          5854 => x"81",
          5855 => x"17",
          5856 => x"d8",
          5857 => x"3d",
          5858 => x"3d",
          5859 => x"52",
          5860 => x"3f",
          5861 => x"08",
          5862 => x"c8",
          5863 => x"38",
          5864 => x"74",
          5865 => x"81",
          5866 => x"38",
          5867 => x"59",
          5868 => x"09",
          5869 => x"e3",
          5870 => x"53",
          5871 => x"08",
          5872 => x"70",
          5873 => x"d3",
          5874 => x"d5",
          5875 => x"17",
          5876 => x"3f",
          5877 => x"a4",
          5878 => x"51",
          5879 => x"86",
          5880 => x"f2",
          5881 => x"17",
          5882 => x"3f",
          5883 => x"52",
          5884 => x"51",
          5885 => x"90",
          5886 => x"84",
          5887 => x"fb",
          5888 => x"17",
          5889 => x"70",
          5890 => x"79",
          5891 => x"52",
          5892 => x"51",
          5893 => x"77",
          5894 => x"80",
          5895 => x"81",
          5896 => x"f9",
          5897 => x"d8",
          5898 => x"2e",
          5899 => x"58",
          5900 => x"c8",
          5901 => x"0d",
          5902 => x"0d",
          5903 => x"9c",
          5904 => x"05",
          5905 => x"80",
          5906 => x"27",
          5907 => x"14",
          5908 => x"29",
          5909 => x"05",
          5910 => x"82",
          5911 => x"87",
          5912 => x"f9",
          5913 => x"7a",
          5914 => x"54",
          5915 => x"27",
          5916 => x"76",
          5917 => x"27",
          5918 => x"ff",
          5919 => x"58",
          5920 => x"80",
          5921 => x"82",
          5922 => x"72",
          5923 => x"38",
          5924 => x"72",
          5925 => x"8e",
          5926 => x"39",
          5927 => x"17",
          5928 => x"a8",
          5929 => x"53",
          5930 => x"fd",
          5931 => x"d8",
          5932 => x"9f",
          5933 => x"ff",
          5934 => x"11",
          5935 => x"70",
          5936 => x"18",
          5937 => x"76",
          5938 => x"53",
          5939 => x"82",
          5940 => x"80",
          5941 => x"83",
          5942 => x"b8",
          5943 => x"88",
          5944 => x"79",
          5945 => x"84",
          5946 => x"58",
          5947 => x"80",
          5948 => x"9f",
          5949 => x"80",
          5950 => x"88",
          5951 => x"08",
          5952 => x"51",
          5953 => x"82",
          5954 => x"80",
          5955 => x"10",
          5956 => x"74",
          5957 => x"51",
          5958 => x"82",
          5959 => x"83",
          5960 => x"58",
          5961 => x"87",
          5962 => x"08",
          5963 => x"51",
          5964 => x"82",
          5965 => x"9b",
          5966 => x"2b",
          5967 => x"74",
          5968 => x"51",
          5969 => x"82",
          5970 => x"f0",
          5971 => x"83",
          5972 => x"77",
          5973 => x"0c",
          5974 => x"04",
          5975 => x"7a",
          5976 => x"58",
          5977 => x"81",
          5978 => x"9e",
          5979 => x"17",
          5980 => x"96",
          5981 => x"53",
          5982 => x"81",
          5983 => x"79",
          5984 => x"72",
          5985 => x"38",
          5986 => x"72",
          5987 => x"b8",
          5988 => x"39",
          5989 => x"17",
          5990 => x"a8",
          5991 => x"53",
          5992 => x"fb",
          5993 => x"d8",
          5994 => x"82",
          5995 => x"81",
          5996 => x"83",
          5997 => x"b8",
          5998 => x"78",
          5999 => x"56",
          6000 => x"76",
          6001 => x"38",
          6002 => x"9f",
          6003 => x"33",
          6004 => x"07",
          6005 => x"74",
          6006 => x"83",
          6007 => x"89",
          6008 => x"08",
          6009 => x"51",
          6010 => x"82",
          6011 => x"59",
          6012 => x"08",
          6013 => x"74",
          6014 => x"16",
          6015 => x"84",
          6016 => x"76",
          6017 => x"88",
          6018 => x"81",
          6019 => x"8f",
          6020 => x"53",
          6021 => x"80",
          6022 => x"88",
          6023 => x"08",
          6024 => x"51",
          6025 => x"82",
          6026 => x"59",
          6027 => x"08",
          6028 => x"77",
          6029 => x"06",
          6030 => x"83",
          6031 => x"05",
          6032 => x"f6",
          6033 => x"39",
          6034 => x"a8",
          6035 => x"52",
          6036 => x"ef",
          6037 => x"c8",
          6038 => x"d8",
          6039 => x"38",
          6040 => x"06",
          6041 => x"83",
          6042 => x"18",
          6043 => x"54",
          6044 => x"f6",
          6045 => x"d8",
          6046 => x"0a",
          6047 => x"52",
          6048 => x"c5",
          6049 => x"83",
          6050 => x"82",
          6051 => x"8a",
          6052 => x"f8",
          6053 => x"7c",
          6054 => x"59",
          6055 => x"81",
          6056 => x"38",
          6057 => x"08",
          6058 => x"73",
          6059 => x"38",
          6060 => x"52",
          6061 => x"a4",
          6062 => x"c8",
          6063 => x"d8",
          6064 => x"f2",
          6065 => x"82",
          6066 => x"39",
          6067 => x"e6",
          6068 => x"c8",
          6069 => x"de",
          6070 => x"78",
          6071 => x"3f",
          6072 => x"08",
          6073 => x"c8",
          6074 => x"80",
          6075 => x"d8",
          6076 => x"2e",
          6077 => x"d8",
          6078 => x"2e",
          6079 => x"53",
          6080 => x"51",
          6081 => x"82",
          6082 => x"c5",
          6083 => x"08",
          6084 => x"18",
          6085 => x"57",
          6086 => x"90",
          6087 => x"94",
          6088 => x"16",
          6089 => x"54",
          6090 => x"34",
          6091 => x"78",
          6092 => x"38",
          6093 => x"82",
          6094 => x"8a",
          6095 => x"f6",
          6096 => x"7e",
          6097 => x"5b",
          6098 => x"38",
          6099 => x"58",
          6100 => x"88",
          6101 => x"08",
          6102 => x"38",
          6103 => x"39",
          6104 => x"51",
          6105 => x"81",
          6106 => x"d8",
          6107 => x"82",
          6108 => x"d8",
          6109 => x"82",
          6110 => x"ff",
          6111 => x"38",
          6112 => x"82",
          6113 => x"26",
          6114 => x"79",
          6115 => x"08",
          6116 => x"73",
          6117 => x"b9",
          6118 => x"2e",
          6119 => x"80",
          6120 => x"1a",
          6121 => x"08",
          6122 => x"38",
          6123 => x"52",
          6124 => x"af",
          6125 => x"82",
          6126 => x"81",
          6127 => x"06",
          6128 => x"d8",
          6129 => x"82",
          6130 => x"09",
          6131 => x"72",
          6132 => x"70",
          6133 => x"d8",
          6134 => x"51",
          6135 => x"73",
          6136 => x"82",
          6137 => x"80",
          6138 => x"90",
          6139 => x"81",
          6140 => x"38",
          6141 => x"08",
          6142 => x"73",
          6143 => x"75",
          6144 => x"77",
          6145 => x"56",
          6146 => x"76",
          6147 => x"82",
          6148 => x"26",
          6149 => x"75",
          6150 => x"f8",
          6151 => x"d8",
          6152 => x"2e",
          6153 => x"59",
          6154 => x"08",
          6155 => x"81",
          6156 => x"82",
          6157 => x"59",
          6158 => x"08",
          6159 => x"70",
          6160 => x"25",
          6161 => x"51",
          6162 => x"73",
          6163 => x"75",
          6164 => x"81",
          6165 => x"38",
          6166 => x"f5",
          6167 => x"75",
          6168 => x"f9",
          6169 => x"d8",
          6170 => x"d8",
          6171 => x"70",
          6172 => x"08",
          6173 => x"51",
          6174 => x"80",
          6175 => x"73",
          6176 => x"38",
          6177 => x"52",
          6178 => x"d0",
          6179 => x"c8",
          6180 => x"a5",
          6181 => x"18",
          6182 => x"08",
          6183 => x"18",
          6184 => x"74",
          6185 => x"38",
          6186 => x"18",
          6187 => x"33",
          6188 => x"73",
          6189 => x"97",
          6190 => x"74",
          6191 => x"38",
          6192 => x"55",
          6193 => x"d8",
          6194 => x"85",
          6195 => x"75",
          6196 => x"d8",
          6197 => x"3d",
          6198 => x"3d",
          6199 => x"52",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"82",
          6203 => x"80",
          6204 => x"52",
          6205 => x"c1",
          6206 => x"c8",
          6207 => x"c8",
          6208 => x"0c",
          6209 => x"53",
          6210 => x"15",
          6211 => x"f2",
          6212 => x"56",
          6213 => x"16",
          6214 => x"22",
          6215 => x"27",
          6216 => x"54",
          6217 => x"76",
          6218 => x"33",
          6219 => x"3f",
          6220 => x"08",
          6221 => x"38",
          6222 => x"76",
          6223 => x"70",
          6224 => x"9f",
          6225 => x"56",
          6226 => x"d8",
          6227 => x"3d",
          6228 => x"3d",
          6229 => x"71",
          6230 => x"57",
          6231 => x"0a",
          6232 => x"38",
          6233 => x"53",
          6234 => x"38",
          6235 => x"0c",
          6236 => x"54",
          6237 => x"75",
          6238 => x"73",
          6239 => x"ac",
          6240 => x"73",
          6241 => x"85",
          6242 => x"0b",
          6243 => x"5a",
          6244 => x"27",
          6245 => x"ac",
          6246 => x"18",
          6247 => x"39",
          6248 => x"70",
          6249 => x"58",
          6250 => x"b2",
          6251 => x"76",
          6252 => x"3f",
          6253 => x"08",
          6254 => x"c8",
          6255 => x"bd",
          6256 => x"82",
          6257 => x"27",
          6258 => x"16",
          6259 => x"c8",
          6260 => x"38",
          6261 => x"39",
          6262 => x"55",
          6263 => x"52",
          6264 => x"d5",
          6265 => x"c8",
          6266 => x"0c",
          6267 => x"0c",
          6268 => x"53",
          6269 => x"80",
          6270 => x"85",
          6271 => x"94",
          6272 => x"2a",
          6273 => x"0c",
          6274 => x"06",
          6275 => x"9c",
          6276 => x"58",
          6277 => x"c8",
          6278 => x"0d",
          6279 => x"0d",
          6280 => x"90",
          6281 => x"05",
          6282 => x"f0",
          6283 => x"27",
          6284 => x"0b",
          6285 => x"98",
          6286 => x"84",
          6287 => x"2e",
          6288 => x"76",
          6289 => x"58",
          6290 => x"38",
          6291 => x"15",
          6292 => x"08",
          6293 => x"38",
          6294 => x"88",
          6295 => x"53",
          6296 => x"81",
          6297 => x"c0",
          6298 => x"22",
          6299 => x"89",
          6300 => x"72",
          6301 => x"74",
          6302 => x"f3",
          6303 => x"d8",
          6304 => x"82",
          6305 => x"82",
          6306 => x"27",
          6307 => x"81",
          6308 => x"c8",
          6309 => x"80",
          6310 => x"16",
          6311 => x"c8",
          6312 => x"ca",
          6313 => x"38",
          6314 => x"0c",
          6315 => x"dd",
          6316 => x"08",
          6317 => x"f9",
          6318 => x"d8",
          6319 => x"87",
          6320 => x"c8",
          6321 => x"80",
          6322 => x"55",
          6323 => x"08",
          6324 => x"38",
          6325 => x"d8",
          6326 => x"2e",
          6327 => x"d8",
          6328 => x"75",
          6329 => x"3f",
          6330 => x"08",
          6331 => x"94",
          6332 => x"52",
          6333 => x"c1",
          6334 => x"c8",
          6335 => x"0c",
          6336 => x"0c",
          6337 => x"05",
          6338 => x"80",
          6339 => x"d8",
          6340 => x"3d",
          6341 => x"3d",
          6342 => x"71",
          6343 => x"57",
          6344 => x"51",
          6345 => x"82",
          6346 => x"54",
          6347 => x"08",
          6348 => x"82",
          6349 => x"56",
          6350 => x"52",
          6351 => x"83",
          6352 => x"c8",
          6353 => x"d8",
          6354 => x"d2",
          6355 => x"c8",
          6356 => x"08",
          6357 => x"54",
          6358 => x"e5",
          6359 => x"06",
          6360 => x"58",
          6361 => x"08",
          6362 => x"38",
          6363 => x"75",
          6364 => x"80",
          6365 => x"81",
          6366 => x"7a",
          6367 => x"06",
          6368 => x"39",
          6369 => x"08",
          6370 => x"76",
          6371 => x"3f",
          6372 => x"08",
          6373 => x"c8",
          6374 => x"ff",
          6375 => x"84",
          6376 => x"06",
          6377 => x"54",
          6378 => x"c8",
          6379 => x"0d",
          6380 => x"0d",
          6381 => x"52",
          6382 => x"3f",
          6383 => x"08",
          6384 => x"06",
          6385 => x"51",
          6386 => x"83",
          6387 => x"06",
          6388 => x"14",
          6389 => x"3f",
          6390 => x"08",
          6391 => x"07",
          6392 => x"d8",
          6393 => x"3d",
          6394 => x"3d",
          6395 => x"70",
          6396 => x"06",
          6397 => x"53",
          6398 => x"af",
          6399 => x"33",
          6400 => x"83",
          6401 => x"06",
          6402 => x"90",
          6403 => x"15",
          6404 => x"3f",
          6405 => x"04",
          6406 => x"75",
          6407 => x"8b",
          6408 => x"2a",
          6409 => x"29",
          6410 => x"81",
          6411 => x"71",
          6412 => x"ff",
          6413 => x"56",
          6414 => x"72",
          6415 => x"82",
          6416 => x"85",
          6417 => x"f2",
          6418 => x"62",
          6419 => x"79",
          6420 => x"81",
          6421 => x"5d",
          6422 => x"80",
          6423 => x"38",
          6424 => x"52",
          6425 => x"db",
          6426 => x"c8",
          6427 => x"d8",
          6428 => x"eb",
          6429 => x"08",
          6430 => x"55",
          6431 => x"84",
          6432 => x"39",
          6433 => x"bf",
          6434 => x"ff",
          6435 => x"72",
          6436 => x"82",
          6437 => x"56",
          6438 => x"2e",
          6439 => x"83",
          6440 => x"82",
          6441 => x"53",
          6442 => x"09",
          6443 => x"38",
          6444 => x"73",
          6445 => x"99",
          6446 => x"c8",
          6447 => x"06",
          6448 => x"88",
          6449 => x"06",
          6450 => x"56",
          6451 => x"87",
          6452 => x"5c",
          6453 => x"76",
          6454 => x"81",
          6455 => x"38",
          6456 => x"70",
          6457 => x"53",
          6458 => x"92",
          6459 => x"33",
          6460 => x"06",
          6461 => x"08",
          6462 => x"56",
          6463 => x"7c",
          6464 => x"06",
          6465 => x"8d",
          6466 => x"7c",
          6467 => x"81",
          6468 => x"38",
          6469 => x"9a",
          6470 => x"e8",
          6471 => x"d8",
          6472 => x"ff",
          6473 => x"72",
          6474 => x"74",
          6475 => x"bf",
          6476 => x"f3",
          6477 => x"81",
          6478 => x"82",
          6479 => x"33",
          6480 => x"e8",
          6481 => x"d8",
          6482 => x"ff",
          6483 => x"77",
          6484 => x"38",
          6485 => x"26",
          6486 => x"73",
          6487 => x"59",
          6488 => x"23",
          6489 => x"8b",
          6490 => x"ff",
          6491 => x"81",
          6492 => x"81",
          6493 => x"77",
          6494 => x"74",
          6495 => x"2a",
          6496 => x"51",
          6497 => x"80",
          6498 => x"73",
          6499 => x"92",
          6500 => x"1a",
          6501 => x"23",
          6502 => x"81",
          6503 => x"53",
          6504 => x"ff",
          6505 => x"9d",
          6506 => x"38",
          6507 => x"e8",
          6508 => x"c8",
          6509 => x"06",
          6510 => x"2e",
          6511 => x"0b",
          6512 => x"a0",
          6513 => x"78",
          6514 => x"3f",
          6515 => x"08",
          6516 => x"c8",
          6517 => x"98",
          6518 => x"84",
          6519 => x"80",
          6520 => x"0c",
          6521 => x"c8",
          6522 => x"0d",
          6523 => x"0d",
          6524 => x"40",
          6525 => x"78",
          6526 => x"3f",
          6527 => x"08",
          6528 => x"c8",
          6529 => x"38",
          6530 => x"5f",
          6531 => x"ac",
          6532 => x"19",
          6533 => x"51",
          6534 => x"82",
          6535 => x"58",
          6536 => x"08",
          6537 => x"9c",
          6538 => x"33",
          6539 => x"86",
          6540 => x"82",
          6541 => x"17",
          6542 => x"70",
          6543 => x"56",
          6544 => x"1a",
          6545 => x"e5",
          6546 => x"38",
          6547 => x"70",
          6548 => x"54",
          6549 => x"8e",
          6550 => x"b2",
          6551 => x"2e",
          6552 => x"81",
          6553 => x"19",
          6554 => x"2a",
          6555 => x"51",
          6556 => x"82",
          6557 => x"86",
          6558 => x"06",
          6559 => x"80",
          6560 => x"8d",
          6561 => x"81",
          6562 => x"90",
          6563 => x"1d",
          6564 => x"5e",
          6565 => x"09",
          6566 => x"b9",
          6567 => x"33",
          6568 => x"2e",
          6569 => x"81",
          6570 => x"1f",
          6571 => x"52",
          6572 => x"3f",
          6573 => x"08",
          6574 => x"06",
          6575 => x"95",
          6576 => x"70",
          6577 => x"29",
          6578 => x"56",
          6579 => x"5a",
          6580 => x"1b",
          6581 => x"51",
          6582 => x"82",
          6583 => x"83",
          6584 => x"56",
          6585 => x"b1",
          6586 => x"fe",
          6587 => x"38",
          6588 => x"df",
          6589 => x"d8",
          6590 => x"10",
          6591 => x"53",
          6592 => x"59",
          6593 => x"a1",
          6594 => x"d8",
          6595 => x"09",
          6596 => x"c1",
          6597 => x"8b",
          6598 => x"ff",
          6599 => x"81",
          6600 => x"81",
          6601 => x"7b",
          6602 => x"38",
          6603 => x"86",
          6604 => x"06",
          6605 => x"79",
          6606 => x"38",
          6607 => x"8b",
          6608 => x"1d",
          6609 => x"54",
          6610 => x"ff",
          6611 => x"ff",
          6612 => x"84",
          6613 => x"54",
          6614 => x"39",
          6615 => x"76",
          6616 => x"3f",
          6617 => x"08",
          6618 => x"54",
          6619 => x"bb",
          6620 => x"33",
          6621 => x"73",
          6622 => x"53",
          6623 => x"9c",
          6624 => x"e5",
          6625 => x"d8",
          6626 => x"2e",
          6627 => x"ff",
          6628 => x"ac",
          6629 => x"52",
          6630 => x"81",
          6631 => x"c8",
          6632 => x"d8",
          6633 => x"2e",
          6634 => x"77",
          6635 => x"0c",
          6636 => x"04",
          6637 => x"64",
          6638 => x"12",
          6639 => x"06",
          6640 => x"86",
          6641 => x"b5",
          6642 => x"1d",
          6643 => x"56",
          6644 => x"80",
          6645 => x"81",
          6646 => x"16",
          6647 => x"55",
          6648 => x"8c",
          6649 => x"70",
          6650 => x"70",
          6651 => x"e4",
          6652 => x"80",
          6653 => x"81",
          6654 => x"80",
          6655 => x"38",
          6656 => x"ab",
          6657 => x"5b",
          6658 => x"7b",
          6659 => x"53",
          6660 => x"51",
          6661 => x"85",
          6662 => x"c6",
          6663 => x"77",
          6664 => x"ff",
          6665 => x"55",
          6666 => x"b4",
          6667 => x"ff",
          6668 => x"19",
          6669 => x"57",
          6670 => x"76",
          6671 => x"81",
          6672 => x"2a",
          6673 => x"51",
          6674 => x"73",
          6675 => x"38",
          6676 => x"a1",
          6677 => x"17",
          6678 => x"25",
          6679 => x"39",
          6680 => x"02",
          6681 => x"05",
          6682 => x"b0",
          6683 => x"54",
          6684 => x"84",
          6685 => x"54",
          6686 => x"ff",
          6687 => x"76",
          6688 => x"58",
          6689 => x"38",
          6690 => x"05",
          6691 => x"fe",
          6692 => x"77",
          6693 => x"78",
          6694 => x"a0",
          6695 => x"74",
          6696 => x"52",
          6697 => x"3f",
          6698 => x"08",
          6699 => x"38",
          6700 => x"74",
          6701 => x"38",
          6702 => x"81",
          6703 => x"77",
          6704 => x"74",
          6705 => x"51",
          6706 => x"94",
          6707 => x"eb",
          6708 => x"15",
          6709 => x"58",
          6710 => x"87",
          6711 => x"81",
          6712 => x"70",
          6713 => x"57",
          6714 => x"87",
          6715 => x"38",
          6716 => x"f9",
          6717 => x"c8",
          6718 => x"81",
          6719 => x"e3",
          6720 => x"84",
          6721 => x"7a",
          6722 => x"82",
          6723 => x"d8",
          6724 => x"82",
          6725 => x"84",
          6726 => x"06",
          6727 => x"02",
          6728 => x"33",
          6729 => x"02",
          6730 => x"33",
          6731 => x"70",
          6732 => x"55",
          6733 => x"73",
          6734 => x"38",
          6735 => x"1d",
          6736 => x"c1",
          6737 => x"c8",
          6738 => x"78",
          6739 => x"f3",
          6740 => x"d8",
          6741 => x"82",
          6742 => x"82",
          6743 => x"19",
          6744 => x"2e",
          6745 => x"78",
          6746 => x"1b",
          6747 => x"53",
          6748 => x"ef",
          6749 => x"d8",
          6750 => x"82",
          6751 => x"81",
          6752 => x"1a",
          6753 => x"3f",
          6754 => x"08",
          6755 => x"5d",
          6756 => x"52",
          6757 => x"ab",
          6758 => x"c8",
          6759 => x"d8",
          6760 => x"d7",
          6761 => x"08",
          6762 => x"7a",
          6763 => x"5a",
          6764 => x"8d",
          6765 => x"0b",
          6766 => x"82",
          6767 => x"8c",
          6768 => x"d8",
          6769 => x"9a",
          6770 => x"df",
          6771 => x"29",
          6772 => x"55",
          6773 => x"ff",
          6774 => x"38",
          6775 => x"70",
          6776 => x"57",
          6777 => x"52",
          6778 => x"17",
          6779 => x"51",
          6780 => x"73",
          6781 => x"ff",
          6782 => x"17",
          6783 => x"27",
          6784 => x"83",
          6785 => x"8b",
          6786 => x"1b",
          6787 => x"54",
          6788 => x"77",
          6789 => x"58",
          6790 => x"81",
          6791 => x"34",
          6792 => x"51",
          6793 => x"82",
          6794 => x"57",
          6795 => x"08",
          6796 => x"ff",
          6797 => x"fe",
          6798 => x"1a",
          6799 => x"51",
          6800 => x"82",
          6801 => x"57",
          6802 => x"08",
          6803 => x"53",
          6804 => x"08",
          6805 => x"08",
          6806 => x"3f",
          6807 => x"1a",
          6808 => x"08",
          6809 => x"3f",
          6810 => x"ab",
          6811 => x"06",
          6812 => x"8c",
          6813 => x"0b",
          6814 => x"76",
          6815 => x"d8",
          6816 => x"3d",
          6817 => x"3d",
          6818 => x"08",
          6819 => x"ac",
          6820 => x"59",
          6821 => x"ff",
          6822 => x"72",
          6823 => x"ed",
          6824 => x"d8",
          6825 => x"82",
          6826 => x"80",
          6827 => x"15",
          6828 => x"51",
          6829 => x"82",
          6830 => x"54",
          6831 => x"08",
          6832 => x"15",
          6833 => x"73",
          6834 => x"83",
          6835 => x"15",
          6836 => x"a2",
          6837 => x"c8",
          6838 => x"51",
          6839 => x"82",
          6840 => x"54",
          6841 => x"08",
          6842 => x"38",
          6843 => x"09",
          6844 => x"38",
          6845 => x"82",
          6846 => x"88",
          6847 => x"f4",
          6848 => x"60",
          6849 => x"59",
          6850 => x"96",
          6851 => x"1c",
          6852 => x"83",
          6853 => x"1c",
          6854 => x"81",
          6855 => x"70",
          6856 => x"05",
          6857 => x"57",
          6858 => x"57",
          6859 => x"81",
          6860 => x"10",
          6861 => x"81",
          6862 => x"53",
          6863 => x"80",
          6864 => x"70",
          6865 => x"06",
          6866 => x"8f",
          6867 => x"38",
          6868 => x"df",
          6869 => x"96",
          6870 => x"79",
          6871 => x"54",
          6872 => x"7a",
          6873 => x"07",
          6874 => x"98",
          6875 => x"c8",
          6876 => x"ff",
          6877 => x"ff",
          6878 => x"38",
          6879 => x"a5",
          6880 => x"2a",
          6881 => x"34",
          6882 => x"34",
          6883 => x"39",
          6884 => x"30",
          6885 => x"80",
          6886 => x"25",
          6887 => x"54",
          6888 => x"85",
          6889 => x"9a",
          6890 => x"34",
          6891 => x"17",
          6892 => x"8c",
          6893 => x"10",
          6894 => x"51",
          6895 => x"fe",
          6896 => x"30",
          6897 => x"70",
          6898 => x"59",
          6899 => x"17",
          6900 => x"80",
          6901 => x"34",
          6902 => x"1a",
          6903 => x"9c",
          6904 => x"70",
          6905 => x"5b",
          6906 => x"a0",
          6907 => x"74",
          6908 => x"81",
          6909 => x"81",
          6910 => x"89",
          6911 => x"70",
          6912 => x"25",
          6913 => x"76",
          6914 => x"38",
          6915 => x"8b",
          6916 => x"70",
          6917 => x"34",
          6918 => x"74",
          6919 => x"05",
          6920 => x"17",
          6921 => x"27",
          6922 => x"77",
          6923 => x"53",
          6924 => x"14",
          6925 => x"33",
          6926 => x"87",
          6927 => x"38",
          6928 => x"19",
          6929 => x"80",
          6930 => x"73",
          6931 => x"55",
          6932 => x"80",
          6933 => x"38",
          6934 => x"19",
          6935 => x"33",
          6936 => x"54",
          6937 => x"26",
          6938 => x"1c",
          6939 => x"33",
          6940 => x"79",
          6941 => x"72",
          6942 => x"85",
          6943 => x"2a",
          6944 => x"06",
          6945 => x"2e",
          6946 => x"15",
          6947 => x"ff",
          6948 => x"74",
          6949 => x"05",
          6950 => x"19",
          6951 => x"19",
          6952 => x"59",
          6953 => x"ff",
          6954 => x"17",
          6955 => x"80",
          6956 => x"34",
          6957 => x"8c",
          6958 => x"53",
          6959 => x"72",
          6960 => x"9c",
          6961 => x"8b",
          6962 => x"19",
          6963 => x"08",
          6964 => x"53",
          6965 => x"82",
          6966 => x"78",
          6967 => x"51",
          6968 => x"82",
          6969 => x"86",
          6970 => x"13",
          6971 => x"3f",
          6972 => x"08",
          6973 => x"8e",
          6974 => x"f0",
          6975 => x"70",
          6976 => x"80",
          6977 => x"51",
          6978 => x"af",
          6979 => x"81",
          6980 => x"dc",
          6981 => x"74",
          6982 => x"38",
          6983 => x"08",
          6984 => x"aa",
          6985 => x"44",
          6986 => x"33",
          6987 => x"73",
          6988 => x"81",
          6989 => x"81",
          6990 => x"dc",
          6991 => x"70",
          6992 => x"07",
          6993 => x"73",
          6994 => x"88",
          6995 => x"70",
          6996 => x"73",
          6997 => x"38",
          6998 => x"ab",
          6999 => x"52",
          7000 => x"ee",
          7001 => x"c8",
          7002 => x"e1",
          7003 => x"7d",
          7004 => x"08",
          7005 => x"59",
          7006 => x"05",
          7007 => x"3f",
          7008 => x"08",
          7009 => x"b1",
          7010 => x"ff",
          7011 => x"c8",
          7012 => x"38",
          7013 => x"82",
          7014 => x"90",
          7015 => x"73",
          7016 => x"19",
          7017 => x"c8",
          7018 => x"ff",
          7019 => x"32",
          7020 => x"73",
          7021 => x"25",
          7022 => x"55",
          7023 => x"38",
          7024 => x"2e",
          7025 => x"80",
          7026 => x"38",
          7027 => x"c9",
          7028 => x"92",
          7029 => x"c8",
          7030 => x"38",
          7031 => x"26",
          7032 => x"78",
          7033 => x"75",
          7034 => x"19",
          7035 => x"39",
          7036 => x"80",
          7037 => x"56",
          7038 => x"af",
          7039 => x"06",
          7040 => x"57",
          7041 => x"32",
          7042 => x"80",
          7043 => x"51",
          7044 => x"dc",
          7045 => x"9f",
          7046 => x"2b",
          7047 => x"2e",
          7048 => x"8c",
          7049 => x"54",
          7050 => x"a5",
          7051 => x"39",
          7052 => x"09",
          7053 => x"c9",
          7054 => x"22",
          7055 => x"2e",
          7056 => x"80",
          7057 => x"22",
          7058 => x"2e",
          7059 => x"b6",
          7060 => x"1a",
          7061 => x"23",
          7062 => x"1f",
          7063 => x"54",
          7064 => x"83",
          7065 => x"73",
          7066 => x"05",
          7067 => x"18",
          7068 => x"27",
          7069 => x"a0",
          7070 => x"ab",
          7071 => x"c4",
          7072 => x"2e",
          7073 => x"10",
          7074 => x"55",
          7075 => x"16",
          7076 => x"32",
          7077 => x"9f",
          7078 => x"53",
          7079 => x"75",
          7080 => x"38",
          7081 => x"ff",
          7082 => x"e0",
          7083 => x"7a",
          7084 => x"80",
          7085 => x"8d",
          7086 => x"85",
          7087 => x"83",
          7088 => x"99",
          7089 => x"22",
          7090 => x"ff",
          7091 => x"5d",
          7092 => x"09",
          7093 => x"38",
          7094 => x"10",
          7095 => x"51",
          7096 => x"a0",
          7097 => x"7c",
          7098 => x"83",
          7099 => x"54",
          7100 => x"09",
          7101 => x"38",
          7102 => x"57",
          7103 => x"aa",
          7104 => x"fe",
          7105 => x"51",
          7106 => x"2e",
          7107 => x"10",
          7108 => x"55",
          7109 => x"78",
          7110 => x"38",
          7111 => x"22",
          7112 => x"ae",
          7113 => x"06",
          7114 => x"53",
          7115 => x"1e",
          7116 => x"3f",
          7117 => x"5c",
          7118 => x"10",
          7119 => x"81",
          7120 => x"54",
          7121 => x"82",
          7122 => x"a0",
          7123 => x"75",
          7124 => x"30",
          7125 => x"51",
          7126 => x"79",
          7127 => x"73",
          7128 => x"38",
          7129 => x"57",
          7130 => x"54",
          7131 => x"78",
          7132 => x"81",
          7133 => x"32",
          7134 => x"72",
          7135 => x"70",
          7136 => x"51",
          7137 => x"80",
          7138 => x"7e",
          7139 => x"ae",
          7140 => x"2e",
          7141 => x"83",
          7142 => x"79",
          7143 => x"38",
          7144 => x"58",
          7145 => x"2b",
          7146 => x"5d",
          7147 => x"39",
          7148 => x"27",
          7149 => x"82",
          7150 => x"b5",
          7151 => x"80",
          7152 => x"82",
          7153 => x"83",
          7154 => x"70",
          7155 => x"81",
          7156 => x"56",
          7157 => x"8c",
          7158 => x"ff",
          7159 => x"e0",
          7160 => x"54",
          7161 => x"27",
          7162 => x"1f",
          7163 => x"26",
          7164 => x"83",
          7165 => x"57",
          7166 => x"7d",
          7167 => x"76",
          7168 => x"55",
          7169 => x"81",
          7170 => x"c3",
          7171 => x"2e",
          7172 => x"52",
          7173 => x"51",
          7174 => x"82",
          7175 => x"80",
          7176 => x"80",
          7177 => x"07",
          7178 => x"39",
          7179 => x"54",
          7180 => x"85",
          7181 => x"07",
          7182 => x"16",
          7183 => x"26",
          7184 => x"81",
          7185 => x"70",
          7186 => x"06",
          7187 => x"7d",
          7188 => x"54",
          7189 => x"81",
          7190 => x"de",
          7191 => x"33",
          7192 => x"e5",
          7193 => x"06",
          7194 => x"0b",
          7195 => x"7e",
          7196 => x"81",
          7197 => x"7b",
          7198 => x"fc",
          7199 => x"8c",
          7200 => x"8c",
          7201 => x"7b",
          7202 => x"73",
          7203 => x"81",
          7204 => x"76",
          7205 => x"76",
          7206 => x"81",
          7207 => x"73",
          7208 => x"81",
          7209 => x"80",
          7210 => x"76",
          7211 => x"7b",
          7212 => x"81",
          7213 => x"73",
          7214 => x"38",
          7215 => x"57",
          7216 => x"34",
          7217 => x"a5",
          7218 => x"c8",
          7219 => x"33",
          7220 => x"d8",
          7221 => x"2e",
          7222 => x"d8",
          7223 => x"2e",
          7224 => x"80",
          7225 => x"85",
          7226 => x"06",
          7227 => x"57",
          7228 => x"80",
          7229 => x"74",
          7230 => x"73",
          7231 => x"ed",
          7232 => x"0b",
          7233 => x"80",
          7234 => x"39",
          7235 => x"54",
          7236 => x"85",
          7237 => x"74",
          7238 => x"81",
          7239 => x"73",
          7240 => x"1e",
          7241 => x"2a",
          7242 => x"51",
          7243 => x"80",
          7244 => x"90",
          7245 => x"ff",
          7246 => x"b8",
          7247 => x"51",
          7248 => x"82",
          7249 => x"88",
          7250 => x"a1",
          7251 => x"d8",
          7252 => x"3d",
          7253 => x"3d",
          7254 => x"ff",
          7255 => x"71",
          7256 => x"5c",
          7257 => x"80",
          7258 => x"38",
          7259 => x"05",
          7260 => x"9f",
          7261 => x"71",
          7262 => x"38",
          7263 => x"71",
          7264 => x"81",
          7265 => x"38",
          7266 => x"11",
          7267 => x"06",
          7268 => x"70",
          7269 => x"38",
          7270 => x"81",
          7271 => x"05",
          7272 => x"76",
          7273 => x"38",
          7274 => x"ca",
          7275 => x"77",
          7276 => x"57",
          7277 => x"05",
          7278 => x"70",
          7279 => x"33",
          7280 => x"53",
          7281 => x"99",
          7282 => x"e0",
          7283 => x"ff",
          7284 => x"ff",
          7285 => x"70",
          7286 => x"38",
          7287 => x"81",
          7288 => x"51",
          7289 => x"9f",
          7290 => x"72",
          7291 => x"81",
          7292 => x"70",
          7293 => x"72",
          7294 => x"32",
          7295 => x"72",
          7296 => x"73",
          7297 => x"53",
          7298 => x"70",
          7299 => x"38",
          7300 => x"19",
          7301 => x"75",
          7302 => x"38",
          7303 => x"83",
          7304 => x"74",
          7305 => x"59",
          7306 => x"39",
          7307 => x"33",
          7308 => x"d8",
          7309 => x"3d",
          7310 => x"3d",
          7311 => x"80",
          7312 => x"34",
          7313 => x"17",
          7314 => x"75",
          7315 => x"3f",
          7316 => x"d8",
          7317 => x"80",
          7318 => x"16",
          7319 => x"3f",
          7320 => x"08",
          7321 => x"06",
          7322 => x"73",
          7323 => x"2e",
          7324 => x"80",
          7325 => x"0b",
          7326 => x"56",
          7327 => x"e9",
          7328 => x"06",
          7329 => x"57",
          7330 => x"32",
          7331 => x"80",
          7332 => x"51",
          7333 => x"8a",
          7334 => x"e8",
          7335 => x"06",
          7336 => x"53",
          7337 => x"52",
          7338 => x"51",
          7339 => x"82",
          7340 => x"55",
          7341 => x"08",
          7342 => x"38",
          7343 => x"ca",
          7344 => x"8a",
          7345 => x"ed",
          7346 => x"c8",
          7347 => x"d8",
          7348 => x"2e",
          7349 => x"55",
          7350 => x"c8",
          7351 => x"0d",
          7352 => x"0d",
          7353 => x"05",
          7354 => x"33",
          7355 => x"75",
          7356 => x"fc",
          7357 => x"d8",
          7358 => x"8b",
          7359 => x"82",
          7360 => x"24",
          7361 => x"82",
          7362 => x"84",
          7363 => x"90",
          7364 => x"55",
          7365 => x"73",
          7366 => x"ee",
          7367 => x"0c",
          7368 => x"06",
          7369 => x"57",
          7370 => x"ae",
          7371 => x"33",
          7372 => x"3f",
          7373 => x"08",
          7374 => x"70",
          7375 => x"55",
          7376 => x"76",
          7377 => x"c0",
          7378 => x"2a",
          7379 => x"51",
          7380 => x"72",
          7381 => x"86",
          7382 => x"74",
          7383 => x"15",
          7384 => x"81",
          7385 => x"c6",
          7386 => x"d8",
          7387 => x"ff",
          7388 => x"06",
          7389 => x"56",
          7390 => x"38",
          7391 => x"8f",
          7392 => x"2a",
          7393 => x"51",
          7394 => x"72",
          7395 => x"80",
          7396 => x"52",
          7397 => x"3f",
          7398 => x"08",
          7399 => x"57",
          7400 => x"09",
          7401 => x"e2",
          7402 => x"74",
          7403 => x"56",
          7404 => x"33",
          7405 => x"72",
          7406 => x"38",
          7407 => x"51",
          7408 => x"82",
          7409 => x"57",
          7410 => x"84",
          7411 => x"ff",
          7412 => x"56",
          7413 => x"25",
          7414 => x"0b",
          7415 => x"56",
          7416 => x"05",
          7417 => x"83",
          7418 => x"2e",
          7419 => x"52",
          7420 => x"c6",
          7421 => x"c8",
          7422 => x"06",
          7423 => x"27",
          7424 => x"16",
          7425 => x"27",
          7426 => x"56",
          7427 => x"84",
          7428 => x"56",
          7429 => x"84",
          7430 => x"c3",
          7431 => x"c9",
          7432 => x"c8",
          7433 => x"ff",
          7434 => x"84",
          7435 => x"81",
          7436 => x"38",
          7437 => x"51",
          7438 => x"82",
          7439 => x"83",
          7440 => x"58",
          7441 => x"80",
          7442 => x"ca",
          7443 => x"d8",
          7444 => x"77",
          7445 => x"80",
          7446 => x"82",
          7447 => x"c8",
          7448 => x"11",
          7449 => x"06",
          7450 => x"8d",
          7451 => x"26",
          7452 => x"74",
          7453 => x"78",
          7454 => x"c5",
          7455 => x"59",
          7456 => x"15",
          7457 => x"2e",
          7458 => x"13",
          7459 => x"72",
          7460 => x"38",
          7461 => x"f2",
          7462 => x"14",
          7463 => x"3f",
          7464 => x"08",
          7465 => x"c8",
          7466 => x"23",
          7467 => x"57",
          7468 => x"83",
          7469 => x"cb",
          7470 => x"ad",
          7471 => x"c8",
          7472 => x"ff",
          7473 => x"8d",
          7474 => x"14",
          7475 => x"3f",
          7476 => x"08",
          7477 => x"14",
          7478 => x"3f",
          7479 => x"08",
          7480 => x"06",
          7481 => x"72",
          7482 => x"9e",
          7483 => x"22",
          7484 => x"84",
          7485 => x"5a",
          7486 => x"83",
          7487 => x"14",
          7488 => x"79",
          7489 => x"dc",
          7490 => x"d8",
          7491 => x"82",
          7492 => x"80",
          7493 => x"38",
          7494 => x"08",
          7495 => x"ff",
          7496 => x"38",
          7497 => x"83",
          7498 => x"83",
          7499 => x"74",
          7500 => x"85",
          7501 => x"89",
          7502 => x"76",
          7503 => x"ca",
          7504 => x"70",
          7505 => x"7b",
          7506 => x"73",
          7507 => x"17",
          7508 => x"b0",
          7509 => x"55",
          7510 => x"09",
          7511 => x"38",
          7512 => x"51",
          7513 => x"82",
          7514 => x"83",
          7515 => x"53",
          7516 => x"82",
          7517 => x"82",
          7518 => x"e4",
          7519 => x"80",
          7520 => x"c8",
          7521 => x"0c",
          7522 => x"53",
          7523 => x"56",
          7524 => x"81",
          7525 => x"13",
          7526 => x"74",
          7527 => x"82",
          7528 => x"74",
          7529 => x"81",
          7530 => x"06",
          7531 => x"83",
          7532 => x"2a",
          7533 => x"72",
          7534 => x"26",
          7535 => x"ff",
          7536 => x"0c",
          7537 => x"15",
          7538 => x"0b",
          7539 => x"76",
          7540 => x"81",
          7541 => x"38",
          7542 => x"51",
          7543 => x"82",
          7544 => x"83",
          7545 => x"53",
          7546 => x"09",
          7547 => x"f9",
          7548 => x"52",
          7549 => x"cb",
          7550 => x"c8",
          7551 => x"38",
          7552 => x"08",
          7553 => x"84",
          7554 => x"c6",
          7555 => x"d8",
          7556 => x"ff",
          7557 => x"72",
          7558 => x"2e",
          7559 => x"80",
          7560 => x"14",
          7561 => x"3f",
          7562 => x"08",
          7563 => x"a4",
          7564 => x"81",
          7565 => x"84",
          7566 => x"c6",
          7567 => x"d8",
          7568 => x"8a",
          7569 => x"2e",
          7570 => x"9d",
          7571 => x"14",
          7572 => x"3f",
          7573 => x"08",
          7574 => x"84",
          7575 => x"c6",
          7576 => x"d8",
          7577 => x"15",
          7578 => x"34",
          7579 => x"22",
          7580 => x"72",
          7581 => x"23",
          7582 => x"23",
          7583 => x"0b",
          7584 => x"80",
          7585 => x"0c",
          7586 => x"82",
          7587 => x"90",
          7588 => x"fb",
          7589 => x"54",
          7590 => x"80",
          7591 => x"73",
          7592 => x"80",
          7593 => x"72",
          7594 => x"80",
          7595 => x"86",
          7596 => x"15",
          7597 => x"71",
          7598 => x"81",
          7599 => x"81",
          7600 => x"ff",
          7601 => x"82",
          7602 => x"81",
          7603 => x"88",
          7604 => x"08",
          7605 => x"39",
          7606 => x"73",
          7607 => x"74",
          7608 => x"0c",
          7609 => x"04",
          7610 => x"02",
          7611 => x"7a",
          7612 => x"fc",
          7613 => x"f4",
          7614 => x"54",
          7615 => x"d8",
          7616 => x"bc",
          7617 => x"c8",
          7618 => x"82",
          7619 => x"70",
          7620 => x"73",
          7621 => x"38",
          7622 => x"78",
          7623 => x"2e",
          7624 => x"74",
          7625 => x"0c",
          7626 => x"80",
          7627 => x"80",
          7628 => x"70",
          7629 => x"51",
          7630 => x"82",
          7631 => x"54",
          7632 => x"c8",
          7633 => x"0d",
          7634 => x"0d",
          7635 => x"05",
          7636 => x"33",
          7637 => x"54",
          7638 => x"84",
          7639 => x"bf",
          7640 => x"99",
          7641 => x"53",
          7642 => x"05",
          7643 => x"f1",
          7644 => x"c8",
          7645 => x"d8",
          7646 => x"a4",
          7647 => x"69",
          7648 => x"70",
          7649 => x"f3",
          7650 => x"c8",
          7651 => x"d8",
          7652 => x"38",
          7653 => x"05",
          7654 => x"2b",
          7655 => x"80",
          7656 => x"86",
          7657 => x"06",
          7658 => x"2e",
          7659 => x"74",
          7660 => x"38",
          7661 => x"09",
          7662 => x"38",
          7663 => x"f4",
          7664 => x"c8",
          7665 => x"39",
          7666 => x"33",
          7667 => x"73",
          7668 => x"77",
          7669 => x"81",
          7670 => x"73",
          7671 => x"38",
          7672 => x"bc",
          7673 => x"07",
          7674 => x"b4",
          7675 => x"2a",
          7676 => x"51",
          7677 => x"2e",
          7678 => x"62",
          7679 => x"d7",
          7680 => x"d8",
          7681 => x"82",
          7682 => x"52",
          7683 => x"51",
          7684 => x"62",
          7685 => x"8b",
          7686 => x"53",
          7687 => x"51",
          7688 => x"80",
          7689 => x"05",
          7690 => x"3f",
          7691 => x"0b",
          7692 => x"75",
          7693 => x"f1",
          7694 => x"11",
          7695 => x"80",
          7696 => x"98",
          7697 => x"51",
          7698 => x"82",
          7699 => x"55",
          7700 => x"08",
          7701 => x"b7",
          7702 => x"c4",
          7703 => x"05",
          7704 => x"2a",
          7705 => x"51",
          7706 => x"80",
          7707 => x"84",
          7708 => x"39",
          7709 => x"70",
          7710 => x"54",
          7711 => x"a9",
          7712 => x"06",
          7713 => x"2e",
          7714 => x"55",
          7715 => x"73",
          7716 => x"c5",
          7717 => x"d8",
          7718 => x"ff",
          7719 => x"0c",
          7720 => x"d8",
          7721 => x"f8",
          7722 => x"2a",
          7723 => x"51",
          7724 => x"2e",
          7725 => x"80",
          7726 => x"7a",
          7727 => x"a0",
          7728 => x"a4",
          7729 => x"53",
          7730 => x"d5",
          7731 => x"d8",
          7732 => x"d8",
          7733 => x"1b",
          7734 => x"05",
          7735 => x"a0",
          7736 => x"c8",
          7737 => x"c8",
          7738 => x"0c",
          7739 => x"56",
          7740 => x"84",
          7741 => x"90",
          7742 => x"0b",
          7743 => x"80",
          7744 => x"0c",
          7745 => x"1a",
          7746 => x"2a",
          7747 => x"51",
          7748 => x"2e",
          7749 => x"82",
          7750 => x"80",
          7751 => x"38",
          7752 => x"08",
          7753 => x"8a",
          7754 => x"89",
          7755 => x"59",
          7756 => x"76",
          7757 => x"c6",
          7758 => x"d8",
          7759 => x"82",
          7760 => x"81",
          7761 => x"82",
          7762 => x"c8",
          7763 => x"09",
          7764 => x"38",
          7765 => x"78",
          7766 => x"30",
          7767 => x"80",
          7768 => x"77",
          7769 => x"38",
          7770 => x"06",
          7771 => x"c3",
          7772 => x"1a",
          7773 => x"38",
          7774 => x"06",
          7775 => x"2e",
          7776 => x"52",
          7777 => x"b1",
          7778 => x"c8",
          7779 => x"82",
          7780 => x"75",
          7781 => x"d8",
          7782 => x"9c",
          7783 => x"39",
          7784 => x"74",
          7785 => x"d8",
          7786 => x"3d",
          7787 => x"3d",
          7788 => x"65",
          7789 => x"5d",
          7790 => x"0c",
          7791 => x"05",
          7792 => x"f9",
          7793 => x"d8",
          7794 => x"82",
          7795 => x"8a",
          7796 => x"33",
          7797 => x"2e",
          7798 => x"56",
          7799 => x"90",
          7800 => x"06",
          7801 => x"74",
          7802 => x"b9",
          7803 => x"82",
          7804 => x"34",
          7805 => x"ad",
          7806 => x"91",
          7807 => x"56",
          7808 => x"8c",
          7809 => x"1a",
          7810 => x"74",
          7811 => x"38",
          7812 => x"80",
          7813 => x"38",
          7814 => x"70",
          7815 => x"56",
          7816 => x"b4",
          7817 => x"11",
          7818 => x"77",
          7819 => x"5b",
          7820 => x"38",
          7821 => x"88",
          7822 => x"8f",
          7823 => x"08",
          7824 => x"c4",
          7825 => x"d8",
          7826 => x"81",
          7827 => x"9f",
          7828 => x"2e",
          7829 => x"74",
          7830 => x"98",
          7831 => x"7e",
          7832 => x"3f",
          7833 => x"08",
          7834 => x"83",
          7835 => x"c8",
          7836 => x"89",
          7837 => x"77",
          7838 => x"d8",
          7839 => x"7f",
          7840 => x"58",
          7841 => x"75",
          7842 => x"75",
          7843 => x"77",
          7844 => x"7c",
          7845 => x"33",
          7846 => x"d4",
          7847 => x"c8",
          7848 => x"38",
          7849 => x"33",
          7850 => x"80",
          7851 => x"b4",
          7852 => x"31",
          7853 => x"27",
          7854 => x"80",
          7855 => x"52",
          7856 => x"77",
          7857 => x"7d",
          7858 => x"be",
          7859 => x"89",
          7860 => x"39",
          7861 => x"0c",
          7862 => x"83",
          7863 => x"80",
          7864 => x"55",
          7865 => x"83",
          7866 => x"9c",
          7867 => x"7e",
          7868 => x"3f",
          7869 => x"08",
          7870 => x"75",
          7871 => x"08",
          7872 => x"1f",
          7873 => x"7c",
          7874 => x"ec",
          7875 => x"31",
          7876 => x"7f",
          7877 => x"94",
          7878 => x"94",
          7879 => x"5c",
          7880 => x"80",
          7881 => x"d8",
          7882 => x"3d",
          7883 => x"3d",
          7884 => x"65",
          7885 => x"5d",
          7886 => x"0c",
          7887 => x"05",
          7888 => x"f6",
          7889 => x"d8",
          7890 => x"82",
          7891 => x"8a",
          7892 => x"33",
          7893 => x"2e",
          7894 => x"56",
          7895 => x"90",
          7896 => x"81",
          7897 => x"06",
          7898 => x"87",
          7899 => x"2e",
          7900 => x"95",
          7901 => x"91",
          7902 => x"56",
          7903 => x"81",
          7904 => x"34",
          7905 => x"94",
          7906 => x"08",
          7907 => x"56",
          7908 => x"84",
          7909 => x"5c",
          7910 => x"82",
          7911 => x"18",
          7912 => x"ff",
          7913 => x"74",
          7914 => x"7e",
          7915 => x"ff",
          7916 => x"2a",
          7917 => x"7a",
          7918 => x"8c",
          7919 => x"08",
          7920 => x"38",
          7921 => x"39",
          7922 => x"52",
          7923 => x"ef",
          7924 => x"c8",
          7925 => x"d8",
          7926 => x"2e",
          7927 => x"74",
          7928 => x"91",
          7929 => x"2e",
          7930 => x"74",
          7931 => x"88",
          7932 => x"38",
          7933 => x"0c",
          7934 => x"15",
          7935 => x"08",
          7936 => x"06",
          7937 => x"51",
          7938 => x"3f",
          7939 => x"08",
          7940 => x"98",
          7941 => x"7e",
          7942 => x"3f",
          7943 => x"08",
          7944 => x"d1",
          7945 => x"c8",
          7946 => x"89",
          7947 => x"78",
          7948 => x"d7",
          7949 => x"7f",
          7950 => x"58",
          7951 => x"75",
          7952 => x"75",
          7953 => x"78",
          7954 => x"7c",
          7955 => x"33",
          7956 => x"86",
          7957 => x"c8",
          7958 => x"38",
          7959 => x"08",
          7960 => x"56",
          7961 => x"9c",
          7962 => x"53",
          7963 => x"77",
          7964 => x"7d",
          7965 => x"16",
          7966 => x"fc",
          7967 => x"80",
          7968 => x"34",
          7969 => x"56",
          7970 => x"8c",
          7971 => x"19",
          7972 => x"38",
          7973 => x"bc",
          7974 => x"d8",
          7975 => x"df",
          7976 => x"b4",
          7977 => x"76",
          7978 => x"94",
          7979 => x"ff",
          7980 => x"71",
          7981 => x"7b",
          7982 => x"38",
          7983 => x"18",
          7984 => x"51",
          7985 => x"3f",
          7986 => x"08",
          7987 => x"75",
          7988 => x"94",
          7989 => x"ff",
          7990 => x"05",
          7991 => x"98",
          7992 => x"81",
          7993 => x"34",
          7994 => x"7e",
          7995 => x"0c",
          7996 => x"1a",
          7997 => x"94",
          7998 => x"1b",
          7999 => x"5e",
          8000 => x"27",
          8001 => x"55",
          8002 => x"0c",
          8003 => x"90",
          8004 => x"c0",
          8005 => x"90",
          8006 => x"56",
          8007 => x"c8",
          8008 => x"0d",
          8009 => x"0d",
          8010 => x"fc",
          8011 => x"52",
          8012 => x"3f",
          8013 => x"08",
          8014 => x"c8",
          8015 => x"38",
          8016 => x"70",
          8017 => x"81",
          8018 => x"55",
          8019 => x"80",
          8020 => x"16",
          8021 => x"51",
          8022 => x"3f",
          8023 => x"08",
          8024 => x"c8",
          8025 => x"38",
          8026 => x"8b",
          8027 => x"07",
          8028 => x"8b",
          8029 => x"16",
          8030 => x"52",
          8031 => x"cc",
          8032 => x"16",
          8033 => x"15",
          8034 => x"bd",
          8035 => x"b2",
          8036 => x"15",
          8037 => x"b1",
          8038 => x"92",
          8039 => x"b8",
          8040 => x"54",
          8041 => x"15",
          8042 => x"ff",
          8043 => x"82",
          8044 => x"90",
          8045 => x"bf",
          8046 => x"73",
          8047 => x"76",
          8048 => x"0c",
          8049 => x"04",
          8050 => x"76",
          8051 => x"fe",
          8052 => x"d8",
          8053 => x"82",
          8054 => x"9c",
          8055 => x"fc",
          8056 => x"51",
          8057 => x"82",
          8058 => x"53",
          8059 => x"08",
          8060 => x"d8",
          8061 => x"0c",
          8062 => x"c8",
          8063 => x"0d",
          8064 => x"0d",
          8065 => x"e6",
          8066 => x"52",
          8067 => x"d8",
          8068 => x"8b",
          8069 => x"c8",
          8070 => x"a4",
          8071 => x"71",
          8072 => x"0c",
          8073 => x"04",
          8074 => x"80",
          8075 => x"cc",
          8076 => x"3d",
          8077 => x"3f",
          8078 => x"08",
          8079 => x"c8",
          8080 => x"38",
          8081 => x"52",
          8082 => x"05",
          8083 => x"3f",
          8084 => x"08",
          8085 => x"c8",
          8086 => x"02",
          8087 => x"33",
          8088 => x"55",
          8089 => x"25",
          8090 => x"7a",
          8091 => x"54",
          8092 => x"a2",
          8093 => x"84",
          8094 => x"06",
          8095 => x"73",
          8096 => x"38",
          8097 => x"70",
          8098 => x"a5",
          8099 => x"c8",
          8100 => x"0c",
          8101 => x"d8",
          8102 => x"2e",
          8103 => x"83",
          8104 => x"74",
          8105 => x"0c",
          8106 => x"04",
          8107 => x"0d",
          8108 => x"08",
          8109 => x"08",
          8110 => x"7a",
          8111 => x"80",
          8112 => x"b4",
          8113 => x"e0",
          8114 => x"95",
          8115 => x"c8",
          8116 => x"d8",
          8117 => x"a1",
          8118 => x"d4",
          8119 => x"7c",
          8120 => x"80",
          8121 => x"55",
          8122 => x"3d",
          8123 => x"80",
          8124 => x"38",
          8125 => x"d3",
          8126 => x"55",
          8127 => x"82",
          8128 => x"57",
          8129 => x"08",
          8130 => x"80",
          8131 => x"52",
          8132 => x"b8",
          8133 => x"d8",
          8134 => x"82",
          8135 => x"82",
          8136 => x"da",
          8137 => x"7b",
          8138 => x"3f",
          8139 => x"08",
          8140 => x"0c",
          8141 => x"51",
          8142 => x"82",
          8143 => x"57",
          8144 => x"08",
          8145 => x"80",
          8146 => x"c9",
          8147 => x"d8",
          8148 => x"82",
          8149 => x"a7",
          8150 => x"3d",
          8151 => x"51",
          8152 => x"73",
          8153 => x"08",
          8154 => x"76",
          8155 => x"c5",
          8156 => x"d8",
          8157 => x"82",
          8158 => x"80",
          8159 => x"76",
          8160 => x"81",
          8161 => x"82",
          8162 => x"39",
          8163 => x"38",
          8164 => x"fd",
          8165 => x"74",
          8166 => x"3f",
          8167 => x"78",
          8168 => x"33",
          8169 => x"56",
          8170 => x"92",
          8171 => x"c6",
          8172 => x"16",
          8173 => x"33",
          8174 => x"73",
          8175 => x"16",
          8176 => x"26",
          8177 => x"75",
          8178 => x"38",
          8179 => x"05",
          8180 => x"80",
          8181 => x"11",
          8182 => x"18",
          8183 => x"58",
          8184 => x"34",
          8185 => x"ff",
          8186 => x"3d",
          8187 => x"58",
          8188 => x"fd",
          8189 => x"7b",
          8190 => x"06",
          8191 => x"18",
          8192 => x"08",
          8193 => x"af",
          8194 => x"0b",
          8195 => x"33",
          8196 => x"82",
          8197 => x"70",
          8198 => x"52",
          8199 => x"56",
          8200 => x"8d",
          8201 => x"70",
          8202 => x"51",
          8203 => x"f5",
          8204 => x"54",
          8205 => x"a7",
          8206 => x"74",
          8207 => x"38",
          8208 => x"73",
          8209 => x"81",
          8210 => x"81",
          8211 => x"39",
          8212 => x"81",
          8213 => x"74",
          8214 => x"81",
          8215 => x"91",
          8216 => x"80",
          8217 => x"18",
          8218 => x"54",
          8219 => x"70",
          8220 => x"34",
          8221 => x"eb",
          8222 => x"34",
          8223 => x"c8",
          8224 => x"3d",
          8225 => x"3d",
          8226 => x"8d",
          8227 => x"54",
          8228 => x"55",
          8229 => x"82",
          8230 => x"53",
          8231 => x"08",
          8232 => x"91",
          8233 => x"72",
          8234 => x"8c",
          8235 => x"73",
          8236 => x"38",
          8237 => x"70",
          8238 => x"81",
          8239 => x"57",
          8240 => x"73",
          8241 => x"08",
          8242 => x"94",
          8243 => x"75",
          8244 => x"9b",
          8245 => x"11",
          8246 => x"2b",
          8247 => x"73",
          8248 => x"38",
          8249 => x"16",
          8250 => x"99",
          8251 => x"c8",
          8252 => x"78",
          8253 => x"55",
          8254 => x"89",
          8255 => x"c8",
          8256 => x"96",
          8257 => x"70",
          8258 => x"94",
          8259 => x"71",
          8260 => x"08",
          8261 => x"53",
          8262 => x"15",
          8263 => x"a7",
          8264 => x"74",
          8265 => x"97",
          8266 => x"c8",
          8267 => x"d8",
          8268 => x"2e",
          8269 => x"82",
          8270 => x"ff",
          8271 => x"38",
          8272 => x"08",
          8273 => x"73",
          8274 => x"73",
          8275 => x"9f",
          8276 => x"27",
          8277 => x"75",
          8278 => x"16",
          8279 => x"17",
          8280 => x"33",
          8281 => x"70",
          8282 => x"55",
          8283 => x"80",
          8284 => x"73",
          8285 => x"ff",
          8286 => x"82",
          8287 => x"54",
          8288 => x"08",
          8289 => x"d8",
          8290 => x"a8",
          8291 => x"74",
          8292 => x"cf",
          8293 => x"c8",
          8294 => x"ff",
          8295 => x"81",
          8296 => x"38",
          8297 => x"9c",
          8298 => x"a7",
          8299 => x"16",
          8300 => x"39",
          8301 => x"16",
          8302 => x"75",
          8303 => x"53",
          8304 => x"ab",
          8305 => x"79",
          8306 => x"ed",
          8307 => x"c8",
          8308 => x"82",
          8309 => x"34",
          8310 => x"c4",
          8311 => x"91",
          8312 => x"53",
          8313 => x"89",
          8314 => x"c8",
          8315 => x"94",
          8316 => x"8c",
          8317 => x"27",
          8318 => x"8c",
          8319 => x"15",
          8320 => x"07",
          8321 => x"16",
          8322 => x"ff",
          8323 => x"80",
          8324 => x"77",
          8325 => x"2e",
          8326 => x"9c",
          8327 => x"53",
          8328 => x"c8",
          8329 => x"0d",
          8330 => x"0d",
          8331 => x"54",
          8332 => x"81",
          8333 => x"53",
          8334 => x"05",
          8335 => x"84",
          8336 => x"9d",
          8337 => x"c8",
          8338 => x"d8",
          8339 => x"eb",
          8340 => x"0c",
          8341 => x"51",
          8342 => x"82",
          8343 => x"55",
          8344 => x"08",
          8345 => x"ab",
          8346 => x"98",
          8347 => x"80",
          8348 => x"38",
          8349 => x"70",
          8350 => x"81",
          8351 => x"57",
          8352 => x"ae",
          8353 => x"08",
          8354 => x"c2",
          8355 => x"d8",
          8356 => x"17",
          8357 => x"86",
          8358 => x"17",
          8359 => x"75",
          8360 => x"ae",
          8361 => x"c8",
          8362 => x"84",
          8363 => x"06",
          8364 => x"55",
          8365 => x"80",
          8366 => x"80",
          8367 => x"54",
          8368 => x"c8",
          8369 => x"0d",
          8370 => x"0d",
          8371 => x"fc",
          8372 => x"52",
          8373 => x"3f",
          8374 => x"08",
          8375 => x"d8",
          8376 => x"0c",
          8377 => x"04",
          8378 => x"77",
          8379 => x"fc",
          8380 => x"53",
          8381 => x"9b",
          8382 => x"c8",
          8383 => x"d8",
          8384 => x"e1",
          8385 => x"38",
          8386 => x"08",
          8387 => x"ff",
          8388 => x"82",
          8389 => x"53",
          8390 => x"82",
          8391 => x"52",
          8392 => x"a3",
          8393 => x"c8",
          8394 => x"d8",
          8395 => x"2e",
          8396 => x"85",
          8397 => x"87",
          8398 => x"c8",
          8399 => x"74",
          8400 => x"cf",
          8401 => x"52",
          8402 => x"bd",
          8403 => x"d8",
          8404 => x"32",
          8405 => x"72",
          8406 => x"70",
          8407 => x"08",
          8408 => x"54",
          8409 => x"d8",
          8410 => x"3d",
          8411 => x"3d",
          8412 => x"80",
          8413 => x"70",
          8414 => x"52",
          8415 => x"3f",
          8416 => x"08",
          8417 => x"c8",
          8418 => x"65",
          8419 => x"d2",
          8420 => x"d8",
          8421 => x"82",
          8422 => x"a0",
          8423 => x"cb",
          8424 => x"98",
          8425 => x"73",
          8426 => x"38",
          8427 => x"39",
          8428 => x"88",
          8429 => x"75",
          8430 => x"3f",
          8431 => x"c8",
          8432 => x"0d",
          8433 => x"0d",
          8434 => x"5c",
          8435 => x"3d",
          8436 => x"93",
          8437 => x"89",
          8438 => x"c8",
          8439 => x"d8",
          8440 => x"82",
          8441 => x"0c",
          8442 => x"11",
          8443 => x"94",
          8444 => x"56",
          8445 => x"74",
          8446 => x"75",
          8447 => x"e6",
          8448 => x"81",
          8449 => x"5b",
          8450 => x"82",
          8451 => x"75",
          8452 => x"73",
          8453 => x"81",
          8454 => x"38",
          8455 => x"57",
          8456 => x"3d",
          8457 => x"ff",
          8458 => x"82",
          8459 => x"ff",
          8460 => x"82",
          8461 => x"81",
          8462 => x"82",
          8463 => x"30",
          8464 => x"c8",
          8465 => x"25",
          8466 => x"19",
          8467 => x"5a",
          8468 => x"08",
          8469 => x"38",
          8470 => x"a8",
          8471 => x"d8",
          8472 => x"58",
          8473 => x"77",
          8474 => x"7d",
          8475 => x"ad",
          8476 => x"d8",
          8477 => x"82",
          8478 => x"80",
          8479 => x"70",
          8480 => x"ff",
          8481 => x"56",
          8482 => x"2e",
          8483 => x"9e",
          8484 => x"51",
          8485 => x"3f",
          8486 => x"08",
          8487 => x"06",
          8488 => x"80",
          8489 => x"19",
          8490 => x"54",
          8491 => x"14",
          8492 => x"cc",
          8493 => x"c8",
          8494 => x"06",
          8495 => x"80",
          8496 => x"19",
          8497 => x"54",
          8498 => x"06",
          8499 => x"79",
          8500 => x"78",
          8501 => x"79",
          8502 => x"84",
          8503 => x"07",
          8504 => x"84",
          8505 => x"82",
          8506 => x"92",
          8507 => x"f9",
          8508 => x"8a",
          8509 => x"53",
          8510 => x"e3",
          8511 => x"d8",
          8512 => x"82",
          8513 => x"81",
          8514 => x"17",
          8515 => x"81",
          8516 => x"17",
          8517 => x"2a",
          8518 => x"51",
          8519 => x"55",
          8520 => x"81",
          8521 => x"17",
          8522 => x"8c",
          8523 => x"81",
          8524 => x"9c",
          8525 => x"c8",
          8526 => x"17",
          8527 => x"51",
          8528 => x"3f",
          8529 => x"08",
          8530 => x"0c",
          8531 => x"39",
          8532 => x"52",
          8533 => x"ae",
          8534 => x"d8",
          8535 => x"2e",
          8536 => x"83",
          8537 => x"82",
          8538 => x"81",
          8539 => x"06",
          8540 => x"56",
          8541 => x"a1",
          8542 => x"82",
          8543 => x"9c",
          8544 => x"95",
          8545 => x"08",
          8546 => x"c8",
          8547 => x"51",
          8548 => x"3f",
          8549 => x"08",
          8550 => x"08",
          8551 => x"90",
          8552 => x"c0",
          8553 => x"90",
          8554 => x"80",
          8555 => x"75",
          8556 => x"75",
          8557 => x"d8",
          8558 => x"3d",
          8559 => x"3d",
          8560 => x"a2",
          8561 => x"05",
          8562 => x"51",
          8563 => x"82",
          8564 => x"55",
          8565 => x"08",
          8566 => x"78",
          8567 => x"08",
          8568 => x"70",
          8569 => x"93",
          8570 => x"c8",
          8571 => x"d8",
          8572 => x"df",
          8573 => x"ff",
          8574 => x"85",
          8575 => x"06",
          8576 => x"86",
          8577 => x"cb",
          8578 => x"2b",
          8579 => x"24",
          8580 => x"02",
          8581 => x"33",
          8582 => x"58",
          8583 => x"76",
          8584 => x"6c",
          8585 => x"ff",
          8586 => x"82",
          8587 => x"74",
          8588 => x"81",
          8589 => x"56",
          8590 => x"80",
          8591 => x"54",
          8592 => x"08",
          8593 => x"2e",
          8594 => x"73",
          8595 => x"c8",
          8596 => x"52",
          8597 => x"52",
          8598 => x"f6",
          8599 => x"c8",
          8600 => x"d8",
          8601 => x"eb",
          8602 => x"c8",
          8603 => x"51",
          8604 => x"3f",
          8605 => x"08",
          8606 => x"c8",
          8607 => x"87",
          8608 => x"39",
          8609 => x"08",
          8610 => x"38",
          8611 => x"08",
          8612 => x"77",
          8613 => x"3f",
          8614 => x"08",
          8615 => x"08",
          8616 => x"d8",
          8617 => x"80",
          8618 => x"55",
          8619 => x"95",
          8620 => x"2e",
          8621 => x"53",
          8622 => x"51",
          8623 => x"3f",
          8624 => x"08",
          8625 => x"38",
          8626 => x"a9",
          8627 => x"d8",
          8628 => x"74",
          8629 => x"0c",
          8630 => x"04",
          8631 => x"82",
          8632 => x"ff",
          8633 => x"9b",
          8634 => x"f5",
          8635 => x"c8",
          8636 => x"d8",
          8637 => x"b7",
          8638 => x"6a",
          8639 => x"70",
          8640 => x"f7",
          8641 => x"c8",
          8642 => x"d8",
          8643 => x"38",
          8644 => x"9b",
          8645 => x"c8",
          8646 => x"09",
          8647 => x"8f",
          8648 => x"df",
          8649 => x"85",
          8650 => x"51",
          8651 => x"74",
          8652 => x"78",
          8653 => x"8a",
          8654 => x"57",
          8655 => x"3f",
          8656 => x"08",
          8657 => x"82",
          8658 => x"83",
          8659 => x"82",
          8660 => x"81",
          8661 => x"06",
          8662 => x"54",
          8663 => x"08",
          8664 => x"81",
          8665 => x"81",
          8666 => x"39",
          8667 => x"38",
          8668 => x"08",
          8669 => x"ff",
          8670 => x"82",
          8671 => x"54",
          8672 => x"08",
          8673 => x"8b",
          8674 => x"b8",
          8675 => x"a5",
          8676 => x"54",
          8677 => x"15",
          8678 => x"90",
          8679 => x"15",
          8680 => x"b2",
          8681 => x"ce",
          8682 => x"a4",
          8683 => x"53",
          8684 => x"53",
          8685 => x"b2",
          8686 => x"78",
          8687 => x"80",
          8688 => x"ff",
          8689 => x"78",
          8690 => x"80",
          8691 => x"7f",
          8692 => x"d8",
          8693 => x"ff",
          8694 => x"78",
          8695 => x"83",
          8696 => x"51",
          8697 => x"3f",
          8698 => x"08",
          8699 => x"c8",
          8700 => x"82",
          8701 => x"52",
          8702 => x"51",
          8703 => x"3f",
          8704 => x"52",
          8705 => x"b7",
          8706 => x"54",
          8707 => x"15",
          8708 => x"81",
          8709 => x"34",
          8710 => x"a6",
          8711 => x"d8",
          8712 => x"8b",
          8713 => x"75",
          8714 => x"ff",
          8715 => x"73",
          8716 => x"0c",
          8717 => x"04",
          8718 => x"ab",
          8719 => x"51",
          8720 => x"82",
          8721 => x"fe",
          8722 => x"ab",
          8723 => x"91",
          8724 => x"c8",
          8725 => x"d8",
          8726 => x"d8",
          8727 => x"ab",
          8728 => x"9e",
          8729 => x"58",
          8730 => x"82",
          8731 => x"55",
          8732 => x"08",
          8733 => x"02",
          8734 => x"33",
          8735 => x"54",
          8736 => x"82",
          8737 => x"53",
          8738 => x"52",
          8739 => x"80",
          8740 => x"a2",
          8741 => x"53",
          8742 => x"3d",
          8743 => x"ff",
          8744 => x"ac",
          8745 => x"73",
          8746 => x"3f",
          8747 => x"08",
          8748 => x"c8",
          8749 => x"63",
          8750 => x"2e",
          8751 => x"88",
          8752 => x"3d",
          8753 => x"38",
          8754 => x"e8",
          8755 => x"c8",
          8756 => x"09",
          8757 => x"bb",
          8758 => x"ff",
          8759 => x"82",
          8760 => x"55",
          8761 => x"08",
          8762 => x"68",
          8763 => x"aa",
          8764 => x"05",
          8765 => x"51",
          8766 => x"3f",
          8767 => x"33",
          8768 => x"8b",
          8769 => x"84",
          8770 => x"06",
          8771 => x"73",
          8772 => x"a0",
          8773 => x"8b",
          8774 => x"54",
          8775 => x"15",
          8776 => x"33",
          8777 => x"70",
          8778 => x"55",
          8779 => x"2e",
          8780 => x"6f",
          8781 => x"e1",
          8782 => x"78",
          8783 => x"f1",
          8784 => x"c8",
          8785 => x"51",
          8786 => x"3f",
          8787 => x"d8",
          8788 => x"2e",
          8789 => x"82",
          8790 => x"52",
          8791 => x"a3",
          8792 => x"d8",
          8793 => x"80",
          8794 => x"58",
          8795 => x"c8",
          8796 => x"38",
          8797 => x"54",
          8798 => x"09",
          8799 => x"38",
          8800 => x"52",
          8801 => x"b4",
          8802 => x"54",
          8803 => x"15",
          8804 => x"82",
          8805 => x"9c",
          8806 => x"c1",
          8807 => x"d8",
          8808 => x"82",
          8809 => x"8c",
          8810 => x"ff",
          8811 => x"82",
          8812 => x"55",
          8813 => x"c8",
          8814 => x"0d",
          8815 => x"0d",
          8816 => x"05",
          8817 => x"05",
          8818 => x"33",
          8819 => x"53",
          8820 => x"05",
          8821 => x"51",
          8822 => x"82",
          8823 => x"55",
          8824 => x"08",
          8825 => x"78",
          8826 => x"96",
          8827 => x"51",
          8828 => x"82",
          8829 => x"55",
          8830 => x"08",
          8831 => x"80",
          8832 => x"81",
          8833 => x"86",
          8834 => x"38",
          8835 => x"61",
          8836 => x"12",
          8837 => x"7a",
          8838 => x"51",
          8839 => x"74",
          8840 => x"78",
          8841 => x"83",
          8842 => x"51",
          8843 => x"3f",
          8844 => x"08",
          8845 => x"d8",
          8846 => x"3d",
          8847 => x"3d",
          8848 => x"82",
          8849 => x"cc",
          8850 => x"3d",
          8851 => x"3f",
          8852 => x"08",
          8853 => x"c8",
          8854 => x"38",
          8855 => x"52",
          8856 => x"05",
          8857 => x"3f",
          8858 => x"08",
          8859 => x"c8",
          8860 => x"02",
          8861 => x"33",
          8862 => x"54",
          8863 => x"a6",
          8864 => x"22",
          8865 => x"71",
          8866 => x"53",
          8867 => x"51",
          8868 => x"3f",
          8869 => x"0b",
          8870 => x"76",
          8871 => x"ea",
          8872 => x"c8",
          8873 => x"82",
          8874 => x"94",
          8875 => x"e9",
          8876 => x"6c",
          8877 => x"53",
          8878 => x"05",
          8879 => x"51",
          8880 => x"82",
          8881 => x"82",
          8882 => x"30",
          8883 => x"c8",
          8884 => x"25",
          8885 => x"79",
          8886 => x"86",
          8887 => x"75",
          8888 => x"73",
          8889 => x"fa",
          8890 => x"80",
          8891 => x"8d",
          8892 => x"54",
          8893 => x"3f",
          8894 => x"08",
          8895 => x"c8",
          8896 => x"38",
          8897 => x"51",
          8898 => x"3f",
          8899 => x"08",
          8900 => x"c8",
          8901 => x"82",
          8902 => x"82",
          8903 => x"65",
          8904 => x"78",
          8905 => x"7b",
          8906 => x"55",
          8907 => x"34",
          8908 => x"8a",
          8909 => x"38",
          8910 => x"1a",
          8911 => x"34",
          8912 => x"9e",
          8913 => x"70",
          8914 => x"51",
          8915 => x"a0",
          8916 => x"8e",
          8917 => x"2e",
          8918 => x"86",
          8919 => x"34",
          8920 => x"30",
          8921 => x"80",
          8922 => x"7a",
          8923 => x"c1",
          8924 => x"2e",
          8925 => x"a4",
          8926 => x"51",
          8927 => x"3f",
          8928 => x"08",
          8929 => x"c8",
          8930 => x"7b",
          8931 => x"55",
          8932 => x"73",
          8933 => x"38",
          8934 => x"73",
          8935 => x"38",
          8936 => x"15",
          8937 => x"ff",
          8938 => x"82",
          8939 => x"7b",
          8940 => x"d8",
          8941 => x"3d",
          8942 => x"3d",
          8943 => x"9c",
          8944 => x"05",
          8945 => x"51",
          8946 => x"82",
          8947 => x"82",
          8948 => x"56",
          8949 => x"c8",
          8950 => x"38",
          8951 => x"52",
          8952 => x"52",
          8953 => x"b3",
          8954 => x"70",
          8955 => x"56",
          8956 => x"81",
          8957 => x"57",
          8958 => x"ff",
          8959 => x"82",
          8960 => x"83",
          8961 => x"80",
          8962 => x"d8",
          8963 => x"95",
          8964 => x"b5",
          8965 => x"c8",
          8966 => x"e8",
          8967 => x"c8",
          8968 => x"ff",
          8969 => x"80",
          8970 => x"74",
          8971 => x"e0",
          8972 => x"b2",
          8973 => x"c8",
          8974 => x"81",
          8975 => x"88",
          8976 => x"26",
          8977 => x"39",
          8978 => x"86",
          8979 => x"81",
          8980 => x"ff",
          8981 => x"38",
          8982 => x"54",
          8983 => x"81",
          8984 => x"81",
          8985 => x"77",
          8986 => x"59",
          8987 => x"6d",
          8988 => x"55",
          8989 => x"26",
          8990 => x"8a",
          8991 => x"86",
          8992 => x"e5",
          8993 => x"38",
          8994 => x"99",
          8995 => x"05",
          8996 => x"70",
          8997 => x"73",
          8998 => x"81",
          8999 => x"ff",
          9000 => x"ed",
          9001 => x"80",
          9002 => x"90",
          9003 => x"55",
          9004 => x"3f",
          9005 => x"08",
          9006 => x"c8",
          9007 => x"38",
          9008 => x"51",
          9009 => x"3f",
          9010 => x"08",
          9011 => x"c8",
          9012 => x"75",
          9013 => x"66",
          9014 => x"34",
          9015 => x"82",
          9016 => x"84",
          9017 => x"06",
          9018 => x"80",
          9019 => x"2e",
          9020 => x"81",
          9021 => x"ff",
          9022 => x"82",
          9023 => x"54",
          9024 => x"08",
          9025 => x"53",
          9026 => x"08",
          9027 => x"ff",
          9028 => x"66",
          9029 => x"8b",
          9030 => x"53",
          9031 => x"51",
          9032 => x"3f",
          9033 => x"0b",
          9034 => x"78",
          9035 => x"da",
          9036 => x"c8",
          9037 => x"55",
          9038 => x"c8",
          9039 => x"0d",
          9040 => x"0d",
          9041 => x"88",
          9042 => x"05",
          9043 => x"fc",
          9044 => x"54",
          9045 => x"d2",
          9046 => x"d8",
          9047 => x"82",
          9048 => x"82",
          9049 => x"1a",
          9050 => x"82",
          9051 => x"80",
          9052 => x"8c",
          9053 => x"78",
          9054 => x"1a",
          9055 => x"2a",
          9056 => x"51",
          9057 => x"90",
          9058 => x"82",
          9059 => x"58",
          9060 => x"81",
          9061 => x"39",
          9062 => x"22",
          9063 => x"70",
          9064 => x"56",
          9065 => x"ab",
          9066 => x"14",
          9067 => x"30",
          9068 => x"9f",
          9069 => x"c8",
          9070 => x"19",
          9071 => x"5a",
          9072 => x"81",
          9073 => x"38",
          9074 => x"77",
          9075 => x"82",
          9076 => x"56",
          9077 => x"74",
          9078 => x"ff",
          9079 => x"81",
          9080 => x"55",
          9081 => x"75",
          9082 => x"82",
          9083 => x"c8",
          9084 => x"ff",
          9085 => x"d8",
          9086 => x"2e",
          9087 => x"82",
          9088 => x"8e",
          9089 => x"56",
          9090 => x"09",
          9091 => x"38",
          9092 => x"59",
          9093 => x"77",
          9094 => x"06",
          9095 => x"87",
          9096 => x"39",
          9097 => x"ba",
          9098 => x"55",
          9099 => x"2e",
          9100 => x"15",
          9101 => x"2e",
          9102 => x"83",
          9103 => x"75",
          9104 => x"7e",
          9105 => x"94",
          9106 => x"c8",
          9107 => x"d8",
          9108 => x"ce",
          9109 => x"16",
          9110 => x"56",
          9111 => x"38",
          9112 => x"19",
          9113 => x"90",
          9114 => x"7d",
          9115 => x"38",
          9116 => x"0c",
          9117 => x"0c",
          9118 => x"80",
          9119 => x"73",
          9120 => x"9c",
          9121 => x"05",
          9122 => x"57",
          9123 => x"26",
          9124 => x"7b",
          9125 => x"0c",
          9126 => x"81",
          9127 => x"84",
          9128 => x"54",
          9129 => x"c8",
          9130 => x"0d",
          9131 => x"0d",
          9132 => x"88",
          9133 => x"05",
          9134 => x"54",
          9135 => x"c5",
          9136 => x"56",
          9137 => x"d8",
          9138 => x"8b",
          9139 => x"d8",
          9140 => x"29",
          9141 => x"05",
          9142 => x"55",
          9143 => x"84",
          9144 => x"34",
          9145 => x"08",
          9146 => x"5f",
          9147 => x"51",
          9148 => x"3f",
          9149 => x"08",
          9150 => x"70",
          9151 => x"57",
          9152 => x"8b",
          9153 => x"82",
          9154 => x"06",
          9155 => x"56",
          9156 => x"38",
          9157 => x"05",
          9158 => x"7e",
          9159 => x"9e",
          9160 => x"c8",
          9161 => x"67",
          9162 => x"2e",
          9163 => x"82",
          9164 => x"8b",
          9165 => x"75",
          9166 => x"80",
          9167 => x"81",
          9168 => x"2e",
          9169 => x"80",
          9170 => x"38",
          9171 => x"0a",
          9172 => x"ff",
          9173 => x"55",
          9174 => x"86",
          9175 => x"8a",
          9176 => x"89",
          9177 => x"2a",
          9178 => x"77",
          9179 => x"59",
          9180 => x"81",
          9181 => x"70",
          9182 => x"07",
          9183 => x"56",
          9184 => x"38",
          9185 => x"05",
          9186 => x"7e",
          9187 => x"ae",
          9188 => x"82",
          9189 => x"8a",
          9190 => x"83",
          9191 => x"06",
          9192 => x"08",
          9193 => x"74",
          9194 => x"41",
          9195 => x"56",
          9196 => x"8a",
          9197 => x"61",
          9198 => x"55",
          9199 => x"27",
          9200 => x"93",
          9201 => x"80",
          9202 => x"38",
          9203 => x"70",
          9204 => x"43",
          9205 => x"95",
          9206 => x"06",
          9207 => x"2e",
          9208 => x"77",
          9209 => x"74",
          9210 => x"83",
          9211 => x"06",
          9212 => x"82",
          9213 => x"2e",
          9214 => x"78",
          9215 => x"2e",
          9216 => x"80",
          9217 => x"ae",
          9218 => x"2a",
          9219 => x"82",
          9220 => x"56",
          9221 => x"2e",
          9222 => x"77",
          9223 => x"82",
          9224 => x"79",
          9225 => x"70",
          9226 => x"5a",
          9227 => x"86",
          9228 => x"27",
          9229 => x"52",
          9230 => x"a6",
          9231 => x"d8",
          9232 => x"29",
          9233 => x"70",
          9234 => x"55",
          9235 => x"0b",
          9236 => x"08",
          9237 => x"05",
          9238 => x"ff",
          9239 => x"27",
          9240 => x"88",
          9241 => x"ae",
          9242 => x"2a",
          9243 => x"82",
          9244 => x"56",
          9245 => x"2e",
          9246 => x"77",
          9247 => x"82",
          9248 => x"79",
          9249 => x"70",
          9250 => x"5a",
          9251 => x"86",
          9252 => x"27",
          9253 => x"52",
          9254 => x"a5",
          9255 => x"d8",
          9256 => x"84",
          9257 => x"d8",
          9258 => x"f5",
          9259 => x"81",
          9260 => x"c8",
          9261 => x"d8",
          9262 => x"71",
          9263 => x"83",
          9264 => x"5e",
          9265 => x"89",
          9266 => x"5c",
          9267 => x"1c",
          9268 => x"05",
          9269 => x"ff",
          9270 => x"70",
          9271 => x"31",
          9272 => x"57",
          9273 => x"83",
          9274 => x"06",
          9275 => x"1c",
          9276 => x"5c",
          9277 => x"1d",
          9278 => x"29",
          9279 => x"31",
          9280 => x"55",
          9281 => x"87",
          9282 => x"7c",
          9283 => x"7a",
          9284 => x"31",
          9285 => x"a4",
          9286 => x"d8",
          9287 => x"7d",
          9288 => x"81",
          9289 => x"82",
          9290 => x"83",
          9291 => x"80",
          9292 => x"87",
          9293 => x"81",
          9294 => x"fd",
          9295 => x"f8",
          9296 => x"2e",
          9297 => x"80",
          9298 => x"ff",
          9299 => x"d8",
          9300 => x"a0",
          9301 => x"38",
          9302 => x"74",
          9303 => x"86",
          9304 => x"fd",
          9305 => x"81",
          9306 => x"80",
          9307 => x"83",
          9308 => x"39",
          9309 => x"08",
          9310 => x"92",
          9311 => x"b8",
          9312 => x"59",
          9313 => x"27",
          9314 => x"86",
          9315 => x"55",
          9316 => x"09",
          9317 => x"38",
          9318 => x"f5",
          9319 => x"38",
          9320 => x"55",
          9321 => x"86",
          9322 => x"80",
          9323 => x"7a",
          9324 => x"e7",
          9325 => x"82",
          9326 => x"7a",
          9327 => x"b8",
          9328 => x"52",
          9329 => x"ff",
          9330 => x"79",
          9331 => x"7b",
          9332 => x"06",
          9333 => x"51",
          9334 => x"3f",
          9335 => x"1c",
          9336 => x"32",
          9337 => x"96",
          9338 => x"06",
          9339 => x"91",
          9340 => x"8f",
          9341 => x"55",
          9342 => x"ff",
          9343 => x"74",
          9344 => x"06",
          9345 => x"51",
          9346 => x"3f",
          9347 => x"52",
          9348 => x"ff",
          9349 => x"f8",
          9350 => x"34",
          9351 => x"1b",
          9352 => x"87",
          9353 => x"52",
          9354 => x"ff",
          9355 => x"60",
          9356 => x"51",
          9357 => x"3f",
          9358 => x"09",
          9359 => x"cb",
          9360 => x"b2",
          9361 => x"c3",
          9362 => x"8e",
          9363 => x"52",
          9364 => x"ff",
          9365 => x"82",
          9366 => x"51",
          9367 => x"3f",
          9368 => x"1b",
          9369 => x"c3",
          9370 => x"b2",
          9371 => x"8e",
          9372 => x"80",
          9373 => x"1c",
          9374 => x"80",
          9375 => x"93",
          9376 => x"98",
          9377 => x"1b",
          9378 => x"82",
          9379 => x"52",
          9380 => x"ff",
          9381 => x"7c",
          9382 => x"06",
          9383 => x"51",
          9384 => x"3f",
          9385 => x"a4",
          9386 => x"0b",
          9387 => x"93",
          9388 => x"ac",
          9389 => x"51",
          9390 => x"3f",
          9391 => x"52",
          9392 => x"70",
          9393 => x"8d",
          9394 => x"54",
          9395 => x"52",
          9396 => x"8a",
          9397 => x"56",
          9398 => x"08",
          9399 => x"7d",
          9400 => x"81",
          9401 => x"38",
          9402 => x"86",
          9403 => x"52",
          9404 => x"89",
          9405 => x"80",
          9406 => x"7a",
          9407 => x"9b",
          9408 => x"85",
          9409 => x"7a",
          9410 => x"bd",
          9411 => x"85",
          9412 => x"83",
          9413 => x"ff",
          9414 => x"ff",
          9415 => x"e8",
          9416 => x"8d",
          9417 => x"52",
          9418 => x"51",
          9419 => x"3f",
          9420 => x"52",
          9421 => x"8c",
          9422 => x"54",
          9423 => x"53",
          9424 => x"51",
          9425 => x"3f",
          9426 => x"16",
          9427 => x"7e",
          9428 => x"86",
          9429 => x"80",
          9430 => x"ff",
          9431 => x"7f",
          9432 => x"7d",
          9433 => x"81",
          9434 => x"f8",
          9435 => x"ff",
          9436 => x"ff",
          9437 => x"51",
          9438 => x"3f",
          9439 => x"88",
          9440 => x"39",
          9441 => x"f8",
          9442 => x"2e",
          9443 => x"55",
          9444 => x"51",
          9445 => x"3f",
          9446 => x"57",
          9447 => x"83",
          9448 => x"76",
          9449 => x"7a",
          9450 => x"ff",
          9451 => x"82",
          9452 => x"82",
          9453 => x"80",
          9454 => x"c8",
          9455 => x"51",
          9456 => x"3f",
          9457 => x"78",
          9458 => x"74",
          9459 => x"18",
          9460 => x"2e",
          9461 => x"79",
          9462 => x"2e",
          9463 => x"55",
          9464 => x"62",
          9465 => x"74",
          9466 => x"75",
          9467 => x"7e",
          9468 => x"e6",
          9469 => x"c8",
          9470 => x"38",
          9471 => x"78",
          9472 => x"74",
          9473 => x"56",
          9474 => x"93",
          9475 => x"66",
          9476 => x"26",
          9477 => x"56",
          9478 => x"83",
          9479 => x"64",
          9480 => x"77",
          9481 => x"84",
          9482 => x"52",
          9483 => x"8b",
          9484 => x"d4",
          9485 => x"51",
          9486 => x"3f",
          9487 => x"55",
          9488 => x"81",
          9489 => x"34",
          9490 => x"16",
          9491 => x"16",
          9492 => x"16",
          9493 => x"05",
          9494 => x"c1",
          9495 => x"fe",
          9496 => x"fe",
          9497 => x"34",
          9498 => x"08",
          9499 => x"07",
          9500 => x"16",
          9501 => x"c8",
          9502 => x"34",
          9503 => x"c6",
          9504 => x"8a",
          9505 => x"52",
          9506 => x"51",
          9507 => x"3f",
          9508 => x"53",
          9509 => x"51",
          9510 => x"3f",
          9511 => x"d8",
          9512 => x"38",
          9513 => x"52",
          9514 => x"88",
          9515 => x"56",
          9516 => x"08",
          9517 => x"39",
          9518 => x"39",
          9519 => x"39",
          9520 => x"08",
          9521 => x"d8",
          9522 => x"3d",
          9523 => x"3d",
          9524 => x"5b",
          9525 => x"60",
          9526 => x"57",
          9527 => x"25",
          9528 => x"3d",
          9529 => x"55",
          9530 => x"15",
          9531 => x"c9",
          9532 => x"81",
          9533 => x"06",
          9534 => x"3d",
          9535 => x"8d",
          9536 => x"74",
          9537 => x"05",
          9538 => x"17",
          9539 => x"2e",
          9540 => x"c9",
          9541 => x"34",
          9542 => x"83",
          9543 => x"74",
          9544 => x"0c",
          9545 => x"04",
          9546 => x"7b",
          9547 => x"b3",
          9548 => x"57",
          9549 => x"09",
          9550 => x"38",
          9551 => x"51",
          9552 => x"17",
          9553 => x"76",
          9554 => x"88",
          9555 => x"17",
          9556 => x"59",
          9557 => x"81",
          9558 => x"76",
          9559 => x"8b",
          9560 => x"54",
          9561 => x"17",
          9562 => x"51",
          9563 => x"79",
          9564 => x"30",
          9565 => x"9f",
          9566 => x"53",
          9567 => x"75",
          9568 => x"81",
          9569 => x"0c",
          9570 => x"04",
          9571 => x"79",
          9572 => x"56",
          9573 => x"24",
          9574 => x"3d",
          9575 => x"74",
          9576 => x"52",
          9577 => x"cb",
          9578 => x"d8",
          9579 => x"38",
          9580 => x"78",
          9581 => x"06",
          9582 => x"16",
          9583 => x"39",
          9584 => x"82",
          9585 => x"89",
          9586 => x"fd",
          9587 => x"54",
          9588 => x"80",
          9589 => x"ff",
          9590 => x"76",
          9591 => x"3d",
          9592 => x"3d",
          9593 => x"e3",
          9594 => x"53",
          9595 => x"53",
          9596 => x"3f",
          9597 => x"51",
          9598 => x"72",
          9599 => x"3f",
          9600 => x"04",
          9601 => x"75",
          9602 => x"9a",
          9603 => x"53",
          9604 => x"80",
          9605 => x"38",
          9606 => x"ff",
          9607 => x"c3",
          9608 => x"ff",
          9609 => x"73",
          9610 => x"09",
          9611 => x"38",
          9612 => x"af",
          9613 => x"94",
          9614 => x"71",
          9615 => x"81",
          9616 => x"ff",
          9617 => x"51",
          9618 => x"26",
          9619 => x"10",
          9620 => x"05",
          9621 => x"51",
          9622 => x"80",
          9623 => x"ff",
          9624 => x"71",
          9625 => x"0c",
          9626 => x"04",
          9627 => x"02",
          9628 => x"02",
          9629 => x"05",
          9630 => x"80",
          9631 => x"ff",
          9632 => x"70",
          9633 => x"71",
          9634 => x"09",
          9635 => x"38",
          9636 => x"26",
          9637 => x"10",
          9638 => x"05",
          9639 => x"51",
          9640 => x"c8",
          9641 => x"0d",
          9642 => x"0d",
          9643 => x"83",
          9644 => x"81",
          9645 => x"83",
          9646 => x"82",
          9647 => x"52",
          9648 => x"27",
          9649 => x"d2",
          9650 => x"70",
          9651 => x"22",
          9652 => x"80",
          9653 => x"26",
          9654 => x"55",
          9655 => x"38",
          9656 => x"05",
          9657 => x"88",
          9658 => x"ff",
          9659 => x"54",
          9660 => x"71",
          9661 => x"d7",
          9662 => x"26",
          9663 => x"73",
          9664 => x"b0",
          9665 => x"70",
          9666 => x"75",
          9667 => x"11",
          9668 => x"51",
          9669 => x"39",
          9670 => x"81",
          9671 => x"31",
          9672 => x"39",
          9673 => x"9f",
          9674 => x"51",
          9675 => x"12",
          9676 => x"e6",
          9677 => x"39",
          9678 => x"8b",
          9679 => x"12",
          9680 => x"c7",
          9681 => x"70",
          9682 => x"06",
          9683 => x"73",
          9684 => x"72",
          9685 => x"fe",
          9686 => x"51",
          9687 => x"c8",
          9688 => x"0d",
          9689 => x"ff",
          9690 => x"00",
          9691 => x"ff",
          9692 => x"ff",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"00",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"69",
          9839 => x"00",
          9840 => x"69",
          9841 => x"6c",
          9842 => x"69",
          9843 => x"00",
          9844 => x"6c",
          9845 => x"00",
          9846 => x"65",
          9847 => x"00",
          9848 => x"63",
          9849 => x"72",
          9850 => x"63",
          9851 => x"00",
          9852 => x"64",
          9853 => x"00",
          9854 => x"64",
          9855 => x"00",
          9856 => x"65",
          9857 => x"65",
          9858 => x"65",
          9859 => x"69",
          9860 => x"69",
          9861 => x"66",
          9862 => x"66",
          9863 => x"61",
          9864 => x"00",
          9865 => x"6d",
          9866 => x"65",
          9867 => x"72",
          9868 => x"65",
          9869 => x"00",
          9870 => x"6e",
          9871 => x"00",
          9872 => x"65",
          9873 => x"00",
          9874 => x"62",
          9875 => x"63",
          9876 => x"62",
          9877 => x"63",
          9878 => x"69",
          9879 => x"00",
          9880 => x"64",
          9881 => x"69",
          9882 => x"45",
          9883 => x"72",
          9884 => x"6e",
          9885 => x"6e",
          9886 => x"65",
          9887 => x"72",
          9888 => x"69",
          9889 => x"6e",
          9890 => x"72",
          9891 => x"79",
          9892 => x"6f",
          9893 => x"6c",
          9894 => x"6f",
          9895 => x"2e",
          9896 => x"6f",
          9897 => x"74",
          9898 => x"6f",
          9899 => x"2e",
          9900 => x"6e",
          9901 => x"69",
          9902 => x"69",
          9903 => x"61",
          9904 => x"00",
          9905 => x"63",
          9906 => x"73",
          9907 => x"6e",
          9908 => x"2e",
          9909 => x"69",
          9910 => x"61",
          9911 => x"61",
          9912 => x"65",
          9913 => x"74",
          9914 => x"00",
          9915 => x"69",
          9916 => x"68",
          9917 => x"6c",
          9918 => x"6e",
          9919 => x"69",
          9920 => x"00",
          9921 => x"44",
          9922 => x"20",
          9923 => x"74",
          9924 => x"72",
          9925 => x"63",
          9926 => x"2e",
          9927 => x"72",
          9928 => x"20",
          9929 => x"62",
          9930 => x"69",
          9931 => x"6e",
          9932 => x"69",
          9933 => x"00",
          9934 => x"69",
          9935 => x"6e",
          9936 => x"65",
          9937 => x"6c",
          9938 => x"00",
          9939 => x"6f",
          9940 => x"6d",
          9941 => x"69",
          9942 => x"20",
          9943 => x"65",
          9944 => x"74",
          9945 => x"66",
          9946 => x"64",
          9947 => x"20",
          9948 => x"6b",
          9949 => x"6f",
          9950 => x"74",
          9951 => x"6f",
          9952 => x"64",
          9953 => x"69",
          9954 => x"75",
          9955 => x"6f",
          9956 => x"61",
          9957 => x"6e",
          9958 => x"6e",
          9959 => x"6c",
          9960 => x"00",
          9961 => x"69",
          9962 => x"69",
          9963 => x"6f",
          9964 => x"64",
          9965 => x"6e",
          9966 => x"66",
          9967 => x"65",
          9968 => x"6d",
          9969 => x"72",
          9970 => x"00",
          9971 => x"6f",
          9972 => x"61",
          9973 => x"6f",
          9974 => x"20",
          9975 => x"65",
          9976 => x"00",
          9977 => x"61",
          9978 => x"65",
          9979 => x"73",
          9980 => x"63",
          9981 => x"65",
          9982 => x"00",
          9983 => x"75",
          9984 => x"73",
          9985 => x"00",
          9986 => x"6e",
          9987 => x"77",
          9988 => x"72",
          9989 => x"2e",
          9990 => x"25",
          9991 => x"62",
          9992 => x"73",
          9993 => x"20",
          9994 => x"25",
          9995 => x"62",
          9996 => x"73",
          9997 => x"63",
          9998 => x"00",
          9999 => x"65",
         10000 => x"00",
         10001 => x"3d",
         10002 => x"6c",
         10003 => x"31",
         10004 => x"38",
         10005 => x"20",
         10006 => x"30",
         10007 => x"2c",
         10008 => x"4f",
         10009 => x"30",
         10010 => x"20",
         10011 => x"6c",
         10012 => x"30",
         10013 => x"0a",
         10014 => x"30",
         10015 => x"00",
         10016 => x"20",
         10017 => x"30",
         10018 => x"00",
         10019 => x"20",
         10020 => x"20",
         10021 => x"00",
         10022 => x"30",
         10023 => x"00",
         10024 => x"20",
         10025 => x"7c",
         10026 => x"00",
         10027 => x"50",
         10028 => x"00",
         10029 => x"2a",
         10030 => x"73",
         10031 => x"00",
         10032 => x"32",
         10033 => x"2f",
         10034 => x"30",
         10035 => x"31",
         10036 => x"00",
         10037 => x"5a",
         10038 => x"20",
         10039 => x"20",
         10040 => x"78",
         10041 => x"73",
         10042 => x"20",
         10043 => x"0a",
         10044 => x"50",
         10045 => x"20",
         10046 => x"65",
         10047 => x"70",
         10048 => x"61",
         10049 => x"65",
         10050 => x"69",
         10051 => x"20",
         10052 => x"65",
         10053 => x"70",
         10054 => x"53",
         10055 => x"6e",
         10056 => x"72",
         10057 => x"00",
         10058 => x"4f",
         10059 => x"20",
         10060 => x"69",
         10061 => x"72",
         10062 => x"74",
         10063 => x"4f",
         10064 => x"20",
         10065 => x"69",
         10066 => x"72",
         10067 => x"74",
         10068 => x"41",
         10069 => x"20",
         10070 => x"69",
         10071 => x"72",
         10072 => x"74",
         10073 => x"41",
         10074 => x"20",
         10075 => x"69",
         10076 => x"72",
         10077 => x"74",
         10078 => x"41",
         10079 => x"20",
         10080 => x"69",
         10081 => x"72",
         10082 => x"74",
         10083 => x"41",
         10084 => x"20",
         10085 => x"69",
         10086 => x"72",
         10087 => x"74",
         10088 => x"65",
         10089 => x"6e",
         10090 => x"70",
         10091 => x"6d",
         10092 => x"2e",
         10093 => x"6e",
         10094 => x"69",
         10095 => x"74",
         10096 => x"72",
         10097 => x"00",
         10098 => x"75",
         10099 => x"78",
         10100 => x"62",
         10101 => x"00",
         10102 => x"70",
         10103 => x"2e",
         10104 => x"00",
         10105 => x"3a",
         10106 => x"61",
         10107 => x"64",
         10108 => x"20",
         10109 => x"74",
         10110 => x"69",
         10111 => x"73",
         10112 => x"61",
         10113 => x"30",
         10114 => x"6c",
         10115 => x"65",
         10116 => x"69",
         10117 => x"61",
         10118 => x"6c",
         10119 => x"00",
         10120 => x"20",
         10121 => x"61",
         10122 => x"69",
         10123 => x"69",
         10124 => x"00",
         10125 => x"6e",
         10126 => x"61",
         10127 => x"65",
         10128 => x"00",
         10129 => x"61",
         10130 => x"64",
         10131 => x"20",
         10132 => x"74",
         10133 => x"69",
         10134 => x"00",
         10135 => x"63",
         10136 => x"0a",
         10137 => x"75",
         10138 => x"6c",
         10139 => x"69",
         10140 => x"2e",
         10141 => x"00",
         10142 => x"6f",
         10143 => x"6e",
         10144 => x"2e",
         10145 => x"6f",
         10146 => x"72",
         10147 => x"2e",
         10148 => x"00",
         10149 => x"30",
         10150 => x"28",
         10151 => x"78",
         10152 => x"25",
         10153 => x"78",
         10154 => x"38",
         10155 => x"00",
         10156 => x"75",
         10157 => x"4d",
         10158 => x"72",
         10159 => x"43",
         10160 => x"6c",
         10161 => x"2e",
         10162 => x"30",
         10163 => x"20",
         10164 => x"58",
         10165 => x"3f",
         10166 => x"30",
         10167 => x"20",
         10168 => x"58",
         10169 => x"30",
         10170 => x"20",
         10171 => x"6c",
         10172 => x"00",
         10173 => x"69",
         10174 => x"6c",
         10175 => x"20",
         10176 => x"65",
         10177 => x"70",
         10178 => x"00",
         10179 => x"6e",
         10180 => x"69",
         10181 => x"69",
         10182 => x"72",
         10183 => x"74",
         10184 => x"69",
         10185 => x"6c",
         10186 => x"75",
         10187 => x"20",
         10188 => x"6f",
         10189 => x"6e",
         10190 => x"69",
         10191 => x"75",
         10192 => x"20",
         10193 => x"6f",
         10194 => x"78",
         10195 => x"74",
         10196 => x"20",
         10197 => x"65",
         10198 => x"25",
         10199 => x"78",
         10200 => x"2e",
         10201 => x"61",
         10202 => x"6e",
         10203 => x"6f",
         10204 => x"40",
         10205 => x"38",
         10206 => x"2e",
         10207 => x"00",
         10208 => x"61",
         10209 => x"72",
         10210 => x"72",
         10211 => x"20",
         10212 => x"65",
         10213 => x"64",
         10214 => x"00",
         10215 => x"65",
         10216 => x"72",
         10217 => x"67",
         10218 => x"70",
         10219 => x"61",
         10220 => x"6e",
         10221 => x"00",
         10222 => x"6f",
         10223 => x"72",
         10224 => x"6f",
         10225 => x"67",
         10226 => x"00",
         10227 => x"50",
         10228 => x"69",
         10229 => x"64",
         10230 => x"73",
         10231 => x"2e",
         10232 => x"00",
         10233 => x"64",
         10234 => x"73",
         10235 => x"00",
         10236 => x"64",
         10237 => x"73",
         10238 => x"61",
         10239 => x"6f",
         10240 => x"6e",
         10241 => x"00",
         10242 => x"75",
         10243 => x"6e",
         10244 => x"2e",
         10245 => x"6e",
         10246 => x"69",
         10247 => x"69",
         10248 => x"72",
         10249 => x"74",
         10250 => x"2e",
         10251 => x"64",
         10252 => x"2f",
         10253 => x"25",
         10254 => x"64",
         10255 => x"2e",
         10256 => x"64",
         10257 => x"6f",
         10258 => x"6f",
         10259 => x"67",
         10260 => x"74",
         10261 => x"00",
         10262 => x"28",
         10263 => x"6d",
         10264 => x"43",
         10265 => x"6e",
         10266 => x"29",
         10267 => x"0a",
         10268 => x"69",
         10269 => x"20",
         10270 => x"6c",
         10271 => x"6e",
         10272 => x"3a",
         10273 => x"20",
         10274 => x"42",
         10275 => x"52",
         10276 => x"20",
         10277 => x"38",
         10278 => x"30",
         10279 => x"2e",
         10280 => x"20",
         10281 => x"44",
         10282 => x"20",
         10283 => x"20",
         10284 => x"38",
         10285 => x"30",
         10286 => x"2e",
         10287 => x"20",
         10288 => x"4e",
         10289 => x"42",
         10290 => x"20",
         10291 => x"38",
         10292 => x"30",
         10293 => x"2e",
         10294 => x"20",
         10295 => x"52",
         10296 => x"20",
         10297 => x"20",
         10298 => x"38",
         10299 => x"30",
         10300 => x"2e",
         10301 => x"20",
         10302 => x"41",
         10303 => x"20",
         10304 => x"20",
         10305 => x"38",
         10306 => x"30",
         10307 => x"2e",
         10308 => x"20",
         10309 => x"44",
         10310 => x"52",
         10311 => x"20",
         10312 => x"76",
         10313 => x"73",
         10314 => x"30",
         10315 => x"2e",
         10316 => x"20",
         10317 => x"49",
         10318 => x"31",
         10319 => x"20",
         10320 => x"6d",
         10321 => x"20",
         10322 => x"30",
         10323 => x"2e",
         10324 => x"20",
         10325 => x"4e",
         10326 => x"43",
         10327 => x"20",
         10328 => x"61",
         10329 => x"6c",
         10330 => x"30",
         10331 => x"2e",
         10332 => x"20",
         10333 => x"49",
         10334 => x"4f",
         10335 => x"42",
         10336 => x"00",
         10337 => x"20",
         10338 => x"42",
         10339 => x"43",
         10340 => x"20",
         10341 => x"4f",
         10342 => x"00",
         10343 => x"20",
         10344 => x"53",
         10345 => x"20",
         10346 => x"50",
         10347 => x"64",
         10348 => x"73",
         10349 => x"3a",
         10350 => x"20",
         10351 => x"50",
         10352 => x"65",
         10353 => x"20",
         10354 => x"74",
         10355 => x"41",
         10356 => x"65",
         10357 => x"3d",
         10358 => x"38",
         10359 => x"00",
         10360 => x"20",
         10361 => x"50",
         10362 => x"65",
         10363 => x"79",
         10364 => x"61",
         10365 => x"41",
         10366 => x"65",
         10367 => x"3d",
         10368 => x"38",
         10369 => x"00",
         10370 => x"20",
         10371 => x"74",
         10372 => x"20",
         10373 => x"72",
         10374 => x"64",
         10375 => x"73",
         10376 => x"20",
         10377 => x"3d",
         10378 => x"38",
         10379 => x"00",
         10380 => x"69",
         10381 => x"00",
         10382 => x"20",
         10383 => x"50",
         10384 => x"64",
         10385 => x"20",
         10386 => x"20",
         10387 => x"20",
         10388 => x"20",
         10389 => x"3d",
         10390 => x"34",
         10391 => x"00",
         10392 => x"20",
         10393 => x"79",
         10394 => x"6d",
         10395 => x"6f",
         10396 => x"46",
         10397 => x"20",
         10398 => x"20",
         10399 => x"3d",
         10400 => x"2e",
         10401 => x"64",
         10402 => x"0a",
         10403 => x"20",
         10404 => x"44",
         10405 => x"20",
         10406 => x"63",
         10407 => x"72",
         10408 => x"20",
         10409 => x"20",
         10410 => x"3d",
         10411 => x"2e",
         10412 => x"64",
         10413 => x"0a",
         10414 => x"20",
         10415 => x"69",
         10416 => x"6f",
         10417 => x"53",
         10418 => x"4d",
         10419 => x"6f",
         10420 => x"46",
         10421 => x"3d",
         10422 => x"2e",
         10423 => x"64",
         10424 => x"0a",
         10425 => x"6d",
         10426 => x"00",
         10427 => x"65",
         10428 => x"6d",
         10429 => x"6c",
         10430 => x"00",
         10431 => x"56",
         10432 => x"56",
         10433 => x"00",
         10434 => x"6e",
         10435 => x"77",
         10436 => x"00",
         10437 => x"00",
         10438 => x"00",
         10439 => x"00",
         10440 => x"00",
         10441 => x"00",
         10442 => x"00",
         10443 => x"00",
         10444 => x"00",
         10445 => x"00",
         10446 => x"00",
         10447 => x"00",
         10448 => x"00",
         10449 => x"00",
         10450 => x"00",
         10451 => x"00",
         10452 => x"00",
         10453 => x"00",
         10454 => x"00",
         10455 => x"00",
         10456 => x"00",
         10457 => x"00",
         10458 => x"00",
         10459 => x"00",
         10460 => x"00",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"00",
         10465 => x"00",
         10466 => x"00",
         10467 => x"00",
         10468 => x"00",
         10469 => x"00",
         10470 => x"00",
         10471 => x"00",
         10472 => x"00",
         10473 => x"00",
         10474 => x"00",
         10475 => x"00",
         10476 => x"00",
         10477 => x"00",
         10478 => x"00",
         10479 => x"00",
         10480 => x"00",
         10481 => x"00",
         10482 => x"00",
         10483 => x"00",
         10484 => x"00",
         10485 => x"00",
         10486 => x"00",
         10487 => x"00",
         10488 => x"00",
         10489 => x"00",
         10490 => x"00",
         10491 => x"00",
         10492 => x"00",
         10493 => x"00",
         10494 => x"00",
         10495 => x"00",
         10496 => x"00",
         10497 => x"00",
         10498 => x"00",
         10499 => x"00",
         10500 => x"00",
         10501 => x"00",
         10502 => x"5b",
         10503 => x"5b",
         10504 => x"5b",
         10505 => x"5b",
         10506 => x"5b",
         10507 => x"5b",
         10508 => x"5b",
         10509 => x"30",
         10510 => x"5b",
         10511 => x"5b",
         10512 => x"5b",
         10513 => x"00",
         10514 => x"00",
         10515 => x"00",
         10516 => x"00",
         10517 => x"00",
         10518 => x"00",
         10519 => x"00",
         10520 => x"00",
         10521 => x"00",
         10522 => x"00",
         10523 => x"00",
         10524 => x"69",
         10525 => x"72",
         10526 => x"69",
         10527 => x"00",
         10528 => x"00",
         10529 => x"30",
         10530 => x"20",
         10531 => x"0a",
         10532 => x"61",
         10533 => x"64",
         10534 => x"20",
         10535 => x"65",
         10536 => x"68",
         10537 => x"69",
         10538 => x"72",
         10539 => x"69",
         10540 => x"74",
         10541 => x"4f",
         10542 => x"00",
         10543 => x"61",
         10544 => x"74",
         10545 => x"65",
         10546 => x"72",
         10547 => x"65",
         10548 => x"73",
         10549 => x"79",
         10550 => x"6c",
         10551 => x"64",
         10552 => x"62",
         10553 => x"67",
         10554 => x"44",
         10555 => x"2a",
         10556 => x"3f",
         10557 => x"00",
         10558 => x"2c",
         10559 => x"5d",
         10560 => x"41",
         10561 => x"41",
         10562 => x"00",
         10563 => x"fe",
         10564 => x"44",
         10565 => x"2e",
         10566 => x"4f",
         10567 => x"4d",
         10568 => x"20",
         10569 => x"54",
         10570 => x"20",
         10571 => x"4f",
         10572 => x"4d",
         10573 => x"20",
         10574 => x"54",
         10575 => x"20",
         10576 => x"00",
         10577 => x"00",
         10578 => x"00",
         10579 => x"00",
         10580 => x"03",
         10581 => x"0e",
         10582 => x"16",
         10583 => x"00",
         10584 => x"9a",
         10585 => x"41",
         10586 => x"45",
         10587 => x"49",
         10588 => x"92",
         10589 => x"4f",
         10590 => x"99",
         10591 => x"9d",
         10592 => x"49",
         10593 => x"a5",
         10594 => x"a9",
         10595 => x"ad",
         10596 => x"b1",
         10597 => x"b5",
         10598 => x"b9",
         10599 => x"bd",
         10600 => x"c1",
         10601 => x"c5",
         10602 => x"c9",
         10603 => x"cd",
         10604 => x"d1",
         10605 => x"d5",
         10606 => x"d9",
         10607 => x"dd",
         10608 => x"e1",
         10609 => x"e5",
         10610 => x"e9",
         10611 => x"ed",
         10612 => x"f1",
         10613 => x"f5",
         10614 => x"f9",
         10615 => x"fd",
         10616 => x"2e",
         10617 => x"5b",
         10618 => x"22",
         10619 => x"3e",
         10620 => x"00",
         10621 => x"01",
         10622 => x"10",
         10623 => x"00",
         10624 => x"00",
         10625 => x"01",
         10626 => x"04",
         10627 => x"10",
         10628 => x"00",
         10629 => x"c7",
         10630 => x"e9",
         10631 => x"e4",
         10632 => x"e5",
         10633 => x"ea",
         10634 => x"e8",
         10635 => x"ee",
         10636 => x"c4",
         10637 => x"c9",
         10638 => x"c6",
         10639 => x"f6",
         10640 => x"fb",
         10641 => x"ff",
         10642 => x"dc",
         10643 => x"a3",
         10644 => x"a7",
         10645 => x"e1",
         10646 => x"f3",
         10647 => x"f1",
         10648 => x"aa",
         10649 => x"bf",
         10650 => x"ac",
         10651 => x"bc",
         10652 => x"ab",
         10653 => x"91",
         10654 => x"93",
         10655 => x"24",
         10656 => x"62",
         10657 => x"55",
         10658 => x"51",
         10659 => x"5d",
         10660 => x"5b",
         10661 => x"14",
         10662 => x"2c",
         10663 => x"00",
         10664 => x"5e",
         10665 => x"5a",
         10666 => x"69",
         10667 => x"60",
         10668 => x"6c",
         10669 => x"68",
         10670 => x"65",
         10671 => x"58",
         10672 => x"53",
         10673 => x"6a",
         10674 => x"0c",
         10675 => x"84",
         10676 => x"90",
         10677 => x"b1",
         10678 => x"93",
         10679 => x"a3",
         10680 => x"b5",
         10681 => x"a6",
         10682 => x"a9",
         10683 => x"1e",
         10684 => x"b5",
         10685 => x"61",
         10686 => x"65",
         10687 => x"20",
         10688 => x"f7",
         10689 => x"b0",
         10690 => x"b7",
         10691 => x"7f",
         10692 => x"a0",
         10693 => x"61",
         10694 => x"e0",
         10695 => x"f8",
         10696 => x"ff",
         10697 => x"78",
         10698 => x"30",
         10699 => x"06",
         10700 => x"10",
         10701 => x"2e",
         10702 => x"06",
         10703 => x"4d",
         10704 => x"81",
         10705 => x"82",
         10706 => x"84",
         10707 => x"87",
         10708 => x"89",
         10709 => x"8b",
         10710 => x"8d",
         10711 => x"8f",
         10712 => x"91",
         10713 => x"93",
         10714 => x"f6",
         10715 => x"97",
         10716 => x"98",
         10717 => x"9b",
         10718 => x"9d",
         10719 => x"9f",
         10720 => x"a0",
         10721 => x"a2",
         10722 => x"a4",
         10723 => x"a7",
         10724 => x"a9",
         10725 => x"ab",
         10726 => x"ac",
         10727 => x"af",
         10728 => x"b1",
         10729 => x"b3",
         10730 => x"b5",
         10731 => x"b7",
         10732 => x"b8",
         10733 => x"bb",
         10734 => x"bc",
         10735 => x"f7",
         10736 => x"c1",
         10737 => x"c3",
         10738 => x"c5",
         10739 => x"c7",
         10740 => x"c7",
         10741 => x"cb",
         10742 => x"cd",
         10743 => x"dd",
         10744 => x"8e",
         10745 => x"12",
         10746 => x"03",
         10747 => x"f4",
         10748 => x"f8",
         10749 => x"22",
         10750 => x"3a",
         10751 => x"65",
         10752 => x"3b",
         10753 => x"66",
         10754 => x"40",
         10755 => x"41",
         10756 => x"0a",
         10757 => x"40",
         10758 => x"86",
         10759 => x"89",
         10760 => x"58",
         10761 => x"5a",
         10762 => x"5c",
         10763 => x"5e",
         10764 => x"93",
         10765 => x"62",
         10766 => x"64",
         10767 => x"66",
         10768 => x"97",
         10769 => x"6a",
         10770 => x"6c",
         10771 => x"6e",
         10772 => x"70",
         10773 => x"9d",
         10774 => x"74",
         10775 => x"76",
         10776 => x"78",
         10777 => x"7a",
         10778 => x"7c",
         10779 => x"7e",
         10780 => x"a6",
         10781 => x"82",
         10782 => x"84",
         10783 => x"86",
         10784 => x"ae",
         10785 => x"b1",
         10786 => x"45",
         10787 => x"8e",
         10788 => x"90",
         10789 => x"b7",
         10790 => x"03",
         10791 => x"fe",
         10792 => x"ac",
         10793 => x"86",
         10794 => x"89",
         10795 => x"b1",
         10796 => x"c2",
         10797 => x"a3",
         10798 => x"c4",
         10799 => x"cc",
         10800 => x"8c",
         10801 => x"8f",
         10802 => x"18",
         10803 => x"0a",
         10804 => x"f3",
         10805 => x"f5",
         10806 => x"f7",
         10807 => x"f9",
         10808 => x"fa",
         10809 => x"20",
         10810 => x"10",
         10811 => x"22",
         10812 => x"36",
         10813 => x"0e",
         10814 => x"01",
         10815 => x"d0",
         10816 => x"61",
         10817 => x"00",
         10818 => x"7d",
         10819 => x"63",
         10820 => x"96",
         10821 => x"5a",
         10822 => x"08",
         10823 => x"06",
         10824 => x"08",
         10825 => x"08",
         10826 => x"06",
         10827 => x"07",
         10828 => x"52",
         10829 => x"54",
         10830 => x"56",
         10831 => x"60",
         10832 => x"70",
         10833 => x"ba",
         10834 => x"c8",
         10835 => x"ca",
         10836 => x"da",
         10837 => x"f8",
         10838 => x"ea",
         10839 => x"fa",
         10840 => x"80",
         10841 => x"90",
         10842 => x"a0",
         10843 => x"b0",
         10844 => x"b8",
         10845 => x"b2",
         10846 => x"cc",
         10847 => x"c3",
         10848 => x"02",
         10849 => x"02",
         10850 => x"01",
         10851 => x"f3",
         10852 => x"fc",
         10853 => x"01",
         10854 => x"70",
         10855 => x"84",
         10856 => x"83",
         10857 => x"1a",
         10858 => x"2f",
         10859 => x"02",
         10860 => x"06",
         10861 => x"02",
         10862 => x"64",
         10863 => x"26",
         10864 => x"1a",
         10865 => x"00",
         10866 => x"00",
         10867 => x"02",
         10868 => x"00",
         10869 => x"00",
         10870 => x"00",
         10871 => x"04",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"14",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"2b",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"30",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"3c",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"3d",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"3f",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"40",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"41",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"42",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"43",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"50",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"51",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"54",
         10924 => x"00",
         10925 => x"00",
         10926 => x"00",
         10927 => x"55",
         10928 => x"00",
         10929 => x"00",
         10930 => x"00",
         10931 => x"79",
         10932 => x"00",
         10933 => x"00",
         10934 => x"00",
         10935 => x"78",
         10936 => x"00",
         10937 => x"00",
         10938 => x"00",
         10939 => x"82",
         10940 => x"00",
         10941 => x"00",
         10942 => x"00",
         10943 => x"83",
         10944 => x"00",
         10945 => x"00",
         10946 => x"00",
         10947 => x"85",
         10948 => x"00",
         10949 => x"00",
         10950 => x"00",
         10951 => x"87",
         10952 => x"00",
         10953 => x"00",
         10954 => x"00",
         10955 => x"8c",
         10956 => x"00",
         10957 => x"00",
         10958 => x"00",
         10959 => x"8d",
         10960 => x"00",
         10961 => x"00",
         10962 => x"00",
         10963 => x"8e",
         10964 => x"00",
         10965 => x"00",
         10966 => x"00",
         10967 => x"8f",
         10968 => x"00",
         10969 => x"00",
         10970 => x"00",
         10971 => x"00",
         10972 => x"00",
         10973 => x"00",
         10974 => x"00",
         10975 => x"01",
         10976 => x"00",
         10977 => x"01",
         10978 => x"81",
         10979 => x"00",
         10980 => x"7f",
         10981 => x"00",
         10982 => x"00",
         10983 => x"00",
         10984 => x"00",
         10985 => x"f5",
         10986 => x"f5",
         10987 => x"f5",
         10988 => x"00",
         10989 => x"01",
         10990 => x"01",
         10991 => x"01",
         10992 => x"00",
         10993 => x"00",
         10994 => x"00",
         10995 => x"00",
         10996 => x"00",
         10997 => x"00",
         10998 => x"00",
         10999 => x"00",
         11000 => x"00",
         11001 => x"00",
         11002 => x"00",
         11003 => x"00",
         11004 => x"00",
         11005 => x"00",
         11006 => x"00",
         11007 => x"00",
         11008 => x"00",
         11009 => x"00",
         11010 => x"00",
         11011 => x"00",
         11012 => x"00",
         11013 => x"00",
         11014 => x"00",
         11015 => x"00",
         11016 => x"00",
         11017 => x"00",
         11018 => x"00",
         11019 => x"00",
         11020 => x"00",
         11021 => x"00",
         11022 => x"00",
         11023 => x"00",
         11024 => x"00",
         11025 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"e4",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"f4",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"e0",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"84",
           393 => x"82",
           394 => x"af",
           395 => x"d8",
           396 => x"80",
           397 => x"d8",
           398 => x"ad",
           399 => x"d4",
           400 => x"90",
           401 => x"d4",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"84",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"84",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"84",
           416 => x"82",
           417 => x"93",
           418 => x"d8",
           419 => x"80",
           420 => x"d8",
           421 => x"c0",
           422 => x"d4",
           423 => x"90",
           424 => x"d4",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"f3",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"d8",
           636 => x"05",
           637 => x"d4",
           638 => x"08",
           639 => x"d4",
           640 => x"08",
           641 => x"ac",
           642 => x"84",
           643 => x"d8",
           644 => x"82",
           645 => x"f8",
           646 => x"d8",
           647 => x"05",
           648 => x"d8",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"d4",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"d4",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"d4",
           668 => x"08",
           669 => x"d8",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"d8",
           674 => x"05",
           675 => x"d4",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"d8",
           681 => x"05",
           682 => x"e9",
           683 => x"d4",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"d4",
           688 => x"0c",
           689 => x"d4",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"d4",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"d8",
           698 => x"05",
           699 => x"71",
           700 => x"d8",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"d8",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"d4",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"d8",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"d4",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"d4",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"d8",
           736 => x"05",
           737 => x"d8",
           738 => x"05",
           739 => x"d8",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"d8",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"d4",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"d8",
           763 => x"05",
           764 => x"d8",
           765 => x"05",
           766 => x"d8",
           767 => x"05",
           768 => x"a3",
           769 => x"c8",
           770 => x"d8",
           771 => x"05",
           772 => x"d4",
           773 => x"08",
           774 => x"c8",
           775 => x"87",
           776 => x"d8",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"d4",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"d4",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"d8",
           797 => x"05",
           798 => x"33",
           799 => x"d8",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"d4",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"d8",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"d8",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"d8",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"d4",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"d8",
           856 => x"05",
           857 => x"d4",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"d4",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"d4",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"d4",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"d4",
           894 => x"0c",
           895 => x"d4",
           896 => x"08",
           897 => x"92",
           898 => x"d8",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"d4",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"d4",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"d4",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"d4",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"d4",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"d4",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"d8",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"d8",
           960 => x"05",
           961 => x"51",
           962 => x"d8",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"d4",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"d8",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"d4",
           983 => x"08",
           984 => x"d8",
           985 => x"c8",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"d4",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"d4",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"d8",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"d4",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"d8",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"d8",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"d8",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"d8",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"d8",
          1055 => x"05",
          1056 => x"d4",
          1057 => x"08",
          1058 => x"d8",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"d8",
          1065 => x"05",
          1066 => x"d4",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"d4",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"d4",
          1082 => x"23",
          1083 => x"88",
          1084 => x"d4",
          1085 => x"23",
          1086 => x"d8",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"d8",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"d8",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"d8",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"d8",
          1111 => x"05",
          1112 => x"d4",
          1113 => x"08",
          1114 => x"d8",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"d8",
          1121 => x"05",
          1122 => x"d4",
          1123 => x"22",
          1124 => x"51",
          1125 => x"d8",
          1126 => x"05",
          1127 => x"d8",
          1128 => x"d4",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"d8",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"d8",
          1142 => x"05",
          1143 => x"d4",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"d4",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"d8",
          1162 => x"05",
          1163 => x"d8",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"d4",
          1177 => x"0c",
          1178 => x"d4",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"d8",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"d4",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"d8",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"d8",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"d8",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"d8",
          1224 => x"05",
          1225 => x"d4",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"d4",
          1235 => x"33",
          1236 => x"70",
          1237 => x"d8",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"d8",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"d4",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"d4",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"d4",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"d8",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"d4",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"d8",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"d8",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"d8",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"d8",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"d4",
          1382 => x"22",
          1383 => x"54",
          1384 => x"d4",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"d4",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"d4",
          1398 => x"08",
          1399 => x"d4",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"d4",
          1408 => x"22",
          1409 => x"53",
          1410 => x"d4",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"d8",
          1416 => x"05",
          1417 => x"d8",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"d4",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"d4",
          1431 => x"22",
          1432 => x"53",
          1433 => x"d4",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"d8",
          1439 => x"05",
          1440 => x"d8",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"d4",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"d8",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"d4",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"d8",
          1468 => x"05",
          1469 => x"54",
          1470 => x"d8",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"d8",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"d4",
          1480 => x"08",
          1481 => x"d4",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"d8",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"d8",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"d4",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"d4",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"d4",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"d4",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"d4",
          1521 => x"08",
          1522 => x"d4",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"c8",
          1527 => x"3d",
          1528 => x"d4",
          1529 => x"d8",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"d4",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"d4",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"f4",
          1556 => x"f4",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"d8",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"ac",
          1568 => x"ac",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"d8",
          1577 => x"05",
          1578 => x"d8",
          1579 => x"05",
          1580 => x"d8",
          1581 => x"05",
          1582 => x"c8",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"d4",
          1586 => x"d8",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"d8",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"d4",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"d4",
          1604 => x"08",
          1605 => x"d8",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"d8",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"d4",
          1626 => x"08",
          1627 => x"d4",
          1628 => x"0c",
          1629 => x"d4",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"d4",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"d4",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"d4",
          1646 => x"d8",
          1647 => x"3d",
          1648 => x"d4",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"d8",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"d4",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"d8",
          1683 => x"05",
          1684 => x"d8",
          1685 => x"05",
          1686 => x"80",
          1687 => x"d8",
          1688 => x"05",
          1689 => x"d4",
          1690 => x"08",
          1691 => x"d4",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"c8",
          1697 => x"a3",
          1698 => x"d4",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"d4",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"d8",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"d8",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"d8",
          1733 => x"05",
          1734 => x"d4",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"d8",
          1744 => x"05",
          1745 => x"33",
          1746 => x"d4",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"d8",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"d4",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"d4",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"d8",
          1778 => x"05",
          1779 => x"d4",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"d4",
          1785 => x"0c",
          1786 => x"d4",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"d4",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"d4",
          1796 => x"0c",
          1797 => x"d4",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"d8",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"d8",
          1809 => x"05",
          1810 => x"d4",
          1811 => x"08",
          1812 => x"d4",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"d4",
          1816 => x"0c",
          1817 => x"d8",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"d4",
          1822 => x"08",
          1823 => x"06",
          1824 => x"d4",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"d8",
          1829 => x"3d",
          1830 => x"d4",
          1831 => x"d8",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"d8",
          1835 => x"05",
          1836 => x"d4",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"d8",
          1842 => x"05",
          1843 => x"82",
          1844 => x"d8",
          1845 => x"05",
          1846 => x"d4",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"d8",
          1862 => x"05",
          1863 => x"d4",
          1864 => x"08",
          1865 => x"d4",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"d4",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"d4",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"d4",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"d4",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"d8",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"d4",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"d4",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"d4",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"d8",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"d4",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"d4",
          1939 => x"08",
          1940 => x"d8",
          1941 => x"05",
          1942 => x"d4",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"c8",
          1947 => x"3d",
          1948 => x"d4",
          1949 => x"d8",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"d8",
          1953 => x"05",
          1954 => x"d4",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"d8",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"d8",
          1963 => x"05",
          1964 => x"70",
          1965 => x"d8",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"d4",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"d8",
          1985 => x"05",
          1986 => x"d4",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"d4",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"d4",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"d4",
          2005 => x"08",
          2006 => x"d8",
          2007 => x"05",
          2008 => x"d4",
          2009 => x"08",
          2010 => x"71",
          2011 => x"d4",
          2012 => x"08",
          2013 => x"d8",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"d4",
          2022 => x"d8",
          2023 => x"3d",
          2024 => x"d4",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"d4",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"d8",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"d4",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"d4",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"d4",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"d4",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"d4",
          2082 => x"08",
          2083 => x"71",
          2084 => x"d8",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"d8",
          2089 => x"05",
          2090 => x"d4",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"d4",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"82",
          2100 => x"f8",
          2101 => x"d8",
          2102 => x"05",
          2103 => x"80",
          2104 => x"d4",
          2105 => x"0c",
          2106 => x"82",
          2107 => x"f8",
          2108 => x"71",
          2109 => x"d4",
          2110 => x"08",
          2111 => x"d8",
          2112 => x"05",
          2113 => x"ff",
          2114 => x"70",
          2115 => x"38",
          2116 => x"08",
          2117 => x"ff",
          2118 => x"d4",
          2119 => x"0c",
          2120 => x"08",
          2121 => x"ff",
          2122 => x"ff",
          2123 => x"d8",
          2124 => x"05",
          2125 => x"82",
          2126 => x"f8",
          2127 => x"d8",
          2128 => x"05",
          2129 => x"d4",
          2130 => x"08",
          2131 => x"d8",
          2132 => x"05",
          2133 => x"d8",
          2134 => x"05",
          2135 => x"c8",
          2136 => x"0d",
          2137 => x"0c",
          2138 => x"d4",
          2139 => x"d8",
          2140 => x"3d",
          2141 => x"d4",
          2142 => x"08",
          2143 => x"08",
          2144 => x"82",
          2145 => x"90",
          2146 => x"2e",
          2147 => x"82",
          2148 => x"90",
          2149 => x"05",
          2150 => x"08",
          2151 => x"82",
          2152 => x"90",
          2153 => x"05",
          2154 => x"08",
          2155 => x"82",
          2156 => x"90",
          2157 => x"2e",
          2158 => x"d8",
          2159 => x"05",
          2160 => x"82",
          2161 => x"fc",
          2162 => x"52",
          2163 => x"82",
          2164 => x"fc",
          2165 => x"05",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"d8",
          2169 => x"05",
          2170 => x"d8",
          2171 => x"84",
          2172 => x"d8",
          2173 => x"82",
          2174 => x"02",
          2175 => x"0c",
          2176 => x"80",
          2177 => x"d4",
          2178 => x"0c",
          2179 => x"08",
          2180 => x"80",
          2181 => x"82",
          2182 => x"88",
          2183 => x"82",
          2184 => x"88",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"82",
          2188 => x"fc",
          2189 => x"38",
          2190 => x"d8",
          2191 => x"05",
          2192 => x"d4",
          2193 => x"08",
          2194 => x"08",
          2195 => x"82",
          2196 => x"8c",
          2197 => x"25",
          2198 => x"d8",
          2199 => x"05",
          2200 => x"d8",
          2201 => x"05",
          2202 => x"82",
          2203 => x"f0",
          2204 => x"d8",
          2205 => x"05",
          2206 => x"81",
          2207 => x"d4",
          2208 => x"0c",
          2209 => x"08",
          2210 => x"82",
          2211 => x"fc",
          2212 => x"53",
          2213 => x"08",
          2214 => x"52",
          2215 => x"08",
          2216 => x"51",
          2217 => x"82",
          2218 => x"70",
          2219 => x"08",
          2220 => x"54",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"f8",
          2225 => x"82",
          2226 => x"f8",
          2227 => x"d8",
          2228 => x"05",
          2229 => x"d8",
          2230 => x"89",
          2231 => x"d8",
          2232 => x"82",
          2233 => x"02",
          2234 => x"0c",
          2235 => x"80",
          2236 => x"d4",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"88",
          2242 => x"82",
          2243 => x"88",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"8c",
          2248 => x"25",
          2249 => x"d8",
          2250 => x"05",
          2251 => x"d8",
          2252 => x"05",
          2253 => x"82",
          2254 => x"8c",
          2255 => x"82",
          2256 => x"88",
          2257 => x"81",
          2258 => x"d8",
          2259 => x"82",
          2260 => x"f8",
          2261 => x"82",
          2262 => x"fc",
          2263 => x"2e",
          2264 => x"d8",
          2265 => x"05",
          2266 => x"d8",
          2267 => x"05",
          2268 => x"d4",
          2269 => x"08",
          2270 => x"c8",
          2271 => x"3d",
          2272 => x"d4",
          2273 => x"d8",
          2274 => x"82",
          2275 => x"fd",
          2276 => x"53",
          2277 => x"08",
          2278 => x"52",
          2279 => x"08",
          2280 => x"51",
          2281 => x"82",
          2282 => x"70",
          2283 => x"0c",
          2284 => x"0d",
          2285 => x"0c",
          2286 => x"d4",
          2287 => x"d8",
          2288 => x"3d",
          2289 => x"82",
          2290 => x"8c",
          2291 => x"82",
          2292 => x"88",
          2293 => x"93",
          2294 => x"c8",
          2295 => x"d8",
          2296 => x"85",
          2297 => x"d8",
          2298 => x"82",
          2299 => x"02",
          2300 => x"0c",
          2301 => x"81",
          2302 => x"d4",
          2303 => x"0c",
          2304 => x"d8",
          2305 => x"05",
          2306 => x"d4",
          2307 => x"08",
          2308 => x"08",
          2309 => x"27",
          2310 => x"d8",
          2311 => x"05",
          2312 => x"ae",
          2313 => x"82",
          2314 => x"8c",
          2315 => x"a2",
          2316 => x"d4",
          2317 => x"08",
          2318 => x"d4",
          2319 => x"0c",
          2320 => x"08",
          2321 => x"10",
          2322 => x"08",
          2323 => x"ff",
          2324 => x"d8",
          2325 => x"05",
          2326 => x"80",
          2327 => x"d8",
          2328 => x"05",
          2329 => x"d4",
          2330 => x"08",
          2331 => x"82",
          2332 => x"88",
          2333 => x"d8",
          2334 => x"05",
          2335 => x"d8",
          2336 => x"05",
          2337 => x"d4",
          2338 => x"08",
          2339 => x"08",
          2340 => x"07",
          2341 => x"08",
          2342 => x"82",
          2343 => x"fc",
          2344 => x"2a",
          2345 => x"08",
          2346 => x"82",
          2347 => x"8c",
          2348 => x"2a",
          2349 => x"08",
          2350 => x"ff",
          2351 => x"d8",
          2352 => x"05",
          2353 => x"93",
          2354 => x"d4",
          2355 => x"08",
          2356 => x"d4",
          2357 => x"0c",
          2358 => x"82",
          2359 => x"f8",
          2360 => x"82",
          2361 => x"f4",
          2362 => x"82",
          2363 => x"f4",
          2364 => x"d8",
          2365 => x"3d",
          2366 => x"d4",
          2367 => x"d8",
          2368 => x"82",
          2369 => x"f7",
          2370 => x"0b",
          2371 => x"08",
          2372 => x"82",
          2373 => x"8c",
          2374 => x"80",
          2375 => x"d8",
          2376 => x"05",
          2377 => x"51",
          2378 => x"53",
          2379 => x"d4",
          2380 => x"34",
          2381 => x"06",
          2382 => x"2e",
          2383 => x"91",
          2384 => x"d4",
          2385 => x"08",
          2386 => x"05",
          2387 => x"ce",
          2388 => x"d4",
          2389 => x"33",
          2390 => x"2e",
          2391 => x"a4",
          2392 => x"82",
          2393 => x"f0",
          2394 => x"d8",
          2395 => x"05",
          2396 => x"81",
          2397 => x"70",
          2398 => x"72",
          2399 => x"d4",
          2400 => x"34",
          2401 => x"08",
          2402 => x"53",
          2403 => x"09",
          2404 => x"dc",
          2405 => x"d4",
          2406 => x"08",
          2407 => x"05",
          2408 => x"08",
          2409 => x"33",
          2410 => x"08",
          2411 => x"82",
          2412 => x"f8",
          2413 => x"d8",
          2414 => x"05",
          2415 => x"d4",
          2416 => x"08",
          2417 => x"b6",
          2418 => x"d4",
          2419 => x"08",
          2420 => x"84",
          2421 => x"39",
          2422 => x"d8",
          2423 => x"05",
          2424 => x"d4",
          2425 => x"08",
          2426 => x"05",
          2427 => x"08",
          2428 => x"33",
          2429 => x"08",
          2430 => x"81",
          2431 => x"0b",
          2432 => x"08",
          2433 => x"82",
          2434 => x"88",
          2435 => x"08",
          2436 => x"0c",
          2437 => x"53",
          2438 => x"d8",
          2439 => x"05",
          2440 => x"39",
          2441 => x"08",
          2442 => x"53",
          2443 => x"8d",
          2444 => x"82",
          2445 => x"ec",
          2446 => x"80",
          2447 => x"d4",
          2448 => x"33",
          2449 => x"27",
          2450 => x"d8",
          2451 => x"05",
          2452 => x"b9",
          2453 => x"8d",
          2454 => x"82",
          2455 => x"ec",
          2456 => x"d8",
          2457 => x"82",
          2458 => x"f4",
          2459 => x"39",
          2460 => x"08",
          2461 => x"53",
          2462 => x"90",
          2463 => x"d4",
          2464 => x"33",
          2465 => x"26",
          2466 => x"39",
          2467 => x"d8",
          2468 => x"05",
          2469 => x"39",
          2470 => x"d8",
          2471 => x"05",
          2472 => x"82",
          2473 => x"fc",
          2474 => x"d8",
          2475 => x"05",
          2476 => x"73",
          2477 => x"38",
          2478 => x"08",
          2479 => x"53",
          2480 => x"27",
          2481 => x"d8",
          2482 => x"05",
          2483 => x"51",
          2484 => x"d8",
          2485 => x"05",
          2486 => x"d4",
          2487 => x"33",
          2488 => x"53",
          2489 => x"d4",
          2490 => x"34",
          2491 => x"08",
          2492 => x"53",
          2493 => x"ad",
          2494 => x"d4",
          2495 => x"33",
          2496 => x"53",
          2497 => x"d4",
          2498 => x"34",
          2499 => x"08",
          2500 => x"53",
          2501 => x"8d",
          2502 => x"82",
          2503 => x"ec",
          2504 => x"98",
          2505 => x"d4",
          2506 => x"33",
          2507 => x"08",
          2508 => x"54",
          2509 => x"26",
          2510 => x"0b",
          2511 => x"08",
          2512 => x"80",
          2513 => x"d8",
          2514 => x"05",
          2515 => x"d8",
          2516 => x"05",
          2517 => x"d8",
          2518 => x"05",
          2519 => x"82",
          2520 => x"fc",
          2521 => x"d8",
          2522 => x"05",
          2523 => x"81",
          2524 => x"70",
          2525 => x"52",
          2526 => x"33",
          2527 => x"08",
          2528 => x"fe",
          2529 => x"d8",
          2530 => x"05",
          2531 => x"80",
          2532 => x"82",
          2533 => x"fc",
          2534 => x"82",
          2535 => x"fc",
          2536 => x"d8",
          2537 => x"05",
          2538 => x"d4",
          2539 => x"08",
          2540 => x"81",
          2541 => x"d4",
          2542 => x"0c",
          2543 => x"08",
          2544 => x"82",
          2545 => x"8b",
          2546 => x"d8",
          2547 => x"82",
          2548 => x"02",
          2549 => x"0c",
          2550 => x"80",
          2551 => x"d4",
          2552 => x"34",
          2553 => x"08",
          2554 => x"53",
          2555 => x"82",
          2556 => x"88",
          2557 => x"08",
          2558 => x"33",
          2559 => x"d8",
          2560 => x"05",
          2561 => x"ff",
          2562 => x"a0",
          2563 => x"06",
          2564 => x"d8",
          2565 => x"05",
          2566 => x"81",
          2567 => x"53",
          2568 => x"d8",
          2569 => x"05",
          2570 => x"ad",
          2571 => x"06",
          2572 => x"0b",
          2573 => x"08",
          2574 => x"82",
          2575 => x"88",
          2576 => x"08",
          2577 => x"0c",
          2578 => x"53",
          2579 => x"d8",
          2580 => x"05",
          2581 => x"d4",
          2582 => x"33",
          2583 => x"2e",
          2584 => x"81",
          2585 => x"d8",
          2586 => x"05",
          2587 => x"81",
          2588 => x"70",
          2589 => x"72",
          2590 => x"d4",
          2591 => x"34",
          2592 => x"08",
          2593 => x"82",
          2594 => x"e8",
          2595 => x"d8",
          2596 => x"05",
          2597 => x"2e",
          2598 => x"d8",
          2599 => x"05",
          2600 => x"2e",
          2601 => x"cd",
          2602 => x"82",
          2603 => x"f4",
          2604 => x"d8",
          2605 => x"05",
          2606 => x"81",
          2607 => x"70",
          2608 => x"72",
          2609 => x"d4",
          2610 => x"34",
          2611 => x"82",
          2612 => x"d4",
          2613 => x"34",
          2614 => x"08",
          2615 => x"70",
          2616 => x"71",
          2617 => x"51",
          2618 => x"82",
          2619 => x"f8",
          2620 => x"fe",
          2621 => x"d4",
          2622 => x"33",
          2623 => x"26",
          2624 => x"0b",
          2625 => x"08",
          2626 => x"83",
          2627 => x"d8",
          2628 => x"05",
          2629 => x"73",
          2630 => x"82",
          2631 => x"f8",
          2632 => x"72",
          2633 => x"38",
          2634 => x"0b",
          2635 => x"08",
          2636 => x"82",
          2637 => x"0b",
          2638 => x"08",
          2639 => x"b2",
          2640 => x"d4",
          2641 => x"33",
          2642 => x"27",
          2643 => x"d8",
          2644 => x"05",
          2645 => x"b9",
          2646 => x"8d",
          2647 => x"82",
          2648 => x"ec",
          2649 => x"a5",
          2650 => x"82",
          2651 => x"f4",
          2652 => x"0b",
          2653 => x"08",
          2654 => x"82",
          2655 => x"f8",
          2656 => x"a0",
          2657 => x"cf",
          2658 => x"d4",
          2659 => x"33",
          2660 => x"73",
          2661 => x"82",
          2662 => x"f8",
          2663 => x"11",
          2664 => x"82",
          2665 => x"f8",
          2666 => x"d8",
          2667 => x"05",
          2668 => x"51",
          2669 => x"d8",
          2670 => x"05",
          2671 => x"d4",
          2672 => x"33",
          2673 => x"27",
          2674 => x"d8",
          2675 => x"05",
          2676 => x"51",
          2677 => x"d8",
          2678 => x"05",
          2679 => x"d4",
          2680 => x"33",
          2681 => x"26",
          2682 => x"0b",
          2683 => x"08",
          2684 => x"81",
          2685 => x"d8",
          2686 => x"05",
          2687 => x"d4",
          2688 => x"33",
          2689 => x"74",
          2690 => x"80",
          2691 => x"d4",
          2692 => x"0c",
          2693 => x"82",
          2694 => x"f4",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"82",
          2698 => x"f8",
          2699 => x"12",
          2700 => x"08",
          2701 => x"82",
          2702 => x"88",
          2703 => x"08",
          2704 => x"0c",
          2705 => x"51",
          2706 => x"72",
          2707 => x"d4",
          2708 => x"34",
          2709 => x"82",
          2710 => x"f0",
          2711 => x"72",
          2712 => x"38",
          2713 => x"08",
          2714 => x"30",
          2715 => x"08",
          2716 => x"82",
          2717 => x"8c",
          2718 => x"d8",
          2719 => x"05",
          2720 => x"53",
          2721 => x"d8",
          2722 => x"05",
          2723 => x"d4",
          2724 => x"08",
          2725 => x"0c",
          2726 => x"82",
          2727 => x"04",
          2728 => x"79",
          2729 => x"56",
          2730 => x"80",
          2731 => x"38",
          2732 => x"08",
          2733 => x"3f",
          2734 => x"08",
          2735 => x"85",
          2736 => x"80",
          2737 => x"33",
          2738 => x"2e",
          2739 => x"86",
          2740 => x"55",
          2741 => x"57",
          2742 => x"82",
          2743 => x"70",
          2744 => x"e6",
          2745 => x"d8",
          2746 => x"74",
          2747 => x"51",
          2748 => x"82",
          2749 => x"8b",
          2750 => x"33",
          2751 => x"2e",
          2752 => x"81",
          2753 => x"ff",
          2754 => x"99",
          2755 => x"38",
          2756 => x"82",
          2757 => x"89",
          2758 => x"ff",
          2759 => x"52",
          2760 => x"81",
          2761 => x"84",
          2762 => x"f4",
          2763 => x"08",
          2764 => x"e4",
          2765 => x"39",
          2766 => x"51",
          2767 => x"82",
          2768 => x"80",
          2769 => x"b5",
          2770 => x"eb",
          2771 => x"a0",
          2772 => x"39",
          2773 => x"51",
          2774 => x"82",
          2775 => x"80",
          2776 => x"b5",
          2777 => x"cf",
          2778 => x"ec",
          2779 => x"39",
          2780 => x"51",
          2781 => x"82",
          2782 => x"bb",
          2783 => x"b8",
          2784 => x"82",
          2785 => x"af",
          2786 => x"f4",
          2787 => x"82",
          2788 => x"a3",
          2789 => x"a4",
          2790 => x"82",
          2791 => x"97",
          2792 => x"cc",
          2793 => x"82",
          2794 => x"8b",
          2795 => x"fc",
          2796 => x"82",
          2797 => x"d8",
          2798 => x"3d",
          2799 => x"3d",
          2800 => x"56",
          2801 => x"e7",
          2802 => x"74",
          2803 => x"e8",
          2804 => x"39",
          2805 => x"74",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"ef",
          2809 => x"d8",
          2810 => x"79",
          2811 => x"82",
          2812 => x"ff",
          2813 => x"87",
          2814 => x"ec",
          2815 => x"02",
          2816 => x"e3",
          2817 => x"57",
          2818 => x"30",
          2819 => x"73",
          2820 => x"59",
          2821 => x"77",
          2822 => x"83",
          2823 => x"74",
          2824 => x"81",
          2825 => x"55",
          2826 => x"81",
          2827 => x"53",
          2828 => x"3d",
          2829 => x"81",
          2830 => x"82",
          2831 => x"57",
          2832 => x"08",
          2833 => x"d8",
          2834 => x"c0",
          2835 => x"82",
          2836 => x"59",
          2837 => x"05",
          2838 => x"53",
          2839 => x"51",
          2840 => x"3f",
          2841 => x"08",
          2842 => x"c8",
          2843 => x"7a",
          2844 => x"2e",
          2845 => x"19",
          2846 => x"59",
          2847 => x"3d",
          2848 => x"81",
          2849 => x"76",
          2850 => x"07",
          2851 => x"30",
          2852 => x"72",
          2853 => x"51",
          2854 => x"2e",
          2855 => x"b8",
          2856 => x"c0",
          2857 => x"52",
          2858 => x"92",
          2859 => x"75",
          2860 => x"0c",
          2861 => x"04",
          2862 => x"7d",
          2863 => x"bb",
          2864 => x"5a",
          2865 => x"53",
          2866 => x"51",
          2867 => x"82",
          2868 => x"80",
          2869 => x"80",
          2870 => x"77",
          2871 => x"38",
          2872 => x"f4",
          2873 => x"f4",
          2874 => x"f4",
          2875 => x"f4",
          2876 => x"82",
          2877 => x"53",
          2878 => x"08",
          2879 => x"c4",
          2880 => x"d7",
          2881 => x"a8",
          2882 => x"61",
          2883 => x"c8",
          2884 => x"7f",
          2885 => x"82",
          2886 => x"59",
          2887 => x"04",
          2888 => x"c8",
          2889 => x"0d",
          2890 => x"0d",
          2891 => x"02",
          2892 => x"cf",
          2893 => x"73",
          2894 => x"5f",
          2895 => x"5e",
          2896 => x"82",
          2897 => x"ff",
          2898 => x"82",
          2899 => x"ff",
          2900 => x"80",
          2901 => x"27",
          2902 => x"7b",
          2903 => x"38",
          2904 => x"a7",
          2905 => x"39",
          2906 => x"72",
          2907 => x"38",
          2908 => x"82",
          2909 => x"ff",
          2910 => x"89",
          2911 => x"90",
          2912 => x"d7",
          2913 => x"55",
          2914 => x"74",
          2915 => x"7a",
          2916 => x"72",
          2917 => x"b8",
          2918 => x"b8",
          2919 => x"39",
          2920 => x"51",
          2921 => x"3f",
          2922 => x"a1",
          2923 => x"53",
          2924 => x"8e",
          2925 => x"52",
          2926 => x"51",
          2927 => x"3f",
          2928 => x"b9",
          2929 => x"b8",
          2930 => x"15",
          2931 => x"ac",
          2932 => x"51",
          2933 => x"fe",
          2934 => x"b9",
          2935 => x"b7",
          2936 => x"55",
          2937 => x"80",
          2938 => x"18",
          2939 => x"53",
          2940 => x"7a",
          2941 => x"81",
          2942 => x"9f",
          2943 => x"38",
          2944 => x"73",
          2945 => x"ff",
          2946 => x"72",
          2947 => x"38",
          2948 => x"26",
          2949 => x"f4",
          2950 => x"73",
          2951 => x"82",
          2952 => x"52",
          2953 => x"8d",
          2954 => x"55",
          2955 => x"82",
          2956 => x"d3",
          2957 => x"18",
          2958 => x"58",
          2959 => x"82",
          2960 => x"98",
          2961 => x"2c",
          2962 => x"a0",
          2963 => x"06",
          2964 => x"ea",
          2965 => x"c8",
          2966 => x"70",
          2967 => x"a0",
          2968 => x"72",
          2969 => x"30",
          2970 => x"73",
          2971 => x"51",
          2972 => x"57",
          2973 => x"73",
          2974 => x"76",
          2975 => x"81",
          2976 => x"80",
          2977 => x"7c",
          2978 => x"78",
          2979 => x"38",
          2980 => x"82",
          2981 => x"8f",
          2982 => x"fc",
          2983 => x"9b",
          2984 => x"b9",
          2985 => x"b9",
          2986 => x"ff",
          2987 => x"82",
          2988 => x"51",
          2989 => x"82",
          2990 => x"82",
          2991 => x"82",
          2992 => x"52",
          2993 => x"51",
          2994 => x"3f",
          2995 => x"84",
          2996 => x"3f",
          2997 => x"04",
          2998 => x"87",
          2999 => x"08",
          3000 => x"3f",
          3001 => x"c3",
          3002 => x"f0",
          3003 => x"3f",
          3004 => x"b7",
          3005 => x"2a",
          3006 => x"51",
          3007 => x"2e",
          3008 => x"51",
          3009 => x"82",
          3010 => x"9d",
          3011 => x"51",
          3012 => x"72",
          3013 => x"81",
          3014 => x"71",
          3015 => x"38",
          3016 => x"87",
          3017 => x"98",
          3018 => x"3f",
          3019 => x"fb",
          3020 => x"2a",
          3021 => x"51",
          3022 => x"2e",
          3023 => x"51",
          3024 => x"82",
          3025 => x"9c",
          3026 => x"51",
          3027 => x"72",
          3028 => x"81",
          3029 => x"71",
          3030 => x"38",
          3031 => x"cb",
          3032 => x"bc",
          3033 => x"3f",
          3034 => x"bf",
          3035 => x"2a",
          3036 => x"51",
          3037 => x"2e",
          3038 => x"51",
          3039 => x"82",
          3040 => x"9c",
          3041 => x"51",
          3042 => x"72",
          3043 => x"81",
          3044 => x"71",
          3045 => x"38",
          3046 => x"8f",
          3047 => x"e4",
          3048 => x"3f",
          3049 => x"83",
          3050 => x"2a",
          3051 => x"51",
          3052 => x"2e",
          3053 => x"51",
          3054 => x"82",
          3055 => x"9c",
          3056 => x"51",
          3057 => x"72",
          3058 => x"81",
          3059 => x"71",
          3060 => x"38",
          3061 => x"d3",
          3062 => x"8c",
          3063 => x"3f",
          3064 => x"c7",
          3065 => x"3f",
          3066 => x"04",
          3067 => x"77",
          3068 => x"a3",
          3069 => x"55",
          3070 => x"52",
          3071 => x"e9",
          3072 => x"82",
          3073 => x"54",
          3074 => x"81",
          3075 => x"c8",
          3076 => x"d8",
          3077 => x"b2",
          3078 => x"c8",
          3079 => x"82",
          3080 => x"07",
          3081 => x"71",
          3082 => x"54",
          3083 => x"82",
          3084 => x"0b",
          3085 => x"c4",
          3086 => x"81",
          3087 => x"06",
          3088 => x"ef",
          3089 => x"52",
          3090 => x"c9",
          3091 => x"d8",
          3092 => x"2e",
          3093 => x"d8",
          3094 => x"cf",
          3095 => x"39",
          3096 => x"51",
          3097 => x"3f",
          3098 => x"0b",
          3099 => x"34",
          3100 => x"d3",
          3101 => x"73",
          3102 => x"81",
          3103 => x"82",
          3104 => x"74",
          3105 => x"ae",
          3106 => x"0b",
          3107 => x"0c",
          3108 => x"04",
          3109 => x"80",
          3110 => x"ef",
          3111 => x"5d",
          3112 => x"51",
          3113 => x"3f",
          3114 => x"08",
          3115 => x"59",
          3116 => x"09",
          3117 => x"38",
          3118 => x"83",
          3119 => x"e4",
          3120 => x"dc",
          3121 => x"53",
          3122 => x"d9",
          3123 => x"8c",
          3124 => x"d8",
          3125 => x"2e",
          3126 => x"bb",
          3127 => x"d7",
          3128 => x"5f",
          3129 => x"a0",
          3130 => x"ef",
          3131 => x"70",
          3132 => x"f8",
          3133 => x"fd",
          3134 => x"3d",
          3135 => x"51",
          3136 => x"82",
          3137 => x"90",
          3138 => x"2c",
          3139 => x"80",
          3140 => x"d4",
          3141 => x"c1",
          3142 => x"38",
          3143 => x"83",
          3144 => x"ab",
          3145 => x"78",
          3146 => x"b3",
          3147 => x"24",
          3148 => x"80",
          3149 => x"38",
          3150 => x"78",
          3151 => x"83",
          3152 => x"2e",
          3153 => x"8e",
          3154 => x"bd",
          3155 => x"38",
          3156 => x"90",
          3157 => x"2e",
          3158 => x"78",
          3159 => x"84",
          3160 => x"39",
          3161 => x"85",
          3162 => x"80",
          3163 => x"bd",
          3164 => x"39",
          3165 => x"2e",
          3166 => x"78",
          3167 => x"b0",
          3168 => x"d0",
          3169 => x"38",
          3170 => x"24",
          3171 => x"80",
          3172 => x"fc",
          3173 => x"c3",
          3174 => x"38",
          3175 => x"78",
          3176 => x"8c",
          3177 => x"80",
          3178 => x"d3",
          3179 => x"39",
          3180 => x"2e",
          3181 => x"78",
          3182 => x"92",
          3183 => x"f8",
          3184 => x"38",
          3185 => x"2e",
          3186 => x"8d",
          3187 => x"81",
          3188 => x"d5",
          3189 => x"85",
          3190 => x"38",
          3191 => x"b4",
          3192 => x"11",
          3193 => x"05",
          3194 => x"3f",
          3195 => x"08",
          3196 => x"bc",
          3197 => x"bf",
          3198 => x"fe",
          3199 => x"ff",
          3200 => x"eb",
          3201 => x"d8",
          3202 => x"2e",
          3203 => x"63",
          3204 => x"80",
          3205 => x"cb",
          3206 => x"02",
          3207 => x"33",
          3208 => x"ce",
          3209 => x"c8",
          3210 => x"06",
          3211 => x"38",
          3212 => x"51",
          3213 => x"81",
          3214 => x"39",
          3215 => x"51",
          3216 => x"b4",
          3217 => x"11",
          3218 => x"05",
          3219 => x"3f",
          3220 => x"08",
          3221 => x"8d",
          3222 => x"80",
          3223 => x"cf",
          3224 => x"80",
          3225 => x"82",
          3226 => x"52",
          3227 => x"51",
          3228 => x"b4",
          3229 => x"11",
          3230 => x"05",
          3231 => x"3f",
          3232 => x"08",
          3233 => x"38",
          3234 => x"fc",
          3235 => x"3d",
          3236 => x"53",
          3237 => x"51",
          3238 => x"82",
          3239 => x"86",
          3240 => x"c8",
          3241 => x"53",
          3242 => x"52",
          3243 => x"b1",
          3244 => x"80",
          3245 => x"53",
          3246 => x"84",
          3247 => x"d9",
          3248 => x"81",
          3249 => x"82",
          3250 => x"81",
          3251 => x"bc",
          3252 => x"92",
          3253 => x"fc",
          3254 => x"3d",
          3255 => x"51",
          3256 => x"82",
          3257 => x"b5",
          3258 => x"05",
          3259 => x"d8",
          3260 => x"82",
          3261 => x"52",
          3262 => x"ff",
          3263 => x"39",
          3264 => x"84",
          3265 => x"9c",
          3266 => x"c8",
          3267 => x"ff",
          3268 => x"5b",
          3269 => x"82",
          3270 => x"b5",
          3271 => x"05",
          3272 => x"a4",
          3273 => x"c8",
          3274 => x"ff",
          3275 => x"59",
          3276 => x"82",
          3277 => x"82",
          3278 => x"80",
          3279 => x"82",
          3280 => x"81",
          3281 => x"78",
          3282 => x"7a",
          3283 => x"3f",
          3284 => x"08",
          3285 => x"8d",
          3286 => x"c8",
          3287 => x"bb",
          3288 => x"39",
          3289 => x"80",
          3290 => x"84",
          3291 => x"df",
          3292 => x"c8",
          3293 => x"fa",
          3294 => x"3d",
          3295 => x"53",
          3296 => x"51",
          3297 => x"82",
          3298 => x"80",
          3299 => x"38",
          3300 => x"f8",
          3301 => x"84",
          3302 => x"b3",
          3303 => x"c8",
          3304 => x"82",
          3305 => x"42",
          3306 => x"51",
          3307 => x"3f",
          3308 => x"5a",
          3309 => x"81",
          3310 => x"59",
          3311 => x"84",
          3312 => x"7a",
          3313 => x"38",
          3314 => x"b4",
          3315 => x"11",
          3316 => x"05",
          3317 => x"3f",
          3318 => x"08",
          3319 => x"85",
          3320 => x"fe",
          3321 => x"ff",
          3322 => x"e7",
          3323 => x"d8",
          3324 => x"2e",
          3325 => x"b4",
          3326 => x"11",
          3327 => x"05",
          3328 => x"3f",
          3329 => x"08",
          3330 => x"d9",
          3331 => x"f8",
          3332 => x"c7",
          3333 => x"79",
          3334 => x"89",
          3335 => x"79",
          3336 => x"5b",
          3337 => x"61",
          3338 => x"eb",
          3339 => x"ff",
          3340 => x"ff",
          3341 => x"e7",
          3342 => x"d8",
          3343 => x"2e",
          3344 => x"b4",
          3345 => x"11",
          3346 => x"05",
          3347 => x"3f",
          3348 => x"08",
          3349 => x"8d",
          3350 => x"fe",
          3351 => x"ff",
          3352 => x"e6",
          3353 => x"d8",
          3354 => x"2e",
          3355 => x"82",
          3356 => x"ff",
          3357 => x"63",
          3358 => x"27",
          3359 => x"70",
          3360 => x"5e",
          3361 => x"7c",
          3362 => x"78",
          3363 => x"79",
          3364 => x"52",
          3365 => x"51",
          3366 => x"3f",
          3367 => x"81",
          3368 => x"d5",
          3369 => x"c9",
          3370 => x"b9",
          3371 => x"ff",
          3372 => x"ff",
          3373 => x"e6",
          3374 => x"d8",
          3375 => x"df",
          3376 => x"b4",
          3377 => x"80",
          3378 => x"82",
          3379 => x"44",
          3380 => x"82",
          3381 => x"59",
          3382 => x"88",
          3383 => x"f4",
          3384 => x"39",
          3385 => x"33",
          3386 => x"2e",
          3387 => x"d6",
          3388 => x"ab",
          3389 => x"b7",
          3390 => x"80",
          3391 => x"82",
          3392 => x"44",
          3393 => x"d7",
          3394 => x"78",
          3395 => x"38",
          3396 => x"08",
          3397 => x"82",
          3398 => x"fc",
          3399 => x"b4",
          3400 => x"11",
          3401 => x"05",
          3402 => x"3f",
          3403 => x"08",
          3404 => x"82",
          3405 => x"59",
          3406 => x"89",
          3407 => x"f0",
          3408 => x"cc",
          3409 => x"b5",
          3410 => x"80",
          3411 => x"82",
          3412 => x"43",
          3413 => x"d7",
          3414 => x"78",
          3415 => x"38",
          3416 => x"08",
          3417 => x"82",
          3418 => x"59",
          3419 => x"88",
          3420 => x"88",
          3421 => x"39",
          3422 => x"33",
          3423 => x"2e",
          3424 => x"d7",
          3425 => x"88",
          3426 => x"9c",
          3427 => x"43",
          3428 => x"f8",
          3429 => x"84",
          3430 => x"b3",
          3431 => x"c8",
          3432 => x"a7",
          3433 => x"5c",
          3434 => x"2e",
          3435 => x"5c",
          3436 => x"70",
          3437 => x"07",
          3438 => x"7f",
          3439 => x"5a",
          3440 => x"2e",
          3441 => x"a0",
          3442 => x"88",
          3443 => x"b0",
          3444 => x"3f",
          3445 => x"54",
          3446 => x"52",
          3447 => x"c9",
          3448 => x"bc",
          3449 => x"39",
          3450 => x"80",
          3451 => x"84",
          3452 => x"db",
          3453 => x"c8",
          3454 => x"f5",
          3455 => x"3d",
          3456 => x"53",
          3457 => x"51",
          3458 => x"82",
          3459 => x"80",
          3460 => x"63",
          3461 => x"cb",
          3462 => x"34",
          3463 => x"44",
          3464 => x"fc",
          3465 => x"84",
          3466 => x"a3",
          3467 => x"c8",
          3468 => x"f5",
          3469 => x"70",
          3470 => x"82",
          3471 => x"ff",
          3472 => x"82",
          3473 => x"53",
          3474 => x"79",
          3475 => x"e0",
          3476 => x"79",
          3477 => x"ae",
          3478 => x"38",
          3479 => x"9f",
          3480 => x"fe",
          3481 => x"ff",
          3482 => x"e2",
          3483 => x"d8",
          3484 => x"2e",
          3485 => x"59",
          3486 => x"05",
          3487 => x"63",
          3488 => x"ff",
          3489 => x"bd",
          3490 => x"da",
          3491 => x"39",
          3492 => x"f4",
          3493 => x"84",
          3494 => x"e2",
          3495 => x"c8",
          3496 => x"f4",
          3497 => x"3d",
          3498 => x"53",
          3499 => x"51",
          3500 => x"82",
          3501 => x"80",
          3502 => x"60",
          3503 => x"05",
          3504 => x"82",
          3505 => x"78",
          3506 => x"fe",
          3507 => x"ff",
          3508 => x"dc",
          3509 => x"d8",
          3510 => x"38",
          3511 => x"60",
          3512 => x"52",
          3513 => x"51",
          3514 => x"3f",
          3515 => x"08",
          3516 => x"52",
          3517 => x"a6",
          3518 => x"45",
          3519 => x"78",
          3520 => x"e1",
          3521 => x"26",
          3522 => x"82",
          3523 => x"39",
          3524 => x"f0",
          3525 => x"84",
          3526 => x"e2",
          3527 => x"c8",
          3528 => x"92",
          3529 => x"02",
          3530 => x"79",
          3531 => x"5b",
          3532 => x"ff",
          3533 => x"bd",
          3534 => x"aa",
          3535 => x"39",
          3536 => x"f4",
          3537 => x"84",
          3538 => x"b2",
          3539 => x"c8",
          3540 => x"f3",
          3541 => x"3d",
          3542 => x"53",
          3543 => x"51",
          3544 => x"82",
          3545 => x"80",
          3546 => x"60",
          3547 => x"59",
          3548 => x"41",
          3549 => x"f0",
          3550 => x"84",
          3551 => x"fe",
          3552 => x"c8",
          3553 => x"f2",
          3554 => x"70",
          3555 => x"82",
          3556 => x"ff",
          3557 => x"82",
          3558 => x"53",
          3559 => x"79",
          3560 => x"8c",
          3561 => x"79",
          3562 => x"ae",
          3563 => x"38",
          3564 => x"9b",
          3565 => x"fe",
          3566 => x"ff",
          3567 => x"da",
          3568 => x"d8",
          3569 => x"2e",
          3570 => x"60",
          3571 => x"60",
          3572 => x"ff",
          3573 => x"bd",
          3574 => x"8a",
          3575 => x"39",
          3576 => x"51",
          3577 => x"82",
          3578 => x"3f",
          3579 => x"82",
          3580 => x"ff",
          3581 => x"a2",
          3582 => x"3f",
          3583 => x"82",
          3584 => x"ff",
          3585 => x"84",
          3586 => x"87",
          3587 => x"0c",
          3588 => x"0b",
          3589 => x"94",
          3590 => x"39",
          3591 => x"51",
          3592 => x"3f",
          3593 => x"0b",
          3594 => x"84",
          3595 => x"83",
          3596 => x"94",
          3597 => x"ad",
          3598 => x"ff",
          3599 => x"ff",
          3600 => x"df",
          3601 => x"d8",
          3602 => x"2e",
          3603 => x"63",
          3604 => x"c8",
          3605 => x"83",
          3606 => x"78",
          3607 => x"ff",
          3608 => x"ff",
          3609 => x"de",
          3610 => x"d8",
          3611 => x"2e",
          3612 => x"63",
          3613 => x"e4",
          3614 => x"df",
          3615 => x"78",
          3616 => x"c8",
          3617 => x"f0",
          3618 => x"d8",
          3619 => x"82",
          3620 => x"ff",
          3621 => x"f0",
          3622 => x"bf",
          3623 => x"be",
          3624 => x"a2",
          3625 => x"bd",
          3626 => x"b8",
          3627 => x"b6",
          3628 => x"ff",
          3629 => x"a8",
          3630 => x"39",
          3631 => x"33",
          3632 => x"2e",
          3633 => x"7d",
          3634 => x"78",
          3635 => x"cf",
          3636 => x"ff",
          3637 => x"83",
          3638 => x"d8",
          3639 => x"81",
          3640 => x"2e",
          3641 => x"82",
          3642 => x"7b",
          3643 => x"38",
          3644 => x"7b",
          3645 => x"38",
          3646 => x"82",
          3647 => x"7a",
          3648 => x"d0",
          3649 => x"82",
          3650 => x"b4",
          3651 => x"05",
          3652 => x"af",
          3653 => x"7a",
          3654 => x"ff",
          3655 => x"ca",
          3656 => x"39",
          3657 => x"bf",
          3658 => x"53",
          3659 => x"52",
          3660 => x"b0",
          3661 => x"a4",
          3662 => x"39",
          3663 => x"53",
          3664 => x"52",
          3665 => x"b0",
          3666 => x"a3",
          3667 => x"d6",
          3668 => x"d8",
          3669 => x"56",
          3670 => x"54",
          3671 => x"53",
          3672 => x"52",
          3673 => x"b0",
          3674 => x"cc",
          3675 => x"c8",
          3676 => x"c8",
          3677 => x"30",
          3678 => x"80",
          3679 => x"5b",
          3680 => x"7b",
          3681 => x"38",
          3682 => x"7a",
          3683 => x"80",
          3684 => x"81",
          3685 => x"ff",
          3686 => x"7b",
          3687 => x"7d",
          3688 => x"81",
          3689 => x"78",
          3690 => x"ff",
          3691 => x"06",
          3692 => x"82",
          3693 => x"ff",
          3694 => x"ee",
          3695 => x"3d",
          3696 => x"82",
          3697 => x"87",
          3698 => x"70",
          3699 => x"87",
          3700 => x"72",
          3701 => x"3f",
          3702 => x"08",
          3703 => x"08",
          3704 => x"84",
          3705 => x"51",
          3706 => x"72",
          3707 => x"08",
          3708 => x"87",
          3709 => x"70",
          3710 => x"87",
          3711 => x"72",
          3712 => x"3f",
          3713 => x"08",
          3714 => x"08",
          3715 => x"84",
          3716 => x"51",
          3717 => x"72",
          3718 => x"08",
          3719 => x"8c",
          3720 => x"87",
          3721 => x"0c",
          3722 => x"0b",
          3723 => x"94",
          3724 => x"c0",
          3725 => x"ac",
          3726 => x"84",
          3727 => x"34",
          3728 => x"f4",
          3729 => x"3d",
          3730 => x"0c",
          3731 => x"82",
          3732 => x"54",
          3733 => x"93",
          3734 => x"c0",
          3735 => x"bb",
          3736 => x"c0",
          3737 => x"ba",
          3738 => x"dd",
          3739 => x"e3",
          3740 => x"e8",
          3741 => x"9c",
          3742 => x"fe",
          3743 => x"52",
          3744 => x"88",
          3745 => x"d8",
          3746 => x"c8",
          3747 => x"06",
          3748 => x"14",
          3749 => x"80",
          3750 => x"71",
          3751 => x"0c",
          3752 => x"04",
          3753 => x"76",
          3754 => x"55",
          3755 => x"54",
          3756 => x"81",
          3757 => x"33",
          3758 => x"2e",
          3759 => x"86",
          3760 => x"53",
          3761 => x"33",
          3762 => x"2e",
          3763 => x"86",
          3764 => x"53",
          3765 => x"52",
          3766 => x"09",
          3767 => x"38",
          3768 => x"12",
          3769 => x"33",
          3770 => x"a2",
          3771 => x"81",
          3772 => x"2e",
          3773 => x"ea",
          3774 => x"81",
          3775 => x"72",
          3776 => x"70",
          3777 => x"38",
          3778 => x"80",
          3779 => x"73",
          3780 => x"72",
          3781 => x"70",
          3782 => x"81",
          3783 => x"81",
          3784 => x"32",
          3785 => x"80",
          3786 => x"51",
          3787 => x"80",
          3788 => x"80",
          3789 => x"05",
          3790 => x"75",
          3791 => x"70",
          3792 => x"0c",
          3793 => x"04",
          3794 => x"76",
          3795 => x"80",
          3796 => x"86",
          3797 => x"52",
          3798 => x"a2",
          3799 => x"c8",
          3800 => x"80",
          3801 => x"74",
          3802 => x"d8",
          3803 => x"3d",
          3804 => x"3d",
          3805 => x"11",
          3806 => x"52",
          3807 => x"70",
          3808 => x"98",
          3809 => x"33",
          3810 => x"82",
          3811 => x"26",
          3812 => x"84",
          3813 => x"83",
          3814 => x"26",
          3815 => x"85",
          3816 => x"84",
          3817 => x"26",
          3818 => x"86",
          3819 => x"85",
          3820 => x"26",
          3821 => x"88",
          3822 => x"86",
          3823 => x"e7",
          3824 => x"38",
          3825 => x"54",
          3826 => x"87",
          3827 => x"cc",
          3828 => x"87",
          3829 => x"0c",
          3830 => x"c0",
          3831 => x"82",
          3832 => x"c0",
          3833 => x"83",
          3834 => x"c0",
          3835 => x"84",
          3836 => x"c0",
          3837 => x"85",
          3838 => x"c0",
          3839 => x"86",
          3840 => x"c0",
          3841 => x"74",
          3842 => x"a4",
          3843 => x"c0",
          3844 => x"80",
          3845 => x"98",
          3846 => x"52",
          3847 => x"c8",
          3848 => x"0d",
          3849 => x"0d",
          3850 => x"c0",
          3851 => x"81",
          3852 => x"c0",
          3853 => x"5e",
          3854 => x"87",
          3855 => x"08",
          3856 => x"1c",
          3857 => x"98",
          3858 => x"79",
          3859 => x"87",
          3860 => x"08",
          3861 => x"1c",
          3862 => x"98",
          3863 => x"79",
          3864 => x"87",
          3865 => x"08",
          3866 => x"1c",
          3867 => x"98",
          3868 => x"7b",
          3869 => x"87",
          3870 => x"08",
          3871 => x"1c",
          3872 => x"0c",
          3873 => x"ff",
          3874 => x"83",
          3875 => x"58",
          3876 => x"57",
          3877 => x"56",
          3878 => x"55",
          3879 => x"54",
          3880 => x"53",
          3881 => x"ff",
          3882 => x"c0",
          3883 => x"9a",
          3884 => x"3d",
          3885 => x"3d",
          3886 => x"05",
          3887 => x"e8",
          3888 => x"ff",
          3889 => x"55",
          3890 => x"84",
          3891 => x"2e",
          3892 => x"c0",
          3893 => x"70",
          3894 => x"2a",
          3895 => x"53",
          3896 => x"80",
          3897 => x"71",
          3898 => x"81",
          3899 => x"70",
          3900 => x"81",
          3901 => x"06",
          3902 => x"80",
          3903 => x"71",
          3904 => x"81",
          3905 => x"70",
          3906 => x"73",
          3907 => x"51",
          3908 => x"80",
          3909 => x"2e",
          3910 => x"c0",
          3911 => x"74",
          3912 => x"82",
          3913 => x"87",
          3914 => x"ff",
          3915 => x"8f",
          3916 => x"30",
          3917 => x"51",
          3918 => x"82",
          3919 => x"83",
          3920 => x"f9",
          3921 => x"a7",
          3922 => x"77",
          3923 => x"81",
          3924 => x"7a",
          3925 => x"eb",
          3926 => x"e8",
          3927 => x"ff",
          3928 => x"87",
          3929 => x"53",
          3930 => x"86",
          3931 => x"94",
          3932 => x"08",
          3933 => x"70",
          3934 => x"56",
          3935 => x"2e",
          3936 => x"91",
          3937 => x"06",
          3938 => x"d7",
          3939 => x"32",
          3940 => x"51",
          3941 => x"2e",
          3942 => x"93",
          3943 => x"06",
          3944 => x"ff",
          3945 => x"81",
          3946 => x"87",
          3947 => x"54",
          3948 => x"86",
          3949 => x"94",
          3950 => x"74",
          3951 => x"82",
          3952 => x"89",
          3953 => x"f9",
          3954 => x"54",
          3955 => x"70",
          3956 => x"53",
          3957 => x"77",
          3958 => x"38",
          3959 => x"06",
          3960 => x"d6",
          3961 => x"81",
          3962 => x"57",
          3963 => x"c0",
          3964 => x"75",
          3965 => x"38",
          3966 => x"94",
          3967 => x"70",
          3968 => x"81",
          3969 => x"52",
          3970 => x"8c",
          3971 => x"2a",
          3972 => x"51",
          3973 => x"38",
          3974 => x"70",
          3975 => x"51",
          3976 => x"8d",
          3977 => x"2a",
          3978 => x"51",
          3979 => x"be",
          3980 => x"ff",
          3981 => x"c0",
          3982 => x"70",
          3983 => x"38",
          3984 => x"90",
          3985 => x"0c",
          3986 => x"33",
          3987 => x"06",
          3988 => x"70",
          3989 => x"76",
          3990 => x"0c",
          3991 => x"04",
          3992 => x"82",
          3993 => x"70",
          3994 => x"54",
          3995 => x"94",
          3996 => x"80",
          3997 => x"87",
          3998 => x"51",
          3999 => x"82",
          4000 => x"06",
          4001 => x"70",
          4002 => x"38",
          4003 => x"06",
          4004 => x"94",
          4005 => x"80",
          4006 => x"87",
          4007 => x"52",
          4008 => x"81",
          4009 => x"d8",
          4010 => x"84",
          4011 => x"ff",
          4012 => x"d8",
          4013 => x"ff",
          4014 => x"c8",
          4015 => x"3d",
          4016 => x"e8",
          4017 => x"ff",
          4018 => x"87",
          4019 => x"52",
          4020 => x"86",
          4021 => x"94",
          4022 => x"08",
          4023 => x"70",
          4024 => x"51",
          4025 => x"70",
          4026 => x"38",
          4027 => x"06",
          4028 => x"94",
          4029 => x"80",
          4030 => x"87",
          4031 => x"52",
          4032 => x"98",
          4033 => x"2c",
          4034 => x"71",
          4035 => x"0c",
          4036 => x"04",
          4037 => x"87",
          4038 => x"08",
          4039 => x"8a",
          4040 => x"70",
          4041 => x"b4",
          4042 => x"9e",
          4043 => x"d6",
          4044 => x"c0",
          4045 => x"82",
          4046 => x"87",
          4047 => x"08",
          4048 => x"0c",
          4049 => x"98",
          4050 => x"f8",
          4051 => x"9e",
          4052 => x"d6",
          4053 => x"c0",
          4054 => x"82",
          4055 => x"87",
          4056 => x"08",
          4057 => x"0c",
          4058 => x"b0",
          4059 => x"88",
          4060 => x"9e",
          4061 => x"d7",
          4062 => x"c0",
          4063 => x"82",
          4064 => x"87",
          4065 => x"08",
          4066 => x"0c",
          4067 => x"c0",
          4068 => x"98",
          4069 => x"9e",
          4070 => x"d7",
          4071 => x"c0",
          4072 => x"51",
          4073 => x"a0",
          4074 => x"9e",
          4075 => x"d7",
          4076 => x"c0",
          4077 => x"82",
          4078 => x"87",
          4079 => x"08",
          4080 => x"0c",
          4081 => x"d7",
          4082 => x"0b",
          4083 => x"90",
          4084 => x"80",
          4085 => x"52",
          4086 => x"2e",
          4087 => x"52",
          4088 => x"b1",
          4089 => x"87",
          4090 => x"08",
          4091 => x"0a",
          4092 => x"52",
          4093 => x"83",
          4094 => x"71",
          4095 => x"34",
          4096 => x"c0",
          4097 => x"70",
          4098 => x"06",
          4099 => x"70",
          4100 => x"38",
          4101 => x"82",
          4102 => x"80",
          4103 => x"9e",
          4104 => x"88",
          4105 => x"51",
          4106 => x"80",
          4107 => x"81",
          4108 => x"d7",
          4109 => x"0b",
          4110 => x"90",
          4111 => x"80",
          4112 => x"52",
          4113 => x"2e",
          4114 => x"52",
          4115 => x"b5",
          4116 => x"87",
          4117 => x"08",
          4118 => x"80",
          4119 => x"52",
          4120 => x"83",
          4121 => x"71",
          4122 => x"34",
          4123 => x"c0",
          4124 => x"70",
          4125 => x"06",
          4126 => x"70",
          4127 => x"38",
          4128 => x"82",
          4129 => x"80",
          4130 => x"9e",
          4131 => x"82",
          4132 => x"51",
          4133 => x"80",
          4134 => x"81",
          4135 => x"d7",
          4136 => x"0b",
          4137 => x"90",
          4138 => x"80",
          4139 => x"52",
          4140 => x"2e",
          4141 => x"52",
          4142 => x"b9",
          4143 => x"87",
          4144 => x"08",
          4145 => x"80",
          4146 => x"52",
          4147 => x"83",
          4148 => x"71",
          4149 => x"34",
          4150 => x"c0",
          4151 => x"70",
          4152 => x"51",
          4153 => x"80",
          4154 => x"81",
          4155 => x"d7",
          4156 => x"c0",
          4157 => x"70",
          4158 => x"70",
          4159 => x"51",
          4160 => x"d7",
          4161 => x"0b",
          4162 => x"90",
          4163 => x"80",
          4164 => x"52",
          4165 => x"83",
          4166 => x"71",
          4167 => x"34",
          4168 => x"90",
          4169 => x"f0",
          4170 => x"2a",
          4171 => x"70",
          4172 => x"34",
          4173 => x"c0",
          4174 => x"70",
          4175 => x"52",
          4176 => x"2e",
          4177 => x"52",
          4178 => x"bf",
          4179 => x"9e",
          4180 => x"87",
          4181 => x"70",
          4182 => x"34",
          4183 => x"04",
          4184 => x"82",
          4185 => x"ff",
          4186 => x"82",
          4187 => x"54",
          4188 => x"89",
          4189 => x"d8",
          4190 => x"df",
          4191 => x"ec",
          4192 => x"e2",
          4193 => x"b2",
          4194 => x"80",
          4195 => x"82",
          4196 => x"82",
          4197 => x"11",
          4198 => x"c1",
          4199 => x"90",
          4200 => x"d7",
          4201 => x"73",
          4202 => x"38",
          4203 => x"08",
          4204 => x"08",
          4205 => x"82",
          4206 => x"ff",
          4207 => x"82",
          4208 => x"54",
          4209 => x"94",
          4210 => x"ec",
          4211 => x"f0",
          4212 => x"52",
          4213 => x"51",
          4214 => x"3f",
          4215 => x"33",
          4216 => x"2e",
          4217 => x"d6",
          4218 => x"d6",
          4219 => x"54",
          4220 => x"d8",
          4221 => x"e3",
          4222 => x"b6",
          4223 => x"80",
          4224 => x"82",
          4225 => x"82",
          4226 => x"11",
          4227 => x"c1",
          4228 => x"8f",
          4229 => x"d7",
          4230 => x"73",
          4231 => x"38",
          4232 => x"33",
          4233 => x"90",
          4234 => x"af",
          4235 => x"bf",
          4236 => x"80",
          4237 => x"82",
          4238 => x"52",
          4239 => x"51",
          4240 => x"3f",
          4241 => x"33",
          4242 => x"2e",
          4243 => x"d7",
          4244 => x"82",
          4245 => x"ff",
          4246 => x"82",
          4247 => x"54",
          4248 => x"89",
          4249 => x"f0",
          4250 => x"fa",
          4251 => x"b3",
          4252 => x"80",
          4253 => x"82",
          4254 => x"ff",
          4255 => x"82",
          4256 => x"54",
          4257 => x"89",
          4258 => x"90",
          4259 => x"d6",
          4260 => x"b9",
          4261 => x"80",
          4262 => x"82",
          4263 => x"ff",
          4264 => x"82",
          4265 => x"54",
          4266 => x"89",
          4267 => x"a4",
          4268 => x"b2",
          4269 => x"ac",
          4270 => x"aa",
          4271 => x"94",
          4272 => x"c3",
          4273 => x"8e",
          4274 => x"d7",
          4275 => x"82",
          4276 => x"ff",
          4277 => x"82",
          4278 => x"52",
          4279 => x"51",
          4280 => x"3f",
          4281 => x"51",
          4282 => x"3f",
          4283 => x"22",
          4284 => x"b8",
          4285 => x"e3",
          4286 => x"a4",
          4287 => x"84",
          4288 => x"51",
          4289 => x"82",
          4290 => x"bd",
          4291 => x"76",
          4292 => x"54",
          4293 => x"08",
          4294 => x"e0",
          4295 => x"bb",
          4296 => x"b7",
          4297 => x"80",
          4298 => x"82",
          4299 => x"56",
          4300 => x"52",
          4301 => x"ce",
          4302 => x"c8",
          4303 => x"c0",
          4304 => x"31",
          4305 => x"d8",
          4306 => x"82",
          4307 => x"ff",
          4308 => x"82",
          4309 => x"54",
          4310 => x"a9",
          4311 => x"ac",
          4312 => x"84",
          4313 => x"51",
          4314 => x"82",
          4315 => x"bd",
          4316 => x"76",
          4317 => x"54",
          4318 => x"08",
          4319 => x"b8",
          4320 => x"d7",
          4321 => x"ff",
          4322 => x"87",
          4323 => x"fe",
          4324 => x"92",
          4325 => x"05",
          4326 => x"26",
          4327 => x"84",
          4328 => x"c4",
          4329 => x"08",
          4330 => x"e4",
          4331 => x"82",
          4332 => x"97",
          4333 => x"f4",
          4334 => x"82",
          4335 => x"8b",
          4336 => x"80",
          4337 => x"82",
          4338 => x"ff",
          4339 => x"84",
          4340 => x"71",
          4341 => x"04",
          4342 => x"87",
          4343 => x"70",
          4344 => x"80",
          4345 => x"74",
          4346 => x"d7",
          4347 => x"0c",
          4348 => x"04",
          4349 => x"87",
          4350 => x"70",
          4351 => x"c4",
          4352 => x"72",
          4353 => x"70",
          4354 => x"08",
          4355 => x"d7",
          4356 => x"0c",
          4357 => x"0d",
          4358 => x"87",
          4359 => x"0c",
          4360 => x"c4",
          4361 => x"96",
          4362 => x"fd",
          4363 => x"98",
          4364 => x"2c",
          4365 => x"70",
          4366 => x"10",
          4367 => x"2b",
          4368 => x"54",
          4369 => x"0b",
          4370 => x"12",
          4371 => x"71",
          4372 => x"38",
          4373 => x"11",
          4374 => x"84",
          4375 => x"33",
          4376 => x"52",
          4377 => x"2e",
          4378 => x"83",
          4379 => x"72",
          4380 => x"0c",
          4381 => x"04",
          4382 => x"79",
          4383 => x"a3",
          4384 => x"33",
          4385 => x"72",
          4386 => x"38",
          4387 => x"08",
          4388 => x"ff",
          4389 => x"82",
          4390 => x"52",
          4391 => x"aa",
          4392 => x"f4",
          4393 => x"88",
          4394 => x"89",
          4395 => x"ff",
          4396 => x"74",
          4397 => x"ff",
          4398 => x"39",
          4399 => x"8a",
          4400 => x"74",
          4401 => x"0d",
          4402 => x"0d",
          4403 => x"05",
          4404 => x"02",
          4405 => x"05",
          4406 => x"a0",
          4407 => x"29",
          4408 => x"05",
          4409 => x"59",
          4410 => x"59",
          4411 => x"86",
          4412 => x"9a",
          4413 => x"d8",
          4414 => x"84",
          4415 => x"c8",
          4416 => x"70",
          4417 => x"5a",
          4418 => x"82",
          4419 => x"75",
          4420 => x"a0",
          4421 => x"29",
          4422 => x"05",
          4423 => x"56",
          4424 => x"2e",
          4425 => x"53",
          4426 => x"51",
          4427 => x"3f",
          4428 => x"33",
          4429 => x"74",
          4430 => x"34",
          4431 => x"06",
          4432 => x"27",
          4433 => x"0b",
          4434 => x"34",
          4435 => x"b6",
          4436 => x"9c",
          4437 => x"80",
          4438 => x"82",
          4439 => x"55",
          4440 => x"8c",
          4441 => x"54",
          4442 => x"52",
          4443 => x"eb",
          4444 => x"d8",
          4445 => x"8a",
          4446 => x"e7",
          4447 => x"9c",
          4448 => x"ef",
          4449 => x"3d",
          4450 => x"3d",
          4451 => x"c8",
          4452 => x"72",
          4453 => x"80",
          4454 => x"71",
          4455 => x"3f",
          4456 => x"ff",
          4457 => x"54",
          4458 => x"25",
          4459 => x"0b",
          4460 => x"34",
          4461 => x"08",
          4462 => x"2e",
          4463 => x"51",
          4464 => x"3f",
          4465 => x"08",
          4466 => x"3f",
          4467 => x"d8",
          4468 => x"3d",
          4469 => x"3d",
          4470 => x"80",
          4471 => x"9c",
          4472 => x"f5",
          4473 => x"d8",
          4474 => x"d3",
          4475 => x"9c",
          4476 => x"f8",
          4477 => x"70",
          4478 => x"9d",
          4479 => x"d8",
          4480 => x"2e",
          4481 => x"51",
          4482 => x"3f",
          4483 => x"08",
          4484 => x"82",
          4485 => x"25",
          4486 => x"d8",
          4487 => x"05",
          4488 => x"55",
          4489 => x"75",
          4490 => x"81",
          4491 => x"84",
          4492 => x"87",
          4493 => x"ff",
          4494 => x"06",
          4495 => x"a6",
          4496 => x"d9",
          4497 => x"3d",
          4498 => x"08",
          4499 => x"70",
          4500 => x"52",
          4501 => x"08",
          4502 => x"ab",
          4503 => x"c8",
          4504 => x"38",
          4505 => x"d8",
          4506 => x"55",
          4507 => x"8b",
          4508 => x"56",
          4509 => x"3f",
          4510 => x"08",
          4511 => x"38",
          4512 => x"af",
          4513 => x"d8",
          4514 => x"18",
          4515 => x"0b",
          4516 => x"08",
          4517 => x"82",
          4518 => x"ff",
          4519 => x"55",
          4520 => x"34",
          4521 => x"30",
          4522 => x"9f",
          4523 => x"55",
          4524 => x"85",
          4525 => x"ac",
          4526 => x"9c",
          4527 => x"08",
          4528 => x"f3",
          4529 => x"d8",
          4530 => x"2e",
          4531 => x"c9",
          4532 => x"86",
          4533 => x"77",
          4534 => x"06",
          4535 => x"52",
          4536 => x"af",
          4537 => x"51",
          4538 => x"3f",
          4539 => x"54",
          4540 => x"08",
          4541 => x"58",
          4542 => x"c8",
          4543 => x"0d",
          4544 => x"0d",
          4545 => x"5c",
          4546 => x"57",
          4547 => x"73",
          4548 => x"81",
          4549 => x"78",
          4550 => x"56",
          4551 => x"98",
          4552 => x"70",
          4553 => x"33",
          4554 => x"73",
          4555 => x"81",
          4556 => x"75",
          4557 => x"38",
          4558 => x"88",
          4559 => x"a4",
          4560 => x"52",
          4561 => x"c0",
          4562 => x"c8",
          4563 => x"52",
          4564 => x"ff",
          4565 => x"82",
          4566 => x"80",
          4567 => x"15",
          4568 => x"81",
          4569 => x"74",
          4570 => x"38",
          4571 => x"e6",
          4572 => x"81",
          4573 => x"3d",
          4574 => x"f8",
          4575 => x"cf",
          4576 => x"c8",
          4577 => x"9a",
          4578 => x"53",
          4579 => x"51",
          4580 => x"82",
          4581 => x"81",
          4582 => x"74",
          4583 => x"54",
          4584 => x"14",
          4585 => x"06",
          4586 => x"74",
          4587 => x"38",
          4588 => x"82",
          4589 => x"8c",
          4590 => x"d3",
          4591 => x"3d",
          4592 => x"08",
          4593 => x"59",
          4594 => x"0b",
          4595 => x"82",
          4596 => x"82",
          4597 => x"55",
          4598 => x"cb",
          4599 => x"d8",
          4600 => x"55",
          4601 => x"81",
          4602 => x"2e",
          4603 => x"81",
          4604 => x"55",
          4605 => x"2e",
          4606 => x"a8",
          4607 => x"3f",
          4608 => x"08",
          4609 => x"0c",
          4610 => x"08",
          4611 => x"92",
          4612 => x"76",
          4613 => x"c8",
          4614 => x"de",
          4615 => x"d8",
          4616 => x"2e",
          4617 => x"c9",
          4618 => x"9f",
          4619 => x"f7",
          4620 => x"c8",
          4621 => x"d8",
          4622 => x"80",
          4623 => x"3d",
          4624 => x"81",
          4625 => x"82",
          4626 => x"56",
          4627 => x"08",
          4628 => x"81",
          4629 => x"38",
          4630 => x"08",
          4631 => x"a8",
          4632 => x"c8",
          4633 => x"0b",
          4634 => x"08",
          4635 => x"82",
          4636 => x"ff",
          4637 => x"55",
          4638 => x"34",
          4639 => x"81",
          4640 => x"75",
          4641 => x"3f",
          4642 => x"81",
          4643 => x"54",
          4644 => x"83",
          4645 => x"74",
          4646 => x"81",
          4647 => x"38",
          4648 => x"82",
          4649 => x"76",
          4650 => x"d8",
          4651 => x"2e",
          4652 => x"d6",
          4653 => x"5d",
          4654 => x"82",
          4655 => x"98",
          4656 => x"2c",
          4657 => x"ff",
          4658 => x"78",
          4659 => x"82",
          4660 => x"70",
          4661 => x"98",
          4662 => x"80",
          4663 => x"2b",
          4664 => x"71",
          4665 => x"70",
          4666 => x"c6",
          4667 => x"08",
          4668 => x"51",
          4669 => x"59",
          4670 => x"5d",
          4671 => x"73",
          4672 => x"e9",
          4673 => x"27",
          4674 => x"81",
          4675 => x"81",
          4676 => x"70",
          4677 => x"55",
          4678 => x"80",
          4679 => x"53",
          4680 => x"51",
          4681 => x"82",
          4682 => x"81",
          4683 => x"73",
          4684 => x"38",
          4685 => x"80",
          4686 => x"b1",
          4687 => x"80",
          4688 => x"80",
          4689 => x"98",
          4690 => x"ff",
          4691 => x"55",
          4692 => x"97",
          4693 => x"74",
          4694 => x"f5",
          4695 => x"d8",
          4696 => x"ff",
          4697 => x"cc",
          4698 => x"80",
          4699 => x"2e",
          4700 => x"81",
          4701 => x"82",
          4702 => x"74",
          4703 => x"98",
          4704 => x"80",
          4705 => x"2b",
          4706 => x"70",
          4707 => x"82",
          4708 => x"94",
          4709 => x"51",
          4710 => x"58",
          4711 => x"77",
          4712 => x"06",
          4713 => x"82",
          4714 => x"08",
          4715 => x"0b",
          4716 => x"34",
          4717 => x"f0",
          4718 => x"39",
          4719 => x"84",
          4720 => x"f0",
          4721 => x"af",
          4722 => x"7d",
          4723 => x"73",
          4724 => x"e1",
          4725 => x"29",
          4726 => x"05",
          4727 => x"04",
          4728 => x"33",
          4729 => x"2e",
          4730 => x"82",
          4731 => x"55",
          4732 => x"ab",
          4733 => x"2b",
          4734 => x"51",
          4735 => x"24",
          4736 => x"1a",
          4737 => x"81",
          4738 => x"81",
          4739 => x"81",
          4740 => x"70",
          4741 => x"f0",
          4742 => x"51",
          4743 => x"82",
          4744 => x"81",
          4745 => x"74",
          4746 => x"34",
          4747 => x"ae",
          4748 => x"34",
          4749 => x"33",
          4750 => x"25",
          4751 => x"14",
          4752 => x"f0",
          4753 => x"f0",
          4754 => x"81",
          4755 => x"81",
          4756 => x"70",
          4757 => x"f0",
          4758 => x"51",
          4759 => x"77",
          4760 => x"82",
          4761 => x"52",
          4762 => x"33",
          4763 => x"9e",
          4764 => x"81",
          4765 => x"81",
          4766 => x"70",
          4767 => x"f0",
          4768 => x"51",
          4769 => x"24",
          4770 => x"f0",
          4771 => x"98",
          4772 => x"2c",
          4773 => x"33",
          4774 => x"56",
          4775 => x"fc",
          4776 => x"f4",
          4777 => x"88",
          4778 => x"89",
          4779 => x"80",
          4780 => x"80",
          4781 => x"98",
          4782 => x"88",
          4783 => x"55",
          4784 => x"de",
          4785 => x"39",
          4786 => x"80",
          4787 => x"34",
          4788 => x"53",
          4789 => x"b8",
          4790 => x"9c",
          4791 => x"39",
          4792 => x"33",
          4793 => x"06",
          4794 => x"80",
          4795 => x"38",
          4796 => x"33",
          4797 => x"73",
          4798 => x"34",
          4799 => x"73",
          4800 => x"34",
          4801 => x"08",
          4802 => x"ff",
          4803 => x"82",
          4804 => x"70",
          4805 => x"98",
          4806 => x"88",
          4807 => x"56",
          4808 => x"25",
          4809 => x"1a",
          4810 => x"33",
          4811 => x"f4",
          4812 => x"73",
          4813 => x"9c",
          4814 => x"81",
          4815 => x"81",
          4816 => x"70",
          4817 => x"f0",
          4818 => x"51",
          4819 => x"24",
          4820 => x"f4",
          4821 => x"a0",
          4822 => x"d9",
          4823 => x"8c",
          4824 => x"2b",
          4825 => x"82",
          4826 => x"57",
          4827 => x"74",
          4828 => x"c1",
          4829 => x"ac",
          4830 => x"51",
          4831 => x"3f",
          4832 => x"0a",
          4833 => x"0a",
          4834 => x"2c",
          4835 => x"33",
          4836 => x"75",
          4837 => x"38",
          4838 => x"82",
          4839 => x"7a",
          4840 => x"74",
          4841 => x"ac",
          4842 => x"51",
          4843 => x"3f",
          4844 => x"52",
          4845 => x"c9",
          4846 => x"c8",
          4847 => x"06",
          4848 => x"38",
          4849 => x"33",
          4850 => x"2e",
          4851 => x"53",
          4852 => x"51",
          4853 => x"84",
          4854 => x"34",
          4855 => x"f0",
          4856 => x"0b",
          4857 => x"34",
          4858 => x"c8",
          4859 => x"0d",
          4860 => x"8c",
          4861 => x"80",
          4862 => x"38",
          4863 => x"08",
          4864 => x"ff",
          4865 => x"82",
          4866 => x"ff",
          4867 => x"82",
          4868 => x"73",
          4869 => x"54",
          4870 => x"f0",
          4871 => x"f0",
          4872 => x"55",
          4873 => x"f9",
          4874 => x"14",
          4875 => x"f0",
          4876 => x"98",
          4877 => x"2c",
          4878 => x"06",
          4879 => x"74",
          4880 => x"38",
          4881 => x"81",
          4882 => x"34",
          4883 => x"08",
          4884 => x"51",
          4885 => x"3f",
          4886 => x"0a",
          4887 => x"0a",
          4888 => x"2c",
          4889 => x"33",
          4890 => x"75",
          4891 => x"38",
          4892 => x"08",
          4893 => x"ff",
          4894 => x"82",
          4895 => x"70",
          4896 => x"98",
          4897 => x"88",
          4898 => x"56",
          4899 => x"24",
          4900 => x"82",
          4901 => x"52",
          4902 => x"9a",
          4903 => x"81",
          4904 => x"81",
          4905 => x"70",
          4906 => x"f0",
          4907 => x"51",
          4908 => x"25",
          4909 => x"fd",
          4910 => x"8c",
          4911 => x"ff",
          4912 => x"88",
          4913 => x"54",
          4914 => x"f7",
          4915 => x"f4",
          4916 => x"81",
          4917 => x"82",
          4918 => x"74",
          4919 => x"52",
          4920 => x"d1",
          4921 => x"8c",
          4922 => x"ff",
          4923 => x"88",
          4924 => x"54",
          4925 => x"d6",
          4926 => x"39",
          4927 => x"53",
          4928 => x"b8",
          4929 => x"f0",
          4930 => x"82",
          4931 => x"80",
          4932 => x"88",
          4933 => x"39",
          4934 => x"82",
          4935 => x"55",
          4936 => x"a6",
          4937 => x"ff",
          4938 => x"82",
          4939 => x"82",
          4940 => x"82",
          4941 => x"81",
          4942 => x"05",
          4943 => x"79",
          4944 => x"a4",
          4945 => x"81",
          4946 => x"84",
          4947 => x"c8",
          4948 => x"08",
          4949 => x"80",
          4950 => x"74",
          4951 => x"a8",
          4952 => x"c8",
          4953 => x"88",
          4954 => x"c8",
          4955 => x"06",
          4956 => x"74",
          4957 => x"ff",
          4958 => x"ff",
          4959 => x"fa",
          4960 => x"55",
          4961 => x"f6",
          4962 => x"51",
          4963 => x"3f",
          4964 => x"93",
          4965 => x"06",
          4966 => x"d7",
          4967 => x"74",
          4968 => x"38",
          4969 => x"a0",
          4970 => x"d8",
          4971 => x"f0",
          4972 => x"d8",
          4973 => x"ff",
          4974 => x"53",
          4975 => x"51",
          4976 => x"3f",
          4977 => x"7a",
          4978 => x"d7",
          4979 => x"08",
          4980 => x"80",
          4981 => x"74",
          4982 => x"ac",
          4983 => x"c8",
          4984 => x"88",
          4985 => x"c8",
          4986 => x"06",
          4987 => x"74",
          4988 => x"ff",
          4989 => x"81",
          4990 => x"81",
          4991 => x"89",
          4992 => x"f0",
          4993 => x"7a",
          4994 => x"8c",
          4995 => x"88",
          4996 => x"51",
          4997 => x"f5",
          4998 => x"f0",
          4999 => x"81",
          5000 => x"f0",
          5001 => x"56",
          5002 => x"27",
          5003 => x"82",
          5004 => x"52",
          5005 => x"73",
          5006 => x"34",
          5007 => x"33",
          5008 => x"96",
          5009 => x"ed",
          5010 => x"8c",
          5011 => x"80",
          5012 => x"38",
          5013 => x"08",
          5014 => x"ff",
          5015 => x"82",
          5016 => x"ff",
          5017 => x"82",
          5018 => x"f4",
          5019 => x"3d",
          5020 => x"80",
          5021 => x"c0",
          5022 => x"0b",
          5023 => x"23",
          5024 => x"80",
          5025 => x"80",
          5026 => x"dd",
          5027 => x"c0",
          5028 => x"58",
          5029 => x"81",
          5030 => x"15",
          5031 => x"c0",
          5032 => x"84",
          5033 => x"85",
          5034 => x"d8",
          5035 => x"77",
          5036 => x"76",
          5037 => x"82",
          5038 => x"82",
          5039 => x"ff",
          5040 => x"80",
          5041 => x"ff",
          5042 => x"88",
          5043 => x"55",
          5044 => x"17",
          5045 => x"17",
          5046 => x"bc",
          5047 => x"29",
          5048 => x"08",
          5049 => x"51",
          5050 => x"82",
          5051 => x"83",
          5052 => x"3d",
          5053 => x"3d",
          5054 => x"81",
          5055 => x"27",
          5056 => x"12",
          5057 => x"11",
          5058 => x"ff",
          5059 => x"51",
          5060 => x"c8",
          5061 => x"0d",
          5062 => x"0d",
          5063 => x"22",
          5064 => x"aa",
          5065 => x"05",
          5066 => x"08",
          5067 => x"71",
          5068 => x"2b",
          5069 => x"33",
          5070 => x"71",
          5071 => x"02",
          5072 => x"05",
          5073 => x"ff",
          5074 => x"70",
          5075 => x"51",
          5076 => x"5b",
          5077 => x"54",
          5078 => x"34",
          5079 => x"34",
          5080 => x"08",
          5081 => x"2a",
          5082 => x"82",
          5083 => x"83",
          5084 => x"d8",
          5085 => x"17",
          5086 => x"12",
          5087 => x"2b",
          5088 => x"2b",
          5089 => x"06",
          5090 => x"52",
          5091 => x"83",
          5092 => x"70",
          5093 => x"54",
          5094 => x"12",
          5095 => x"ff",
          5096 => x"83",
          5097 => x"d8",
          5098 => x"56",
          5099 => x"72",
          5100 => x"89",
          5101 => x"fb",
          5102 => x"d8",
          5103 => x"84",
          5104 => x"22",
          5105 => x"72",
          5106 => x"33",
          5107 => x"71",
          5108 => x"83",
          5109 => x"5b",
          5110 => x"52",
          5111 => x"12",
          5112 => x"33",
          5113 => x"07",
          5114 => x"54",
          5115 => x"70",
          5116 => x"73",
          5117 => x"82",
          5118 => x"70",
          5119 => x"33",
          5120 => x"71",
          5121 => x"83",
          5122 => x"59",
          5123 => x"05",
          5124 => x"87",
          5125 => x"88",
          5126 => x"88",
          5127 => x"56",
          5128 => x"13",
          5129 => x"13",
          5130 => x"c0",
          5131 => x"33",
          5132 => x"71",
          5133 => x"70",
          5134 => x"06",
          5135 => x"53",
          5136 => x"53",
          5137 => x"70",
          5138 => x"87",
          5139 => x"fa",
          5140 => x"a2",
          5141 => x"d8",
          5142 => x"83",
          5143 => x"70",
          5144 => x"33",
          5145 => x"07",
          5146 => x"15",
          5147 => x"12",
          5148 => x"2b",
          5149 => x"07",
          5150 => x"55",
          5151 => x"57",
          5152 => x"80",
          5153 => x"38",
          5154 => x"ab",
          5155 => x"c0",
          5156 => x"70",
          5157 => x"33",
          5158 => x"71",
          5159 => x"74",
          5160 => x"81",
          5161 => x"88",
          5162 => x"83",
          5163 => x"f8",
          5164 => x"54",
          5165 => x"58",
          5166 => x"74",
          5167 => x"52",
          5168 => x"34",
          5169 => x"34",
          5170 => x"08",
          5171 => x"33",
          5172 => x"71",
          5173 => x"83",
          5174 => x"59",
          5175 => x"05",
          5176 => x"12",
          5177 => x"2b",
          5178 => x"ff",
          5179 => x"88",
          5180 => x"52",
          5181 => x"74",
          5182 => x"15",
          5183 => x"0d",
          5184 => x"0d",
          5185 => x"08",
          5186 => x"9e",
          5187 => x"83",
          5188 => x"82",
          5189 => x"12",
          5190 => x"2b",
          5191 => x"07",
          5192 => x"52",
          5193 => x"05",
          5194 => x"13",
          5195 => x"2b",
          5196 => x"05",
          5197 => x"71",
          5198 => x"2a",
          5199 => x"53",
          5200 => x"34",
          5201 => x"34",
          5202 => x"08",
          5203 => x"33",
          5204 => x"71",
          5205 => x"83",
          5206 => x"59",
          5207 => x"05",
          5208 => x"83",
          5209 => x"88",
          5210 => x"88",
          5211 => x"56",
          5212 => x"13",
          5213 => x"13",
          5214 => x"c0",
          5215 => x"11",
          5216 => x"33",
          5217 => x"07",
          5218 => x"0c",
          5219 => x"3d",
          5220 => x"3d",
          5221 => x"d8",
          5222 => x"83",
          5223 => x"ff",
          5224 => x"53",
          5225 => x"a7",
          5226 => x"c0",
          5227 => x"2b",
          5228 => x"11",
          5229 => x"33",
          5230 => x"71",
          5231 => x"75",
          5232 => x"81",
          5233 => x"98",
          5234 => x"2b",
          5235 => x"40",
          5236 => x"58",
          5237 => x"72",
          5238 => x"38",
          5239 => x"52",
          5240 => x"9d",
          5241 => x"39",
          5242 => x"85",
          5243 => x"8b",
          5244 => x"2b",
          5245 => x"79",
          5246 => x"51",
          5247 => x"76",
          5248 => x"75",
          5249 => x"56",
          5250 => x"34",
          5251 => x"08",
          5252 => x"12",
          5253 => x"33",
          5254 => x"07",
          5255 => x"54",
          5256 => x"53",
          5257 => x"34",
          5258 => x"34",
          5259 => x"08",
          5260 => x"0b",
          5261 => x"80",
          5262 => x"34",
          5263 => x"08",
          5264 => x"14",
          5265 => x"14",
          5266 => x"c0",
          5267 => x"33",
          5268 => x"71",
          5269 => x"70",
          5270 => x"07",
          5271 => x"53",
          5272 => x"54",
          5273 => x"72",
          5274 => x"8b",
          5275 => x"ff",
          5276 => x"52",
          5277 => x"08",
          5278 => x"f2",
          5279 => x"2e",
          5280 => x"51",
          5281 => x"83",
          5282 => x"f5",
          5283 => x"7e",
          5284 => x"e2",
          5285 => x"c8",
          5286 => x"ff",
          5287 => x"c0",
          5288 => x"33",
          5289 => x"71",
          5290 => x"70",
          5291 => x"58",
          5292 => x"ff",
          5293 => x"2e",
          5294 => x"75",
          5295 => x"70",
          5296 => x"33",
          5297 => x"07",
          5298 => x"ff",
          5299 => x"70",
          5300 => x"06",
          5301 => x"52",
          5302 => x"59",
          5303 => x"27",
          5304 => x"80",
          5305 => x"75",
          5306 => x"84",
          5307 => x"16",
          5308 => x"2b",
          5309 => x"75",
          5310 => x"81",
          5311 => x"85",
          5312 => x"59",
          5313 => x"83",
          5314 => x"c0",
          5315 => x"33",
          5316 => x"71",
          5317 => x"70",
          5318 => x"06",
          5319 => x"56",
          5320 => x"75",
          5321 => x"81",
          5322 => x"79",
          5323 => x"cc",
          5324 => x"74",
          5325 => x"c4",
          5326 => x"2e",
          5327 => x"89",
          5328 => x"f8",
          5329 => x"ac",
          5330 => x"80",
          5331 => x"75",
          5332 => x"3f",
          5333 => x"08",
          5334 => x"11",
          5335 => x"33",
          5336 => x"71",
          5337 => x"53",
          5338 => x"74",
          5339 => x"70",
          5340 => x"06",
          5341 => x"5c",
          5342 => x"78",
          5343 => x"76",
          5344 => x"57",
          5345 => x"34",
          5346 => x"08",
          5347 => x"71",
          5348 => x"86",
          5349 => x"12",
          5350 => x"2b",
          5351 => x"2a",
          5352 => x"53",
          5353 => x"73",
          5354 => x"75",
          5355 => x"82",
          5356 => x"70",
          5357 => x"33",
          5358 => x"71",
          5359 => x"83",
          5360 => x"5d",
          5361 => x"05",
          5362 => x"15",
          5363 => x"15",
          5364 => x"c0",
          5365 => x"71",
          5366 => x"33",
          5367 => x"71",
          5368 => x"70",
          5369 => x"5a",
          5370 => x"54",
          5371 => x"34",
          5372 => x"34",
          5373 => x"08",
          5374 => x"54",
          5375 => x"c8",
          5376 => x"0d",
          5377 => x"0d",
          5378 => x"d8",
          5379 => x"38",
          5380 => x"71",
          5381 => x"2e",
          5382 => x"51",
          5383 => x"82",
          5384 => x"53",
          5385 => x"c8",
          5386 => x"0d",
          5387 => x"0d",
          5388 => x"5c",
          5389 => x"40",
          5390 => x"08",
          5391 => x"81",
          5392 => x"f4",
          5393 => x"8e",
          5394 => x"ff",
          5395 => x"d8",
          5396 => x"83",
          5397 => x"8b",
          5398 => x"fc",
          5399 => x"54",
          5400 => x"7e",
          5401 => x"3f",
          5402 => x"08",
          5403 => x"06",
          5404 => x"08",
          5405 => x"83",
          5406 => x"ff",
          5407 => x"83",
          5408 => x"70",
          5409 => x"33",
          5410 => x"07",
          5411 => x"70",
          5412 => x"06",
          5413 => x"fc",
          5414 => x"29",
          5415 => x"81",
          5416 => x"88",
          5417 => x"90",
          5418 => x"4e",
          5419 => x"52",
          5420 => x"41",
          5421 => x"5b",
          5422 => x"8f",
          5423 => x"ff",
          5424 => x"31",
          5425 => x"ff",
          5426 => x"82",
          5427 => x"17",
          5428 => x"2b",
          5429 => x"29",
          5430 => x"81",
          5431 => x"98",
          5432 => x"2b",
          5433 => x"45",
          5434 => x"73",
          5435 => x"38",
          5436 => x"70",
          5437 => x"06",
          5438 => x"7b",
          5439 => x"38",
          5440 => x"73",
          5441 => x"81",
          5442 => x"78",
          5443 => x"3f",
          5444 => x"ff",
          5445 => x"e5",
          5446 => x"38",
          5447 => x"89",
          5448 => x"f6",
          5449 => x"a5",
          5450 => x"55",
          5451 => x"80",
          5452 => x"1d",
          5453 => x"83",
          5454 => x"88",
          5455 => x"57",
          5456 => x"3f",
          5457 => x"51",
          5458 => x"82",
          5459 => x"83",
          5460 => x"7e",
          5461 => x"70",
          5462 => x"d8",
          5463 => x"84",
          5464 => x"59",
          5465 => x"3f",
          5466 => x"08",
          5467 => x"75",
          5468 => x"06",
          5469 => x"85",
          5470 => x"54",
          5471 => x"80",
          5472 => x"51",
          5473 => x"82",
          5474 => x"1d",
          5475 => x"83",
          5476 => x"88",
          5477 => x"43",
          5478 => x"3f",
          5479 => x"51",
          5480 => x"82",
          5481 => x"83",
          5482 => x"7e",
          5483 => x"70",
          5484 => x"d8",
          5485 => x"84",
          5486 => x"59",
          5487 => x"3f",
          5488 => x"08",
          5489 => x"60",
          5490 => x"55",
          5491 => x"ff",
          5492 => x"a9",
          5493 => x"52",
          5494 => x"3f",
          5495 => x"08",
          5496 => x"c8",
          5497 => x"93",
          5498 => x"73",
          5499 => x"c8",
          5500 => x"91",
          5501 => x"51",
          5502 => x"7a",
          5503 => x"27",
          5504 => x"53",
          5505 => x"51",
          5506 => x"7a",
          5507 => x"82",
          5508 => x"05",
          5509 => x"f6",
          5510 => x"54",
          5511 => x"c8",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"70",
          5515 => x"d5",
          5516 => x"c8",
          5517 => x"d8",
          5518 => x"2e",
          5519 => x"53",
          5520 => x"d8",
          5521 => x"ff",
          5522 => x"74",
          5523 => x"0c",
          5524 => x"04",
          5525 => x"02",
          5526 => x"51",
          5527 => x"72",
          5528 => x"82",
          5529 => x"33",
          5530 => x"d8",
          5531 => x"3d",
          5532 => x"3d",
          5533 => x"05",
          5534 => x"05",
          5535 => x"56",
          5536 => x"72",
          5537 => x"e0",
          5538 => x"2b",
          5539 => x"8c",
          5540 => x"88",
          5541 => x"2e",
          5542 => x"88",
          5543 => x"0c",
          5544 => x"8c",
          5545 => x"71",
          5546 => x"87",
          5547 => x"0c",
          5548 => x"08",
          5549 => x"51",
          5550 => x"2e",
          5551 => x"c0",
          5552 => x"51",
          5553 => x"71",
          5554 => x"80",
          5555 => x"92",
          5556 => x"98",
          5557 => x"70",
          5558 => x"38",
          5559 => x"c4",
          5560 => x"d8",
          5561 => x"51",
          5562 => x"c8",
          5563 => x"0d",
          5564 => x"0d",
          5565 => x"02",
          5566 => x"05",
          5567 => x"58",
          5568 => x"52",
          5569 => x"3f",
          5570 => x"08",
          5571 => x"54",
          5572 => x"be",
          5573 => x"75",
          5574 => x"c0",
          5575 => x"87",
          5576 => x"12",
          5577 => x"84",
          5578 => x"40",
          5579 => x"85",
          5580 => x"98",
          5581 => x"7d",
          5582 => x"0c",
          5583 => x"85",
          5584 => x"06",
          5585 => x"71",
          5586 => x"38",
          5587 => x"71",
          5588 => x"05",
          5589 => x"19",
          5590 => x"a2",
          5591 => x"71",
          5592 => x"38",
          5593 => x"83",
          5594 => x"38",
          5595 => x"8a",
          5596 => x"98",
          5597 => x"71",
          5598 => x"c0",
          5599 => x"52",
          5600 => x"87",
          5601 => x"80",
          5602 => x"81",
          5603 => x"c0",
          5604 => x"53",
          5605 => x"82",
          5606 => x"71",
          5607 => x"1a",
          5608 => x"84",
          5609 => x"19",
          5610 => x"06",
          5611 => x"79",
          5612 => x"38",
          5613 => x"80",
          5614 => x"87",
          5615 => x"26",
          5616 => x"73",
          5617 => x"06",
          5618 => x"2e",
          5619 => x"52",
          5620 => x"82",
          5621 => x"8f",
          5622 => x"f3",
          5623 => x"62",
          5624 => x"05",
          5625 => x"57",
          5626 => x"83",
          5627 => x"52",
          5628 => x"3f",
          5629 => x"08",
          5630 => x"54",
          5631 => x"2e",
          5632 => x"81",
          5633 => x"74",
          5634 => x"c0",
          5635 => x"87",
          5636 => x"12",
          5637 => x"84",
          5638 => x"5f",
          5639 => x"0b",
          5640 => x"8c",
          5641 => x"0c",
          5642 => x"80",
          5643 => x"70",
          5644 => x"81",
          5645 => x"54",
          5646 => x"8c",
          5647 => x"81",
          5648 => x"7c",
          5649 => x"58",
          5650 => x"70",
          5651 => x"52",
          5652 => x"8a",
          5653 => x"98",
          5654 => x"71",
          5655 => x"c0",
          5656 => x"52",
          5657 => x"87",
          5658 => x"80",
          5659 => x"81",
          5660 => x"c0",
          5661 => x"53",
          5662 => x"82",
          5663 => x"71",
          5664 => x"19",
          5665 => x"81",
          5666 => x"ff",
          5667 => x"19",
          5668 => x"78",
          5669 => x"38",
          5670 => x"80",
          5671 => x"87",
          5672 => x"26",
          5673 => x"73",
          5674 => x"06",
          5675 => x"2e",
          5676 => x"52",
          5677 => x"82",
          5678 => x"8f",
          5679 => x"fa",
          5680 => x"02",
          5681 => x"05",
          5682 => x"05",
          5683 => x"71",
          5684 => x"57",
          5685 => x"82",
          5686 => x"81",
          5687 => x"54",
          5688 => x"38",
          5689 => x"c0",
          5690 => x"81",
          5691 => x"2e",
          5692 => x"71",
          5693 => x"38",
          5694 => x"87",
          5695 => x"11",
          5696 => x"80",
          5697 => x"80",
          5698 => x"83",
          5699 => x"38",
          5700 => x"72",
          5701 => x"2a",
          5702 => x"51",
          5703 => x"80",
          5704 => x"87",
          5705 => x"08",
          5706 => x"38",
          5707 => x"8c",
          5708 => x"96",
          5709 => x"0c",
          5710 => x"8c",
          5711 => x"08",
          5712 => x"51",
          5713 => x"38",
          5714 => x"56",
          5715 => x"80",
          5716 => x"85",
          5717 => x"77",
          5718 => x"83",
          5719 => x"75",
          5720 => x"d8",
          5721 => x"3d",
          5722 => x"3d",
          5723 => x"11",
          5724 => x"71",
          5725 => x"82",
          5726 => x"53",
          5727 => x"0d",
          5728 => x"0d",
          5729 => x"33",
          5730 => x"71",
          5731 => x"88",
          5732 => x"14",
          5733 => x"07",
          5734 => x"33",
          5735 => x"d8",
          5736 => x"53",
          5737 => x"52",
          5738 => x"04",
          5739 => x"73",
          5740 => x"92",
          5741 => x"52",
          5742 => x"81",
          5743 => x"70",
          5744 => x"70",
          5745 => x"3d",
          5746 => x"3d",
          5747 => x"52",
          5748 => x"70",
          5749 => x"34",
          5750 => x"51",
          5751 => x"81",
          5752 => x"70",
          5753 => x"70",
          5754 => x"05",
          5755 => x"88",
          5756 => x"72",
          5757 => x"0d",
          5758 => x"0d",
          5759 => x"54",
          5760 => x"80",
          5761 => x"71",
          5762 => x"53",
          5763 => x"81",
          5764 => x"ff",
          5765 => x"39",
          5766 => x"04",
          5767 => x"75",
          5768 => x"52",
          5769 => x"70",
          5770 => x"34",
          5771 => x"70",
          5772 => x"3d",
          5773 => x"3d",
          5774 => x"79",
          5775 => x"74",
          5776 => x"56",
          5777 => x"81",
          5778 => x"71",
          5779 => x"16",
          5780 => x"52",
          5781 => x"86",
          5782 => x"2e",
          5783 => x"82",
          5784 => x"86",
          5785 => x"fe",
          5786 => x"76",
          5787 => x"39",
          5788 => x"8a",
          5789 => x"51",
          5790 => x"71",
          5791 => x"33",
          5792 => x"0c",
          5793 => x"04",
          5794 => x"d8",
          5795 => x"fb",
          5796 => x"70",
          5797 => x"81",
          5798 => x"70",
          5799 => x"56",
          5800 => x"55",
          5801 => x"08",
          5802 => x"80",
          5803 => x"83",
          5804 => x"51",
          5805 => x"3f",
          5806 => x"08",
          5807 => x"06",
          5808 => x"2e",
          5809 => x"76",
          5810 => x"74",
          5811 => x"0c",
          5812 => x"04",
          5813 => x"7b",
          5814 => x"83",
          5815 => x"5a",
          5816 => x"80",
          5817 => x"54",
          5818 => x"53",
          5819 => x"53",
          5820 => x"52",
          5821 => x"3f",
          5822 => x"08",
          5823 => x"81",
          5824 => x"82",
          5825 => x"83",
          5826 => x"16",
          5827 => x"18",
          5828 => x"18",
          5829 => x"58",
          5830 => x"9f",
          5831 => x"33",
          5832 => x"2e",
          5833 => x"93",
          5834 => x"76",
          5835 => x"52",
          5836 => x"51",
          5837 => x"83",
          5838 => x"79",
          5839 => x"0c",
          5840 => x"04",
          5841 => x"78",
          5842 => x"80",
          5843 => x"17",
          5844 => x"38",
          5845 => x"fc",
          5846 => x"c8",
          5847 => x"d8",
          5848 => x"38",
          5849 => x"53",
          5850 => x"81",
          5851 => x"f7",
          5852 => x"d8",
          5853 => x"2e",
          5854 => x"55",
          5855 => x"b4",
          5856 => x"82",
          5857 => x"88",
          5858 => x"f8",
          5859 => x"70",
          5860 => x"c0",
          5861 => x"c8",
          5862 => x"d8",
          5863 => x"91",
          5864 => x"55",
          5865 => x"09",
          5866 => x"f0",
          5867 => x"33",
          5868 => x"2e",
          5869 => x"80",
          5870 => x"80",
          5871 => x"c8",
          5872 => x"17",
          5873 => x"fc",
          5874 => x"d4",
          5875 => x"b6",
          5876 => x"d8",
          5877 => x"85",
          5878 => x"75",
          5879 => x"3f",
          5880 => x"e4",
          5881 => x"9c",
          5882 => x"de",
          5883 => x"08",
          5884 => x"17",
          5885 => x"3f",
          5886 => x"52",
          5887 => x"51",
          5888 => x"a4",
          5889 => x"05",
          5890 => x"0c",
          5891 => x"75",
          5892 => x"33",
          5893 => x"3f",
          5894 => x"34",
          5895 => x"52",
          5896 => x"51",
          5897 => x"82",
          5898 => x"80",
          5899 => x"81",
          5900 => x"d8",
          5901 => x"3d",
          5902 => x"3d",
          5903 => x"1a",
          5904 => x"fe",
          5905 => x"54",
          5906 => x"73",
          5907 => x"8a",
          5908 => x"71",
          5909 => x"08",
          5910 => x"75",
          5911 => x"0c",
          5912 => x"04",
          5913 => x"7a",
          5914 => x"56",
          5915 => x"77",
          5916 => x"38",
          5917 => x"08",
          5918 => x"38",
          5919 => x"54",
          5920 => x"2e",
          5921 => x"72",
          5922 => x"38",
          5923 => x"8d",
          5924 => x"39",
          5925 => x"81",
          5926 => x"b6",
          5927 => x"2a",
          5928 => x"2a",
          5929 => x"05",
          5930 => x"55",
          5931 => x"82",
          5932 => x"81",
          5933 => x"83",
          5934 => x"b8",
          5935 => x"17",
          5936 => x"a8",
          5937 => x"55",
          5938 => x"57",
          5939 => x"3f",
          5940 => x"08",
          5941 => x"74",
          5942 => x"14",
          5943 => x"70",
          5944 => x"07",
          5945 => x"71",
          5946 => x"52",
          5947 => x"72",
          5948 => x"75",
          5949 => x"58",
          5950 => x"76",
          5951 => x"15",
          5952 => x"73",
          5953 => x"3f",
          5954 => x"08",
          5955 => x"76",
          5956 => x"06",
          5957 => x"05",
          5958 => x"3f",
          5959 => x"08",
          5960 => x"06",
          5961 => x"76",
          5962 => x"15",
          5963 => x"73",
          5964 => x"3f",
          5965 => x"08",
          5966 => x"82",
          5967 => x"06",
          5968 => x"05",
          5969 => x"3f",
          5970 => x"08",
          5971 => x"58",
          5972 => x"58",
          5973 => x"c8",
          5974 => x"0d",
          5975 => x"0d",
          5976 => x"5a",
          5977 => x"59",
          5978 => x"82",
          5979 => x"9c",
          5980 => x"82",
          5981 => x"33",
          5982 => x"2e",
          5983 => x"72",
          5984 => x"38",
          5985 => x"8d",
          5986 => x"39",
          5987 => x"81",
          5988 => x"f7",
          5989 => x"2a",
          5990 => x"2a",
          5991 => x"05",
          5992 => x"55",
          5993 => x"82",
          5994 => x"59",
          5995 => x"08",
          5996 => x"74",
          5997 => x"16",
          5998 => x"16",
          5999 => x"59",
          6000 => x"53",
          6001 => x"8f",
          6002 => x"2b",
          6003 => x"74",
          6004 => x"71",
          6005 => x"72",
          6006 => x"0b",
          6007 => x"74",
          6008 => x"17",
          6009 => x"75",
          6010 => x"3f",
          6011 => x"08",
          6012 => x"c8",
          6013 => x"38",
          6014 => x"06",
          6015 => x"78",
          6016 => x"54",
          6017 => x"77",
          6018 => x"33",
          6019 => x"71",
          6020 => x"51",
          6021 => x"34",
          6022 => x"76",
          6023 => x"17",
          6024 => x"75",
          6025 => x"3f",
          6026 => x"08",
          6027 => x"c8",
          6028 => x"38",
          6029 => x"ff",
          6030 => x"10",
          6031 => x"76",
          6032 => x"51",
          6033 => x"be",
          6034 => x"2a",
          6035 => x"05",
          6036 => x"f9",
          6037 => x"d8",
          6038 => x"82",
          6039 => x"ab",
          6040 => x"0a",
          6041 => x"2b",
          6042 => x"70",
          6043 => x"70",
          6044 => x"54",
          6045 => x"82",
          6046 => x"8f",
          6047 => x"07",
          6048 => x"f6",
          6049 => x"0b",
          6050 => x"78",
          6051 => x"0c",
          6052 => x"04",
          6053 => x"7a",
          6054 => x"08",
          6055 => x"59",
          6056 => x"a4",
          6057 => x"17",
          6058 => x"38",
          6059 => x"aa",
          6060 => x"73",
          6061 => x"fd",
          6062 => x"d8",
          6063 => x"82",
          6064 => x"80",
          6065 => x"39",
          6066 => x"eb",
          6067 => x"80",
          6068 => x"d8",
          6069 => x"80",
          6070 => x"52",
          6071 => x"84",
          6072 => x"c8",
          6073 => x"d8",
          6074 => x"2e",
          6075 => x"82",
          6076 => x"81",
          6077 => x"82",
          6078 => x"ff",
          6079 => x"80",
          6080 => x"75",
          6081 => x"3f",
          6082 => x"08",
          6083 => x"16",
          6084 => x"94",
          6085 => x"55",
          6086 => x"27",
          6087 => x"15",
          6088 => x"84",
          6089 => x"07",
          6090 => x"17",
          6091 => x"76",
          6092 => x"a6",
          6093 => x"73",
          6094 => x"0c",
          6095 => x"04",
          6096 => x"7c",
          6097 => x"59",
          6098 => x"95",
          6099 => x"08",
          6100 => x"2e",
          6101 => x"17",
          6102 => x"b2",
          6103 => x"ae",
          6104 => x"7a",
          6105 => x"3f",
          6106 => x"82",
          6107 => x"27",
          6108 => x"82",
          6109 => x"55",
          6110 => x"08",
          6111 => x"d2",
          6112 => x"08",
          6113 => x"08",
          6114 => x"38",
          6115 => x"17",
          6116 => x"54",
          6117 => x"82",
          6118 => x"7a",
          6119 => x"06",
          6120 => x"81",
          6121 => x"17",
          6122 => x"83",
          6123 => x"75",
          6124 => x"f9",
          6125 => x"59",
          6126 => x"08",
          6127 => x"81",
          6128 => x"82",
          6129 => x"59",
          6130 => x"08",
          6131 => x"70",
          6132 => x"25",
          6133 => x"82",
          6134 => x"54",
          6135 => x"55",
          6136 => x"38",
          6137 => x"08",
          6138 => x"38",
          6139 => x"54",
          6140 => x"90",
          6141 => x"18",
          6142 => x"38",
          6143 => x"39",
          6144 => x"38",
          6145 => x"16",
          6146 => x"08",
          6147 => x"38",
          6148 => x"78",
          6149 => x"38",
          6150 => x"51",
          6151 => x"82",
          6152 => x"80",
          6153 => x"80",
          6154 => x"c8",
          6155 => x"09",
          6156 => x"38",
          6157 => x"08",
          6158 => x"c8",
          6159 => x"30",
          6160 => x"80",
          6161 => x"07",
          6162 => x"55",
          6163 => x"38",
          6164 => x"09",
          6165 => x"ae",
          6166 => x"80",
          6167 => x"53",
          6168 => x"51",
          6169 => x"82",
          6170 => x"82",
          6171 => x"30",
          6172 => x"c8",
          6173 => x"25",
          6174 => x"79",
          6175 => x"38",
          6176 => x"8f",
          6177 => x"79",
          6178 => x"f9",
          6179 => x"d8",
          6180 => x"74",
          6181 => x"90",
          6182 => x"17",
          6183 => x"94",
          6184 => x"54",
          6185 => x"86",
          6186 => x"94",
          6187 => x"17",
          6188 => x"54",
          6189 => x"34",
          6190 => x"56",
          6191 => x"90",
          6192 => x"80",
          6193 => x"82",
          6194 => x"55",
          6195 => x"56",
          6196 => x"82",
          6197 => x"8c",
          6198 => x"f8",
          6199 => x"70",
          6200 => x"f0",
          6201 => x"c8",
          6202 => x"56",
          6203 => x"08",
          6204 => x"7b",
          6205 => x"f6",
          6206 => x"d8",
          6207 => x"d8",
          6208 => x"17",
          6209 => x"80",
          6210 => x"b8",
          6211 => x"57",
          6212 => x"77",
          6213 => x"81",
          6214 => x"15",
          6215 => x"78",
          6216 => x"81",
          6217 => x"53",
          6218 => x"15",
          6219 => x"ab",
          6220 => x"c8",
          6221 => x"df",
          6222 => x"22",
          6223 => x"30",
          6224 => x"70",
          6225 => x"51",
          6226 => x"82",
          6227 => x"8a",
          6228 => x"f8",
          6229 => x"7c",
          6230 => x"56",
          6231 => x"80",
          6232 => x"f1",
          6233 => x"06",
          6234 => x"e9",
          6235 => x"18",
          6236 => x"08",
          6237 => x"38",
          6238 => x"82",
          6239 => x"38",
          6240 => x"54",
          6241 => x"74",
          6242 => x"82",
          6243 => x"22",
          6244 => x"79",
          6245 => x"38",
          6246 => x"98",
          6247 => x"cd",
          6248 => x"22",
          6249 => x"54",
          6250 => x"26",
          6251 => x"52",
          6252 => x"b0",
          6253 => x"c8",
          6254 => x"d8",
          6255 => x"2e",
          6256 => x"0b",
          6257 => x"08",
          6258 => x"9c",
          6259 => x"d8",
          6260 => x"85",
          6261 => x"bd",
          6262 => x"31",
          6263 => x"73",
          6264 => x"f4",
          6265 => x"d8",
          6266 => x"18",
          6267 => x"18",
          6268 => x"08",
          6269 => x"72",
          6270 => x"38",
          6271 => x"58",
          6272 => x"89",
          6273 => x"18",
          6274 => x"ff",
          6275 => x"05",
          6276 => x"80",
          6277 => x"d8",
          6278 => x"3d",
          6279 => x"3d",
          6280 => x"08",
          6281 => x"a0",
          6282 => x"54",
          6283 => x"77",
          6284 => x"80",
          6285 => x"0c",
          6286 => x"53",
          6287 => x"80",
          6288 => x"38",
          6289 => x"06",
          6290 => x"b5",
          6291 => x"98",
          6292 => x"14",
          6293 => x"92",
          6294 => x"2a",
          6295 => x"56",
          6296 => x"26",
          6297 => x"80",
          6298 => x"16",
          6299 => x"77",
          6300 => x"53",
          6301 => x"38",
          6302 => x"51",
          6303 => x"82",
          6304 => x"53",
          6305 => x"0b",
          6306 => x"08",
          6307 => x"38",
          6308 => x"d8",
          6309 => x"2e",
          6310 => x"9c",
          6311 => x"d8",
          6312 => x"80",
          6313 => x"8a",
          6314 => x"15",
          6315 => x"80",
          6316 => x"14",
          6317 => x"51",
          6318 => x"82",
          6319 => x"53",
          6320 => x"d8",
          6321 => x"2e",
          6322 => x"82",
          6323 => x"c8",
          6324 => x"ba",
          6325 => x"82",
          6326 => x"ff",
          6327 => x"82",
          6328 => x"52",
          6329 => x"f3",
          6330 => x"c8",
          6331 => x"72",
          6332 => x"72",
          6333 => x"f2",
          6334 => x"d8",
          6335 => x"15",
          6336 => x"15",
          6337 => x"b8",
          6338 => x"0c",
          6339 => x"82",
          6340 => x"8a",
          6341 => x"f7",
          6342 => x"7d",
          6343 => x"5b",
          6344 => x"76",
          6345 => x"3f",
          6346 => x"08",
          6347 => x"c8",
          6348 => x"38",
          6349 => x"08",
          6350 => x"08",
          6351 => x"f0",
          6352 => x"d8",
          6353 => x"82",
          6354 => x"80",
          6355 => x"d8",
          6356 => x"18",
          6357 => x"51",
          6358 => x"81",
          6359 => x"81",
          6360 => x"81",
          6361 => x"c8",
          6362 => x"83",
          6363 => x"77",
          6364 => x"72",
          6365 => x"38",
          6366 => x"75",
          6367 => x"81",
          6368 => x"a5",
          6369 => x"c8",
          6370 => x"52",
          6371 => x"8e",
          6372 => x"c8",
          6373 => x"d8",
          6374 => x"2e",
          6375 => x"73",
          6376 => x"81",
          6377 => x"87",
          6378 => x"d8",
          6379 => x"3d",
          6380 => x"3d",
          6381 => x"11",
          6382 => x"ae",
          6383 => x"c8",
          6384 => x"ff",
          6385 => x"33",
          6386 => x"71",
          6387 => x"81",
          6388 => x"94",
          6389 => x"92",
          6390 => x"c8",
          6391 => x"73",
          6392 => x"82",
          6393 => x"85",
          6394 => x"fc",
          6395 => x"79",
          6396 => x"ff",
          6397 => x"12",
          6398 => x"eb",
          6399 => x"70",
          6400 => x"72",
          6401 => x"81",
          6402 => x"73",
          6403 => x"94",
          6404 => x"98",
          6405 => x"0d",
          6406 => x"0d",
          6407 => x"51",
          6408 => x"81",
          6409 => x"80",
          6410 => x"70",
          6411 => x"33",
          6412 => x"81",
          6413 => x"16",
          6414 => x"51",
          6415 => x"70",
          6416 => x"0c",
          6417 => x"04",
          6418 => x"60",
          6419 => x"84",
          6420 => x"5b",
          6421 => x"5d",
          6422 => x"08",
          6423 => x"80",
          6424 => x"08",
          6425 => x"ed",
          6426 => x"d8",
          6427 => x"82",
          6428 => x"82",
          6429 => x"19",
          6430 => x"55",
          6431 => x"38",
          6432 => x"dc",
          6433 => x"33",
          6434 => x"81",
          6435 => x"53",
          6436 => x"34",
          6437 => x"08",
          6438 => x"e5",
          6439 => x"06",
          6440 => x"56",
          6441 => x"08",
          6442 => x"2e",
          6443 => x"83",
          6444 => x"75",
          6445 => x"72",
          6446 => x"d8",
          6447 => x"df",
          6448 => x"72",
          6449 => x"81",
          6450 => x"81",
          6451 => x"2e",
          6452 => x"ff",
          6453 => x"39",
          6454 => x"09",
          6455 => x"ca",
          6456 => x"2a",
          6457 => x"51",
          6458 => x"2e",
          6459 => x"15",
          6460 => x"bf",
          6461 => x"1c",
          6462 => x"0c",
          6463 => x"73",
          6464 => x"81",
          6465 => x"38",
          6466 => x"53",
          6467 => x"09",
          6468 => x"8f",
          6469 => x"08",
          6470 => x"5a",
          6471 => x"82",
          6472 => x"83",
          6473 => x"53",
          6474 => x"38",
          6475 => x"81",
          6476 => x"29",
          6477 => x"54",
          6478 => x"58",
          6479 => x"17",
          6480 => x"51",
          6481 => x"82",
          6482 => x"83",
          6483 => x"56",
          6484 => x"96",
          6485 => x"fe",
          6486 => x"38",
          6487 => x"76",
          6488 => x"73",
          6489 => x"54",
          6490 => x"83",
          6491 => x"09",
          6492 => x"38",
          6493 => x"8c",
          6494 => x"38",
          6495 => x"86",
          6496 => x"06",
          6497 => x"72",
          6498 => x"38",
          6499 => x"26",
          6500 => x"10",
          6501 => x"73",
          6502 => x"70",
          6503 => x"51",
          6504 => x"81",
          6505 => x"5c",
          6506 => x"93",
          6507 => x"fc",
          6508 => x"d8",
          6509 => x"ff",
          6510 => x"7d",
          6511 => x"ff",
          6512 => x"0c",
          6513 => x"52",
          6514 => x"d2",
          6515 => x"c8",
          6516 => x"d8",
          6517 => x"38",
          6518 => x"fd",
          6519 => x"39",
          6520 => x"1a",
          6521 => x"d8",
          6522 => x"3d",
          6523 => x"3d",
          6524 => x"08",
          6525 => x"52",
          6526 => x"d7",
          6527 => x"c8",
          6528 => x"d8",
          6529 => x"a4",
          6530 => x"70",
          6531 => x"0b",
          6532 => x"98",
          6533 => x"7e",
          6534 => x"3f",
          6535 => x"08",
          6536 => x"c8",
          6537 => x"38",
          6538 => x"70",
          6539 => x"75",
          6540 => x"58",
          6541 => x"8b",
          6542 => x"06",
          6543 => x"06",
          6544 => x"86",
          6545 => x"81",
          6546 => x"c3",
          6547 => x"2a",
          6548 => x"51",
          6549 => x"2e",
          6550 => x"82",
          6551 => x"8f",
          6552 => x"06",
          6553 => x"ab",
          6554 => x"86",
          6555 => x"06",
          6556 => x"73",
          6557 => x"75",
          6558 => x"81",
          6559 => x"73",
          6560 => x"38",
          6561 => x"76",
          6562 => x"70",
          6563 => x"ac",
          6564 => x"5d",
          6565 => x"2e",
          6566 => x"81",
          6567 => x"17",
          6568 => x"76",
          6569 => x"06",
          6570 => x"8c",
          6571 => x"18",
          6572 => x"b6",
          6573 => x"c8",
          6574 => x"ff",
          6575 => x"81",
          6576 => x"33",
          6577 => x"8d",
          6578 => x"59",
          6579 => x"5c",
          6580 => x"d0",
          6581 => x"05",
          6582 => x"3f",
          6583 => x"08",
          6584 => x"06",
          6585 => x"2e",
          6586 => x"81",
          6587 => x"e6",
          6588 => x"80",
          6589 => x"82",
          6590 => x"78",
          6591 => x"22",
          6592 => x"19",
          6593 => x"df",
          6594 => x"82",
          6595 => x"2e",
          6596 => x"80",
          6597 => x"5a",
          6598 => x"83",
          6599 => x"09",
          6600 => x"38",
          6601 => x"8c",
          6602 => x"a5",
          6603 => x"70",
          6604 => x"81",
          6605 => x"57",
          6606 => x"90",
          6607 => x"2e",
          6608 => x"10",
          6609 => x"51",
          6610 => x"38",
          6611 => x"81",
          6612 => x"54",
          6613 => x"ff",
          6614 => x"bb",
          6615 => x"38",
          6616 => x"b5",
          6617 => x"c8",
          6618 => x"06",
          6619 => x"2e",
          6620 => x"19",
          6621 => x"54",
          6622 => x"8b",
          6623 => x"52",
          6624 => x"51",
          6625 => x"82",
          6626 => x"80",
          6627 => x"81",
          6628 => x"0b",
          6629 => x"80",
          6630 => x"f5",
          6631 => x"d8",
          6632 => x"82",
          6633 => x"80",
          6634 => x"38",
          6635 => x"c8",
          6636 => x"0d",
          6637 => x"0d",
          6638 => x"ab",
          6639 => x"a0",
          6640 => x"5a",
          6641 => x"85",
          6642 => x"8c",
          6643 => x"22",
          6644 => x"73",
          6645 => x"38",
          6646 => x"10",
          6647 => x"51",
          6648 => x"39",
          6649 => x"1a",
          6650 => x"3d",
          6651 => x"59",
          6652 => x"02",
          6653 => x"33",
          6654 => x"73",
          6655 => x"a8",
          6656 => x"0b",
          6657 => x"81",
          6658 => x"08",
          6659 => x"8b",
          6660 => x"78",
          6661 => x"3f",
          6662 => x"80",
          6663 => x"56",
          6664 => x"83",
          6665 => x"55",
          6666 => x"2e",
          6667 => x"83",
          6668 => x"82",
          6669 => x"8f",
          6670 => x"06",
          6671 => x"75",
          6672 => x"90",
          6673 => x"06",
          6674 => x"56",
          6675 => x"87",
          6676 => x"a0",
          6677 => x"ff",
          6678 => x"80",
          6679 => x"c0",
          6680 => x"87",
          6681 => x"bf",
          6682 => x"74",
          6683 => x"06",
          6684 => x"27",
          6685 => x"14",
          6686 => x"34",
          6687 => x"18",
          6688 => x"57",
          6689 => x"e3",
          6690 => x"ec",
          6691 => x"80",
          6692 => x"80",
          6693 => x"38",
          6694 => x"73",
          6695 => x"38",
          6696 => x"33",
          6697 => x"e0",
          6698 => x"c8",
          6699 => x"8c",
          6700 => x"54",
          6701 => x"94",
          6702 => x"55",
          6703 => x"74",
          6704 => x"38",
          6705 => x"33",
          6706 => x"39",
          6707 => x"05",
          6708 => x"78",
          6709 => x"56",
          6710 => x"76",
          6711 => x"38",
          6712 => x"15",
          6713 => x"55",
          6714 => x"34",
          6715 => x"e3",
          6716 => x"f9",
          6717 => x"d8",
          6718 => x"38",
          6719 => x"80",
          6720 => x"fe",
          6721 => x"55",
          6722 => x"2e",
          6723 => x"82",
          6724 => x"55",
          6725 => x"08",
          6726 => x"81",
          6727 => x"38",
          6728 => x"05",
          6729 => x"34",
          6730 => x"05",
          6731 => x"2a",
          6732 => x"51",
          6733 => x"59",
          6734 => x"90",
          6735 => x"8c",
          6736 => x"f4",
          6737 => x"d8",
          6738 => x"59",
          6739 => x"51",
          6740 => x"82",
          6741 => x"57",
          6742 => x"08",
          6743 => x"ff",
          6744 => x"80",
          6745 => x"38",
          6746 => x"90",
          6747 => x"31",
          6748 => x"51",
          6749 => x"82",
          6750 => x"57",
          6751 => x"08",
          6752 => x"a0",
          6753 => x"91",
          6754 => x"c8",
          6755 => x"06",
          6756 => x"08",
          6757 => x"e3",
          6758 => x"d8",
          6759 => x"82",
          6760 => x"81",
          6761 => x"1c",
          6762 => x"08",
          6763 => x"06",
          6764 => x"7c",
          6765 => x"8f",
          6766 => x"34",
          6767 => x"08",
          6768 => x"82",
          6769 => x"52",
          6770 => x"df",
          6771 => x"8d",
          6772 => x"77",
          6773 => x"83",
          6774 => x"8b",
          6775 => x"1b",
          6776 => x"17",
          6777 => x"73",
          6778 => x"d0",
          6779 => x"05",
          6780 => x"3f",
          6781 => x"83",
          6782 => x"81",
          6783 => x"77",
          6784 => x"73",
          6785 => x"2e",
          6786 => x"10",
          6787 => x"51",
          6788 => x"38",
          6789 => x"07",
          6790 => x"34",
          6791 => x"1d",
          6792 => x"79",
          6793 => x"3f",
          6794 => x"08",
          6795 => x"c8",
          6796 => x"38",
          6797 => x"78",
          6798 => x"98",
          6799 => x"7b",
          6800 => x"3f",
          6801 => x"08",
          6802 => x"c8",
          6803 => x"a0",
          6804 => x"c8",
          6805 => x"1a",
          6806 => x"c0",
          6807 => x"a0",
          6808 => x"1a",
          6809 => x"91",
          6810 => x"08",
          6811 => x"98",
          6812 => x"73",
          6813 => x"81",
          6814 => x"34",
          6815 => x"82",
          6816 => x"94",
          6817 => x"fa",
          6818 => x"70",
          6819 => x"08",
          6820 => x"56",
          6821 => x"72",
          6822 => x"38",
          6823 => x"51",
          6824 => x"82",
          6825 => x"54",
          6826 => x"08",
          6827 => x"98",
          6828 => x"75",
          6829 => x"3f",
          6830 => x"08",
          6831 => x"c8",
          6832 => x"9c",
          6833 => x"e5",
          6834 => x"0b",
          6835 => x"90",
          6836 => x"27",
          6837 => x"d8",
          6838 => x"74",
          6839 => x"3f",
          6840 => x"08",
          6841 => x"c8",
          6842 => x"c3",
          6843 => x"2e",
          6844 => x"83",
          6845 => x"73",
          6846 => x"0c",
          6847 => x"04",
          6848 => x"7e",
          6849 => x"5f",
          6850 => x"0b",
          6851 => x"98",
          6852 => x"2e",
          6853 => x"ac",
          6854 => x"2e",
          6855 => x"80",
          6856 => x"8c",
          6857 => x"22",
          6858 => x"5c",
          6859 => x"2e",
          6860 => x"78",
          6861 => x"22",
          6862 => x"56",
          6863 => x"38",
          6864 => x"15",
          6865 => x"ff",
          6866 => x"72",
          6867 => x"86",
          6868 => x"80",
          6869 => x"18",
          6870 => x"ff",
          6871 => x"5b",
          6872 => x"52",
          6873 => x"75",
          6874 => x"d5",
          6875 => x"d8",
          6876 => x"ff",
          6877 => x"81",
          6878 => x"95",
          6879 => x"27",
          6880 => x"88",
          6881 => x"7a",
          6882 => x"15",
          6883 => x"9f",
          6884 => x"76",
          6885 => x"07",
          6886 => x"80",
          6887 => x"54",
          6888 => x"2e",
          6889 => x"57",
          6890 => x"7a",
          6891 => x"74",
          6892 => x"5b",
          6893 => x"79",
          6894 => x"22",
          6895 => x"72",
          6896 => x"7a",
          6897 => x"25",
          6898 => x"06",
          6899 => x"77",
          6900 => x"53",
          6901 => x"14",
          6902 => x"89",
          6903 => x"57",
          6904 => x"19",
          6905 => x"1b",
          6906 => x"74",
          6907 => x"38",
          6908 => x"09",
          6909 => x"38",
          6910 => x"78",
          6911 => x"30",
          6912 => x"80",
          6913 => x"54",
          6914 => x"90",
          6915 => x"2e",
          6916 => x"76",
          6917 => x"58",
          6918 => x"57",
          6919 => x"81",
          6920 => x"81",
          6921 => x"79",
          6922 => x"38",
          6923 => x"05",
          6924 => x"81",
          6925 => x"18",
          6926 => x"81",
          6927 => x"8b",
          6928 => x"96",
          6929 => x"57",
          6930 => x"72",
          6931 => x"33",
          6932 => x"72",
          6933 => x"d3",
          6934 => x"89",
          6935 => x"73",
          6936 => x"11",
          6937 => x"99",
          6938 => x"9c",
          6939 => x"11",
          6940 => x"88",
          6941 => x"38",
          6942 => x"53",
          6943 => x"83",
          6944 => x"81",
          6945 => x"80",
          6946 => x"a0",
          6947 => x"ff",
          6948 => x"53",
          6949 => x"81",
          6950 => x"81",
          6951 => x"81",
          6952 => x"56",
          6953 => x"72",
          6954 => x"77",
          6955 => x"53",
          6956 => x"14",
          6957 => x"08",
          6958 => x"51",
          6959 => x"38",
          6960 => x"34",
          6961 => x"53",
          6962 => x"88",
          6963 => x"1c",
          6964 => x"52",
          6965 => x"3f",
          6966 => x"08",
          6967 => x"13",
          6968 => x"3f",
          6969 => x"08",
          6970 => x"98",
          6971 => x"fa",
          6972 => x"c8",
          6973 => x"23",
          6974 => x"04",
          6975 => x"62",
          6976 => x"5e",
          6977 => x"33",
          6978 => x"73",
          6979 => x"38",
          6980 => x"80",
          6981 => x"38",
          6982 => x"8d",
          6983 => x"05",
          6984 => x"0c",
          6985 => x"15",
          6986 => x"70",
          6987 => x"56",
          6988 => x"09",
          6989 => x"38",
          6990 => x"80",
          6991 => x"30",
          6992 => x"78",
          6993 => x"54",
          6994 => x"73",
          6995 => x"63",
          6996 => x"54",
          6997 => x"96",
          6998 => x"0b",
          6999 => x"80",
          7000 => x"e7",
          7001 => x"d8",
          7002 => x"87",
          7003 => x"41",
          7004 => x"11",
          7005 => x"80",
          7006 => x"fc",
          7007 => x"8f",
          7008 => x"c8",
          7009 => x"82",
          7010 => x"ff",
          7011 => x"d8",
          7012 => x"92",
          7013 => x"1a",
          7014 => x"08",
          7015 => x"55",
          7016 => x"81",
          7017 => x"d8",
          7018 => x"ff",
          7019 => x"af",
          7020 => x"9f",
          7021 => x"80",
          7022 => x"51",
          7023 => x"b4",
          7024 => x"dc",
          7025 => x"75",
          7026 => x"91",
          7027 => x"82",
          7028 => x"d9",
          7029 => x"d8",
          7030 => x"de",
          7031 => x"fe",
          7032 => x"38",
          7033 => x"54",
          7034 => x"81",
          7035 => x"89",
          7036 => x"41",
          7037 => x"33",
          7038 => x"73",
          7039 => x"81",
          7040 => x"81",
          7041 => x"dc",
          7042 => x"70",
          7043 => x"07",
          7044 => x"73",
          7045 => x"44",
          7046 => x"82",
          7047 => x"81",
          7048 => x"06",
          7049 => x"22",
          7050 => x"2e",
          7051 => x"d2",
          7052 => x"2e",
          7053 => x"80",
          7054 => x"1a",
          7055 => x"ae",
          7056 => x"06",
          7057 => x"79",
          7058 => x"ae",
          7059 => x"06",
          7060 => x"10",
          7061 => x"74",
          7062 => x"a0",
          7063 => x"ae",
          7064 => x"26",
          7065 => x"54",
          7066 => x"81",
          7067 => x"81",
          7068 => x"78",
          7069 => x"76",
          7070 => x"73",
          7071 => x"84",
          7072 => x"80",
          7073 => x"78",
          7074 => x"05",
          7075 => x"fe",
          7076 => x"a0",
          7077 => x"70",
          7078 => x"51",
          7079 => x"54",
          7080 => x"84",
          7081 => x"38",
          7082 => x"78",
          7083 => x"19",
          7084 => x"56",
          7085 => x"78",
          7086 => x"56",
          7087 => x"76",
          7088 => x"83",
          7089 => x"7a",
          7090 => x"ff",
          7091 => x"56",
          7092 => x"2e",
          7093 => x"93",
          7094 => x"70",
          7095 => x"22",
          7096 => x"73",
          7097 => x"38",
          7098 => x"74",
          7099 => x"06",
          7100 => x"2e",
          7101 => x"85",
          7102 => x"07",
          7103 => x"2e",
          7104 => x"16",
          7105 => x"22",
          7106 => x"ae",
          7107 => x"78",
          7108 => x"05",
          7109 => x"59",
          7110 => x"8f",
          7111 => x"70",
          7112 => x"73",
          7113 => x"81",
          7114 => x"8b",
          7115 => x"a0",
          7116 => x"e8",
          7117 => x"59",
          7118 => x"7c",
          7119 => x"22",
          7120 => x"57",
          7121 => x"2e",
          7122 => x"75",
          7123 => x"38",
          7124 => x"70",
          7125 => x"25",
          7126 => x"7c",
          7127 => x"38",
          7128 => x"89",
          7129 => x"07",
          7130 => x"80",
          7131 => x"7e",
          7132 => x"38",
          7133 => x"79",
          7134 => x"70",
          7135 => x"25",
          7136 => x"51",
          7137 => x"73",
          7138 => x"38",
          7139 => x"fe",
          7140 => x"79",
          7141 => x"76",
          7142 => x"7c",
          7143 => x"be",
          7144 => x"88",
          7145 => x"82",
          7146 => x"06",
          7147 => x"8b",
          7148 => x"76",
          7149 => x"76",
          7150 => x"83",
          7151 => x"51",
          7152 => x"3f",
          7153 => x"08",
          7154 => x"06",
          7155 => x"70",
          7156 => x"55",
          7157 => x"2e",
          7158 => x"80",
          7159 => x"ca",
          7160 => x"57",
          7161 => x"76",
          7162 => x"ff",
          7163 => x"78",
          7164 => x"76",
          7165 => x"59",
          7166 => x"39",
          7167 => x"05",
          7168 => x"55",
          7169 => x"34",
          7170 => x"80",
          7171 => x"80",
          7172 => x"75",
          7173 => x"f8",
          7174 => x"3f",
          7175 => x"08",
          7176 => x"38",
          7177 => x"83",
          7178 => x"a4",
          7179 => x"16",
          7180 => x"26",
          7181 => x"82",
          7182 => x"9f",
          7183 => x"99",
          7184 => x"7b",
          7185 => x"17",
          7186 => x"ff",
          7187 => x"5c",
          7188 => x"05",
          7189 => x"34",
          7190 => x"fd",
          7191 => x"1e",
          7192 => x"81",
          7193 => x"81",
          7194 => x"85",
          7195 => x"34",
          7196 => x"09",
          7197 => x"38",
          7198 => x"81",
          7199 => x"7b",
          7200 => x"73",
          7201 => x"38",
          7202 => x"54",
          7203 => x"09",
          7204 => x"38",
          7205 => x"57",
          7206 => x"70",
          7207 => x"54",
          7208 => x"7b",
          7209 => x"73",
          7210 => x"38",
          7211 => x"57",
          7212 => x"70",
          7213 => x"54",
          7214 => x"85",
          7215 => x"07",
          7216 => x"1f",
          7217 => x"ea",
          7218 => x"d8",
          7219 => x"1f",
          7220 => x"82",
          7221 => x"80",
          7222 => x"82",
          7223 => x"84",
          7224 => x"06",
          7225 => x"74",
          7226 => x"81",
          7227 => x"2a",
          7228 => x"73",
          7229 => x"38",
          7230 => x"54",
          7231 => x"f8",
          7232 => x"80",
          7233 => x"34",
          7234 => x"c2",
          7235 => x"06",
          7236 => x"38",
          7237 => x"39",
          7238 => x"70",
          7239 => x"54",
          7240 => x"86",
          7241 => x"84",
          7242 => x"06",
          7243 => x"73",
          7244 => x"38",
          7245 => x"83",
          7246 => x"05",
          7247 => x"7f",
          7248 => x"3f",
          7249 => x"08",
          7250 => x"f8",
          7251 => x"82",
          7252 => x"92",
          7253 => x"f6",
          7254 => x"5b",
          7255 => x"70",
          7256 => x"59",
          7257 => x"73",
          7258 => x"c6",
          7259 => x"81",
          7260 => x"70",
          7261 => x"52",
          7262 => x"8d",
          7263 => x"38",
          7264 => x"09",
          7265 => x"a5",
          7266 => x"d0",
          7267 => x"ff",
          7268 => x"53",
          7269 => x"91",
          7270 => x"73",
          7271 => x"d0",
          7272 => x"71",
          7273 => x"f7",
          7274 => x"82",
          7275 => x"55",
          7276 => x"55",
          7277 => x"81",
          7278 => x"74",
          7279 => x"56",
          7280 => x"12",
          7281 => x"70",
          7282 => x"38",
          7283 => x"81",
          7284 => x"51",
          7285 => x"51",
          7286 => x"89",
          7287 => x"70",
          7288 => x"53",
          7289 => x"70",
          7290 => x"51",
          7291 => x"09",
          7292 => x"38",
          7293 => x"38",
          7294 => x"77",
          7295 => x"70",
          7296 => x"2a",
          7297 => x"07",
          7298 => x"51",
          7299 => x"8f",
          7300 => x"84",
          7301 => x"83",
          7302 => x"94",
          7303 => x"74",
          7304 => x"38",
          7305 => x"0c",
          7306 => x"86",
          7307 => x"a4",
          7308 => x"82",
          7309 => x"8c",
          7310 => x"fa",
          7311 => x"56",
          7312 => x"17",
          7313 => x"b4",
          7314 => x"52",
          7315 => x"f4",
          7316 => x"82",
          7317 => x"81",
          7318 => x"b6",
          7319 => x"8a",
          7320 => x"c8",
          7321 => x"ff",
          7322 => x"55",
          7323 => x"d5",
          7324 => x"06",
          7325 => x"80",
          7326 => x"33",
          7327 => x"81",
          7328 => x"81",
          7329 => x"81",
          7330 => x"eb",
          7331 => x"70",
          7332 => x"07",
          7333 => x"73",
          7334 => x"81",
          7335 => x"81",
          7336 => x"83",
          7337 => x"80",
          7338 => x"16",
          7339 => x"3f",
          7340 => x"08",
          7341 => x"c8",
          7342 => x"9d",
          7343 => x"82",
          7344 => x"81",
          7345 => x"ce",
          7346 => x"d8",
          7347 => x"82",
          7348 => x"80",
          7349 => x"82",
          7350 => x"d8",
          7351 => x"3d",
          7352 => x"3d",
          7353 => x"84",
          7354 => x"05",
          7355 => x"80",
          7356 => x"51",
          7357 => x"82",
          7358 => x"58",
          7359 => x"0b",
          7360 => x"08",
          7361 => x"38",
          7362 => x"08",
          7363 => x"f0",
          7364 => x"08",
          7365 => x"56",
          7366 => x"86",
          7367 => x"75",
          7368 => x"fe",
          7369 => x"54",
          7370 => x"2e",
          7371 => x"14",
          7372 => x"a0",
          7373 => x"c8",
          7374 => x"06",
          7375 => x"54",
          7376 => x"38",
          7377 => x"86",
          7378 => x"82",
          7379 => x"06",
          7380 => x"56",
          7381 => x"38",
          7382 => x"80",
          7383 => x"81",
          7384 => x"52",
          7385 => x"51",
          7386 => x"82",
          7387 => x"81",
          7388 => x"81",
          7389 => x"83",
          7390 => x"8f",
          7391 => x"2e",
          7392 => x"82",
          7393 => x"06",
          7394 => x"56",
          7395 => x"38",
          7396 => x"74",
          7397 => x"a3",
          7398 => x"c8",
          7399 => x"06",
          7400 => x"2e",
          7401 => x"80",
          7402 => x"3d",
          7403 => x"83",
          7404 => x"15",
          7405 => x"53",
          7406 => x"8d",
          7407 => x"15",
          7408 => x"3f",
          7409 => x"08",
          7410 => x"70",
          7411 => x"0c",
          7412 => x"16",
          7413 => x"80",
          7414 => x"80",
          7415 => x"54",
          7416 => x"84",
          7417 => x"5b",
          7418 => x"80",
          7419 => x"7a",
          7420 => x"fc",
          7421 => x"d8",
          7422 => x"ff",
          7423 => x"77",
          7424 => x"81",
          7425 => x"76",
          7426 => x"81",
          7427 => x"2e",
          7428 => x"8d",
          7429 => x"26",
          7430 => x"80",
          7431 => x"ca",
          7432 => x"d8",
          7433 => x"ff",
          7434 => x"72",
          7435 => x"09",
          7436 => x"d7",
          7437 => x"14",
          7438 => x"3f",
          7439 => x"08",
          7440 => x"06",
          7441 => x"38",
          7442 => x"51",
          7443 => x"82",
          7444 => x"58",
          7445 => x"0c",
          7446 => x"33",
          7447 => x"80",
          7448 => x"ff",
          7449 => x"ff",
          7450 => x"55",
          7451 => x"81",
          7452 => x"38",
          7453 => x"06",
          7454 => x"80",
          7455 => x"52",
          7456 => x"8a",
          7457 => x"80",
          7458 => x"ff",
          7459 => x"53",
          7460 => x"86",
          7461 => x"83",
          7462 => x"c9",
          7463 => x"ca",
          7464 => x"c8",
          7465 => x"d8",
          7466 => x"15",
          7467 => x"06",
          7468 => x"76",
          7469 => x"80",
          7470 => x"c9",
          7471 => x"d8",
          7472 => x"ff",
          7473 => x"74",
          7474 => x"d8",
          7475 => x"b1",
          7476 => x"c8",
          7477 => x"c6",
          7478 => x"8e",
          7479 => x"c8",
          7480 => x"ff",
          7481 => x"56",
          7482 => x"83",
          7483 => x"14",
          7484 => x"71",
          7485 => x"5a",
          7486 => x"26",
          7487 => x"8a",
          7488 => x"74",
          7489 => x"fe",
          7490 => x"82",
          7491 => x"55",
          7492 => x"08",
          7493 => x"f3",
          7494 => x"c8",
          7495 => x"ff",
          7496 => x"83",
          7497 => x"74",
          7498 => x"26",
          7499 => x"57",
          7500 => x"26",
          7501 => x"57",
          7502 => x"56",
          7503 => x"82",
          7504 => x"15",
          7505 => x"0c",
          7506 => x"0c",
          7507 => x"a8",
          7508 => x"1d",
          7509 => x"54",
          7510 => x"2e",
          7511 => x"af",
          7512 => x"14",
          7513 => x"3f",
          7514 => x"08",
          7515 => x"06",
          7516 => x"72",
          7517 => x"79",
          7518 => x"80",
          7519 => x"c8",
          7520 => x"d8",
          7521 => x"15",
          7522 => x"2b",
          7523 => x"8d",
          7524 => x"2e",
          7525 => x"77",
          7526 => x"0c",
          7527 => x"76",
          7528 => x"38",
          7529 => x"70",
          7530 => x"81",
          7531 => x"53",
          7532 => x"89",
          7533 => x"56",
          7534 => x"08",
          7535 => x"38",
          7536 => x"15",
          7537 => x"90",
          7538 => x"80",
          7539 => x"34",
          7540 => x"09",
          7541 => x"92",
          7542 => x"14",
          7543 => x"3f",
          7544 => x"08",
          7545 => x"06",
          7546 => x"2e",
          7547 => x"80",
          7548 => x"1b",
          7549 => x"ca",
          7550 => x"d8",
          7551 => x"ea",
          7552 => x"c8",
          7553 => x"34",
          7554 => x"51",
          7555 => x"82",
          7556 => x"83",
          7557 => x"53",
          7558 => x"d5",
          7559 => x"06",
          7560 => x"b8",
          7561 => x"d9",
          7562 => x"c8",
          7563 => x"85",
          7564 => x"09",
          7565 => x"38",
          7566 => x"51",
          7567 => x"82",
          7568 => x"86",
          7569 => x"f2",
          7570 => x"06",
          7571 => x"a0",
          7572 => x"ad",
          7573 => x"c8",
          7574 => x"0c",
          7575 => x"51",
          7576 => x"82",
          7577 => x"90",
          7578 => x"74",
          7579 => x"a0",
          7580 => x"53",
          7581 => x"a0",
          7582 => x"15",
          7583 => x"a8",
          7584 => x"0c",
          7585 => x"15",
          7586 => x"75",
          7587 => x"0c",
          7588 => x"04",
          7589 => x"77",
          7590 => x"73",
          7591 => x"38",
          7592 => x"72",
          7593 => x"38",
          7594 => x"71",
          7595 => x"38",
          7596 => x"84",
          7597 => x"52",
          7598 => x"09",
          7599 => x"38",
          7600 => x"51",
          7601 => x"3f",
          7602 => x"08",
          7603 => x"71",
          7604 => x"74",
          7605 => x"83",
          7606 => x"78",
          7607 => x"52",
          7608 => x"c8",
          7609 => x"0d",
          7610 => x"0d",
          7611 => x"33",
          7612 => x"3d",
          7613 => x"56",
          7614 => x"8b",
          7615 => x"82",
          7616 => x"24",
          7617 => x"d8",
          7618 => x"29",
          7619 => x"05",
          7620 => x"55",
          7621 => x"84",
          7622 => x"34",
          7623 => x"80",
          7624 => x"80",
          7625 => x"75",
          7626 => x"75",
          7627 => x"38",
          7628 => x"3d",
          7629 => x"05",
          7630 => x"3f",
          7631 => x"08",
          7632 => x"d8",
          7633 => x"3d",
          7634 => x"3d",
          7635 => x"84",
          7636 => x"05",
          7637 => x"89",
          7638 => x"2e",
          7639 => x"77",
          7640 => x"54",
          7641 => x"05",
          7642 => x"84",
          7643 => x"f6",
          7644 => x"d8",
          7645 => x"82",
          7646 => x"84",
          7647 => x"5c",
          7648 => x"3d",
          7649 => x"ea",
          7650 => x"d8",
          7651 => x"82",
          7652 => x"92",
          7653 => x"d7",
          7654 => x"98",
          7655 => x"73",
          7656 => x"38",
          7657 => x"9c",
          7658 => x"80",
          7659 => x"38",
          7660 => x"95",
          7661 => x"2e",
          7662 => x"aa",
          7663 => x"df",
          7664 => x"d8",
          7665 => x"9e",
          7666 => x"05",
          7667 => x"54",
          7668 => x"38",
          7669 => x"70",
          7670 => x"54",
          7671 => x"8e",
          7672 => x"83",
          7673 => x"88",
          7674 => x"83",
          7675 => x"83",
          7676 => x"06",
          7677 => x"80",
          7678 => x"38",
          7679 => x"51",
          7680 => x"82",
          7681 => x"56",
          7682 => x"0a",
          7683 => x"05",
          7684 => x"3f",
          7685 => x"0b",
          7686 => x"80",
          7687 => x"7a",
          7688 => x"3f",
          7689 => x"9c",
          7690 => x"9e",
          7691 => x"81",
          7692 => x"34",
          7693 => x"80",
          7694 => x"b4",
          7695 => x"54",
          7696 => x"52",
          7697 => x"05",
          7698 => x"3f",
          7699 => x"08",
          7700 => x"c8",
          7701 => x"38",
          7702 => x"82",
          7703 => x"b2",
          7704 => x"84",
          7705 => x"06",
          7706 => x"73",
          7707 => x"38",
          7708 => x"ad",
          7709 => x"2a",
          7710 => x"51",
          7711 => x"2e",
          7712 => x"81",
          7713 => x"80",
          7714 => x"87",
          7715 => x"39",
          7716 => x"51",
          7717 => x"82",
          7718 => x"7b",
          7719 => x"12",
          7720 => x"82",
          7721 => x"81",
          7722 => x"83",
          7723 => x"06",
          7724 => x"80",
          7725 => x"77",
          7726 => x"58",
          7727 => x"08",
          7728 => x"63",
          7729 => x"63",
          7730 => x"57",
          7731 => x"82",
          7732 => x"82",
          7733 => x"88",
          7734 => x"9c",
          7735 => x"c1",
          7736 => x"d8",
          7737 => x"d8",
          7738 => x"1b",
          7739 => x"0c",
          7740 => x"22",
          7741 => x"77",
          7742 => x"80",
          7743 => x"34",
          7744 => x"1a",
          7745 => x"94",
          7746 => x"85",
          7747 => x"06",
          7748 => x"80",
          7749 => x"38",
          7750 => x"08",
          7751 => x"84",
          7752 => x"c8",
          7753 => x"0c",
          7754 => x"70",
          7755 => x"52",
          7756 => x"39",
          7757 => x"51",
          7758 => x"82",
          7759 => x"57",
          7760 => x"08",
          7761 => x"38",
          7762 => x"d8",
          7763 => x"2e",
          7764 => x"83",
          7765 => x"75",
          7766 => x"74",
          7767 => x"07",
          7768 => x"54",
          7769 => x"8a",
          7770 => x"75",
          7771 => x"73",
          7772 => x"98",
          7773 => x"a9",
          7774 => x"ff",
          7775 => x"80",
          7776 => x"76",
          7777 => x"c5",
          7778 => x"d8",
          7779 => x"38",
          7780 => x"39",
          7781 => x"82",
          7782 => x"05",
          7783 => x"84",
          7784 => x"0c",
          7785 => x"82",
          7786 => x"98",
          7787 => x"f2",
          7788 => x"63",
          7789 => x"40",
          7790 => x"7e",
          7791 => x"fc",
          7792 => x"51",
          7793 => x"82",
          7794 => x"55",
          7795 => x"08",
          7796 => x"19",
          7797 => x"80",
          7798 => x"74",
          7799 => x"39",
          7800 => x"81",
          7801 => x"56",
          7802 => x"82",
          7803 => x"39",
          7804 => x"1a",
          7805 => x"82",
          7806 => x"0b",
          7807 => x"81",
          7808 => x"39",
          7809 => x"94",
          7810 => x"55",
          7811 => x"83",
          7812 => x"7b",
          7813 => x"8c",
          7814 => x"08",
          7815 => x"06",
          7816 => x"81",
          7817 => x"8a",
          7818 => x"05",
          7819 => x"06",
          7820 => x"a8",
          7821 => x"38",
          7822 => x"55",
          7823 => x"19",
          7824 => x"51",
          7825 => x"82",
          7826 => x"55",
          7827 => x"ff",
          7828 => x"ff",
          7829 => x"38",
          7830 => x"0c",
          7831 => x"52",
          7832 => x"d6",
          7833 => x"c8",
          7834 => x"ff",
          7835 => x"d8",
          7836 => x"7c",
          7837 => x"57",
          7838 => x"80",
          7839 => x"1a",
          7840 => x"22",
          7841 => x"75",
          7842 => x"38",
          7843 => x"58",
          7844 => x"53",
          7845 => x"1b",
          7846 => x"b8",
          7847 => x"d8",
          7848 => x"d6",
          7849 => x"11",
          7850 => x"74",
          7851 => x"38",
          7852 => x"77",
          7853 => x"78",
          7854 => x"84",
          7855 => x"16",
          7856 => x"08",
          7857 => x"2b",
          7858 => x"ff",
          7859 => x"77",
          7860 => x"ba",
          7861 => x"1a",
          7862 => x"08",
          7863 => x"84",
          7864 => x"57",
          7865 => x"27",
          7866 => x"56",
          7867 => x"52",
          7868 => x"d0",
          7869 => x"c8",
          7870 => x"38",
          7871 => x"19",
          7872 => x"06",
          7873 => x"52",
          7874 => x"bd",
          7875 => x"76",
          7876 => x"17",
          7877 => x"1e",
          7878 => x"18",
          7879 => x"5e",
          7880 => x"39",
          7881 => x"82",
          7882 => x"90",
          7883 => x"f2",
          7884 => x"63",
          7885 => x"40",
          7886 => x"7e",
          7887 => x"fc",
          7888 => x"51",
          7889 => x"82",
          7890 => x"55",
          7891 => x"08",
          7892 => x"18",
          7893 => x"80",
          7894 => x"74",
          7895 => x"39",
          7896 => x"70",
          7897 => x"81",
          7898 => x"56",
          7899 => x"80",
          7900 => x"38",
          7901 => x"0b",
          7902 => x"82",
          7903 => x"39",
          7904 => x"19",
          7905 => x"83",
          7906 => x"18",
          7907 => x"56",
          7908 => x"27",
          7909 => x"09",
          7910 => x"2e",
          7911 => x"94",
          7912 => x"83",
          7913 => x"56",
          7914 => x"38",
          7915 => x"22",
          7916 => x"89",
          7917 => x"55",
          7918 => x"75",
          7919 => x"18",
          7920 => x"9c",
          7921 => x"85",
          7922 => x"08",
          7923 => x"c6",
          7924 => x"d8",
          7925 => x"82",
          7926 => x"80",
          7927 => x"38",
          7928 => x"ff",
          7929 => x"ff",
          7930 => x"38",
          7931 => x"0c",
          7932 => x"85",
          7933 => x"19",
          7934 => x"b4",
          7935 => x"19",
          7936 => x"81",
          7937 => x"74",
          7938 => x"c8",
          7939 => x"c8",
          7940 => x"38",
          7941 => x"52",
          7942 => x"9e",
          7943 => x"c8",
          7944 => x"fe",
          7945 => x"d8",
          7946 => x"7c",
          7947 => x"57",
          7948 => x"80",
          7949 => x"1b",
          7950 => x"22",
          7951 => x"75",
          7952 => x"38",
          7953 => x"59",
          7954 => x"53",
          7955 => x"1a",
          7956 => x"b7",
          7957 => x"d8",
          7958 => x"a4",
          7959 => x"11",
          7960 => x"56",
          7961 => x"27",
          7962 => x"80",
          7963 => x"08",
          7964 => x"2b",
          7965 => x"b8",
          7966 => x"ba",
          7967 => x"55",
          7968 => x"16",
          7969 => x"2b",
          7970 => x"39",
          7971 => x"94",
          7972 => x"94",
          7973 => x"ff",
          7974 => x"82",
          7975 => x"fd",
          7976 => x"77",
          7977 => x"55",
          7978 => x"0c",
          7979 => x"83",
          7980 => x"80",
          7981 => x"55",
          7982 => x"83",
          7983 => x"9c",
          7984 => x"7e",
          7985 => x"fc",
          7986 => x"c8",
          7987 => x"38",
          7988 => x"52",
          7989 => x"83",
          7990 => x"b8",
          7991 => x"ba",
          7992 => x"55",
          7993 => x"16",
          7994 => x"31",
          7995 => x"7f",
          7996 => x"94",
          7997 => x"70",
          7998 => x"8c",
          7999 => x"58",
          8000 => x"76",
          8001 => x"75",
          8002 => x"19",
          8003 => x"39",
          8004 => x"80",
          8005 => x"74",
          8006 => x"80",
          8007 => x"d8",
          8008 => x"3d",
          8009 => x"3d",
          8010 => x"3d",
          8011 => x"70",
          8012 => x"e0",
          8013 => x"c8",
          8014 => x"d8",
          8015 => x"80",
          8016 => x"33",
          8017 => x"70",
          8018 => x"55",
          8019 => x"2e",
          8020 => x"a0",
          8021 => x"78",
          8022 => x"e8",
          8023 => x"c8",
          8024 => x"d8",
          8025 => x"d8",
          8026 => x"08",
          8027 => x"a0",
          8028 => x"73",
          8029 => x"88",
          8030 => x"74",
          8031 => x"51",
          8032 => x"8c",
          8033 => x"9c",
          8034 => x"b8",
          8035 => x"88",
          8036 => x"96",
          8037 => x"b8",
          8038 => x"52",
          8039 => x"ff",
          8040 => x"78",
          8041 => x"83",
          8042 => x"51",
          8043 => x"3f",
          8044 => x"08",
          8045 => x"81",
          8046 => x"57",
          8047 => x"34",
          8048 => x"c8",
          8049 => x"0d",
          8050 => x"0d",
          8051 => x"54",
          8052 => x"82",
          8053 => x"53",
          8054 => x"08",
          8055 => x"3d",
          8056 => x"73",
          8057 => x"3f",
          8058 => x"08",
          8059 => x"c8",
          8060 => x"82",
          8061 => x"74",
          8062 => x"d8",
          8063 => x"3d",
          8064 => x"3d",
          8065 => x"51",
          8066 => x"8b",
          8067 => x"82",
          8068 => x"24",
          8069 => x"d8",
          8070 => x"f0",
          8071 => x"52",
          8072 => x"c8",
          8073 => x"0d",
          8074 => x"0d",
          8075 => x"3d",
          8076 => x"95",
          8077 => x"aa",
          8078 => x"c8",
          8079 => x"d8",
          8080 => x"e0",
          8081 => x"64",
          8082 => x"d0",
          8083 => x"ac",
          8084 => x"c8",
          8085 => x"d8",
          8086 => x"38",
          8087 => x"05",
          8088 => x"2b",
          8089 => x"80",
          8090 => x"76",
          8091 => x"0c",
          8092 => x"02",
          8093 => x"70",
          8094 => x"81",
          8095 => x"56",
          8096 => x"9e",
          8097 => x"53",
          8098 => x"ca",
          8099 => x"d8",
          8100 => x"15",
          8101 => x"82",
          8102 => x"84",
          8103 => x"06",
          8104 => x"55",
          8105 => x"c8",
          8106 => x"0d",
          8107 => x"3d",
          8108 => x"3d",
          8109 => x"3d",
          8110 => x"80",
          8111 => x"53",
          8112 => x"fd",
          8113 => x"80",
          8114 => x"e8",
          8115 => x"d8",
          8116 => x"82",
          8117 => x"83",
          8118 => x"80",
          8119 => x"7a",
          8120 => x"08",
          8121 => x"0c",
          8122 => x"d5",
          8123 => x"73",
          8124 => x"83",
          8125 => x"80",
          8126 => x"52",
          8127 => x"3f",
          8128 => x"08",
          8129 => x"c8",
          8130 => x"38",
          8131 => x"08",
          8132 => x"ff",
          8133 => x"82",
          8134 => x"57",
          8135 => x"08",
          8136 => x"80",
          8137 => x"52",
          8138 => x"86",
          8139 => x"c8",
          8140 => x"3d",
          8141 => x"74",
          8142 => x"3f",
          8143 => x"08",
          8144 => x"c8",
          8145 => x"38",
          8146 => x"51",
          8147 => x"82",
          8148 => x"57",
          8149 => x"08",
          8150 => x"da",
          8151 => x"7b",
          8152 => x"3f",
          8153 => x"c8",
          8154 => x"38",
          8155 => x"51",
          8156 => x"82",
          8157 => x"57",
          8158 => x"08",
          8159 => x"38",
          8160 => x"09",
          8161 => x"38",
          8162 => x"ee",
          8163 => x"ea",
          8164 => x"3d",
          8165 => x"52",
          8166 => x"e4",
          8167 => x"3d",
          8168 => x"11",
          8169 => x"5a",
          8170 => x"2e",
          8171 => x"80",
          8172 => x"81",
          8173 => x"70",
          8174 => x"56",
          8175 => x"81",
          8176 => x"78",
          8177 => x"38",
          8178 => x"9c",
          8179 => x"82",
          8180 => x"18",
          8181 => x"08",
          8182 => x"ff",
          8183 => x"55",
          8184 => x"74",
          8185 => x"38",
          8186 => x"e1",
          8187 => x"55",
          8188 => x"34",
          8189 => x"77",
          8190 => x"81",
          8191 => x"ff",
          8192 => x"3d",
          8193 => x"58",
          8194 => x"80",
          8195 => x"a4",
          8196 => x"29",
          8197 => x"05",
          8198 => x"33",
          8199 => x"56",
          8200 => x"2e",
          8201 => x"16",
          8202 => x"33",
          8203 => x"73",
          8204 => x"16",
          8205 => x"26",
          8206 => x"55",
          8207 => x"91",
          8208 => x"54",
          8209 => x"70",
          8210 => x"34",
          8211 => x"ec",
          8212 => x"70",
          8213 => x"34",
          8214 => x"09",
          8215 => x"38",
          8216 => x"39",
          8217 => x"08",
          8218 => x"59",
          8219 => x"7a",
          8220 => x"5c",
          8221 => x"26",
          8222 => x"7a",
          8223 => x"d8",
          8224 => x"df",
          8225 => x"f7",
          8226 => x"7d",
          8227 => x"05",
          8228 => x"57",
          8229 => x"3f",
          8230 => x"08",
          8231 => x"c8",
          8232 => x"38",
          8233 => x"53",
          8234 => x"38",
          8235 => x"54",
          8236 => x"92",
          8237 => x"33",
          8238 => x"70",
          8239 => x"54",
          8240 => x"38",
          8241 => x"15",
          8242 => x"70",
          8243 => x"58",
          8244 => x"82",
          8245 => x"8a",
          8246 => x"89",
          8247 => x"53",
          8248 => x"b7",
          8249 => x"ff",
          8250 => x"c5",
          8251 => x"d8",
          8252 => x"15",
          8253 => x"53",
          8254 => x"c5",
          8255 => x"d8",
          8256 => x"26",
          8257 => x"30",
          8258 => x"70",
          8259 => x"77",
          8260 => x"18",
          8261 => x"51",
          8262 => x"88",
          8263 => x"73",
          8264 => x"52",
          8265 => x"bc",
          8266 => x"d8",
          8267 => x"82",
          8268 => x"81",
          8269 => x"38",
          8270 => x"08",
          8271 => x"9e",
          8272 => x"c8",
          8273 => x"0c",
          8274 => x"0c",
          8275 => x"81",
          8276 => x"76",
          8277 => x"38",
          8278 => x"94",
          8279 => x"94",
          8280 => x"16",
          8281 => x"2a",
          8282 => x"51",
          8283 => x"72",
          8284 => x"38",
          8285 => x"51",
          8286 => x"3f",
          8287 => x"08",
          8288 => x"c8",
          8289 => x"82",
          8290 => x"56",
          8291 => x"52",
          8292 => x"b5",
          8293 => x"d8",
          8294 => x"73",
          8295 => x"38",
          8296 => x"b0",
          8297 => x"73",
          8298 => x"27",
          8299 => x"98",
          8300 => x"9e",
          8301 => x"08",
          8302 => x"0c",
          8303 => x"06",
          8304 => x"2e",
          8305 => x"52",
          8306 => x"b4",
          8307 => x"d8",
          8308 => x"38",
          8309 => x"16",
          8310 => x"80",
          8311 => x"0b",
          8312 => x"81",
          8313 => x"75",
          8314 => x"d8",
          8315 => x"58",
          8316 => x"54",
          8317 => x"74",
          8318 => x"73",
          8319 => x"90",
          8320 => x"c0",
          8321 => x"90",
          8322 => x"83",
          8323 => x"72",
          8324 => x"38",
          8325 => x"08",
          8326 => x"77",
          8327 => x"80",
          8328 => x"d8",
          8329 => x"3d",
          8330 => x"3d",
          8331 => x"89",
          8332 => x"2e",
          8333 => x"80",
          8334 => x"fc",
          8335 => x"3d",
          8336 => x"e1",
          8337 => x"d8",
          8338 => x"82",
          8339 => x"80",
          8340 => x"76",
          8341 => x"75",
          8342 => x"3f",
          8343 => x"08",
          8344 => x"c8",
          8345 => x"38",
          8346 => x"70",
          8347 => x"57",
          8348 => x"a2",
          8349 => x"33",
          8350 => x"70",
          8351 => x"55",
          8352 => x"2e",
          8353 => x"16",
          8354 => x"51",
          8355 => x"82",
          8356 => x"88",
          8357 => x"54",
          8358 => x"84",
          8359 => x"52",
          8360 => x"bd",
          8361 => x"d8",
          8362 => x"74",
          8363 => x"81",
          8364 => x"85",
          8365 => x"74",
          8366 => x"38",
          8367 => x"74",
          8368 => x"d8",
          8369 => x"3d",
          8370 => x"3d",
          8371 => x"3d",
          8372 => x"70",
          8373 => x"bc",
          8374 => x"c8",
          8375 => x"82",
          8376 => x"73",
          8377 => x"0d",
          8378 => x"0d",
          8379 => x"3d",
          8380 => x"71",
          8381 => x"e7",
          8382 => x"d8",
          8383 => x"82",
          8384 => x"80",
          8385 => x"94",
          8386 => x"c8",
          8387 => x"51",
          8388 => x"3f",
          8389 => x"08",
          8390 => x"39",
          8391 => x"08",
          8392 => x"c2",
          8393 => x"d8",
          8394 => x"82",
          8395 => x"84",
          8396 => x"06",
          8397 => x"53",
          8398 => x"d8",
          8399 => x"38",
          8400 => x"51",
          8401 => x"72",
          8402 => x"ff",
          8403 => x"82",
          8404 => x"84",
          8405 => x"70",
          8406 => x"2c",
          8407 => x"c8",
          8408 => x"51",
          8409 => x"82",
          8410 => x"87",
          8411 => x"ed",
          8412 => x"57",
          8413 => x"3d",
          8414 => x"3d",
          8415 => x"e2",
          8416 => x"c8",
          8417 => x"d8",
          8418 => x"38",
          8419 => x"51",
          8420 => x"82",
          8421 => x"55",
          8422 => x"08",
          8423 => x"80",
          8424 => x"70",
          8425 => x"58",
          8426 => x"85",
          8427 => x"8d",
          8428 => x"2e",
          8429 => x"52",
          8430 => x"c4",
          8431 => x"d8",
          8432 => x"3d",
          8433 => x"3d",
          8434 => x"55",
          8435 => x"92",
          8436 => x"52",
          8437 => x"de",
          8438 => x"d8",
          8439 => x"82",
          8440 => x"82",
          8441 => x"74",
          8442 => x"9c",
          8443 => x"11",
          8444 => x"59",
          8445 => x"75",
          8446 => x"38",
          8447 => x"81",
          8448 => x"5b",
          8449 => x"82",
          8450 => x"39",
          8451 => x"08",
          8452 => x"59",
          8453 => x"09",
          8454 => x"c0",
          8455 => x"5f",
          8456 => x"92",
          8457 => x"51",
          8458 => x"3f",
          8459 => x"08",
          8460 => x"38",
          8461 => x"08",
          8462 => x"38",
          8463 => x"08",
          8464 => x"d8",
          8465 => x"80",
          8466 => x"81",
          8467 => x"59",
          8468 => x"14",
          8469 => x"c9",
          8470 => x"39",
          8471 => x"82",
          8472 => x"57",
          8473 => x"38",
          8474 => x"18",
          8475 => x"ff",
          8476 => x"82",
          8477 => x"5b",
          8478 => x"08",
          8479 => x"7c",
          8480 => x"12",
          8481 => x"52",
          8482 => x"82",
          8483 => x"06",
          8484 => x"14",
          8485 => x"d2",
          8486 => x"c8",
          8487 => x"ff",
          8488 => x"70",
          8489 => x"82",
          8490 => x"51",
          8491 => x"b8",
          8492 => x"a9",
          8493 => x"d8",
          8494 => x"0a",
          8495 => x"70",
          8496 => x"84",
          8497 => x"51",
          8498 => x"ff",
          8499 => x"56",
          8500 => x"38",
          8501 => x"7c",
          8502 => x"0c",
          8503 => x"81",
          8504 => x"74",
          8505 => x"7a",
          8506 => x"0c",
          8507 => x"04",
          8508 => x"79",
          8509 => x"05",
          8510 => x"57",
          8511 => x"82",
          8512 => x"56",
          8513 => x"08",
          8514 => x"91",
          8515 => x"75",
          8516 => x"90",
          8517 => x"81",
          8518 => x"06",
          8519 => x"87",
          8520 => x"2e",
          8521 => x"94",
          8522 => x"73",
          8523 => x"27",
          8524 => x"73",
          8525 => x"d8",
          8526 => x"88",
          8527 => x"76",
          8528 => x"d0",
          8529 => x"c8",
          8530 => x"19",
          8531 => x"ca",
          8532 => x"08",
          8533 => x"ff",
          8534 => x"82",
          8535 => x"ff",
          8536 => x"06",
          8537 => x"56",
          8538 => x"08",
          8539 => x"81",
          8540 => x"82",
          8541 => x"75",
          8542 => x"54",
          8543 => x"08",
          8544 => x"27",
          8545 => x"17",
          8546 => x"d8",
          8547 => x"76",
          8548 => x"80",
          8549 => x"c8",
          8550 => x"17",
          8551 => x"0c",
          8552 => x"80",
          8553 => x"73",
          8554 => x"75",
          8555 => x"38",
          8556 => x"34",
          8557 => x"82",
          8558 => x"89",
          8559 => x"e0",
          8560 => x"53",
          8561 => x"9c",
          8562 => x"3d",
          8563 => x"3f",
          8564 => x"08",
          8565 => x"c8",
          8566 => x"38",
          8567 => x"3d",
          8568 => x"3d",
          8569 => x"ce",
          8570 => x"d8",
          8571 => x"82",
          8572 => x"81",
          8573 => x"80",
          8574 => x"70",
          8575 => x"81",
          8576 => x"56",
          8577 => x"81",
          8578 => x"98",
          8579 => x"74",
          8580 => x"38",
          8581 => x"05",
          8582 => x"06",
          8583 => x"55",
          8584 => x"38",
          8585 => x"51",
          8586 => x"3f",
          8587 => x"08",
          8588 => x"70",
          8589 => x"55",
          8590 => x"2e",
          8591 => x"78",
          8592 => x"c8",
          8593 => x"08",
          8594 => x"38",
          8595 => x"d8",
          8596 => x"76",
          8597 => x"70",
          8598 => x"b5",
          8599 => x"d8",
          8600 => x"82",
          8601 => x"80",
          8602 => x"d8",
          8603 => x"73",
          8604 => x"d4",
          8605 => x"c8",
          8606 => x"d8",
          8607 => x"38",
          8608 => x"d0",
          8609 => x"c8",
          8610 => x"88",
          8611 => x"c8",
          8612 => x"38",
          8613 => x"ef",
          8614 => x"c8",
          8615 => x"c8",
          8616 => x"82",
          8617 => x"07",
          8618 => x"55",
          8619 => x"2e",
          8620 => x"80",
          8621 => x"80",
          8622 => x"77",
          8623 => x"d4",
          8624 => x"c8",
          8625 => x"8c",
          8626 => x"ff",
          8627 => x"82",
          8628 => x"55",
          8629 => x"c8",
          8630 => x"0d",
          8631 => x"0d",
          8632 => x"3d",
          8633 => x"52",
          8634 => x"d7",
          8635 => x"d8",
          8636 => x"82",
          8637 => x"82",
          8638 => x"5e",
          8639 => x"3d",
          8640 => x"cb",
          8641 => x"d8",
          8642 => x"82",
          8643 => x"86",
          8644 => x"82",
          8645 => x"d8",
          8646 => x"2e",
          8647 => x"82",
          8648 => x"80",
          8649 => x"70",
          8650 => x"06",
          8651 => x"54",
          8652 => x"38",
          8653 => x"52",
          8654 => x"52",
          8655 => x"80",
          8656 => x"c8",
          8657 => x"56",
          8658 => x"08",
          8659 => x"54",
          8660 => x"08",
          8661 => x"81",
          8662 => x"82",
          8663 => x"c8",
          8664 => x"09",
          8665 => x"38",
          8666 => x"ba",
          8667 => x"b6",
          8668 => x"c8",
          8669 => x"51",
          8670 => x"3f",
          8671 => x"08",
          8672 => x"c8",
          8673 => x"38",
          8674 => x"52",
          8675 => x"ff",
          8676 => x"78",
          8677 => x"b8",
          8678 => x"54",
          8679 => x"c3",
          8680 => x"88",
          8681 => x"80",
          8682 => x"ff",
          8683 => x"75",
          8684 => x"11",
          8685 => x"b8",
          8686 => x"53",
          8687 => x"53",
          8688 => x"51",
          8689 => x"3f",
          8690 => x"0b",
          8691 => x"34",
          8692 => x"80",
          8693 => x"51",
          8694 => x"3f",
          8695 => x"0b",
          8696 => x"77",
          8697 => x"cd",
          8698 => x"c8",
          8699 => x"d8",
          8700 => x"38",
          8701 => x"0a",
          8702 => x"05",
          8703 => x"ca",
          8704 => x"64",
          8705 => x"ff",
          8706 => x"64",
          8707 => x"8b",
          8708 => x"54",
          8709 => x"15",
          8710 => x"ff",
          8711 => x"82",
          8712 => x"54",
          8713 => x"53",
          8714 => x"51",
          8715 => x"3f",
          8716 => x"c8",
          8717 => x"0d",
          8718 => x"0d",
          8719 => x"05",
          8720 => x"3f",
          8721 => x"3d",
          8722 => x"52",
          8723 => x"d5",
          8724 => x"d8",
          8725 => x"82",
          8726 => x"82",
          8727 => x"4e",
          8728 => x"52",
          8729 => x"52",
          8730 => x"3f",
          8731 => x"08",
          8732 => x"c8",
          8733 => x"38",
          8734 => x"05",
          8735 => x"06",
          8736 => x"73",
          8737 => x"a0",
          8738 => x"08",
          8739 => x"ff",
          8740 => x"ff",
          8741 => x"b0",
          8742 => x"92",
          8743 => x"54",
          8744 => x"3f",
          8745 => x"52",
          8746 => x"d0",
          8747 => x"c8",
          8748 => x"d8",
          8749 => x"38",
          8750 => x"08",
          8751 => x"06",
          8752 => x"a3",
          8753 => x"92",
          8754 => x"81",
          8755 => x"d8",
          8756 => x"2e",
          8757 => x"81",
          8758 => x"51",
          8759 => x"3f",
          8760 => x"08",
          8761 => x"c8",
          8762 => x"38",
          8763 => x"53",
          8764 => x"8d",
          8765 => x"16",
          8766 => x"fd",
          8767 => x"05",
          8768 => x"34",
          8769 => x"70",
          8770 => x"81",
          8771 => x"55",
          8772 => x"74",
          8773 => x"73",
          8774 => x"78",
          8775 => x"83",
          8776 => x"16",
          8777 => x"2a",
          8778 => x"51",
          8779 => x"80",
          8780 => x"38",
          8781 => x"80",
          8782 => x"52",
          8783 => x"b4",
          8784 => x"d8",
          8785 => x"78",
          8786 => x"ee",
          8787 => x"82",
          8788 => x"80",
          8789 => x"38",
          8790 => x"08",
          8791 => x"ff",
          8792 => x"82",
          8793 => x"79",
          8794 => x"58",
          8795 => x"d8",
          8796 => x"c1",
          8797 => x"33",
          8798 => x"2e",
          8799 => x"9a",
          8800 => x"75",
          8801 => x"ff",
          8802 => x"78",
          8803 => x"83",
          8804 => x"39",
          8805 => x"08",
          8806 => x"51",
          8807 => x"82",
          8808 => x"55",
          8809 => x"08",
          8810 => x"51",
          8811 => x"3f",
          8812 => x"08",
          8813 => x"d8",
          8814 => x"3d",
          8815 => x"3d",
          8816 => x"df",
          8817 => x"84",
          8818 => x"05",
          8819 => x"82",
          8820 => x"cc",
          8821 => x"3d",
          8822 => x"3f",
          8823 => x"08",
          8824 => x"c8",
          8825 => x"38",
          8826 => x"52",
          8827 => x"05",
          8828 => x"3f",
          8829 => x"08",
          8830 => x"c8",
          8831 => x"02",
          8832 => x"33",
          8833 => x"54",
          8834 => x"aa",
          8835 => x"06",
          8836 => x"8b",
          8837 => x"06",
          8838 => x"07",
          8839 => x"56",
          8840 => x"34",
          8841 => x"0b",
          8842 => x"78",
          8843 => x"db",
          8844 => x"c8",
          8845 => x"82",
          8846 => x"96",
          8847 => x"ee",
          8848 => x"56",
          8849 => x"3d",
          8850 => x"95",
          8851 => x"92",
          8852 => x"c8",
          8853 => x"d8",
          8854 => x"cb",
          8855 => x"64",
          8856 => x"d0",
          8857 => x"94",
          8858 => x"c8",
          8859 => x"d8",
          8860 => x"38",
          8861 => x"05",
          8862 => x"06",
          8863 => x"73",
          8864 => x"16",
          8865 => x"22",
          8866 => x"07",
          8867 => x"1f",
          8868 => x"b6",
          8869 => x"81",
          8870 => x"34",
          8871 => x"a1",
          8872 => x"d8",
          8873 => x"74",
          8874 => x"0c",
          8875 => x"04",
          8876 => x"6a",
          8877 => x"80",
          8878 => x"cc",
          8879 => x"3d",
          8880 => x"3f",
          8881 => x"08",
          8882 => x"08",
          8883 => x"d8",
          8884 => x"80",
          8885 => x"57",
          8886 => x"81",
          8887 => x"70",
          8888 => x"55",
          8889 => x"80",
          8890 => x"5d",
          8891 => x"52",
          8892 => x"52",
          8893 => x"db",
          8894 => x"c8",
          8895 => x"d8",
          8896 => x"d2",
          8897 => x"73",
          8898 => x"bc",
          8899 => x"c8",
          8900 => x"d8",
          8901 => x"38",
          8902 => x"08",
          8903 => x"08",
          8904 => x"56",
          8905 => x"19",
          8906 => x"59",
          8907 => x"74",
          8908 => x"56",
          8909 => x"ec",
          8910 => x"75",
          8911 => x"74",
          8912 => x"2e",
          8913 => x"16",
          8914 => x"33",
          8915 => x"73",
          8916 => x"38",
          8917 => x"84",
          8918 => x"06",
          8919 => x"7a",
          8920 => x"76",
          8921 => x"07",
          8922 => x"54",
          8923 => x"80",
          8924 => x"80",
          8925 => x"7b",
          8926 => x"53",
          8927 => x"c4",
          8928 => x"c8",
          8929 => x"d8",
          8930 => x"38",
          8931 => x"55",
          8932 => x"56",
          8933 => x"8b",
          8934 => x"56",
          8935 => x"83",
          8936 => x"75",
          8937 => x"51",
          8938 => x"3f",
          8939 => x"08",
          8940 => x"82",
          8941 => x"99",
          8942 => x"e6",
          8943 => x"53",
          8944 => x"b4",
          8945 => x"3d",
          8946 => x"3f",
          8947 => x"08",
          8948 => x"08",
          8949 => x"d8",
          8950 => x"dd",
          8951 => x"a0",
          8952 => x"70",
          8953 => x"9c",
          8954 => x"6d",
          8955 => x"55",
          8956 => x"27",
          8957 => x"77",
          8958 => x"51",
          8959 => x"3f",
          8960 => x"08",
          8961 => x"26",
          8962 => x"82",
          8963 => x"51",
          8964 => x"83",
          8965 => x"d8",
          8966 => x"93",
          8967 => x"d8",
          8968 => x"ff",
          8969 => x"74",
          8970 => x"38",
          8971 => x"cb",
          8972 => x"9c",
          8973 => x"d8",
          8974 => x"38",
          8975 => x"27",
          8976 => x"89",
          8977 => x"8b",
          8978 => x"27",
          8979 => x"55",
          8980 => x"81",
          8981 => x"8f",
          8982 => x"2a",
          8983 => x"70",
          8984 => x"34",
          8985 => x"74",
          8986 => x"05",
          8987 => x"16",
          8988 => x"51",
          8989 => x"9f",
          8990 => x"38",
          8991 => x"54",
          8992 => x"81",
          8993 => x"b1",
          8994 => x"2e",
          8995 => x"a3",
          8996 => x"15",
          8997 => x"54",
          8998 => x"09",
          8999 => x"38",
          9000 => x"75",
          9001 => x"40",
          9002 => x"52",
          9003 => x"52",
          9004 => x"9f",
          9005 => x"c8",
          9006 => x"d8",
          9007 => x"f7",
          9008 => x"74",
          9009 => x"80",
          9010 => x"c8",
          9011 => x"d8",
          9012 => x"38",
          9013 => x"38",
          9014 => x"74",
          9015 => x"39",
          9016 => x"08",
          9017 => x"81",
          9018 => x"38",
          9019 => x"74",
          9020 => x"38",
          9021 => x"51",
          9022 => x"3f",
          9023 => x"08",
          9024 => x"c8",
          9025 => x"a0",
          9026 => x"c8",
          9027 => x"51",
          9028 => x"3f",
          9029 => x"0b",
          9030 => x"8b",
          9031 => x"66",
          9032 => x"d5",
          9033 => x"81",
          9034 => x"34",
          9035 => x"9c",
          9036 => x"d8",
          9037 => x"73",
          9038 => x"d8",
          9039 => x"3d",
          9040 => x"3d",
          9041 => x"02",
          9042 => x"cb",
          9043 => x"3d",
          9044 => x"72",
          9045 => x"5a",
          9046 => x"82",
          9047 => x"58",
          9048 => x"08",
          9049 => x"91",
          9050 => x"77",
          9051 => x"7c",
          9052 => x"38",
          9053 => x"59",
          9054 => x"90",
          9055 => x"81",
          9056 => x"06",
          9057 => x"73",
          9058 => x"54",
          9059 => x"82",
          9060 => x"39",
          9061 => x"8b",
          9062 => x"11",
          9063 => x"2b",
          9064 => x"54",
          9065 => x"fe",
          9066 => x"ff",
          9067 => x"70",
          9068 => x"07",
          9069 => x"d8",
          9070 => x"90",
          9071 => x"40",
          9072 => x"55",
          9073 => x"88",
          9074 => x"08",
          9075 => x"38",
          9076 => x"77",
          9077 => x"56",
          9078 => x"51",
          9079 => x"3f",
          9080 => x"55",
          9081 => x"08",
          9082 => x"38",
          9083 => x"d8",
          9084 => x"2e",
          9085 => x"82",
          9086 => x"ff",
          9087 => x"38",
          9088 => x"08",
          9089 => x"16",
          9090 => x"2e",
          9091 => x"87",
          9092 => x"74",
          9093 => x"74",
          9094 => x"81",
          9095 => x"38",
          9096 => x"ff",
          9097 => x"2e",
          9098 => x"7b",
          9099 => x"80",
          9100 => x"81",
          9101 => x"81",
          9102 => x"06",
          9103 => x"56",
          9104 => x"52",
          9105 => x"9e",
          9106 => x"d8",
          9107 => x"82",
          9108 => x"80",
          9109 => x"81",
          9110 => x"56",
          9111 => x"d3",
          9112 => x"ff",
          9113 => x"7c",
          9114 => x"55",
          9115 => x"b3",
          9116 => x"1b",
          9117 => x"1b",
          9118 => x"33",
          9119 => x"54",
          9120 => x"34",
          9121 => x"fe",
          9122 => x"08",
          9123 => x"74",
          9124 => x"75",
          9125 => x"16",
          9126 => x"33",
          9127 => x"73",
          9128 => x"77",
          9129 => x"d8",
          9130 => x"3d",
          9131 => x"3d",
          9132 => x"02",
          9133 => x"eb",
          9134 => x"3d",
          9135 => x"59",
          9136 => x"8b",
          9137 => x"82",
          9138 => x"24",
          9139 => x"82",
          9140 => x"84",
          9141 => x"90",
          9142 => x"51",
          9143 => x"2e",
          9144 => x"75",
          9145 => x"c8",
          9146 => x"06",
          9147 => x"7e",
          9148 => x"fe",
          9149 => x"c8",
          9150 => x"06",
          9151 => x"56",
          9152 => x"74",
          9153 => x"76",
          9154 => x"81",
          9155 => x"8a",
          9156 => x"b2",
          9157 => x"fc",
          9158 => x"52",
          9159 => x"93",
          9160 => x"d8",
          9161 => x"38",
          9162 => x"80",
          9163 => x"74",
          9164 => x"26",
          9165 => x"15",
          9166 => x"74",
          9167 => x"38",
          9168 => x"80",
          9169 => x"84",
          9170 => x"92",
          9171 => x"80",
          9172 => x"38",
          9173 => x"06",
          9174 => x"2e",
          9175 => x"56",
          9176 => x"78",
          9177 => x"89",
          9178 => x"2b",
          9179 => x"43",
          9180 => x"38",
          9181 => x"30",
          9182 => x"77",
          9183 => x"91",
          9184 => x"c2",
          9185 => x"f8",
          9186 => x"52",
          9187 => x"92",
          9188 => x"56",
          9189 => x"08",
          9190 => x"77",
          9191 => x"77",
          9192 => x"c8",
          9193 => x"45",
          9194 => x"bf",
          9195 => x"8e",
          9196 => x"26",
          9197 => x"74",
          9198 => x"48",
          9199 => x"75",
          9200 => x"38",
          9201 => x"81",
          9202 => x"fa",
          9203 => x"2a",
          9204 => x"56",
          9205 => x"2e",
          9206 => x"87",
          9207 => x"82",
          9208 => x"38",
          9209 => x"55",
          9210 => x"83",
          9211 => x"81",
          9212 => x"56",
          9213 => x"80",
          9214 => x"38",
          9215 => x"83",
          9216 => x"06",
          9217 => x"78",
          9218 => x"91",
          9219 => x"0b",
          9220 => x"22",
          9221 => x"80",
          9222 => x"74",
          9223 => x"38",
          9224 => x"56",
          9225 => x"17",
          9226 => x"57",
          9227 => x"2e",
          9228 => x"75",
          9229 => x"79",
          9230 => x"fe",
          9231 => x"82",
          9232 => x"84",
          9233 => x"05",
          9234 => x"5e",
          9235 => x"80",
          9236 => x"c8",
          9237 => x"8a",
          9238 => x"fd",
          9239 => x"75",
          9240 => x"38",
          9241 => x"78",
          9242 => x"8c",
          9243 => x"0b",
          9244 => x"22",
          9245 => x"80",
          9246 => x"74",
          9247 => x"38",
          9248 => x"56",
          9249 => x"17",
          9250 => x"57",
          9251 => x"2e",
          9252 => x"75",
          9253 => x"79",
          9254 => x"fe",
          9255 => x"82",
          9256 => x"10",
          9257 => x"82",
          9258 => x"9f",
          9259 => x"38",
          9260 => x"d8",
          9261 => x"82",
          9262 => x"05",
          9263 => x"2a",
          9264 => x"56",
          9265 => x"17",
          9266 => x"81",
          9267 => x"60",
          9268 => x"65",
          9269 => x"12",
          9270 => x"30",
          9271 => x"74",
          9272 => x"59",
          9273 => x"7d",
          9274 => x"81",
          9275 => x"76",
          9276 => x"41",
          9277 => x"76",
          9278 => x"90",
          9279 => x"62",
          9280 => x"51",
          9281 => x"26",
          9282 => x"75",
          9283 => x"31",
          9284 => x"65",
          9285 => x"fe",
          9286 => x"82",
          9287 => x"58",
          9288 => x"09",
          9289 => x"38",
          9290 => x"08",
          9291 => x"26",
          9292 => x"78",
          9293 => x"79",
          9294 => x"78",
          9295 => x"86",
          9296 => x"82",
          9297 => x"06",
          9298 => x"83",
          9299 => x"82",
          9300 => x"27",
          9301 => x"8f",
          9302 => x"55",
          9303 => x"26",
          9304 => x"59",
          9305 => x"62",
          9306 => x"74",
          9307 => x"38",
          9308 => x"88",
          9309 => x"c8",
          9310 => x"26",
          9311 => x"86",
          9312 => x"1a",
          9313 => x"79",
          9314 => x"38",
          9315 => x"80",
          9316 => x"2e",
          9317 => x"83",
          9318 => x"9f",
          9319 => x"8b",
          9320 => x"06",
          9321 => x"74",
          9322 => x"84",
          9323 => x"52",
          9324 => x"90",
          9325 => x"53",
          9326 => x"52",
          9327 => x"90",
          9328 => x"80",
          9329 => x"51",
          9330 => x"3f",
          9331 => x"34",
          9332 => x"ff",
          9333 => x"1b",
          9334 => x"d0",
          9335 => x"90",
          9336 => x"83",
          9337 => x"70",
          9338 => x"80",
          9339 => x"55",
          9340 => x"ff",
          9341 => x"66",
          9342 => x"ff",
          9343 => x"38",
          9344 => x"ff",
          9345 => x"1b",
          9346 => x"a0",
          9347 => x"74",
          9348 => x"51",
          9349 => x"3f",
          9350 => x"1c",
          9351 => x"98",
          9352 => x"8f",
          9353 => x"ff",
          9354 => x"51",
          9355 => x"3f",
          9356 => x"1b",
          9357 => x"92",
          9358 => x"2e",
          9359 => x"80",
          9360 => x"88",
          9361 => x"80",
          9362 => x"ff",
          9363 => x"7c",
          9364 => x"51",
          9365 => x"3f",
          9366 => x"1b",
          9367 => x"ea",
          9368 => x"b0",
          9369 => x"8e",
          9370 => x"52",
          9371 => x"ff",
          9372 => x"ff",
          9373 => x"c0",
          9374 => x"0b",
          9375 => x"34",
          9376 => x"ca",
          9377 => x"c7",
          9378 => x"39",
          9379 => x"0a",
          9380 => x"51",
          9381 => x"3f",
          9382 => x"ff",
          9383 => x"1b",
          9384 => x"88",
          9385 => x"0b",
          9386 => x"a9",
          9387 => x"34",
          9388 => x"ca",
          9389 => x"1b",
          9390 => x"bd",
          9391 => x"d5",
          9392 => x"1b",
          9393 => x"ff",
          9394 => x"81",
          9395 => x"7a",
          9396 => x"ff",
          9397 => x"81",
          9398 => x"c8",
          9399 => x"38",
          9400 => x"09",
          9401 => x"ee",
          9402 => x"60",
          9403 => x"7a",
          9404 => x"ff",
          9405 => x"84",
          9406 => x"52",
          9407 => x"8e",
          9408 => x"8b",
          9409 => x"52",
          9410 => x"8d",
          9411 => x"8a",
          9412 => x"52",
          9413 => x"51",
          9414 => x"3f",
          9415 => x"83",
          9416 => x"ff",
          9417 => x"82",
          9418 => x"1b",
          9419 => x"9a",
          9420 => x"d5",
          9421 => x"ff",
          9422 => x"75",
          9423 => x"05",
          9424 => x"7e",
          9425 => x"93",
          9426 => x"60",
          9427 => x"52",
          9428 => x"89",
          9429 => x"53",
          9430 => x"51",
          9431 => x"3f",
          9432 => x"58",
          9433 => x"09",
          9434 => x"38",
          9435 => x"51",
          9436 => x"3f",
          9437 => x"1b",
          9438 => x"ce",
          9439 => x"52",
          9440 => x"91",
          9441 => x"ff",
          9442 => x"81",
          9443 => x"f8",
          9444 => x"7a",
          9445 => x"b2",
          9446 => x"61",
          9447 => x"26",
          9448 => x"57",
          9449 => x"53",
          9450 => x"51",
          9451 => x"3f",
          9452 => x"08",
          9453 => x"84",
          9454 => x"d8",
          9455 => x"7a",
          9456 => x"d8",
          9457 => x"75",
          9458 => x"56",
          9459 => x"81",
          9460 => x"80",
          9461 => x"38",
          9462 => x"83",
          9463 => x"63",
          9464 => x"74",
          9465 => x"38",
          9466 => x"54",
          9467 => x"52",
          9468 => x"87",
          9469 => x"d8",
          9470 => x"c1",
          9471 => x"75",
          9472 => x"56",
          9473 => x"8c",
          9474 => x"2e",
          9475 => x"56",
          9476 => x"ff",
          9477 => x"84",
          9478 => x"2e",
          9479 => x"56",
          9480 => x"58",
          9481 => x"38",
          9482 => x"77",
          9483 => x"ff",
          9484 => x"82",
          9485 => x"78",
          9486 => x"f0",
          9487 => x"1b",
          9488 => x"34",
          9489 => x"16",
          9490 => x"82",
          9491 => x"83",
          9492 => x"84",
          9493 => x"67",
          9494 => x"fd",
          9495 => x"51",
          9496 => x"3f",
          9497 => x"16",
          9498 => x"c8",
          9499 => x"bf",
          9500 => x"86",
          9501 => x"d8",
          9502 => x"16",
          9503 => x"83",
          9504 => x"ff",
          9505 => x"66",
          9506 => x"1b",
          9507 => x"ba",
          9508 => x"77",
          9509 => x"7e",
          9510 => x"bf",
          9511 => x"82",
          9512 => x"a2",
          9513 => x"80",
          9514 => x"ff",
          9515 => x"81",
          9516 => x"c8",
          9517 => x"89",
          9518 => x"8a",
          9519 => x"86",
          9520 => x"c8",
          9521 => x"82",
          9522 => x"99",
          9523 => x"f5",
          9524 => x"60",
          9525 => x"79",
          9526 => x"5a",
          9527 => x"78",
          9528 => x"8d",
          9529 => x"55",
          9530 => x"fc",
          9531 => x"51",
          9532 => x"7a",
          9533 => x"81",
          9534 => x"8c",
          9535 => x"74",
          9536 => x"38",
          9537 => x"81",
          9538 => x"81",
          9539 => x"8a",
          9540 => x"06",
          9541 => x"76",
          9542 => x"76",
          9543 => x"55",
          9544 => x"c8",
          9545 => x"0d",
          9546 => x"0d",
          9547 => x"05",
          9548 => x"59",
          9549 => x"2e",
          9550 => x"87",
          9551 => x"76",
          9552 => x"84",
          9553 => x"80",
          9554 => x"38",
          9555 => x"77",
          9556 => x"56",
          9557 => x"34",
          9558 => x"bb",
          9559 => x"38",
          9560 => x"05",
          9561 => x"8c",
          9562 => x"08",
          9563 => x"3f",
          9564 => x"70",
          9565 => x"07",
          9566 => x"30",
          9567 => x"56",
          9568 => x"0c",
          9569 => x"18",
          9570 => x"0d",
          9571 => x"0d",
          9572 => x"08",
          9573 => x"75",
          9574 => x"89",
          9575 => x"54",
          9576 => x"16",
          9577 => x"51",
          9578 => x"82",
          9579 => x"91",
          9580 => x"08",
          9581 => x"81",
          9582 => x"88",
          9583 => x"83",
          9584 => x"74",
          9585 => x"0c",
          9586 => x"04",
          9587 => x"75",
          9588 => x"53",
          9589 => x"51",
          9590 => x"3f",
          9591 => x"85",
          9592 => x"ea",
          9593 => x"80",
          9594 => x"6a",
          9595 => x"70",
          9596 => x"d8",
          9597 => x"72",
          9598 => x"3f",
          9599 => x"8d",
          9600 => x"0d",
          9601 => x"0d",
          9602 => x"05",
          9603 => x"55",
          9604 => x"72",
          9605 => x"8a",
          9606 => x"ff",
          9607 => x"80",
          9608 => x"ff",
          9609 => x"51",
          9610 => x"2e",
          9611 => x"b4",
          9612 => x"2e",
          9613 => x"cc",
          9614 => x"72",
          9615 => x"38",
          9616 => x"83",
          9617 => x"53",
          9618 => x"ff",
          9619 => x"71",
          9620 => x"94",
          9621 => x"51",
          9622 => x"81",
          9623 => x"81",
          9624 => x"51",
          9625 => x"c8",
          9626 => x"0d",
          9627 => x"0d",
          9628 => x"22",
          9629 => x"96",
          9630 => x"51",
          9631 => x"80",
          9632 => x"38",
          9633 => x"39",
          9634 => x"2e",
          9635 => x"91",
          9636 => x"ff",
          9637 => x"70",
          9638 => x"94",
          9639 => x"54",
          9640 => x"d8",
          9641 => x"3d",
          9642 => x"3d",
          9643 => x"70",
          9644 => x"26",
          9645 => x"70",
          9646 => x"06",
          9647 => x"57",
          9648 => x"72",
          9649 => x"82",
          9650 => x"75",
          9651 => x"57",
          9652 => x"70",
          9653 => x"75",
          9654 => x"52",
          9655 => x"fb",
          9656 => x"82",
          9657 => x"70",
          9658 => x"81",
          9659 => x"18",
          9660 => x"53",
          9661 => x"80",
          9662 => x"88",
          9663 => x"38",
          9664 => x"82",
          9665 => x"51",
          9666 => x"71",
          9667 => x"76",
          9668 => x"54",
          9669 => x"c3",
          9670 => x"31",
          9671 => x"71",
          9672 => x"a4",
          9673 => x"51",
          9674 => x"12",
          9675 => x"d0",
          9676 => x"39",
          9677 => x"90",
          9678 => x"51",
          9679 => x"b0",
          9680 => x"39",
          9681 => x"51",
          9682 => x"ff",
          9683 => x"39",
          9684 => x"38",
          9685 => x"56",
          9686 => x"71",
          9687 => x"d8",
          9688 => x"3d",
          9689 => x"00",
          9690 => x"ff",
          9691 => x"ff",
          9692 => x"ff",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"00",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"00",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"00",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"00",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
          9825 => x"00",
          9826 => x"00",
          9827 => x"00",
          9828 => x"00",
          9829 => x"00",
          9830 => x"00",
          9831 => x"00",
          9832 => x"00",
          9833 => x"00",
          9834 => x"00",
          9835 => x"00",
          9836 => x"00",
          9837 => x"00",
          9838 => x"64",
          9839 => x"74",
          9840 => x"64",
          9841 => x"74",
          9842 => x"66",
          9843 => x"74",
          9844 => x"66",
          9845 => x"64",
          9846 => x"66",
          9847 => x"63",
          9848 => x"6d",
          9849 => x"61",
          9850 => x"6d",
          9851 => x"79",
          9852 => x"6d",
          9853 => x"66",
          9854 => x"6d",
          9855 => x"70",
          9856 => x"6d",
          9857 => x"6d",
          9858 => x"6d",
          9859 => x"68",
          9860 => x"68",
          9861 => x"68",
          9862 => x"68",
          9863 => x"63",
          9864 => x"00",
          9865 => x"6a",
          9866 => x"72",
          9867 => x"61",
          9868 => x"72",
          9869 => x"74",
          9870 => x"69",
          9871 => x"00",
          9872 => x"74",
          9873 => x"00",
          9874 => x"74",
          9875 => x"69",
          9876 => x"6d",
          9877 => x"69",
          9878 => x"6b",
          9879 => x"00",
          9880 => x"65",
          9881 => x"44",
          9882 => x"20",
          9883 => x"6f",
          9884 => x"49",
          9885 => x"72",
          9886 => x"20",
          9887 => x"6f",
          9888 => x"44",
          9889 => x"20",
          9890 => x"20",
          9891 => x"64",
          9892 => x"4e",
          9893 => x"69",
          9894 => x"66",
          9895 => x"64",
          9896 => x"4e",
          9897 => x"61",
          9898 => x"66",
          9899 => x"64",
          9900 => x"49",
          9901 => x"6c",
          9902 => x"66",
          9903 => x"6e",
          9904 => x"2e",
          9905 => x"41",
          9906 => x"73",
          9907 => x"65",
          9908 => x"64",
          9909 => x"46",
          9910 => x"20",
          9911 => x"65",
          9912 => x"20",
          9913 => x"73",
          9914 => x"00",
          9915 => x"46",
          9916 => x"20",
          9917 => x"64",
          9918 => x"69",
          9919 => x"6c",
          9920 => x"00",
          9921 => x"53",
          9922 => x"73",
          9923 => x"69",
          9924 => x"70",
          9925 => x"65",
          9926 => x"64",
          9927 => x"44",
          9928 => x"65",
          9929 => x"6d",
          9930 => x"20",
          9931 => x"69",
          9932 => x"6c",
          9933 => x"00",
          9934 => x"44",
          9935 => x"20",
          9936 => x"20",
          9937 => x"62",
          9938 => x"2e",
          9939 => x"4e",
          9940 => x"6f",
          9941 => x"74",
          9942 => x"65",
          9943 => x"6c",
          9944 => x"73",
          9945 => x"20",
          9946 => x"6e",
          9947 => x"6e",
          9948 => x"73",
          9949 => x"46",
          9950 => x"61",
          9951 => x"62",
          9952 => x"65",
          9953 => x"54",
          9954 => x"6f",
          9955 => x"20",
          9956 => x"72",
          9957 => x"6f",
          9958 => x"61",
          9959 => x"6c",
          9960 => x"2e",
          9961 => x"46",
          9962 => x"20",
          9963 => x"6c",
          9964 => x"65",
          9965 => x"49",
          9966 => x"66",
          9967 => x"69",
          9968 => x"20",
          9969 => x"6f",
          9970 => x"00",
          9971 => x"54",
          9972 => x"6d",
          9973 => x"20",
          9974 => x"6e",
          9975 => x"6c",
          9976 => x"00",
          9977 => x"50",
          9978 => x"6d",
          9979 => x"72",
          9980 => x"6e",
          9981 => x"72",
          9982 => x"2e",
          9983 => x"53",
          9984 => x"65",
          9985 => x"00",
          9986 => x"55",
          9987 => x"6f",
          9988 => x"65",
          9989 => x"72",
          9990 => x"0a",
          9991 => x"20",
          9992 => x"65",
          9993 => x"73",
          9994 => x"20",
          9995 => x"20",
          9996 => x"65",
          9997 => x"65",
          9998 => x"00",
          9999 => x"72",
         10000 => x"00",
         10001 => x"30",
         10002 => x"38",
         10003 => x"20",
         10004 => x"30",
         10005 => x"2c",
         10006 => x"25",
         10007 => x"78",
         10008 => x"49",
         10009 => x"25",
         10010 => x"78",
         10011 => x"38",
         10012 => x"25",
         10013 => x"78",
         10014 => x"25",
         10015 => x"58",
         10016 => x"3a",
         10017 => x"25",
         10018 => x"00",
         10019 => x"20",
         10020 => x"20",
         10021 => x"00",
         10022 => x"25",
         10023 => x"00",
         10024 => x"20",
         10025 => x"20",
         10026 => x"7c",
         10027 => x"5a",
         10028 => x"41",
         10029 => x"0a",
         10030 => x"25",
         10031 => x"00",
         10032 => x"30",
         10033 => x"35",
         10034 => x"32",
         10035 => x"76",
         10036 => x"32",
         10037 => x"20",
         10038 => x"2c",
         10039 => x"76",
         10040 => x"32",
         10041 => x"25",
         10042 => x"73",
         10043 => x"0a",
         10044 => x"5a",
         10045 => x"41",
         10046 => x"74",
         10047 => x"75",
         10048 => x"48",
         10049 => x"6c",
         10050 => x"54",
         10051 => x"72",
         10052 => x"74",
         10053 => x"75",
         10054 => x"50",
         10055 => x"69",
         10056 => x"72",
         10057 => x"74",
         10058 => x"49",
         10059 => x"4c",
         10060 => x"20",
         10061 => x"65",
         10062 => x"70",
         10063 => x"49",
         10064 => x"4c",
         10065 => x"20",
         10066 => x"65",
         10067 => x"70",
         10068 => x"55",
         10069 => x"30",
         10070 => x"20",
         10071 => x"65",
         10072 => x"70",
         10073 => x"55",
         10074 => x"30",
         10075 => x"20",
         10076 => x"65",
         10077 => x"70",
         10078 => x"55",
         10079 => x"31",
         10080 => x"20",
         10081 => x"65",
         10082 => x"70",
         10083 => x"55",
         10084 => x"31",
         10085 => x"20",
         10086 => x"65",
         10087 => x"70",
         10088 => x"53",
         10089 => x"69",
         10090 => x"75",
         10091 => x"69",
         10092 => x"2e",
         10093 => x"45",
         10094 => x"6c",
         10095 => x"20",
         10096 => x"65",
         10097 => x"2e",
         10098 => x"61",
         10099 => x"65",
         10100 => x"2e",
         10101 => x"00",
         10102 => x"7a",
         10103 => x"61",
         10104 => x"74",
         10105 => x"30",
         10106 => x"46",
         10107 => x"65",
         10108 => x"6f",
         10109 => x"69",
         10110 => x"6c",
         10111 => x"20",
         10112 => x"63",
         10113 => x"20",
         10114 => x"70",
         10115 => x"73",
         10116 => x"6e",
         10117 => x"6d",
         10118 => x"61",
         10119 => x"2e",
         10120 => x"2a",
         10121 => x"42",
         10122 => x"64",
         10123 => x"20",
         10124 => x"00",
         10125 => x"49",
         10126 => x"69",
         10127 => x"73",
         10128 => x"00",
         10129 => x"46",
         10130 => x"65",
         10131 => x"6f",
         10132 => x"69",
         10133 => x"6c",
         10134 => x"2e",
         10135 => x"72",
         10136 => x"64",
         10137 => x"25",
         10138 => x"43",
         10139 => x"72",
         10140 => x"2e",
         10141 => x"00",
         10142 => x"43",
         10143 => x"69",
         10144 => x"2e",
         10145 => x"43",
         10146 => x"61",
         10147 => x"67",
         10148 => x"00",
         10149 => x"25",
         10150 => x"78",
         10151 => x"38",
         10152 => x"3e",
         10153 => x"6c",
         10154 => x"30",
         10155 => x"0a",
         10156 => x"44",
         10157 => x"20",
         10158 => x"6f",
         10159 => x"0a",
         10160 => x"70",
         10161 => x"65",
         10162 => x"25",
         10163 => x"58",
         10164 => x"32",
         10165 => x"3f",
         10166 => x"25",
         10167 => x"58",
         10168 => x"34",
         10169 => x"25",
         10170 => x"58",
         10171 => x"38",
         10172 => x"00",
         10173 => x"44",
         10174 => x"62",
         10175 => x"67",
         10176 => x"74",
         10177 => x"75",
         10178 => x"00",
         10179 => x"45",
         10180 => x"6c",
         10181 => x"20",
         10182 => x"65",
         10183 => x"70",
         10184 => x"44",
         10185 => x"62",
         10186 => x"20",
         10187 => x"74",
         10188 => x"66",
         10189 => x"45",
         10190 => x"6c",
         10191 => x"20",
         10192 => x"74",
         10193 => x"66",
         10194 => x"45",
         10195 => x"75",
         10196 => x"67",
         10197 => x"64",
         10198 => x"20",
         10199 => x"6c",
         10200 => x"2e",
         10201 => x"43",
         10202 => x"69",
         10203 => x"63",
         10204 => x"20",
         10205 => x"30",
         10206 => x"20",
         10207 => x"0a",
         10208 => x"43",
         10209 => x"20",
         10210 => x"75",
         10211 => x"64",
         10212 => x"64",
         10213 => x"25",
         10214 => x"0a",
         10215 => x"52",
         10216 => x"61",
         10217 => x"6e",
         10218 => x"70",
         10219 => x"63",
         10220 => x"6f",
         10221 => x"2e",
         10222 => x"43",
         10223 => x"20",
         10224 => x"6f",
         10225 => x"6e",
         10226 => x"2e",
         10227 => x"5a",
         10228 => x"62",
         10229 => x"25",
         10230 => x"25",
         10231 => x"73",
         10232 => x"00",
         10233 => x"25",
         10234 => x"25",
         10235 => x"73",
         10236 => x"25",
         10237 => x"25",
         10238 => x"42",
         10239 => x"63",
         10240 => x"61",
         10241 => x"00",
         10242 => x"52",
         10243 => x"69",
         10244 => x"2e",
         10245 => x"45",
         10246 => x"6c",
         10247 => x"20",
         10248 => x"65",
         10249 => x"70",
         10250 => x"2e",
         10251 => x"25",
         10252 => x"64",
         10253 => x"20",
         10254 => x"25",
         10255 => x"64",
         10256 => x"25",
         10257 => x"53",
         10258 => x"43",
         10259 => x"69",
         10260 => x"61",
         10261 => x"6e",
         10262 => x"20",
         10263 => x"6f",
         10264 => x"6f",
         10265 => x"6f",
         10266 => x"67",
         10267 => x"3a",
         10268 => x"76",
         10269 => x"73",
         10270 => x"70",
         10271 => x"65",
         10272 => x"64",
         10273 => x"20",
         10274 => x"57",
         10275 => x"44",
         10276 => x"20",
         10277 => x"30",
         10278 => x"25",
         10279 => x"29",
         10280 => x"20",
         10281 => x"53",
         10282 => x"4d",
         10283 => x"20",
         10284 => x"30",
         10285 => x"25",
         10286 => x"29",
         10287 => x"20",
         10288 => x"49",
         10289 => x"20",
         10290 => x"4d",
         10291 => x"30",
         10292 => x"25",
         10293 => x"29",
         10294 => x"20",
         10295 => x"42",
         10296 => x"20",
         10297 => x"20",
         10298 => x"30",
         10299 => x"25",
         10300 => x"29",
         10301 => x"20",
         10302 => x"52",
         10303 => x"20",
         10304 => x"20",
         10305 => x"30",
         10306 => x"25",
         10307 => x"29",
         10308 => x"20",
         10309 => x"53",
         10310 => x"41",
         10311 => x"20",
         10312 => x"65",
         10313 => x"65",
         10314 => x"25",
         10315 => x"29",
         10316 => x"20",
         10317 => x"54",
         10318 => x"52",
         10319 => x"20",
         10320 => x"69",
         10321 => x"73",
         10322 => x"25",
         10323 => x"29",
         10324 => x"20",
         10325 => x"49",
         10326 => x"20",
         10327 => x"4c",
         10328 => x"68",
         10329 => x"65",
         10330 => x"25",
         10331 => x"29",
         10332 => x"20",
         10333 => x"57",
         10334 => x"42",
         10335 => x"20",
         10336 => x"00",
         10337 => x"20",
         10338 => x"57",
         10339 => x"32",
         10340 => x"20",
         10341 => x"49",
         10342 => x"4c",
         10343 => x"20",
         10344 => x"50",
         10345 => x"20",
         10346 => x"53",
         10347 => x"41",
         10348 => x"65",
         10349 => x"73",
         10350 => x"20",
         10351 => x"43",
         10352 => x"52",
         10353 => x"74",
         10354 => x"63",
         10355 => x"20",
         10356 => x"72",
         10357 => x"20",
         10358 => x"30",
         10359 => x"00",
         10360 => x"20",
         10361 => x"43",
         10362 => x"4d",
         10363 => x"72",
         10364 => x"74",
         10365 => x"20",
         10366 => x"72",
         10367 => x"20",
         10368 => x"30",
         10369 => x"00",
         10370 => x"20",
         10371 => x"53",
         10372 => x"6b",
         10373 => x"61",
         10374 => x"41",
         10375 => x"65",
         10376 => x"20",
         10377 => x"20",
         10378 => x"30",
         10379 => x"00",
         10380 => x"4d",
         10381 => x"3a",
         10382 => x"20",
         10383 => x"5a",
         10384 => x"49",
         10385 => x"20",
         10386 => x"20",
         10387 => x"20",
         10388 => x"20",
         10389 => x"20",
         10390 => x"30",
         10391 => x"00",
         10392 => x"20",
         10393 => x"53",
         10394 => x"65",
         10395 => x"6c",
         10396 => x"20",
         10397 => x"71",
         10398 => x"20",
         10399 => x"20",
         10400 => x"64",
         10401 => x"34",
         10402 => x"7a",
         10403 => x"20",
         10404 => x"53",
         10405 => x"4d",
         10406 => x"6f",
         10407 => x"46",
         10408 => x"20",
         10409 => x"20",
         10410 => x"20",
         10411 => x"64",
         10412 => x"34",
         10413 => x"7a",
         10414 => x"20",
         10415 => x"57",
         10416 => x"62",
         10417 => x"20",
         10418 => x"41",
         10419 => x"6c",
         10420 => x"20",
         10421 => x"71",
         10422 => x"64",
         10423 => x"34",
         10424 => x"7a",
         10425 => x"53",
         10426 => x"6c",
         10427 => x"4d",
         10428 => x"75",
         10429 => x"46",
         10430 => x"00",
         10431 => x"45",
         10432 => x"45",
         10433 => x"00",
         10434 => x"55",
         10435 => x"6f",
         10436 => x"00",
         10437 => x"01",
         10438 => x"00",
         10439 => x"00",
         10440 => x"01",
         10441 => x"00",
         10442 => x"00",
         10443 => x"01",
         10444 => x"00",
         10445 => x"00",
         10446 => x"01",
         10447 => x"00",
         10448 => x"00",
         10449 => x"01",
         10450 => x"00",
         10451 => x"00",
         10452 => x"01",
         10453 => x"00",
         10454 => x"00",
         10455 => x"01",
         10456 => x"00",
         10457 => x"00",
         10458 => x"01",
         10459 => x"00",
         10460 => x"00",
         10461 => x"01",
         10462 => x"00",
         10463 => x"00",
         10464 => x"01",
         10465 => x"00",
         10466 => x"00",
         10467 => x"01",
         10468 => x"00",
         10469 => x"00",
         10470 => x"04",
         10471 => x"00",
         10472 => x"00",
         10473 => x"04",
         10474 => x"00",
         10475 => x"00",
         10476 => x"04",
         10477 => x"00",
         10478 => x"00",
         10479 => x"03",
         10480 => x"00",
         10481 => x"00",
         10482 => x"04",
         10483 => x"00",
         10484 => x"00",
         10485 => x"04",
         10486 => x"00",
         10487 => x"00",
         10488 => x"04",
         10489 => x"00",
         10490 => x"00",
         10491 => x"03",
         10492 => x"00",
         10493 => x"00",
         10494 => x"03",
         10495 => x"00",
         10496 => x"00",
         10497 => x"03",
         10498 => x"00",
         10499 => x"00",
         10500 => x"03",
         10501 => x"00",
         10502 => x"1b",
         10503 => x"1b",
         10504 => x"1b",
         10505 => x"1b",
         10506 => x"1b",
         10507 => x"1b",
         10508 => x"1b",
         10509 => x"1b",
         10510 => x"1b",
         10511 => x"1b",
         10512 => x"1b",
         10513 => x"10",
         10514 => x"0e",
         10515 => x"0d",
         10516 => x"0b",
         10517 => x"08",
         10518 => x"06",
         10519 => x"05",
         10520 => x"04",
         10521 => x"03",
         10522 => x"02",
         10523 => x"01",
         10524 => x"68",
         10525 => x"6f",
         10526 => x"68",
         10527 => x"00",
         10528 => x"21",
         10529 => x"25",
         10530 => x"75",
         10531 => x"73",
         10532 => x"46",
         10533 => x"65",
         10534 => x"6f",
         10535 => x"73",
         10536 => x"74",
         10537 => x"68",
         10538 => x"6f",
         10539 => x"66",
         10540 => x"20",
         10541 => x"45",
         10542 => x"00",
         10543 => x"43",
         10544 => x"6f",
         10545 => x"70",
         10546 => x"63",
         10547 => x"74",
         10548 => x"69",
         10549 => x"72",
         10550 => x"69",
         10551 => x"20",
         10552 => x"61",
         10553 => x"6e",
         10554 => x"53",
         10555 => x"22",
         10556 => x"3e",
         10557 => x"00",
         10558 => x"2b",
         10559 => x"5b",
         10560 => x"46",
         10561 => x"46",
         10562 => x"32",
         10563 => x"eb",
         10564 => x"53",
         10565 => x"35",
         10566 => x"4e",
         10567 => x"41",
         10568 => x"20",
         10569 => x"41",
         10570 => x"20",
         10571 => x"4e",
         10572 => x"41",
         10573 => x"20",
         10574 => x"41",
         10575 => x"20",
         10576 => x"00",
         10577 => x"00",
         10578 => x"00",
         10579 => x"00",
         10580 => x"01",
         10581 => x"09",
         10582 => x"14",
         10583 => x"1e",
         10584 => x"80",
         10585 => x"8e",
         10586 => x"45",
         10587 => x"49",
         10588 => x"90",
         10589 => x"99",
         10590 => x"59",
         10591 => x"9c",
         10592 => x"41",
         10593 => x"a5",
         10594 => x"a8",
         10595 => x"ac",
         10596 => x"b0",
         10597 => x"b4",
         10598 => x"b8",
         10599 => x"bc",
         10600 => x"c0",
         10601 => x"c4",
         10602 => x"c8",
         10603 => x"cc",
         10604 => x"d0",
         10605 => x"d4",
         10606 => x"d8",
         10607 => x"dc",
         10608 => x"e0",
         10609 => x"e4",
         10610 => x"e8",
         10611 => x"ec",
         10612 => x"f0",
         10613 => x"f4",
         10614 => x"f8",
         10615 => x"fc",
         10616 => x"2b",
         10617 => x"3d",
         10618 => x"5c",
         10619 => x"3c",
         10620 => x"7f",
         10621 => x"00",
         10622 => x"00",
         10623 => x"01",
         10624 => x"00",
         10625 => x"00",
         10626 => x"00",
         10627 => x"00",
         10628 => x"00",
         10629 => x"00",
         10630 => x"00",
         10631 => x"00",
         10632 => x"00",
         10633 => x"00",
         10634 => x"00",
         10635 => x"00",
         10636 => x"00",
         10637 => x"00",
         10638 => x"00",
         10639 => x"00",
         10640 => x"00",
         10641 => x"00",
         10642 => x"00",
         10643 => x"00",
         10644 => x"20",
         10645 => x"00",
         10646 => x"00",
         10647 => x"00",
         10648 => x"00",
         10649 => x"00",
         10650 => x"00",
         10651 => x"00",
         10652 => x"00",
         10653 => x"25",
         10654 => x"25",
         10655 => x"25",
         10656 => x"25",
         10657 => x"25",
         10658 => x"25",
         10659 => x"25",
         10660 => x"25",
         10661 => x"25",
         10662 => x"25",
         10663 => x"25",
         10664 => x"25",
         10665 => x"25",
         10666 => x"25",
         10667 => x"25",
         10668 => x"25",
         10669 => x"25",
         10670 => x"25",
         10671 => x"25",
         10672 => x"25",
         10673 => x"25",
         10674 => x"25",
         10675 => x"25",
         10676 => x"25",
         10677 => x"03",
         10678 => x"03",
         10679 => x"03",
         10680 => x"00",
         10681 => x"03",
         10682 => x"03",
         10683 => x"22",
         10684 => x"03",
         10685 => x"22",
         10686 => x"22",
         10687 => x"23",
         10688 => x"00",
         10689 => x"00",
         10690 => x"00",
         10691 => x"20",
         10692 => x"25",
         10693 => x"00",
         10694 => x"00",
         10695 => x"00",
         10696 => x"00",
         10697 => x"01",
         10698 => x"01",
         10699 => x"01",
         10700 => x"01",
         10701 => x"01",
         10702 => x"01",
         10703 => x"00",
         10704 => x"01",
         10705 => x"01",
         10706 => x"01",
         10707 => x"01",
         10708 => x"01",
         10709 => x"01",
         10710 => x"01",
         10711 => x"01",
         10712 => x"01",
         10713 => x"01",
         10714 => x"01",
         10715 => x"01",
         10716 => x"01",
         10717 => x"01",
         10718 => x"01",
         10719 => x"01",
         10720 => x"01",
         10721 => x"01",
         10722 => x"01",
         10723 => x"01",
         10724 => x"01",
         10725 => x"01",
         10726 => x"01",
         10727 => x"01",
         10728 => x"01",
         10729 => x"01",
         10730 => x"01",
         10731 => x"01",
         10732 => x"01",
         10733 => x"01",
         10734 => x"01",
         10735 => x"01",
         10736 => x"01",
         10737 => x"01",
         10738 => x"01",
         10739 => x"01",
         10740 => x"01",
         10741 => x"01",
         10742 => x"01",
         10743 => x"01",
         10744 => x"01",
         10745 => x"01",
         10746 => x"00",
         10747 => x"01",
         10748 => x"01",
         10749 => x"02",
         10750 => x"02",
         10751 => x"2c",
         10752 => x"02",
         10753 => x"2c",
         10754 => x"02",
         10755 => x"02",
         10756 => x"01",
         10757 => x"00",
         10758 => x"01",
         10759 => x"01",
         10760 => x"02",
         10761 => x"02",
         10762 => x"02",
         10763 => x"02",
         10764 => x"01",
         10765 => x"02",
         10766 => x"02",
         10767 => x"02",
         10768 => x"01",
         10769 => x"02",
         10770 => x"02",
         10771 => x"02",
         10772 => x"02",
         10773 => x"01",
         10774 => x"02",
         10775 => x"02",
         10776 => x"02",
         10777 => x"02",
         10778 => x"02",
         10779 => x"02",
         10780 => x"01",
         10781 => x"02",
         10782 => x"02",
         10783 => x"02",
         10784 => x"01",
         10785 => x"01",
         10786 => x"02",
         10787 => x"02",
         10788 => x"02",
         10789 => x"01",
         10790 => x"00",
         10791 => x"03",
         10792 => x"03",
         10793 => x"03",
         10794 => x"03",
         10795 => x"03",
         10796 => x"03",
         10797 => x"03",
         10798 => x"03",
         10799 => x"03",
         10800 => x"03",
         10801 => x"03",
         10802 => x"01",
         10803 => x"00",
         10804 => x"03",
         10805 => x"03",
         10806 => x"03",
         10807 => x"03",
         10808 => x"03",
         10809 => x"03",
         10810 => x"07",
         10811 => x"01",
         10812 => x"01",
         10813 => x"01",
         10814 => x"00",
         10815 => x"04",
         10816 => x"05",
         10817 => x"00",
         10818 => x"1d",
         10819 => x"2c",
         10820 => x"01",
         10821 => x"01",
         10822 => x"06",
         10823 => x"06",
         10824 => x"06",
         10825 => x"06",
         10826 => x"06",
         10827 => x"00",
         10828 => x"1f",
         10829 => x"1f",
         10830 => x"1f",
         10831 => x"1f",
         10832 => x"1f",
         10833 => x"1f",
         10834 => x"1f",
         10835 => x"1f",
         10836 => x"1f",
         10837 => x"1f",
         10838 => x"1f",
         10839 => x"1f",
         10840 => x"1f",
         10841 => x"1f",
         10842 => x"1f",
         10843 => x"1f",
         10844 => x"1f",
         10845 => x"1f",
         10846 => x"1f",
         10847 => x"1f",
         10848 => x"06",
         10849 => x"06",
         10850 => x"00",
         10851 => x"1f",
         10852 => x"1f",
         10853 => x"00",
         10854 => x"21",
         10855 => x"21",
         10856 => x"21",
         10857 => x"05",
         10858 => x"04",
         10859 => x"01",
         10860 => x"01",
         10861 => x"01",
         10862 => x"01",
         10863 => x"08",
         10864 => x"03",
         10865 => x"00",
         10866 => x"00",
         10867 => x"01",
         10868 => x"00",
         10869 => x"00",
         10870 => x"00",
         10871 => x"01",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"01",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"01",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"01",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"01",
         10888 => x"00",
         10889 => x"00",
         10890 => x"00",
         10891 => x"01",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"01",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"01",
         10900 => x"00",
         10901 => x"00",
         10902 => x"00",
         10903 => x"01",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"01",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"01",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"01",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"01",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"01",
         10924 => x"00",
         10925 => x"00",
         10926 => x"00",
         10927 => x"01",
         10928 => x"00",
         10929 => x"00",
         10930 => x"00",
         10931 => x"01",
         10932 => x"00",
         10933 => x"00",
         10934 => x"00",
         10935 => x"01",
         10936 => x"00",
         10937 => x"00",
         10938 => x"00",
         10939 => x"01",
         10940 => x"00",
         10941 => x"00",
         10942 => x"00",
         10943 => x"01",
         10944 => x"00",
         10945 => x"00",
         10946 => x"00",
         10947 => x"01",
         10948 => x"00",
         10949 => x"00",
         10950 => x"00",
         10951 => x"01",
         10952 => x"00",
         10953 => x"00",
         10954 => x"00",
         10955 => x"01",
         10956 => x"00",
         10957 => x"00",
         10958 => x"00",
         10959 => x"01",
         10960 => x"00",
         10961 => x"00",
         10962 => x"00",
         10963 => x"01",
         10964 => x"00",
         10965 => x"00",
         10966 => x"00",
         10967 => x"01",
         10968 => x"00",
         10969 => x"00",
         10970 => x"00",
         10971 => x"00",
         10972 => x"00",
         10973 => x"00",
         10974 => x"00",
         10975 => x"00",
         10976 => x"00",
         10977 => x"00",
         10978 => x"00",
         10979 => x"01",
         10980 => x"01",
         10981 => x"00",
         10982 => x"00",
         10983 => x"00",
         10984 => x"00",
         10985 => x"05",
         10986 => x"05",
         10987 => x"05",
         10988 => x"00",
         10989 => x"01",
         10990 => x"01",
         10991 => x"01",
         10992 => x"01",
         10993 => x"00",
         10994 => x"00",
         10995 => x"00",
         10996 => x"00",
         10997 => x"00",
         10998 => x"00",
         10999 => x"00",
         11000 => x"00",
         11001 => x"00",
         11002 => x"00",
         11003 => x"00",
         11004 => x"00",
         11005 => x"00",
         11006 => x"00",
         11007 => x"00",
         11008 => x"00",
         11009 => x"00",
         11010 => x"00",
         11011 => x"00",
         11012 => x"00",
         11013 => x"00",
         11014 => x"00",
         11015 => x"00",
         11016 => x"00",
         11017 => x"00",
         11018 => x"01",
         11019 => x"00",
         11020 => x"01",
         11021 => x"00",
         11022 => x"02",
         11023 => x"00",
         11024 => x"00",
         11025 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
