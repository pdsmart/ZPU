-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPort32-64BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPort32-64BootBRAM;

architecture arch of DualPort32-64BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"80",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"ad",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"c5",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"c7",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8e",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"8f",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"90",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"91",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"92",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"f0",
           386 => x"c0",
           387 => x"f0",
           388 => x"90",
           389 => x"f0",
           390 => x"2d",
           391 => x"08",
           392 => x"04",
           393 => x"0c",
           394 => x"82",
           395 => x"84",
           396 => x"82",
           397 => x"af",
           398 => x"d5",
           399 => x"80",
           400 => x"d5",
           401 => x"ad",
           402 => x"f0",
           403 => x"90",
           404 => x"f0",
           405 => x"2d",
           406 => x"08",
           407 => x"04",
           408 => x"0c",
           409 => x"2d",
           410 => x"08",
           411 => x"04",
           412 => x"0c",
           413 => x"2d",
           414 => x"08",
           415 => x"04",
           416 => x"0c",
           417 => x"82",
           418 => x"84",
           419 => x"82",
           420 => x"96",
           421 => x"d5",
           422 => x"80",
           423 => x"d5",
           424 => x"cd",
           425 => x"f0",
           426 => x"90",
           427 => x"f0",
           428 => x"ea",
           429 => x"f0",
           430 => x"90",
           431 => x"f0",
           432 => x"c8",
           433 => x"f0",
           434 => x"90",
           435 => x"f0",
           436 => x"85",
           437 => x"f0",
           438 => x"90",
           439 => x"f0",
           440 => x"fc",
           441 => x"f0",
           442 => x"90",
           443 => x"f0",
           444 => x"af",
           445 => x"f0",
           446 => x"90",
           447 => x"f0",
           448 => x"d7",
           449 => x"f0",
           450 => x"90",
           451 => x"f0",
           452 => x"d7",
           453 => x"f0",
           454 => x"90",
           455 => x"f0",
           456 => x"bc",
           457 => x"f0",
           458 => x"90",
           459 => x"f0",
           460 => x"bc",
           461 => x"f0",
           462 => x"90",
           463 => x"f0",
           464 => x"95",
           465 => x"f0",
           466 => x"90",
           467 => x"f0",
           468 => x"fe",
           469 => x"f0",
           470 => x"90",
           471 => x"f0",
           472 => x"b4",
           473 => x"f0",
           474 => x"90",
           475 => x"f0",
           476 => x"b8",
           477 => x"f0",
           478 => x"90",
           479 => x"f0",
           480 => x"d8",
           481 => x"f0",
           482 => x"90",
           483 => x"f0",
           484 => x"f7",
           485 => x"f0",
           486 => x"90",
           487 => x"f0",
           488 => x"eb",
           489 => x"f0",
           490 => x"90",
           491 => x"f0",
           492 => x"cd",
           493 => x"f0",
           494 => x"90",
           495 => x"f0",
           496 => x"c7",
           497 => x"f0",
           498 => x"90",
           499 => x"f0",
           500 => x"fd",
           501 => x"f0",
           502 => x"90",
           503 => x"f0",
           504 => x"cc",
           505 => x"f0",
           506 => x"90",
           507 => x"f0",
           508 => x"cd",
           509 => x"f0",
           510 => x"90",
           511 => x"f0",
           512 => x"b7",
           513 => x"f0",
           514 => x"90",
           515 => x"f0",
           516 => x"90",
           517 => x"f0",
           518 => x"90",
           519 => x"f0",
           520 => x"bb",
           521 => x"f0",
           522 => x"90",
           523 => x"f0",
           524 => x"d4",
           525 => x"f0",
           526 => x"90",
           527 => x"f0",
           528 => x"be",
           529 => x"f0",
           530 => x"90",
           531 => x"f0",
           532 => x"c9",
           533 => x"f0",
           534 => x"90",
           535 => x"f0",
           536 => x"d0",
           537 => x"f0",
           538 => x"90",
           539 => x"f0",
           540 => x"f6",
           541 => x"f0",
           542 => x"90",
           543 => x"f0",
           544 => x"bc",
           545 => x"f0",
           546 => x"90",
           547 => x"f0",
           548 => x"99",
           549 => x"f0",
           550 => x"90",
           551 => x"f0",
           552 => x"85",
           553 => x"f0",
           554 => x"90",
           555 => x"f0",
           556 => x"bb",
           557 => x"f0",
           558 => x"90",
           559 => x"f0",
           560 => x"a5",
           561 => x"f0",
           562 => x"90",
           563 => x"f0",
           564 => x"89",
           565 => x"f0",
           566 => x"90",
           567 => x"f0",
           568 => x"ae",
           569 => x"f0",
           570 => x"90",
           571 => x"f0",
           572 => x"d2",
           573 => x"f0",
           574 => x"90",
           575 => x"f0",
           576 => x"b5",
           577 => x"f0",
           578 => x"90",
           579 => x"f0",
           580 => x"bf",
           581 => x"f0",
           582 => x"90",
           583 => x"f0",
           584 => x"cf",
           585 => x"f0",
           586 => x"90",
           587 => x"f0",
           588 => x"f7",
           589 => x"f0",
           590 => x"90",
           591 => x"f0",
           592 => x"ef",
           593 => x"f0",
           594 => x"90",
           595 => x"f0",
           596 => x"b9",
           597 => x"f0",
           598 => x"90",
           599 => x"00",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"00",
           609 => x"ff",
           610 => x"06",
           611 => x"83",
           612 => x"10",
           613 => x"fc",
           614 => x"51",
           615 => x"80",
           616 => x"ff",
           617 => x"06",
           618 => x"52",
           619 => x"0a",
           620 => x"38",
           621 => x"51",
           622 => x"e4",
           623 => x"d0",
           624 => x"80",
           625 => x"05",
           626 => x"0b",
           627 => x"04",
           628 => x"80",
           629 => x"00",
           630 => x"08",
           631 => x"f0",
           632 => x"0d",
           633 => x"08",
           634 => x"82",
           635 => x"fc",
           636 => x"d5",
           637 => x"05",
           638 => x"d5",
           639 => x"05",
           640 => x"f1",
           641 => x"54",
           642 => x"82",
           643 => x"70",
           644 => x"08",
           645 => x"82",
           646 => x"f8",
           647 => x"82",
           648 => x"51",
           649 => x"0d",
           650 => x"0c",
           651 => x"f0",
           652 => x"d5",
           653 => x"3d",
           654 => x"f0",
           655 => x"08",
           656 => x"70",
           657 => x"81",
           658 => x"51",
           659 => x"38",
           660 => x"d5",
           661 => x"05",
           662 => x"38",
           663 => x"0b",
           664 => x"08",
           665 => x"81",
           666 => x"d5",
           667 => x"05",
           668 => x"82",
           669 => x"8c",
           670 => x"0b",
           671 => x"08",
           672 => x"82",
           673 => x"88",
           674 => x"d5",
           675 => x"05",
           676 => x"f0",
           677 => x"08",
           678 => x"f6",
           679 => x"82",
           680 => x"8c",
           681 => x"80",
           682 => x"d5",
           683 => x"05",
           684 => x"90",
           685 => x"e4",
           686 => x"d5",
           687 => x"05",
           688 => x"d5",
           689 => x"05",
           690 => x"09",
           691 => x"38",
           692 => x"d5",
           693 => x"05",
           694 => x"39",
           695 => x"08",
           696 => x"82",
           697 => x"f8",
           698 => x"53",
           699 => x"82",
           700 => x"8c",
           701 => x"05",
           702 => x"08",
           703 => x"82",
           704 => x"fc",
           705 => x"05",
           706 => x"08",
           707 => x"ff",
           708 => x"d5",
           709 => x"05",
           710 => x"72",
           711 => x"f0",
           712 => x"08",
           713 => x"f0",
           714 => x"0c",
           715 => x"f0",
           716 => x"08",
           717 => x"0c",
           718 => x"82",
           719 => x"04",
           720 => x"08",
           721 => x"f0",
           722 => x"0d",
           723 => x"d5",
           724 => x"05",
           725 => x"f0",
           726 => x"08",
           727 => x"08",
           728 => x"fe",
           729 => x"d5",
           730 => x"05",
           731 => x"f0",
           732 => x"70",
           733 => x"08",
           734 => x"82",
           735 => x"fc",
           736 => x"82",
           737 => x"8c",
           738 => x"82",
           739 => x"e0",
           740 => x"51",
           741 => x"3f",
           742 => x"08",
           743 => x"f0",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"88",
           748 => x"51",
           749 => x"34",
           750 => x"08",
           751 => x"70",
           752 => x"0c",
           753 => x"0d",
           754 => x"0c",
           755 => x"f0",
           756 => x"d5",
           757 => x"3d",
           758 => x"f0",
           759 => x"70",
           760 => x"08",
           761 => x"82",
           762 => x"fc",
           763 => x"82",
           764 => x"8c",
           765 => x"82",
           766 => x"88",
           767 => x"54",
           768 => x"d5",
           769 => x"82",
           770 => x"f8",
           771 => x"d5",
           772 => x"05",
           773 => x"d5",
           774 => x"54",
           775 => x"82",
           776 => x"04",
           777 => x"08",
           778 => x"f0",
           779 => x"0d",
           780 => x"d5",
           781 => x"05",
           782 => x"f0",
           783 => x"08",
           784 => x"8c",
           785 => x"d5",
           786 => x"05",
           787 => x"33",
           788 => x"70",
           789 => x"81",
           790 => x"51",
           791 => x"80",
           792 => x"ff",
           793 => x"f0",
           794 => x"0c",
           795 => x"82",
           796 => x"8c",
           797 => x"72",
           798 => x"82",
           799 => x"f8",
           800 => x"81",
           801 => x"72",
           802 => x"fa",
           803 => x"f0",
           804 => x"08",
           805 => x"d5",
           806 => x"05",
           807 => x"f0",
           808 => x"22",
           809 => x"51",
           810 => x"2e",
           811 => x"82",
           812 => x"f8",
           813 => x"af",
           814 => x"fc",
           815 => x"f0",
           816 => x"33",
           817 => x"26",
           818 => x"82",
           819 => x"f8",
           820 => x"72",
           821 => x"81",
           822 => x"38",
           823 => x"08",
           824 => x"70",
           825 => x"98",
           826 => x"53",
           827 => x"82",
           828 => x"e4",
           829 => x"83",
           830 => x"32",
           831 => x"51",
           832 => x"72",
           833 => x"38",
           834 => x"08",
           835 => x"70",
           836 => x"51",
           837 => x"d5",
           838 => x"05",
           839 => x"39",
           840 => x"08",
           841 => x"70",
           842 => x"98",
           843 => x"83",
           844 => x"73",
           845 => x"51",
           846 => x"53",
           847 => x"f0",
           848 => x"34",
           849 => x"08",
           850 => x"54",
           851 => x"08",
           852 => x"70",
           853 => x"51",
           854 => x"82",
           855 => x"e8",
           856 => x"d5",
           857 => x"05",
           858 => x"2b",
           859 => x"51",
           860 => x"80",
           861 => x"80",
           862 => x"d5",
           863 => x"05",
           864 => x"f0",
           865 => x"22",
           866 => x"70",
           867 => x"51",
           868 => x"db",
           869 => x"f0",
           870 => x"33",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"d5",
           876 => x"05",
           877 => x"39",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"9d",
           883 => x"f0",
           884 => x"33",
           885 => x"70",
           886 => x"51",
           887 => x"38",
           888 => x"d5",
           889 => x"05",
           890 => x"f0",
           891 => x"33",
           892 => x"d5",
           893 => x"05",
           894 => x"d5",
           895 => x"05",
           896 => x"26",
           897 => x"82",
           898 => x"c4",
           899 => x"82",
           900 => x"8c",
           901 => x"51",
           902 => x"72",
           903 => x"f0",
           904 => x"22",
           905 => x"51",
           906 => x"d5",
           907 => x"05",
           908 => x"f0",
           909 => x"22",
           910 => x"51",
           911 => x"d5",
           912 => x"05",
           913 => x"39",
           914 => x"08",
           915 => x"70",
           916 => x"51",
           917 => x"d5",
           918 => x"05",
           919 => x"39",
           920 => x"08",
           921 => x"70",
           922 => x"51",
           923 => x"d5",
           924 => x"05",
           925 => x"39",
           926 => x"08",
           927 => x"70",
           928 => x"53",
           929 => x"f0",
           930 => x"23",
           931 => x"d5",
           932 => x"05",
           933 => x"39",
           934 => x"08",
           935 => x"70",
           936 => x"53",
           937 => x"f0",
           938 => x"23",
           939 => x"bf",
           940 => x"f0",
           941 => x"34",
           942 => x"08",
           943 => x"ff",
           944 => x"72",
           945 => x"08",
           946 => x"80",
           947 => x"d5",
           948 => x"05",
           949 => x"39",
           950 => x"08",
           951 => x"82",
           952 => x"90",
           953 => x"05",
           954 => x"08",
           955 => x"70",
           956 => x"72",
           957 => x"08",
           958 => x"82",
           959 => x"ec",
           960 => x"11",
           961 => x"82",
           962 => x"ec",
           963 => x"ef",
           964 => x"f0",
           965 => x"08",
           966 => x"08",
           967 => x"84",
           968 => x"f0",
           969 => x"0c",
           970 => x"d5",
           971 => x"05",
           972 => x"f0",
           973 => x"22",
           974 => x"70",
           975 => x"51",
           976 => x"80",
           977 => x"82",
           978 => x"e8",
           979 => x"98",
           980 => x"98",
           981 => x"d5",
           982 => x"05",
           983 => x"a4",
           984 => x"d5",
           985 => x"72",
           986 => x"08",
           987 => x"99",
           988 => x"f0",
           989 => x"08",
           990 => x"3f",
           991 => x"08",
           992 => x"d5",
           993 => x"05",
           994 => x"f0",
           995 => x"22",
           996 => x"f0",
           997 => x"22",
           998 => x"54",
           999 => x"d5",
          1000 => x"05",
          1001 => x"39",
          1002 => x"08",
          1003 => x"82",
          1004 => x"90",
          1005 => x"05",
          1006 => x"08",
          1007 => x"70",
          1008 => x"f0",
          1009 => x"0c",
          1010 => x"08",
          1011 => x"70",
          1012 => x"81",
          1013 => x"51",
          1014 => x"2e",
          1015 => x"d5",
          1016 => x"05",
          1017 => x"2b",
          1018 => x"2c",
          1019 => x"f0",
          1020 => x"08",
          1021 => x"ec",
          1022 => x"e4",
          1023 => x"82",
          1024 => x"f4",
          1025 => x"39",
          1026 => x"08",
          1027 => x"51",
          1028 => x"82",
          1029 => x"53",
          1030 => x"f0",
          1031 => x"23",
          1032 => x"08",
          1033 => x"53",
          1034 => x"08",
          1035 => x"73",
          1036 => x"54",
          1037 => x"f0",
          1038 => x"23",
          1039 => x"82",
          1040 => x"e4",
          1041 => x"82",
          1042 => x"06",
          1043 => x"72",
          1044 => x"38",
          1045 => x"08",
          1046 => x"82",
          1047 => x"90",
          1048 => x"05",
          1049 => x"08",
          1050 => x"70",
          1051 => x"f0",
          1052 => x"0c",
          1053 => x"82",
          1054 => x"90",
          1055 => x"d5",
          1056 => x"05",
          1057 => x"82",
          1058 => x"90",
          1059 => x"08",
          1060 => x"08",
          1061 => x"53",
          1062 => x"08",
          1063 => x"82",
          1064 => x"fc",
          1065 => x"d5",
          1066 => x"05",
          1067 => x"a4",
          1068 => x"f0",
          1069 => x"22",
          1070 => x"51",
          1071 => x"d5",
          1072 => x"05",
          1073 => x"f0",
          1074 => x"08",
          1075 => x"f0",
          1076 => x"0c",
          1077 => x"08",
          1078 => x"70",
          1079 => x"51",
          1080 => x"d5",
          1081 => x"05",
          1082 => x"39",
          1083 => x"d5",
          1084 => x"05",
          1085 => x"82",
          1086 => x"e4",
          1087 => x"80",
          1088 => x"53",
          1089 => x"f0",
          1090 => x"23",
          1091 => x"82",
          1092 => x"f8",
          1093 => x"0b",
          1094 => x"08",
          1095 => x"82",
          1096 => x"e4",
          1097 => x"82",
          1098 => x"06",
          1099 => x"72",
          1100 => x"38",
          1101 => x"08",
          1102 => x"82",
          1103 => x"90",
          1104 => x"05",
          1105 => x"08",
          1106 => x"70",
          1107 => x"f0",
          1108 => x"0c",
          1109 => x"82",
          1110 => x"90",
          1111 => x"d5",
          1112 => x"05",
          1113 => x"82",
          1114 => x"90",
          1115 => x"08",
          1116 => x"08",
          1117 => x"53",
          1118 => x"08",
          1119 => x"82",
          1120 => x"fc",
          1121 => x"d5",
          1122 => x"05",
          1123 => x"06",
          1124 => x"82",
          1125 => x"e4",
          1126 => x"d5",
          1127 => x"d5",
          1128 => x"05",
          1129 => x"f0",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"55",
          1135 => x"54",
          1136 => x"3f",
          1137 => x"08",
          1138 => x"34",
          1139 => x"08",
          1140 => x"82",
          1141 => x"d4",
          1142 => x"d5",
          1143 => x"05",
          1144 => x"51",
          1145 => x"27",
          1146 => x"d5",
          1147 => x"05",
          1148 => x"33",
          1149 => x"f0",
          1150 => x"33",
          1151 => x"11",
          1152 => x"72",
          1153 => x"08",
          1154 => x"97",
          1155 => x"f0",
          1156 => x"08",
          1157 => x"b0",
          1158 => x"72",
          1159 => x"08",
          1160 => x"82",
          1161 => x"d4",
          1162 => x"82",
          1163 => x"d0",
          1164 => x"34",
          1165 => x"08",
          1166 => x"81",
          1167 => x"f0",
          1168 => x"0c",
          1169 => x"08",
          1170 => x"70",
          1171 => x"f0",
          1172 => x"08",
          1173 => x"d6",
          1174 => x"e4",
          1175 => x"d5",
          1176 => x"05",
          1177 => x"d5",
          1178 => x"05",
          1179 => x"84",
          1180 => x"39",
          1181 => x"08",
          1182 => x"82",
          1183 => x"55",
          1184 => x"70",
          1185 => x"53",
          1186 => x"f0",
          1187 => x"34",
          1188 => x"08",
          1189 => x"70",
          1190 => x"53",
          1191 => x"94",
          1192 => x"f0",
          1193 => x"22",
          1194 => x"53",
          1195 => x"f0",
          1196 => x"23",
          1197 => x"08",
          1198 => x"70",
          1199 => x"81",
          1200 => x"53",
          1201 => x"80",
          1202 => x"d5",
          1203 => x"05",
          1204 => x"2b",
          1205 => x"08",
          1206 => x"82",
          1207 => x"cc",
          1208 => x"2c",
          1209 => x"08",
          1210 => x"82",
          1211 => x"f4",
          1212 => x"53",
          1213 => x"09",
          1214 => x"38",
          1215 => x"08",
          1216 => x"fe",
          1217 => x"82",
          1218 => x"c8",
          1219 => x"39",
          1220 => x"08",
          1221 => x"ff",
          1222 => x"82",
          1223 => x"c8",
          1224 => x"d5",
          1225 => x"05",
          1226 => x"f0",
          1227 => x"23",
          1228 => x"08",
          1229 => x"70",
          1230 => x"81",
          1231 => x"53",
          1232 => x"80",
          1233 => x"d5",
          1234 => x"05",
          1235 => x"2b",
          1236 => x"82",
          1237 => x"fc",
          1238 => x"51",
          1239 => x"74",
          1240 => x"82",
          1241 => x"e4",
          1242 => x"f7",
          1243 => x"72",
          1244 => x"08",
          1245 => x"9d",
          1246 => x"f0",
          1247 => x"33",
          1248 => x"f0",
          1249 => x"33",
          1250 => x"54",
          1251 => x"d5",
          1252 => x"05",
          1253 => x"f0",
          1254 => x"22",
          1255 => x"70",
          1256 => x"51",
          1257 => x"2e",
          1258 => x"d5",
          1259 => x"05",
          1260 => x"2b",
          1261 => x"70",
          1262 => x"88",
          1263 => x"51",
          1264 => x"54",
          1265 => x"08",
          1266 => x"70",
          1267 => x"53",
          1268 => x"f0",
          1269 => x"23",
          1270 => x"d5",
          1271 => x"05",
          1272 => x"2b",
          1273 => x"70",
          1274 => x"88",
          1275 => x"51",
          1276 => x"54",
          1277 => x"08",
          1278 => x"70",
          1279 => x"53",
          1280 => x"f0",
          1281 => x"23",
          1282 => x"08",
          1283 => x"70",
          1284 => x"51",
          1285 => x"38",
          1286 => x"08",
          1287 => x"ff",
          1288 => x"72",
          1289 => x"08",
          1290 => x"73",
          1291 => x"90",
          1292 => x"80",
          1293 => x"38",
          1294 => x"08",
          1295 => x"52",
          1296 => x"ee",
          1297 => x"82",
          1298 => x"e4",
          1299 => x"81",
          1300 => x"06",
          1301 => x"72",
          1302 => x"38",
          1303 => x"08",
          1304 => x"52",
          1305 => x"ca",
          1306 => x"39",
          1307 => x"08",
          1308 => x"70",
          1309 => x"81",
          1310 => x"53",
          1311 => x"90",
          1312 => x"f0",
          1313 => x"08",
          1314 => x"8a",
          1315 => x"39",
          1316 => x"08",
          1317 => x"70",
          1318 => x"81",
          1319 => x"53",
          1320 => x"8e",
          1321 => x"f0",
          1322 => x"08",
          1323 => x"8a",
          1324 => x"d5",
          1325 => x"05",
          1326 => x"2a",
          1327 => x"51",
          1328 => x"80",
          1329 => x"82",
          1330 => x"88",
          1331 => x"b0",
          1332 => x"3f",
          1333 => x"08",
          1334 => x"53",
          1335 => x"09",
          1336 => x"38",
          1337 => x"08",
          1338 => x"52",
          1339 => x"08",
          1340 => x"51",
          1341 => x"82",
          1342 => x"e4",
          1343 => x"88",
          1344 => x"06",
          1345 => x"72",
          1346 => x"38",
          1347 => x"08",
          1348 => x"ff",
          1349 => x"72",
          1350 => x"08",
          1351 => x"73",
          1352 => x"90",
          1353 => x"80",
          1354 => x"38",
          1355 => x"08",
          1356 => x"52",
          1357 => x"fa",
          1358 => x"82",
          1359 => x"e4",
          1360 => x"83",
          1361 => x"06",
          1362 => x"72",
          1363 => x"38",
          1364 => x"08",
          1365 => x"ff",
          1366 => x"72",
          1367 => x"08",
          1368 => x"73",
          1369 => x"98",
          1370 => x"80",
          1371 => x"38",
          1372 => x"08",
          1373 => x"52",
          1374 => x"b6",
          1375 => x"82",
          1376 => x"e4",
          1377 => x"87",
          1378 => x"06",
          1379 => x"72",
          1380 => x"d5",
          1381 => x"05",
          1382 => x"54",
          1383 => x"d5",
          1384 => x"05",
          1385 => x"2b",
          1386 => x"51",
          1387 => x"25",
          1388 => x"d5",
          1389 => x"05",
          1390 => x"51",
          1391 => x"d2",
          1392 => x"f0",
          1393 => x"33",
          1394 => x"e3",
          1395 => x"06",
          1396 => x"d5",
          1397 => x"05",
          1398 => x"d5",
          1399 => x"05",
          1400 => x"ce",
          1401 => x"39",
          1402 => x"08",
          1403 => x"53",
          1404 => x"2e",
          1405 => x"80",
          1406 => x"d5",
          1407 => x"05",
          1408 => x"51",
          1409 => x"d5",
          1410 => x"05",
          1411 => x"ff",
          1412 => x"72",
          1413 => x"2e",
          1414 => x"82",
          1415 => x"88",
          1416 => x"82",
          1417 => x"fc",
          1418 => x"33",
          1419 => x"f0",
          1420 => x"08",
          1421 => x"d5",
          1422 => x"05",
          1423 => x"f2",
          1424 => x"39",
          1425 => x"08",
          1426 => x"53",
          1427 => x"2e",
          1428 => x"80",
          1429 => x"d5",
          1430 => x"05",
          1431 => x"51",
          1432 => x"d5",
          1433 => x"05",
          1434 => x"ff",
          1435 => x"72",
          1436 => x"2e",
          1437 => x"82",
          1438 => x"88",
          1439 => x"82",
          1440 => x"fc",
          1441 => x"33",
          1442 => x"a6",
          1443 => x"f0",
          1444 => x"08",
          1445 => x"d5",
          1446 => x"05",
          1447 => x"39",
          1448 => x"08",
          1449 => x"82",
          1450 => x"a9",
          1451 => x"f0",
          1452 => x"08",
          1453 => x"f0",
          1454 => x"08",
          1455 => x"d5",
          1456 => x"05",
          1457 => x"f0",
          1458 => x"08",
          1459 => x"53",
          1460 => x"cc",
          1461 => x"f0",
          1462 => x"22",
          1463 => x"70",
          1464 => x"51",
          1465 => x"2e",
          1466 => x"82",
          1467 => x"ec",
          1468 => x"11",
          1469 => x"82",
          1470 => x"ec",
          1471 => x"90",
          1472 => x"2c",
          1473 => x"73",
          1474 => x"82",
          1475 => x"88",
          1476 => x"a0",
          1477 => x"3f",
          1478 => x"d5",
          1479 => x"05",
          1480 => x"d5",
          1481 => x"05",
          1482 => x"86",
          1483 => x"82",
          1484 => x"e4",
          1485 => x"b7",
          1486 => x"f0",
          1487 => x"33",
          1488 => x"2e",
          1489 => x"a8",
          1490 => x"82",
          1491 => x"e4",
          1492 => x"0b",
          1493 => x"08",
          1494 => x"80",
          1495 => x"f0",
          1496 => x"34",
          1497 => x"d5",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"52",
          1502 => x"08",
          1503 => x"51",
          1504 => x"e9",
          1505 => x"d5",
          1506 => x"05",
          1507 => x"08",
          1508 => x"f0",
          1509 => x"0c",
          1510 => x"d5",
          1511 => x"05",
          1512 => x"e4",
          1513 => x"0d",
          1514 => x"0c",
          1515 => x"f0",
          1516 => x"d5",
          1517 => x"3d",
          1518 => x"c4",
          1519 => x"d5",
          1520 => x"05",
          1521 => x"d5",
          1522 => x"05",
          1523 => x"dd",
          1524 => x"e4",
          1525 => x"d5",
          1526 => x"85",
          1527 => x"d5",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"80",
          1532 => x"f0",
          1533 => x"0c",
          1534 => x"08",
          1535 => x"70",
          1536 => x"81",
          1537 => x"06",
          1538 => x"51",
          1539 => x"2e",
          1540 => x"0b",
          1541 => x"08",
          1542 => x"81",
          1543 => x"d5",
          1544 => x"05",
          1545 => x"33",
          1546 => x"08",
          1547 => x"81",
          1548 => x"f0",
          1549 => x"0c",
          1550 => x"d5",
          1551 => x"05",
          1552 => x"ff",
          1553 => x"80",
          1554 => x"82",
          1555 => x"82",
          1556 => x"53",
          1557 => x"08",
          1558 => x"52",
          1559 => x"51",
          1560 => x"82",
          1561 => x"53",
          1562 => x"ff",
          1563 => x"0b",
          1564 => x"08",
          1565 => x"ff",
          1566 => x"f1",
          1567 => x"f1",
          1568 => x"53",
          1569 => x"13",
          1570 => x"2d",
          1571 => x"08",
          1572 => x"2e",
          1573 => x"0b",
          1574 => x"08",
          1575 => x"82",
          1576 => x"f8",
          1577 => x"82",
          1578 => x"f4",
          1579 => x"82",
          1580 => x"f4",
          1581 => x"d5",
          1582 => x"3d",
          1583 => x"f0",
          1584 => x"d5",
          1585 => x"82",
          1586 => x"fb",
          1587 => x"0b",
          1588 => x"08",
          1589 => x"82",
          1590 => x"8c",
          1591 => x"11",
          1592 => x"2a",
          1593 => x"70",
          1594 => x"51",
          1595 => x"72",
          1596 => x"38",
          1597 => x"d5",
          1598 => x"05",
          1599 => x"39",
          1600 => x"08",
          1601 => x"53",
          1602 => x"d5",
          1603 => x"05",
          1604 => x"82",
          1605 => x"88",
          1606 => x"72",
          1607 => x"08",
          1608 => x"72",
          1609 => x"53",
          1610 => x"b6",
          1611 => x"f0",
          1612 => x"08",
          1613 => x"08",
          1614 => x"53",
          1615 => x"08",
          1616 => x"52",
          1617 => x"51",
          1618 => x"82",
          1619 => x"53",
          1620 => x"ff",
          1621 => x"0b",
          1622 => x"08",
          1623 => x"ff",
          1624 => x"d5",
          1625 => x"05",
          1626 => x"d5",
          1627 => x"05",
          1628 => x"d5",
          1629 => x"05",
          1630 => x"e4",
          1631 => x"0d",
          1632 => x"0c",
          1633 => x"f0",
          1634 => x"d5",
          1635 => x"3d",
          1636 => x"c8",
          1637 => x"d5",
          1638 => x"05",
          1639 => x"3f",
          1640 => x"08",
          1641 => x"e4",
          1642 => x"3d",
          1643 => x"f0",
          1644 => x"d5",
          1645 => x"82",
          1646 => x"fb",
          1647 => x"d5",
          1648 => x"05",
          1649 => x"33",
          1650 => x"70",
          1651 => x"81",
          1652 => x"51",
          1653 => x"80",
          1654 => x"ff",
          1655 => x"f0",
          1656 => x"0c",
          1657 => x"82",
          1658 => x"8c",
          1659 => x"11",
          1660 => x"2a",
          1661 => x"51",
          1662 => x"72",
          1663 => x"db",
          1664 => x"f0",
          1665 => x"08",
          1666 => x"08",
          1667 => x"54",
          1668 => x"08",
          1669 => x"25",
          1670 => x"d5",
          1671 => x"05",
          1672 => x"70",
          1673 => x"08",
          1674 => x"52",
          1675 => x"72",
          1676 => x"08",
          1677 => x"0c",
          1678 => x"08",
          1679 => x"8c",
          1680 => x"05",
          1681 => x"82",
          1682 => x"88",
          1683 => x"82",
          1684 => x"fc",
          1685 => x"53",
          1686 => x"82",
          1687 => x"8c",
          1688 => x"d5",
          1689 => x"05",
          1690 => x"d5",
          1691 => x"05",
          1692 => x"ff",
          1693 => x"12",
          1694 => x"54",
          1695 => x"d5",
          1696 => x"72",
          1697 => x"d5",
          1698 => x"05",
          1699 => x"08",
          1700 => x"12",
          1701 => x"f0",
          1702 => x"08",
          1703 => x"f0",
          1704 => x"0c",
          1705 => x"39",
          1706 => x"d5",
          1707 => x"05",
          1708 => x"f0",
          1709 => x"08",
          1710 => x"0c",
          1711 => x"82",
          1712 => x"04",
          1713 => x"08",
          1714 => x"f0",
          1715 => x"0d",
          1716 => x"08",
          1717 => x"85",
          1718 => x"81",
          1719 => x"06",
          1720 => x"52",
          1721 => x"8d",
          1722 => x"82",
          1723 => x"f8",
          1724 => x"94",
          1725 => x"f0",
          1726 => x"08",
          1727 => x"70",
          1728 => x"81",
          1729 => x"51",
          1730 => x"2e",
          1731 => x"82",
          1732 => x"88",
          1733 => x"d5",
          1734 => x"05",
          1735 => x"85",
          1736 => x"ff",
          1737 => x"52",
          1738 => x"34",
          1739 => x"08",
          1740 => x"8c",
          1741 => x"05",
          1742 => x"82",
          1743 => x"88",
          1744 => x"11",
          1745 => x"d5",
          1746 => x"05",
          1747 => x"52",
          1748 => x"82",
          1749 => x"88",
          1750 => x"11",
          1751 => x"2a",
          1752 => x"51",
          1753 => x"71",
          1754 => x"d7",
          1755 => x"f0",
          1756 => x"08",
          1757 => x"33",
          1758 => x"08",
          1759 => x"51",
          1760 => x"f0",
          1761 => x"08",
          1762 => x"d5",
          1763 => x"05",
          1764 => x"f0",
          1765 => x"08",
          1766 => x"12",
          1767 => x"07",
          1768 => x"85",
          1769 => x"0b",
          1770 => x"08",
          1771 => x"81",
          1772 => x"d5",
          1773 => x"05",
          1774 => x"81",
          1775 => x"52",
          1776 => x"82",
          1777 => x"88",
          1778 => x"d5",
          1779 => x"05",
          1780 => x"11",
          1781 => x"71",
          1782 => x"e4",
          1783 => x"d5",
          1784 => x"05",
          1785 => x"d5",
          1786 => x"05",
          1787 => x"80",
          1788 => x"d5",
          1789 => x"05",
          1790 => x"f0",
          1791 => x"0c",
          1792 => x"08",
          1793 => x"85",
          1794 => x"d5",
          1795 => x"05",
          1796 => x"d5",
          1797 => x"05",
          1798 => x"09",
          1799 => x"38",
          1800 => x"08",
          1801 => x"90",
          1802 => x"82",
          1803 => x"ec",
          1804 => x"39",
          1805 => x"08",
          1806 => x"a0",
          1807 => x"82",
          1808 => x"ec",
          1809 => x"d5",
          1810 => x"05",
          1811 => x"d5",
          1812 => x"05",
          1813 => x"34",
          1814 => x"d5",
          1815 => x"05",
          1816 => x"82",
          1817 => x"88",
          1818 => x"11",
          1819 => x"8c",
          1820 => x"d5",
          1821 => x"05",
          1822 => x"ff",
          1823 => x"d5",
          1824 => x"05",
          1825 => x"52",
          1826 => x"08",
          1827 => x"82",
          1828 => x"89",
          1829 => x"d5",
          1830 => x"82",
          1831 => x"02",
          1832 => x"0c",
          1833 => x"82",
          1834 => x"88",
          1835 => x"d5",
          1836 => x"05",
          1837 => x"f0",
          1838 => x"08",
          1839 => x"08",
          1840 => x"82",
          1841 => x"90",
          1842 => x"2e",
          1843 => x"82",
          1844 => x"f8",
          1845 => x"d5",
          1846 => x"05",
          1847 => x"ac",
          1848 => x"f0",
          1849 => x"08",
          1850 => x"08",
          1851 => x"05",
          1852 => x"f0",
          1853 => x"08",
          1854 => x"90",
          1855 => x"f0",
          1856 => x"08",
          1857 => x"08",
          1858 => x"05",
          1859 => x"08",
          1860 => x"82",
          1861 => x"f8",
          1862 => x"d5",
          1863 => x"05",
          1864 => x"d5",
          1865 => x"05",
          1866 => x"f0",
          1867 => x"08",
          1868 => x"d5",
          1869 => x"05",
          1870 => x"f0",
          1871 => x"08",
          1872 => x"d5",
          1873 => x"05",
          1874 => x"f0",
          1875 => x"08",
          1876 => x"9c",
          1877 => x"f0",
          1878 => x"08",
          1879 => x"d5",
          1880 => x"05",
          1881 => x"f0",
          1882 => x"08",
          1883 => x"d5",
          1884 => x"05",
          1885 => x"f0",
          1886 => x"08",
          1887 => x"08",
          1888 => x"53",
          1889 => x"71",
          1890 => x"39",
          1891 => x"08",
          1892 => x"81",
          1893 => x"f0",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"f0",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"80",
          1901 => x"82",
          1902 => x"f8",
          1903 => x"70",
          1904 => x"f0",
          1905 => x"08",
          1906 => x"d5",
          1907 => x"05",
          1908 => x"f0",
          1909 => x"08",
          1910 => x"71",
          1911 => x"f0",
          1912 => x"08",
          1913 => x"d5",
          1914 => x"05",
          1915 => x"39",
          1916 => x"08",
          1917 => x"70",
          1918 => x"0c",
          1919 => x"0d",
          1920 => x"0c",
          1921 => x"f0",
          1922 => x"d5",
          1923 => x"3d",
          1924 => x"f0",
          1925 => x"08",
          1926 => x"08",
          1927 => x"82",
          1928 => x"fc",
          1929 => x"71",
          1930 => x"f0",
          1931 => x"08",
          1932 => x"d5",
          1933 => x"05",
          1934 => x"ff",
          1935 => x"70",
          1936 => x"38",
          1937 => x"d5",
          1938 => x"05",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"d5",
          1942 => x"05",
          1943 => x"f0",
          1944 => x"08",
          1945 => x"d5",
          1946 => x"84",
          1947 => x"d5",
          1948 => x"82",
          1949 => x"02",
          1950 => x"0c",
          1951 => x"82",
          1952 => x"88",
          1953 => x"d5",
          1954 => x"05",
          1955 => x"f0",
          1956 => x"08",
          1957 => x"82",
          1958 => x"8c",
          1959 => x"05",
          1960 => x"08",
          1961 => x"82",
          1962 => x"fc",
          1963 => x"51",
          1964 => x"82",
          1965 => x"fc",
          1966 => x"05",
          1967 => x"08",
          1968 => x"70",
          1969 => x"51",
          1970 => x"84",
          1971 => x"39",
          1972 => x"08",
          1973 => x"70",
          1974 => x"0c",
          1975 => x"0d",
          1976 => x"0c",
          1977 => x"f0",
          1978 => x"d5",
          1979 => x"3d",
          1980 => x"f0",
          1981 => x"08",
          1982 => x"08",
          1983 => x"82",
          1984 => x"8c",
          1985 => x"d5",
          1986 => x"05",
          1987 => x"f0",
          1988 => x"08",
          1989 => x"e5",
          1990 => x"f0",
          1991 => x"08",
          1992 => x"d5",
          1993 => x"05",
          1994 => x"f0",
          1995 => x"08",
          1996 => x"d5",
          1997 => x"05",
          1998 => x"f0",
          1999 => x"08",
          2000 => x"38",
          2001 => x"08",
          2002 => x"51",
          2003 => x"d5",
          2004 => x"05",
          2005 => x"82",
          2006 => x"f8",
          2007 => x"d5",
          2008 => x"05",
          2009 => x"71",
          2010 => x"d5",
          2011 => x"05",
          2012 => x"82",
          2013 => x"fc",
          2014 => x"ad",
          2015 => x"f0",
          2016 => x"08",
          2017 => x"e4",
          2018 => x"3d",
          2019 => x"f0",
          2020 => x"d5",
          2021 => x"82",
          2022 => x"fd",
          2023 => x"d5",
          2024 => x"05",
          2025 => x"81",
          2026 => x"d5",
          2027 => x"05",
          2028 => x"33",
          2029 => x"08",
          2030 => x"81",
          2031 => x"f0",
          2032 => x"0c",
          2033 => x"08",
          2034 => x"70",
          2035 => x"ff",
          2036 => x"54",
          2037 => x"2e",
          2038 => x"ce",
          2039 => x"f0",
          2040 => x"08",
          2041 => x"82",
          2042 => x"88",
          2043 => x"05",
          2044 => x"08",
          2045 => x"70",
          2046 => x"51",
          2047 => x"38",
          2048 => x"d5",
          2049 => x"05",
          2050 => x"39",
          2051 => x"08",
          2052 => x"ff",
          2053 => x"f0",
          2054 => x"0c",
          2055 => x"08",
          2056 => x"80",
          2057 => x"ff",
          2058 => x"d5",
          2059 => x"05",
          2060 => x"80",
          2061 => x"d5",
          2062 => x"05",
          2063 => x"52",
          2064 => x"38",
          2065 => x"d5",
          2066 => x"05",
          2067 => x"39",
          2068 => x"08",
          2069 => x"ff",
          2070 => x"f0",
          2071 => x"0c",
          2072 => x"08",
          2073 => x"70",
          2074 => x"70",
          2075 => x"0b",
          2076 => x"08",
          2077 => x"ae",
          2078 => x"f0",
          2079 => x"08",
          2080 => x"d5",
          2081 => x"05",
          2082 => x"72",
          2083 => x"82",
          2084 => x"fc",
          2085 => x"55",
          2086 => x"8a",
          2087 => x"82",
          2088 => x"fc",
          2089 => x"d5",
          2090 => x"05",
          2091 => x"e4",
          2092 => x"0d",
          2093 => x"0c",
          2094 => x"f0",
          2095 => x"d5",
          2096 => x"3d",
          2097 => x"f0",
          2098 => x"08",
          2099 => x"f0",
          2100 => x"08",
          2101 => x"3f",
          2102 => x"08",
          2103 => x"f0",
          2104 => x"0c",
          2105 => x"08",
          2106 => x"81",
          2107 => x"51",
          2108 => x"db",
          2109 => x"e4",
          2110 => x"d5",
          2111 => x"05",
          2112 => x"d5",
          2113 => x"05",
          2114 => x"80",
          2115 => x"f0",
          2116 => x"0c",
          2117 => x"d5",
          2118 => x"05",
          2119 => x"f0",
          2120 => x"08",
          2121 => x"74",
          2122 => x"f0",
          2123 => x"08",
          2124 => x"f0",
          2125 => x"08",
          2126 => x"f0",
          2127 => x"08",
          2128 => x"3f",
          2129 => x"08",
          2130 => x"f0",
          2131 => x"0c",
          2132 => x"f0",
          2133 => x"08",
          2134 => x"0c",
          2135 => x"82",
          2136 => x"04",
          2137 => x"08",
          2138 => x"f0",
          2139 => x"0d",
          2140 => x"08",
          2141 => x"82",
          2142 => x"f8",
          2143 => x"d5",
          2144 => x"05",
          2145 => x"80",
          2146 => x"f0",
          2147 => x"0c",
          2148 => x"82",
          2149 => x"f8",
          2150 => x"71",
          2151 => x"f0",
          2152 => x"08",
          2153 => x"d5",
          2154 => x"05",
          2155 => x"ff",
          2156 => x"70",
          2157 => x"38",
          2158 => x"08",
          2159 => x"ff",
          2160 => x"f0",
          2161 => x"0c",
          2162 => x"08",
          2163 => x"ff",
          2164 => x"ff",
          2165 => x"d5",
          2166 => x"05",
          2167 => x"82",
          2168 => x"f8",
          2169 => x"d5",
          2170 => x"05",
          2171 => x"f0",
          2172 => x"08",
          2173 => x"d5",
          2174 => x"05",
          2175 => x"d5",
          2176 => x"05",
          2177 => x"e4",
          2178 => x"0d",
          2179 => x"0c",
          2180 => x"f0",
          2181 => x"d5",
          2182 => x"3d",
          2183 => x"f0",
          2184 => x"08",
          2185 => x"08",
          2186 => x"82",
          2187 => x"90",
          2188 => x"2e",
          2189 => x"82",
          2190 => x"90",
          2191 => x"05",
          2192 => x"08",
          2193 => x"82",
          2194 => x"90",
          2195 => x"05",
          2196 => x"08",
          2197 => x"82",
          2198 => x"90",
          2199 => x"2e",
          2200 => x"d5",
          2201 => x"05",
          2202 => x"82",
          2203 => x"fc",
          2204 => x"52",
          2205 => x"82",
          2206 => x"fc",
          2207 => x"05",
          2208 => x"08",
          2209 => x"ff",
          2210 => x"d5",
          2211 => x"05",
          2212 => x"d5",
          2213 => x"84",
          2214 => x"d5",
          2215 => x"82",
          2216 => x"02",
          2217 => x"0c",
          2218 => x"80",
          2219 => x"f0",
          2220 => x"0c",
          2221 => x"08",
          2222 => x"80",
          2223 => x"82",
          2224 => x"88",
          2225 => x"82",
          2226 => x"88",
          2227 => x"0b",
          2228 => x"08",
          2229 => x"82",
          2230 => x"fc",
          2231 => x"38",
          2232 => x"d5",
          2233 => x"05",
          2234 => x"f0",
          2235 => x"08",
          2236 => x"08",
          2237 => x"82",
          2238 => x"8c",
          2239 => x"25",
          2240 => x"d5",
          2241 => x"05",
          2242 => x"d5",
          2243 => x"05",
          2244 => x"82",
          2245 => x"f0",
          2246 => x"d5",
          2247 => x"05",
          2248 => x"81",
          2249 => x"f0",
          2250 => x"0c",
          2251 => x"08",
          2252 => x"82",
          2253 => x"fc",
          2254 => x"53",
          2255 => x"08",
          2256 => x"52",
          2257 => x"08",
          2258 => x"51",
          2259 => x"82",
          2260 => x"70",
          2261 => x"08",
          2262 => x"54",
          2263 => x"08",
          2264 => x"80",
          2265 => x"82",
          2266 => x"f8",
          2267 => x"82",
          2268 => x"f8",
          2269 => x"d5",
          2270 => x"05",
          2271 => x"d5",
          2272 => x"89",
          2273 => x"d5",
          2274 => x"82",
          2275 => x"02",
          2276 => x"0c",
          2277 => x"80",
          2278 => x"f0",
          2279 => x"0c",
          2280 => x"08",
          2281 => x"80",
          2282 => x"82",
          2283 => x"88",
          2284 => x"82",
          2285 => x"88",
          2286 => x"0b",
          2287 => x"08",
          2288 => x"82",
          2289 => x"8c",
          2290 => x"25",
          2291 => x"d5",
          2292 => x"05",
          2293 => x"d5",
          2294 => x"05",
          2295 => x"82",
          2296 => x"8c",
          2297 => x"82",
          2298 => x"88",
          2299 => x"81",
          2300 => x"d5",
          2301 => x"82",
          2302 => x"f8",
          2303 => x"82",
          2304 => x"fc",
          2305 => x"2e",
          2306 => x"d5",
          2307 => x"05",
          2308 => x"d5",
          2309 => x"05",
          2310 => x"f0",
          2311 => x"08",
          2312 => x"e4",
          2313 => x"3d",
          2314 => x"f0",
          2315 => x"d5",
          2316 => x"82",
          2317 => x"fd",
          2318 => x"53",
          2319 => x"08",
          2320 => x"52",
          2321 => x"08",
          2322 => x"51",
          2323 => x"82",
          2324 => x"70",
          2325 => x"0c",
          2326 => x"0d",
          2327 => x"0c",
          2328 => x"f0",
          2329 => x"d5",
          2330 => x"3d",
          2331 => x"82",
          2332 => x"8c",
          2333 => x"82",
          2334 => x"88",
          2335 => x"93",
          2336 => x"e4",
          2337 => x"d5",
          2338 => x"85",
          2339 => x"d5",
          2340 => x"82",
          2341 => x"02",
          2342 => x"0c",
          2343 => x"81",
          2344 => x"f0",
          2345 => x"0c",
          2346 => x"d5",
          2347 => x"05",
          2348 => x"f0",
          2349 => x"08",
          2350 => x"08",
          2351 => x"27",
          2352 => x"d5",
          2353 => x"05",
          2354 => x"ae",
          2355 => x"82",
          2356 => x"8c",
          2357 => x"a2",
          2358 => x"f0",
          2359 => x"08",
          2360 => x"f0",
          2361 => x"0c",
          2362 => x"08",
          2363 => x"10",
          2364 => x"08",
          2365 => x"ff",
          2366 => x"d5",
          2367 => x"05",
          2368 => x"80",
          2369 => x"d5",
          2370 => x"05",
          2371 => x"f0",
          2372 => x"08",
          2373 => x"82",
          2374 => x"88",
          2375 => x"d5",
          2376 => x"05",
          2377 => x"d5",
          2378 => x"05",
          2379 => x"f0",
          2380 => x"08",
          2381 => x"08",
          2382 => x"07",
          2383 => x"08",
          2384 => x"82",
          2385 => x"fc",
          2386 => x"2a",
          2387 => x"08",
          2388 => x"82",
          2389 => x"8c",
          2390 => x"2a",
          2391 => x"08",
          2392 => x"ff",
          2393 => x"d5",
          2394 => x"05",
          2395 => x"93",
          2396 => x"f0",
          2397 => x"08",
          2398 => x"f0",
          2399 => x"0c",
          2400 => x"82",
          2401 => x"f8",
          2402 => x"82",
          2403 => x"f4",
          2404 => x"82",
          2405 => x"f4",
          2406 => x"d5",
          2407 => x"3d",
          2408 => x"f0",
          2409 => x"d5",
          2410 => x"82",
          2411 => x"f7",
          2412 => x"0b",
          2413 => x"08",
          2414 => x"82",
          2415 => x"8c",
          2416 => x"80",
          2417 => x"d5",
          2418 => x"05",
          2419 => x"51",
          2420 => x"53",
          2421 => x"f0",
          2422 => x"34",
          2423 => x"06",
          2424 => x"2e",
          2425 => x"91",
          2426 => x"f0",
          2427 => x"08",
          2428 => x"05",
          2429 => x"ce",
          2430 => x"f0",
          2431 => x"33",
          2432 => x"2e",
          2433 => x"a4",
          2434 => x"82",
          2435 => x"f0",
          2436 => x"d5",
          2437 => x"05",
          2438 => x"81",
          2439 => x"70",
          2440 => x"72",
          2441 => x"f0",
          2442 => x"34",
          2443 => x"08",
          2444 => x"53",
          2445 => x"09",
          2446 => x"dc",
          2447 => x"f0",
          2448 => x"08",
          2449 => x"05",
          2450 => x"08",
          2451 => x"33",
          2452 => x"08",
          2453 => x"82",
          2454 => x"f8",
          2455 => x"d5",
          2456 => x"05",
          2457 => x"f0",
          2458 => x"08",
          2459 => x"b6",
          2460 => x"f0",
          2461 => x"08",
          2462 => x"84",
          2463 => x"39",
          2464 => x"d5",
          2465 => x"05",
          2466 => x"f0",
          2467 => x"08",
          2468 => x"05",
          2469 => x"08",
          2470 => x"33",
          2471 => x"08",
          2472 => x"81",
          2473 => x"0b",
          2474 => x"08",
          2475 => x"82",
          2476 => x"88",
          2477 => x"08",
          2478 => x"0c",
          2479 => x"53",
          2480 => x"d5",
          2481 => x"05",
          2482 => x"39",
          2483 => x"08",
          2484 => x"53",
          2485 => x"8d",
          2486 => x"82",
          2487 => x"ec",
          2488 => x"80",
          2489 => x"f0",
          2490 => x"33",
          2491 => x"27",
          2492 => x"d5",
          2493 => x"05",
          2494 => x"b9",
          2495 => x"8d",
          2496 => x"82",
          2497 => x"ec",
          2498 => x"d8",
          2499 => x"82",
          2500 => x"f4",
          2501 => x"39",
          2502 => x"08",
          2503 => x"53",
          2504 => x"90",
          2505 => x"f0",
          2506 => x"33",
          2507 => x"26",
          2508 => x"39",
          2509 => x"d5",
          2510 => x"05",
          2511 => x"39",
          2512 => x"d5",
          2513 => x"05",
          2514 => x"82",
          2515 => x"fc",
          2516 => x"d5",
          2517 => x"05",
          2518 => x"73",
          2519 => x"38",
          2520 => x"08",
          2521 => x"53",
          2522 => x"27",
          2523 => x"d5",
          2524 => x"05",
          2525 => x"51",
          2526 => x"d5",
          2527 => x"05",
          2528 => x"f0",
          2529 => x"33",
          2530 => x"53",
          2531 => x"f0",
          2532 => x"34",
          2533 => x"08",
          2534 => x"53",
          2535 => x"ad",
          2536 => x"f0",
          2537 => x"33",
          2538 => x"53",
          2539 => x"f0",
          2540 => x"34",
          2541 => x"08",
          2542 => x"53",
          2543 => x"8d",
          2544 => x"82",
          2545 => x"ec",
          2546 => x"98",
          2547 => x"f0",
          2548 => x"33",
          2549 => x"08",
          2550 => x"54",
          2551 => x"26",
          2552 => x"0b",
          2553 => x"08",
          2554 => x"80",
          2555 => x"d5",
          2556 => x"05",
          2557 => x"d5",
          2558 => x"05",
          2559 => x"d5",
          2560 => x"05",
          2561 => x"82",
          2562 => x"fc",
          2563 => x"d5",
          2564 => x"05",
          2565 => x"81",
          2566 => x"70",
          2567 => x"52",
          2568 => x"33",
          2569 => x"08",
          2570 => x"fe",
          2571 => x"d5",
          2572 => x"05",
          2573 => x"80",
          2574 => x"82",
          2575 => x"fc",
          2576 => x"82",
          2577 => x"fc",
          2578 => x"d5",
          2579 => x"05",
          2580 => x"f0",
          2581 => x"08",
          2582 => x"81",
          2583 => x"f0",
          2584 => x"0c",
          2585 => x"08",
          2586 => x"82",
          2587 => x"8b",
          2588 => x"d5",
          2589 => x"82",
          2590 => x"02",
          2591 => x"0c",
          2592 => x"80",
          2593 => x"f0",
          2594 => x"34",
          2595 => x"08",
          2596 => x"53",
          2597 => x"82",
          2598 => x"88",
          2599 => x"08",
          2600 => x"33",
          2601 => x"d5",
          2602 => x"05",
          2603 => x"ff",
          2604 => x"a0",
          2605 => x"06",
          2606 => x"d5",
          2607 => x"05",
          2608 => x"81",
          2609 => x"53",
          2610 => x"d5",
          2611 => x"05",
          2612 => x"ad",
          2613 => x"06",
          2614 => x"0b",
          2615 => x"08",
          2616 => x"82",
          2617 => x"88",
          2618 => x"08",
          2619 => x"0c",
          2620 => x"53",
          2621 => x"d5",
          2622 => x"05",
          2623 => x"f0",
          2624 => x"33",
          2625 => x"2e",
          2626 => x"81",
          2627 => x"d5",
          2628 => x"05",
          2629 => x"81",
          2630 => x"70",
          2631 => x"72",
          2632 => x"f0",
          2633 => x"34",
          2634 => x"08",
          2635 => x"82",
          2636 => x"e8",
          2637 => x"d5",
          2638 => x"05",
          2639 => x"2e",
          2640 => x"d5",
          2641 => x"05",
          2642 => x"2e",
          2643 => x"cd",
          2644 => x"82",
          2645 => x"f4",
          2646 => x"d5",
          2647 => x"05",
          2648 => x"81",
          2649 => x"70",
          2650 => x"72",
          2651 => x"f0",
          2652 => x"34",
          2653 => x"82",
          2654 => x"f0",
          2655 => x"34",
          2656 => x"08",
          2657 => x"70",
          2658 => x"71",
          2659 => x"51",
          2660 => x"82",
          2661 => x"f8",
          2662 => x"fe",
          2663 => x"f0",
          2664 => x"33",
          2665 => x"26",
          2666 => x"0b",
          2667 => x"08",
          2668 => x"83",
          2669 => x"d5",
          2670 => x"05",
          2671 => x"73",
          2672 => x"82",
          2673 => x"f8",
          2674 => x"72",
          2675 => x"38",
          2676 => x"0b",
          2677 => x"08",
          2678 => x"82",
          2679 => x"0b",
          2680 => x"08",
          2681 => x"b2",
          2682 => x"f0",
          2683 => x"33",
          2684 => x"27",
          2685 => x"d5",
          2686 => x"05",
          2687 => x"b9",
          2688 => x"8d",
          2689 => x"82",
          2690 => x"ec",
          2691 => x"a5",
          2692 => x"82",
          2693 => x"f4",
          2694 => x"0b",
          2695 => x"08",
          2696 => x"82",
          2697 => x"f8",
          2698 => x"a0",
          2699 => x"cf",
          2700 => x"f0",
          2701 => x"33",
          2702 => x"73",
          2703 => x"82",
          2704 => x"f8",
          2705 => x"11",
          2706 => x"82",
          2707 => x"f8",
          2708 => x"d5",
          2709 => x"05",
          2710 => x"51",
          2711 => x"d5",
          2712 => x"05",
          2713 => x"f0",
          2714 => x"33",
          2715 => x"27",
          2716 => x"d5",
          2717 => x"05",
          2718 => x"51",
          2719 => x"d5",
          2720 => x"05",
          2721 => x"f0",
          2722 => x"33",
          2723 => x"26",
          2724 => x"0b",
          2725 => x"08",
          2726 => x"81",
          2727 => x"d5",
          2728 => x"05",
          2729 => x"f0",
          2730 => x"33",
          2731 => x"74",
          2732 => x"80",
          2733 => x"f0",
          2734 => x"0c",
          2735 => x"82",
          2736 => x"f4",
          2737 => x"82",
          2738 => x"fc",
          2739 => x"82",
          2740 => x"f8",
          2741 => x"12",
          2742 => x"08",
          2743 => x"82",
          2744 => x"88",
          2745 => x"08",
          2746 => x"0c",
          2747 => x"51",
          2748 => x"72",
          2749 => x"f0",
          2750 => x"34",
          2751 => x"82",
          2752 => x"f0",
          2753 => x"72",
          2754 => x"38",
          2755 => x"08",
          2756 => x"30",
          2757 => x"08",
          2758 => x"82",
          2759 => x"8c",
          2760 => x"d5",
          2761 => x"05",
          2762 => x"53",
          2763 => x"d5",
          2764 => x"05",
          2765 => x"f0",
          2766 => x"08",
          2767 => x"0c",
          2768 => x"82",
          2769 => x"04",
          2770 => x"7a",
          2771 => x"56",
          2772 => x"80",
          2773 => x"38",
          2774 => x"15",
          2775 => x"16",
          2776 => x"d2",
          2777 => x"54",
          2778 => x"09",
          2779 => x"38",
          2780 => x"f1",
          2781 => x"76",
          2782 => x"d0",
          2783 => x"08",
          2784 => x"81",
          2785 => x"e4",
          2786 => x"e4",
          2787 => x"53",
          2788 => x"58",
          2789 => x"82",
          2790 => x"8b",
          2791 => x"33",
          2792 => x"2e",
          2793 => x"81",
          2794 => x"ff",
          2795 => x"99",
          2796 => x"38",
          2797 => x"82",
          2798 => x"8a",
          2799 => x"ff",
          2800 => x"52",
          2801 => x"81",
          2802 => x"84",
          2803 => x"ac",
          2804 => x"08",
          2805 => x"9c",
          2806 => x"39",
          2807 => x"51",
          2808 => x"82",
          2809 => x"80",
          2810 => x"b3",
          2811 => x"eb",
          2812 => x"d8",
          2813 => x"39",
          2814 => x"51",
          2815 => x"82",
          2816 => x"80",
          2817 => x"b4",
          2818 => x"cf",
          2819 => x"a4",
          2820 => x"39",
          2821 => x"51",
          2822 => x"82",
          2823 => x"bb",
          2824 => x"f0",
          2825 => x"82",
          2826 => x"af",
          2827 => x"ac",
          2828 => x"82",
          2829 => x"a3",
          2830 => x"dc",
          2831 => x"82",
          2832 => x"97",
          2833 => x"84",
          2834 => x"82",
          2835 => x"8b",
          2836 => x"b4",
          2837 => x"82",
          2838 => x"d7",
          2839 => x"3d",
          2840 => x"3d",
          2841 => x"56",
          2842 => x"e7",
          2843 => x"74",
          2844 => x"e8",
          2845 => x"39",
          2846 => x"74",
          2847 => x"3f",
          2848 => x"08",
          2849 => x"ef",
          2850 => x"d5",
          2851 => x"79",
          2852 => x"82",
          2853 => x"ff",
          2854 => x"87",
          2855 => x"ec",
          2856 => x"02",
          2857 => x"e3",
          2858 => x"57",
          2859 => x"30",
          2860 => x"73",
          2861 => x"59",
          2862 => x"77",
          2863 => x"83",
          2864 => x"74",
          2865 => x"81",
          2866 => x"55",
          2867 => x"81",
          2868 => x"53",
          2869 => x"3d",
          2870 => x"81",
          2871 => x"82",
          2872 => x"57",
          2873 => x"08",
          2874 => x"d5",
          2875 => x"c0",
          2876 => x"82",
          2877 => x"59",
          2878 => x"05",
          2879 => x"53",
          2880 => x"51",
          2881 => x"3f",
          2882 => x"08",
          2883 => x"e4",
          2884 => x"7a",
          2885 => x"2e",
          2886 => x"19",
          2887 => x"59",
          2888 => x"3d",
          2889 => x"81",
          2890 => x"76",
          2891 => x"07",
          2892 => x"30",
          2893 => x"72",
          2894 => x"51",
          2895 => x"2e",
          2896 => x"b6",
          2897 => x"c0",
          2898 => x"52",
          2899 => x"92",
          2900 => x"75",
          2901 => x"0c",
          2902 => x"04",
          2903 => x"7c",
          2904 => x"b7",
          2905 => x"59",
          2906 => x"53",
          2907 => x"51",
          2908 => x"82",
          2909 => x"a8",
          2910 => x"2e",
          2911 => x"81",
          2912 => x"9c",
          2913 => x"c4",
          2914 => x"60",
          2915 => x"e4",
          2916 => x"7e",
          2917 => x"82",
          2918 => x"58",
          2919 => x"04",
          2920 => x"e4",
          2921 => x"0d",
          2922 => x"0d",
          2923 => x"02",
          2924 => x"cf",
          2925 => x"73",
          2926 => x"5f",
          2927 => x"5e",
          2928 => x"82",
          2929 => x"ff",
          2930 => x"82",
          2931 => x"ff",
          2932 => x"80",
          2933 => x"27",
          2934 => x"7b",
          2935 => x"38",
          2936 => x"a7",
          2937 => x"39",
          2938 => x"72",
          2939 => x"38",
          2940 => x"82",
          2941 => x"ff",
          2942 => x"89",
          2943 => x"94",
          2944 => x"d4",
          2945 => x"55",
          2946 => x"74",
          2947 => x"7a",
          2948 => x"72",
          2949 => x"b6",
          2950 => x"b7",
          2951 => x"39",
          2952 => x"51",
          2953 => x"3f",
          2954 => x"a1",
          2955 => x"53",
          2956 => x"8e",
          2957 => x"52",
          2958 => x"51",
          2959 => x"3f",
          2960 => x"b7",
          2961 => x"b7",
          2962 => x"15",
          2963 => x"c8",
          2964 => x"51",
          2965 => x"fe",
          2966 => x"b7",
          2967 => x"b6",
          2968 => x"55",
          2969 => x"80",
          2970 => x"18",
          2971 => x"53",
          2972 => x"7a",
          2973 => x"81",
          2974 => x"9f",
          2975 => x"38",
          2976 => x"73",
          2977 => x"ff",
          2978 => x"72",
          2979 => x"38",
          2980 => x"26",
          2981 => x"f1",
          2982 => x"73",
          2983 => x"82",
          2984 => x"52",
          2985 => x"8a",
          2986 => x"55",
          2987 => x"82",
          2988 => x"d2",
          2989 => x"18",
          2990 => x"58",
          2991 => x"82",
          2992 => x"98",
          2993 => x"2c",
          2994 => x"a0",
          2995 => x"06",
          2996 => x"f4",
          2997 => x"e4",
          2998 => x"70",
          2999 => x"a0",
          3000 => x"72",
          3001 => x"30",
          3002 => x"73",
          3003 => x"51",
          3004 => x"57",
          3005 => x"73",
          3006 => x"76",
          3007 => x"81",
          3008 => x"80",
          3009 => x"7c",
          3010 => x"78",
          3011 => x"38",
          3012 => x"82",
          3013 => x"8f",
          3014 => x"fc",
          3015 => x"9b",
          3016 => x"b7",
          3017 => x"b7",
          3018 => x"ff",
          3019 => x"82",
          3020 => x"51",
          3021 => x"82",
          3022 => x"82",
          3023 => x"82",
          3024 => x"52",
          3025 => x"51",
          3026 => x"3f",
          3027 => x"84",
          3028 => x"3f",
          3029 => x"04",
          3030 => x"87",
          3031 => x"08",
          3032 => x"3f",
          3033 => x"cd",
          3034 => x"f0",
          3035 => x"3f",
          3036 => x"c1",
          3037 => x"2a",
          3038 => x"51",
          3039 => x"2e",
          3040 => x"51",
          3041 => x"82",
          3042 => x"99",
          3043 => x"51",
          3044 => x"72",
          3045 => x"81",
          3046 => x"71",
          3047 => x"38",
          3048 => x"91",
          3049 => x"98",
          3050 => x"3f",
          3051 => x"85",
          3052 => x"2a",
          3053 => x"51",
          3054 => x"2e",
          3055 => x"51",
          3056 => x"82",
          3057 => x"99",
          3058 => x"51",
          3059 => x"72",
          3060 => x"81",
          3061 => x"71",
          3062 => x"38",
          3063 => x"d5",
          3064 => x"bc",
          3065 => x"3f",
          3066 => x"c9",
          3067 => x"2a",
          3068 => x"51",
          3069 => x"2e",
          3070 => x"51",
          3071 => x"82",
          3072 => x"98",
          3073 => x"51",
          3074 => x"72",
          3075 => x"81",
          3076 => x"71",
          3077 => x"38",
          3078 => x"99",
          3079 => x"e4",
          3080 => x"3f",
          3081 => x"8d",
          3082 => x"2a",
          3083 => x"51",
          3084 => x"2e",
          3085 => x"51",
          3086 => x"82",
          3087 => x"98",
          3088 => x"51",
          3089 => x"72",
          3090 => x"81",
          3091 => x"71",
          3092 => x"38",
          3093 => x"dd",
          3094 => x"8c",
          3095 => x"3f",
          3096 => x"d1",
          3097 => x"3f",
          3098 => x"04",
          3099 => x"77",
          3100 => x"a3",
          3101 => x"55",
          3102 => x"52",
          3103 => x"91",
          3104 => x"82",
          3105 => x"54",
          3106 => x"81",
          3107 => x"c8",
          3108 => x"f4",
          3109 => x"bf",
          3110 => x"e4",
          3111 => x"82",
          3112 => x"07",
          3113 => x"71",
          3114 => x"54",
          3115 => x"82",
          3116 => x"0b",
          3117 => x"d8",
          3118 => x"81",
          3119 => x"06",
          3120 => x"ec",
          3121 => x"52",
          3122 => x"c6",
          3123 => x"d5",
          3124 => x"2e",
          3125 => x"d5",
          3126 => x"ce",
          3127 => x"39",
          3128 => x"51",
          3129 => x"3f",
          3130 => x"0b",
          3131 => x"34",
          3132 => x"d0",
          3133 => x"73",
          3134 => x"81",
          3135 => x"82",
          3136 => x"74",
          3137 => x"a9",
          3138 => x"0b",
          3139 => x"0c",
          3140 => x"04",
          3141 => x"80",
          3142 => x"ff",
          3143 => x"f0",
          3144 => x"52",
          3145 => x"c7",
          3146 => x"d5",
          3147 => x"ff",
          3148 => x"7e",
          3149 => x"06",
          3150 => x"3d",
          3151 => x"82",
          3152 => x"78",
          3153 => x"3f",
          3154 => x"52",
          3155 => x"51",
          3156 => x"3f",
          3157 => x"08",
          3158 => x"38",
          3159 => x"51",
          3160 => x"81",
          3161 => x"82",
          3162 => x"ff",
          3163 => x"97",
          3164 => x"5a",
          3165 => x"79",
          3166 => x"3f",
          3167 => x"84",
          3168 => x"c4",
          3169 => x"e4",
          3170 => x"70",
          3171 => x"59",
          3172 => x"2e",
          3173 => x"78",
          3174 => x"b2",
          3175 => x"2e",
          3176 => x"78",
          3177 => x"38",
          3178 => x"ff",
          3179 => x"bc",
          3180 => x"38",
          3181 => x"78",
          3182 => x"83",
          3183 => x"80",
          3184 => x"cd",
          3185 => x"2e",
          3186 => x"8a",
          3187 => x"80",
          3188 => x"db",
          3189 => x"f9",
          3190 => x"78",
          3191 => x"88",
          3192 => x"80",
          3193 => x"a3",
          3194 => x"39",
          3195 => x"2e",
          3196 => x"78",
          3197 => x"8b",
          3198 => x"82",
          3199 => x"38",
          3200 => x"78",
          3201 => x"89",
          3202 => x"80",
          3203 => x"ff",
          3204 => x"ff",
          3205 => x"ec",
          3206 => x"d5",
          3207 => x"2e",
          3208 => x"b5",
          3209 => x"11",
          3210 => x"05",
          3211 => x"3f",
          3212 => x"08",
          3213 => x"af",
          3214 => x"fe",
          3215 => x"ff",
          3216 => x"ec",
          3217 => x"d5",
          3218 => x"38",
          3219 => x"08",
          3220 => x"a4",
          3221 => x"80",
          3222 => x"5c",
          3223 => x"27",
          3224 => x"62",
          3225 => x"70",
          3226 => x"0c",
          3227 => x"f5",
          3228 => x"39",
          3229 => x"80",
          3230 => x"84",
          3231 => x"f7",
          3232 => x"e4",
          3233 => x"fd",
          3234 => x"3d",
          3235 => x"53",
          3236 => x"51",
          3237 => x"82",
          3238 => x"80",
          3239 => x"38",
          3240 => x"f8",
          3241 => x"84",
          3242 => x"cb",
          3243 => x"e4",
          3244 => x"fd",
          3245 => x"ba",
          3246 => x"ae",
          3247 => x"5a",
          3248 => x"81",
          3249 => x"59",
          3250 => x"05",
          3251 => x"34",
          3252 => x"43",
          3253 => x"3d",
          3254 => x"53",
          3255 => x"51",
          3256 => x"82",
          3257 => x"80",
          3258 => x"38",
          3259 => x"fc",
          3260 => x"84",
          3261 => x"ff",
          3262 => x"e4",
          3263 => x"fc",
          3264 => x"3d",
          3265 => x"53",
          3266 => x"51",
          3267 => x"82",
          3268 => x"80",
          3269 => x"38",
          3270 => x"51",
          3271 => x"3f",
          3272 => x"64",
          3273 => x"62",
          3274 => x"33",
          3275 => x"78",
          3276 => x"38",
          3277 => x"54",
          3278 => x"79",
          3279 => x"d0",
          3280 => x"94",
          3281 => x"63",
          3282 => x"5a",
          3283 => x"51",
          3284 => x"fc",
          3285 => x"3d",
          3286 => x"53",
          3287 => x"51",
          3288 => x"82",
          3289 => x"80",
          3290 => x"d4",
          3291 => x"78",
          3292 => x"38",
          3293 => x"08",
          3294 => x"39",
          3295 => x"33",
          3296 => x"2e",
          3297 => x"d4",
          3298 => x"bc",
          3299 => x"ca",
          3300 => x"80",
          3301 => x"82",
          3302 => x"45",
          3303 => x"d4",
          3304 => x"78",
          3305 => x"38",
          3306 => x"08",
          3307 => x"82",
          3308 => x"59",
          3309 => x"88",
          3310 => x"a0",
          3311 => x"39",
          3312 => x"08",
          3313 => x"45",
          3314 => x"fc",
          3315 => x"84",
          3316 => x"a3",
          3317 => x"e4",
          3318 => x"38",
          3319 => x"33",
          3320 => x"2e",
          3321 => x"d4",
          3322 => x"80",
          3323 => x"d4",
          3324 => x"78",
          3325 => x"38",
          3326 => x"08",
          3327 => x"82",
          3328 => x"59",
          3329 => x"88",
          3330 => x"94",
          3331 => x"39",
          3332 => x"33",
          3333 => x"2e",
          3334 => x"d4",
          3335 => x"99",
          3336 => x"c6",
          3337 => x"80",
          3338 => x"82",
          3339 => x"44",
          3340 => x"d4",
          3341 => x"05",
          3342 => x"fe",
          3343 => x"ff",
          3344 => x"e8",
          3345 => x"d5",
          3346 => x"2e",
          3347 => x"63",
          3348 => x"88",
          3349 => x"81",
          3350 => x"32",
          3351 => x"72",
          3352 => x"70",
          3353 => x"51",
          3354 => x"80",
          3355 => x"7a",
          3356 => x"38",
          3357 => x"ba",
          3358 => x"e7",
          3359 => x"64",
          3360 => x"63",
          3361 => x"f2",
          3362 => x"ba",
          3363 => x"b1",
          3364 => x"ff",
          3365 => x"ff",
          3366 => x"e7",
          3367 => x"d5",
          3368 => x"2e",
          3369 => x"b5",
          3370 => x"11",
          3371 => x"05",
          3372 => x"3f",
          3373 => x"08",
          3374 => x"38",
          3375 => x"80",
          3376 => x"79",
          3377 => x"05",
          3378 => x"fe",
          3379 => x"ff",
          3380 => x"e7",
          3381 => x"d5",
          3382 => x"38",
          3383 => x"64",
          3384 => x"52",
          3385 => x"51",
          3386 => x"3f",
          3387 => x"08",
          3388 => x"52",
          3389 => x"aa",
          3390 => x"46",
          3391 => x"78",
          3392 => x"e3",
          3393 => x"27",
          3394 => x"3d",
          3395 => x"53",
          3396 => x"51",
          3397 => x"82",
          3398 => x"80",
          3399 => x"64",
          3400 => x"cf",
          3401 => x"34",
          3402 => x"45",
          3403 => x"82",
          3404 => x"c5",
          3405 => x"a7",
          3406 => x"fe",
          3407 => x"ff",
          3408 => x"e0",
          3409 => x"d5",
          3410 => x"2e",
          3411 => x"b5",
          3412 => x"11",
          3413 => x"05",
          3414 => x"3f",
          3415 => x"08",
          3416 => x"38",
          3417 => x"80",
          3418 => x"79",
          3419 => x"5b",
          3420 => x"b5",
          3421 => x"11",
          3422 => x"05",
          3423 => x"3f",
          3424 => x"08",
          3425 => x"df",
          3426 => x"22",
          3427 => x"bb",
          3428 => x"a8",
          3429 => x"f1",
          3430 => x"80",
          3431 => x"51",
          3432 => x"3f",
          3433 => x"33",
          3434 => x"2e",
          3435 => x"78",
          3436 => x"38",
          3437 => x"42",
          3438 => x"3d",
          3439 => x"53",
          3440 => x"51",
          3441 => x"82",
          3442 => x"80",
          3443 => x"61",
          3444 => x"c2",
          3445 => x"70",
          3446 => x"23",
          3447 => x"a9",
          3448 => x"90",
          3449 => x"3f",
          3450 => x"b5",
          3451 => x"11",
          3452 => x"05",
          3453 => x"3f",
          3454 => x"08",
          3455 => x"e7",
          3456 => x"fe",
          3457 => x"ff",
          3458 => x"df",
          3459 => x"d5",
          3460 => x"2e",
          3461 => x"61",
          3462 => x"61",
          3463 => x"b5",
          3464 => x"11",
          3465 => x"05",
          3466 => x"3f",
          3467 => x"08",
          3468 => x"b3",
          3469 => x"08",
          3470 => x"bb",
          3471 => x"a7",
          3472 => x"f1",
          3473 => x"80",
          3474 => x"51",
          3475 => x"3f",
          3476 => x"33",
          3477 => x"2e",
          3478 => x"9f",
          3479 => x"38",
          3480 => x"f0",
          3481 => x"84",
          3482 => x"ba",
          3483 => x"e4",
          3484 => x"8d",
          3485 => x"71",
          3486 => x"84",
          3487 => x"b5",
          3488 => x"90",
          3489 => x"3f",
          3490 => x"b5",
          3491 => x"11",
          3492 => x"05",
          3493 => x"3f",
          3494 => x"08",
          3495 => x"c7",
          3496 => x"82",
          3497 => x"ff",
          3498 => x"64",
          3499 => x"b5",
          3500 => x"11",
          3501 => x"05",
          3502 => x"3f",
          3503 => x"08",
          3504 => x"a3",
          3505 => x"82",
          3506 => x"ff",
          3507 => x"64",
          3508 => x"82",
          3509 => x"80",
          3510 => x"38",
          3511 => x"08",
          3512 => x"e8",
          3513 => x"f0",
          3514 => x"39",
          3515 => x"51",
          3516 => x"ff",
          3517 => x"f4",
          3518 => x"bc",
          3519 => x"e3",
          3520 => x"ff",
          3521 => x"e2",
          3522 => x"39",
          3523 => x"59",
          3524 => x"f4",
          3525 => x"f8",
          3526 => x"d3",
          3527 => x"d5",
          3528 => x"82",
          3529 => x"80",
          3530 => x"38",
          3531 => x"08",
          3532 => x"ff",
          3533 => x"83",
          3534 => x"d5",
          3535 => x"7f",
          3536 => x"78",
          3537 => x"d2",
          3538 => x"e4",
          3539 => x"b5",
          3540 => x"e4",
          3541 => x"81",
          3542 => x"5b",
          3543 => x"b2",
          3544 => x"24",
          3545 => x"81",
          3546 => x"80",
          3547 => x"83",
          3548 => x"80",
          3549 => x"bc",
          3550 => x"55",
          3551 => x"54",
          3552 => x"bc",
          3553 => x"3d",
          3554 => x"51",
          3555 => x"3f",
          3556 => x"52",
          3557 => x"b0",
          3558 => x"d7",
          3559 => x"7b",
          3560 => x"b8",
          3561 => x"82",
          3562 => x"b5",
          3563 => x"05",
          3564 => x"8c",
          3565 => x"7b",
          3566 => x"82",
          3567 => x"b5",
          3568 => x"05",
          3569 => x"f8",
          3570 => x"80",
          3571 => x"94",
          3572 => x"65",
          3573 => x"84",
          3574 => x"84",
          3575 => x"b5",
          3576 => x"05",
          3577 => x"3f",
          3578 => x"08",
          3579 => x"08",
          3580 => x"70",
          3581 => x"25",
          3582 => x"5f",
          3583 => x"83",
          3584 => x"81",
          3585 => x"06",
          3586 => x"2e",
          3587 => x"1b",
          3588 => x"06",
          3589 => x"fe",
          3590 => x"81",
          3591 => x"32",
          3592 => x"89",
          3593 => x"2e",
          3594 => x"89",
          3595 => x"e0",
          3596 => x"af",
          3597 => x"b1",
          3598 => x"ab",
          3599 => x"f0",
          3600 => x"9f",
          3601 => x"39",
          3602 => x"80",
          3603 => x"94",
          3604 => x"94",
          3605 => x"54",
          3606 => x"80",
          3607 => x"d7",
          3608 => x"d5",
          3609 => x"2b",
          3610 => x"53",
          3611 => x"52",
          3612 => x"ba",
          3613 => x"d5",
          3614 => x"75",
          3615 => x"94",
          3616 => x"54",
          3617 => x"80",
          3618 => x"d7",
          3619 => x"d5",
          3620 => x"2b",
          3621 => x"53",
          3622 => x"52",
          3623 => x"8e",
          3624 => x"d5",
          3625 => x"75",
          3626 => x"83",
          3627 => x"94",
          3628 => x"80",
          3629 => x"c0",
          3630 => x"80",
          3631 => x"80",
          3632 => x"83",
          3633 => x"99",
          3634 => x"5c",
          3635 => x"0b",
          3636 => x"88",
          3637 => x"72",
          3638 => x"c8",
          3639 => x"be",
          3640 => x"3f",
          3641 => x"51",
          3642 => x"3f",
          3643 => x"51",
          3644 => x"3f",
          3645 => x"51",
          3646 => x"81",
          3647 => x"3f",
          3648 => x"80",
          3649 => x"0d",
          3650 => x"53",
          3651 => x"52",
          3652 => x"82",
          3653 => x"81",
          3654 => x"07",
          3655 => x"52",
          3656 => x"e8",
          3657 => x"d5",
          3658 => x"3d",
          3659 => x"3d",
          3660 => x"08",
          3661 => x"73",
          3662 => x"74",
          3663 => x"38",
          3664 => x"70",
          3665 => x"81",
          3666 => x"81",
          3667 => x"39",
          3668 => x"70",
          3669 => x"81",
          3670 => x"81",
          3671 => x"54",
          3672 => x"81",
          3673 => x"06",
          3674 => x"39",
          3675 => x"80",
          3676 => x"54",
          3677 => x"83",
          3678 => x"70",
          3679 => x"38",
          3680 => x"98",
          3681 => x"52",
          3682 => x"52",
          3683 => x"2e",
          3684 => x"54",
          3685 => x"84",
          3686 => x"38",
          3687 => x"52",
          3688 => x"2e",
          3689 => x"83",
          3690 => x"70",
          3691 => x"30",
          3692 => x"76",
          3693 => x"51",
          3694 => x"88",
          3695 => x"70",
          3696 => x"34",
          3697 => x"72",
          3698 => x"d5",
          3699 => x"3d",
          3700 => x"3d",
          3701 => x"72",
          3702 => x"91",
          3703 => x"fc",
          3704 => x"51",
          3705 => x"82",
          3706 => x"85",
          3707 => x"83",
          3708 => x"72",
          3709 => x"0c",
          3710 => x"04",
          3711 => x"76",
          3712 => x"ff",
          3713 => x"81",
          3714 => x"26",
          3715 => x"83",
          3716 => x"05",
          3717 => x"70",
          3718 => x"8a",
          3719 => x"33",
          3720 => x"70",
          3721 => x"fe",
          3722 => x"33",
          3723 => x"70",
          3724 => x"f2",
          3725 => x"33",
          3726 => x"70",
          3727 => x"e6",
          3728 => x"22",
          3729 => x"74",
          3730 => x"80",
          3731 => x"13",
          3732 => x"52",
          3733 => x"26",
          3734 => x"81",
          3735 => x"98",
          3736 => x"22",
          3737 => x"bc",
          3738 => x"33",
          3739 => x"b8",
          3740 => x"33",
          3741 => x"b4",
          3742 => x"33",
          3743 => x"b0",
          3744 => x"33",
          3745 => x"ac",
          3746 => x"33",
          3747 => x"a8",
          3748 => x"c0",
          3749 => x"73",
          3750 => x"a0",
          3751 => x"87",
          3752 => x"0c",
          3753 => x"82",
          3754 => x"86",
          3755 => x"f3",
          3756 => x"5b",
          3757 => x"9c",
          3758 => x"0c",
          3759 => x"bc",
          3760 => x"7b",
          3761 => x"98",
          3762 => x"79",
          3763 => x"87",
          3764 => x"08",
          3765 => x"1c",
          3766 => x"98",
          3767 => x"79",
          3768 => x"87",
          3769 => x"08",
          3770 => x"1c",
          3771 => x"98",
          3772 => x"79",
          3773 => x"87",
          3774 => x"08",
          3775 => x"1c",
          3776 => x"98",
          3777 => x"79",
          3778 => x"80",
          3779 => x"83",
          3780 => x"59",
          3781 => x"ff",
          3782 => x"1b",
          3783 => x"1b",
          3784 => x"1b",
          3785 => x"1b",
          3786 => x"1b",
          3787 => x"83",
          3788 => x"52",
          3789 => x"51",
          3790 => x"3f",
          3791 => x"04",
          3792 => x"02",
          3793 => x"82",
          3794 => x"70",
          3795 => x"58",
          3796 => x"c0",
          3797 => x"75",
          3798 => x"38",
          3799 => x"94",
          3800 => x"70",
          3801 => x"81",
          3802 => x"52",
          3803 => x"8c",
          3804 => x"2a",
          3805 => x"51",
          3806 => x"38",
          3807 => x"70",
          3808 => x"51",
          3809 => x"8d",
          3810 => x"2a",
          3811 => x"51",
          3812 => x"be",
          3813 => x"ff",
          3814 => x"c0",
          3815 => x"70",
          3816 => x"38",
          3817 => x"90",
          3818 => x"0c",
          3819 => x"e4",
          3820 => x"0d",
          3821 => x"0d",
          3822 => x"33",
          3823 => x"9f",
          3824 => x"52",
          3825 => x"fc",
          3826 => x"0d",
          3827 => x"0d",
          3828 => x"33",
          3829 => x"2e",
          3830 => x"87",
          3831 => x"8d",
          3832 => x"82",
          3833 => x"70",
          3834 => x"58",
          3835 => x"94",
          3836 => x"80",
          3837 => x"87",
          3838 => x"53",
          3839 => x"96",
          3840 => x"06",
          3841 => x"72",
          3842 => x"38",
          3843 => x"70",
          3844 => x"53",
          3845 => x"74",
          3846 => x"81",
          3847 => x"72",
          3848 => x"38",
          3849 => x"70",
          3850 => x"53",
          3851 => x"38",
          3852 => x"06",
          3853 => x"94",
          3854 => x"80",
          3855 => x"87",
          3856 => x"54",
          3857 => x"80",
          3858 => x"e4",
          3859 => x"0d",
          3860 => x"0d",
          3861 => x"74",
          3862 => x"ff",
          3863 => x"57",
          3864 => x"80",
          3865 => x"81",
          3866 => x"15",
          3867 => x"33",
          3868 => x"06",
          3869 => x"58",
          3870 => x"84",
          3871 => x"2e",
          3872 => x"c0",
          3873 => x"70",
          3874 => x"2a",
          3875 => x"53",
          3876 => x"80",
          3877 => x"71",
          3878 => x"81",
          3879 => x"70",
          3880 => x"81",
          3881 => x"06",
          3882 => x"80",
          3883 => x"71",
          3884 => x"81",
          3885 => x"70",
          3886 => x"74",
          3887 => x"51",
          3888 => x"80",
          3889 => x"2e",
          3890 => x"c0",
          3891 => x"77",
          3892 => x"17",
          3893 => x"81",
          3894 => x"53",
          3895 => x"86",
          3896 => x"d5",
          3897 => x"3d",
          3898 => x"3d",
          3899 => x"fc",
          3900 => x"ff",
          3901 => x"87",
          3902 => x"51",
          3903 => x"86",
          3904 => x"94",
          3905 => x"08",
          3906 => x"70",
          3907 => x"51",
          3908 => x"2e",
          3909 => x"81",
          3910 => x"87",
          3911 => x"52",
          3912 => x"86",
          3913 => x"94",
          3914 => x"08",
          3915 => x"06",
          3916 => x"0c",
          3917 => x"0d",
          3918 => x"3f",
          3919 => x"08",
          3920 => x"82",
          3921 => x"04",
          3922 => x"82",
          3923 => x"70",
          3924 => x"52",
          3925 => x"94",
          3926 => x"80",
          3927 => x"87",
          3928 => x"52",
          3929 => x"82",
          3930 => x"06",
          3931 => x"ff",
          3932 => x"2e",
          3933 => x"81",
          3934 => x"87",
          3935 => x"52",
          3936 => x"86",
          3937 => x"94",
          3938 => x"08",
          3939 => x"70",
          3940 => x"53",
          3941 => x"d5",
          3942 => x"3d",
          3943 => x"3d",
          3944 => x"9e",
          3945 => x"9c",
          3946 => x"51",
          3947 => x"2e",
          3948 => x"87",
          3949 => x"08",
          3950 => x"0c",
          3951 => x"a8",
          3952 => x"84",
          3953 => x"9e",
          3954 => x"d4",
          3955 => x"c0",
          3956 => x"82",
          3957 => x"87",
          3958 => x"08",
          3959 => x"0c",
          3960 => x"a0",
          3961 => x"94",
          3962 => x"9e",
          3963 => x"d4",
          3964 => x"c0",
          3965 => x"82",
          3966 => x"87",
          3967 => x"08",
          3968 => x"0c",
          3969 => x"b8",
          3970 => x"a4",
          3971 => x"9e",
          3972 => x"d4",
          3973 => x"c0",
          3974 => x"82",
          3975 => x"87",
          3976 => x"08",
          3977 => x"0c",
          3978 => x"80",
          3979 => x"82",
          3980 => x"87",
          3981 => x"08",
          3982 => x"0c",
          3983 => x"88",
          3984 => x"bc",
          3985 => x"9e",
          3986 => x"d4",
          3987 => x"0b",
          3988 => x"34",
          3989 => x"c0",
          3990 => x"70",
          3991 => x"06",
          3992 => x"70",
          3993 => x"38",
          3994 => x"82",
          3995 => x"80",
          3996 => x"9e",
          3997 => x"88",
          3998 => x"51",
          3999 => x"80",
          4000 => x"81",
          4001 => x"d4",
          4002 => x"0b",
          4003 => x"90",
          4004 => x"80",
          4005 => x"52",
          4006 => x"2e",
          4007 => x"52",
          4008 => x"c7",
          4009 => x"87",
          4010 => x"08",
          4011 => x"80",
          4012 => x"52",
          4013 => x"83",
          4014 => x"71",
          4015 => x"34",
          4016 => x"c0",
          4017 => x"70",
          4018 => x"06",
          4019 => x"70",
          4020 => x"38",
          4021 => x"82",
          4022 => x"80",
          4023 => x"9e",
          4024 => x"90",
          4025 => x"51",
          4026 => x"80",
          4027 => x"81",
          4028 => x"d4",
          4029 => x"0b",
          4030 => x"90",
          4031 => x"80",
          4032 => x"52",
          4033 => x"2e",
          4034 => x"52",
          4035 => x"cb",
          4036 => x"87",
          4037 => x"08",
          4038 => x"80",
          4039 => x"52",
          4040 => x"83",
          4041 => x"71",
          4042 => x"34",
          4043 => x"c0",
          4044 => x"70",
          4045 => x"06",
          4046 => x"70",
          4047 => x"38",
          4048 => x"82",
          4049 => x"80",
          4050 => x"9e",
          4051 => x"80",
          4052 => x"51",
          4053 => x"80",
          4054 => x"81",
          4055 => x"d4",
          4056 => x"0b",
          4057 => x"90",
          4058 => x"80",
          4059 => x"52",
          4060 => x"83",
          4061 => x"71",
          4062 => x"34",
          4063 => x"90",
          4064 => x"80",
          4065 => x"2a",
          4066 => x"70",
          4067 => x"34",
          4068 => x"c0",
          4069 => x"70",
          4070 => x"51",
          4071 => x"80",
          4072 => x"81",
          4073 => x"d4",
          4074 => x"c0",
          4075 => x"70",
          4076 => x"70",
          4077 => x"51",
          4078 => x"d4",
          4079 => x"0b",
          4080 => x"90",
          4081 => x"06",
          4082 => x"70",
          4083 => x"38",
          4084 => x"82",
          4085 => x"87",
          4086 => x"08",
          4087 => x"51",
          4088 => x"d4",
          4089 => x"3d",
          4090 => x"3d",
          4091 => x"d8",
          4092 => x"e4",
          4093 => x"c4",
          4094 => x"80",
          4095 => x"82",
          4096 => x"ff",
          4097 => x"82",
          4098 => x"ff",
          4099 => x"82",
          4100 => x"54",
          4101 => x"94",
          4102 => x"a0",
          4103 => x"a4",
          4104 => x"52",
          4105 => x"51",
          4106 => x"3f",
          4107 => x"33",
          4108 => x"2e",
          4109 => x"d4",
          4110 => x"d4",
          4111 => x"54",
          4112 => x"b4",
          4113 => x"90",
          4114 => x"c8",
          4115 => x"80",
          4116 => x"82",
          4117 => x"82",
          4118 => x"11",
          4119 => x"be",
          4120 => x"92",
          4121 => x"d4",
          4122 => x"73",
          4123 => x"38",
          4124 => x"08",
          4125 => x"08",
          4126 => x"82",
          4127 => x"ff",
          4128 => x"82",
          4129 => x"54",
          4130 => x"94",
          4131 => x"90",
          4132 => x"94",
          4133 => x"52",
          4134 => x"51",
          4135 => x"3f",
          4136 => x"33",
          4137 => x"2e",
          4138 => x"d4",
          4139 => x"82",
          4140 => x"ff",
          4141 => x"82",
          4142 => x"54",
          4143 => x"8e",
          4144 => x"d4",
          4145 => x"bf",
          4146 => x"92",
          4147 => x"d4",
          4148 => x"73",
          4149 => x"38",
          4150 => x"33",
          4151 => x"e4",
          4152 => x"f4",
          4153 => x"c5",
          4154 => x"80",
          4155 => x"82",
          4156 => x"ff",
          4157 => x"82",
          4158 => x"54",
          4159 => x"89",
          4160 => x"98",
          4161 => x"db",
          4162 => x"cc",
          4163 => x"80",
          4164 => x"82",
          4165 => x"ff",
          4166 => x"82",
          4167 => x"54",
          4168 => x"89",
          4169 => x"b0",
          4170 => x"b7",
          4171 => x"ce",
          4172 => x"80",
          4173 => x"82",
          4174 => x"ff",
          4175 => x"82",
          4176 => x"ff",
          4177 => x"82",
          4178 => x"52",
          4179 => x"51",
          4180 => x"3f",
          4181 => x"08",
          4182 => x"f4",
          4183 => x"f8",
          4184 => x"b0",
          4185 => x"c1",
          4186 => x"90",
          4187 => x"c1",
          4188 => x"ac",
          4189 => x"d4",
          4190 => x"82",
          4191 => x"ff",
          4192 => x"82",
          4193 => x"56",
          4194 => x"52",
          4195 => x"9e",
          4196 => x"e4",
          4197 => x"c0",
          4198 => x"31",
          4199 => x"d5",
          4200 => x"82",
          4201 => x"ff",
          4202 => x"82",
          4203 => x"54",
          4204 => x"a9",
          4205 => x"bc",
          4206 => x"84",
          4207 => x"51",
          4208 => x"82",
          4209 => x"bd",
          4210 => x"76",
          4211 => x"54",
          4212 => x"08",
          4213 => x"a0",
          4214 => x"fc",
          4215 => x"c6",
          4216 => x"80",
          4217 => x"82",
          4218 => x"56",
          4219 => x"52",
          4220 => x"ba",
          4221 => x"e4",
          4222 => x"c0",
          4223 => x"31",
          4224 => x"d5",
          4225 => x"82",
          4226 => x"ff",
          4227 => x"8a",
          4228 => x"f1",
          4229 => x"0d",
          4230 => x"0d",
          4231 => x"33",
          4232 => x"71",
          4233 => x"38",
          4234 => x"82",
          4235 => x"52",
          4236 => x"82",
          4237 => x"9d",
          4238 => x"80",
          4239 => x"82",
          4240 => x"91",
          4241 => x"90",
          4242 => x"82",
          4243 => x"85",
          4244 => x"9c",
          4245 => x"80",
          4246 => x"0d",
          4247 => x"80",
          4248 => x"0b",
          4249 => x"84",
          4250 => x"d4",
          4251 => x"c0",
          4252 => x"04",
          4253 => x"76",
          4254 => x"98",
          4255 => x"2b",
          4256 => x"72",
          4257 => x"82",
          4258 => x"51",
          4259 => x"80",
          4260 => x"a8",
          4261 => x"53",
          4262 => x"9c",
          4263 => x"a4",
          4264 => x"02",
          4265 => x"05",
          4266 => x"52",
          4267 => x"72",
          4268 => x"06",
          4269 => x"53",
          4270 => x"e4",
          4271 => x"0d",
          4272 => x"0d",
          4273 => x"05",
          4274 => x"71",
          4275 => x"54",
          4276 => x"b1",
          4277 => x"c8",
          4278 => x"51",
          4279 => x"3f",
          4280 => x"08",
          4281 => x"ff",
          4282 => x"82",
          4283 => x"52",
          4284 => x"ad",
          4285 => x"33",
          4286 => x"72",
          4287 => x"81",
          4288 => x"cc",
          4289 => x"ff",
          4290 => x"74",
          4291 => x"3d",
          4292 => x"3d",
          4293 => x"84",
          4294 => x"33",
          4295 => x"bb",
          4296 => x"d5",
          4297 => x"84",
          4298 => x"dc",
          4299 => x"51",
          4300 => x"58",
          4301 => x"2e",
          4302 => x"51",
          4303 => x"82",
          4304 => x"70",
          4305 => x"d4",
          4306 => x"19",
          4307 => x"56",
          4308 => x"3f",
          4309 => x"08",
          4310 => x"d5",
          4311 => x"84",
          4312 => x"dc",
          4313 => x"51",
          4314 => x"80",
          4315 => x"75",
          4316 => x"74",
          4317 => x"ed",
          4318 => x"b4",
          4319 => x"55",
          4320 => x"b4",
          4321 => x"ff",
          4322 => x"75",
          4323 => x"80",
          4324 => x"b4",
          4325 => x"2e",
          4326 => x"d5",
          4327 => x"75",
          4328 => x"38",
          4329 => x"33",
          4330 => x"38",
          4331 => x"05",
          4332 => x"78",
          4333 => x"80",
          4334 => x"82",
          4335 => x"52",
          4336 => x"a2",
          4337 => x"d5",
          4338 => x"80",
          4339 => x"8c",
          4340 => x"fd",
          4341 => x"d4",
          4342 => x"54",
          4343 => x"71",
          4344 => x"38",
          4345 => x"d1",
          4346 => x"0c",
          4347 => x"14",
          4348 => x"80",
          4349 => x"80",
          4350 => x"b4",
          4351 => x"b0",
          4352 => x"80",
          4353 => x"71",
          4354 => x"cb",
          4355 => x"b0",
          4356 => x"a5",
          4357 => x"82",
          4358 => x"85",
          4359 => x"dc",
          4360 => x"57",
          4361 => x"d5",
          4362 => x"80",
          4363 => x"82",
          4364 => x"80",
          4365 => x"d5",
          4366 => x"80",
          4367 => x"3d",
          4368 => x"81",
          4369 => x"82",
          4370 => x"80",
          4371 => x"75",
          4372 => x"b1",
          4373 => x"e4",
          4374 => x"0b",
          4375 => x"08",
          4376 => x"82",
          4377 => x"ff",
          4378 => x"55",
          4379 => x"34",
          4380 => x"52",
          4381 => x"c6",
          4382 => x"ff",
          4383 => x"74",
          4384 => x"81",
          4385 => x"38",
          4386 => x"04",
          4387 => x"aa",
          4388 => x"3d",
          4389 => x"81",
          4390 => x"80",
          4391 => x"b0",
          4392 => x"f4",
          4393 => x"d5",
          4394 => x"95",
          4395 => x"82",
          4396 => x"54",
          4397 => x"52",
          4398 => x"52",
          4399 => x"c5",
          4400 => x"e4",
          4401 => x"a5",
          4402 => x"ff",
          4403 => x"82",
          4404 => x"81",
          4405 => x"80",
          4406 => x"e4",
          4407 => x"38",
          4408 => x"08",
          4409 => x"17",
          4410 => x"74",
          4411 => x"70",
          4412 => x"07",
          4413 => x"55",
          4414 => x"2e",
          4415 => x"ff",
          4416 => x"d5",
          4417 => x"11",
          4418 => x"80",
          4419 => x"82",
          4420 => x"80",
          4421 => x"82",
          4422 => x"ff",
          4423 => x"78",
          4424 => x"81",
          4425 => x"75",
          4426 => x"ff",
          4427 => x"79",
          4428 => x"d1",
          4429 => x"08",
          4430 => x"e4",
          4431 => x"80",
          4432 => x"d5",
          4433 => x"3d",
          4434 => x"3d",
          4435 => x"71",
          4436 => x"33",
          4437 => x"58",
          4438 => x"09",
          4439 => x"38",
          4440 => x"05",
          4441 => x"27",
          4442 => x"17",
          4443 => x"71",
          4444 => x"55",
          4445 => x"09",
          4446 => x"38",
          4447 => x"ea",
          4448 => x"73",
          4449 => x"d5",
          4450 => x"08",
          4451 => x"b0",
          4452 => x"d5",
          4453 => x"79",
          4454 => x"51",
          4455 => x"3f",
          4456 => x"08",
          4457 => x"84",
          4458 => x"74",
          4459 => x"38",
          4460 => x"88",
          4461 => x"fc",
          4462 => x"39",
          4463 => x"8c",
          4464 => x"53",
          4465 => x"c5",
          4466 => x"d5",
          4467 => x"2e",
          4468 => x"1b",
          4469 => x"77",
          4470 => x"3f",
          4471 => x"08",
          4472 => x"55",
          4473 => x"74",
          4474 => x"81",
          4475 => x"ff",
          4476 => x"82",
          4477 => x"8b",
          4478 => x"73",
          4479 => x"0c",
          4480 => x"04",
          4481 => x"b0",
          4482 => x"3d",
          4483 => x"08",
          4484 => x"80",
          4485 => x"34",
          4486 => x"33",
          4487 => x"08",
          4488 => x"81",
          4489 => x"82",
          4490 => x"55",
          4491 => x"38",
          4492 => x"80",
          4493 => x"38",
          4494 => x"06",
          4495 => x"80",
          4496 => x"38",
          4497 => x"87",
          4498 => x"e4",
          4499 => x"b0",
          4500 => x"e4",
          4501 => x"81",
          4502 => x"53",
          4503 => x"d5",
          4504 => x"80",
          4505 => x"82",
          4506 => x"80",
          4507 => x"82",
          4508 => x"ff",
          4509 => x"80",
          4510 => x"d5",
          4511 => x"82",
          4512 => x"53",
          4513 => x"90",
          4514 => x"54",
          4515 => x"3f",
          4516 => x"08",
          4517 => x"e4",
          4518 => x"09",
          4519 => x"d0",
          4520 => x"e4",
          4521 => x"ae",
          4522 => x"d5",
          4523 => x"80",
          4524 => x"e4",
          4525 => x"38",
          4526 => x"08",
          4527 => x"17",
          4528 => x"74",
          4529 => x"74",
          4530 => x"52",
          4531 => x"c2",
          4532 => x"70",
          4533 => x"5c",
          4534 => x"27",
          4535 => x"5b",
          4536 => x"09",
          4537 => x"97",
          4538 => x"75",
          4539 => x"34",
          4540 => x"82",
          4541 => x"80",
          4542 => x"f9",
          4543 => x"3d",
          4544 => x"3f",
          4545 => x"08",
          4546 => x"98",
          4547 => x"78",
          4548 => x"38",
          4549 => x"06",
          4550 => x"33",
          4551 => x"70",
          4552 => x"ed",
          4553 => x"98",
          4554 => x"2c",
          4555 => x"05",
          4556 => x"82",
          4557 => x"70",
          4558 => x"33",
          4559 => x"51",
          4560 => x"59",
          4561 => x"56",
          4562 => x"80",
          4563 => x"74",
          4564 => x"74",
          4565 => x"29",
          4566 => x"05",
          4567 => x"51",
          4568 => x"24",
          4569 => x"76",
          4570 => x"77",
          4571 => x"3f",
          4572 => x"08",
          4573 => x"54",
          4574 => x"d7",
          4575 => x"ed",
          4576 => x"56",
          4577 => x"81",
          4578 => x"81",
          4579 => x"70",
          4580 => x"81",
          4581 => x"51",
          4582 => x"26",
          4583 => x"53",
          4584 => x"51",
          4585 => x"82",
          4586 => x"81",
          4587 => x"73",
          4588 => x"39",
          4589 => x"80",
          4590 => x"38",
          4591 => x"74",
          4592 => x"34",
          4593 => x"70",
          4594 => x"ed",
          4595 => x"98",
          4596 => x"2c",
          4597 => x"70",
          4598 => x"c3",
          4599 => x"5e",
          4600 => x"57",
          4601 => x"74",
          4602 => x"81",
          4603 => x"38",
          4604 => x"14",
          4605 => x"80",
          4606 => x"a0",
          4607 => x"82",
          4608 => x"92",
          4609 => x"ed",
          4610 => x"82",
          4611 => x"78",
          4612 => x"75",
          4613 => x"54",
          4614 => x"fd",
          4615 => x"84",
          4616 => x"90",
          4617 => x"08",
          4618 => x"a8",
          4619 => x"7e",
          4620 => x"38",
          4621 => x"33",
          4622 => x"27",
          4623 => x"98",
          4624 => x"2c",
          4625 => x"75",
          4626 => x"74",
          4627 => x"33",
          4628 => x"74",
          4629 => x"29",
          4630 => x"05",
          4631 => x"82",
          4632 => x"56",
          4633 => x"39",
          4634 => x"33",
          4635 => x"54",
          4636 => x"a8",
          4637 => x"54",
          4638 => x"74",
          4639 => x"a4",
          4640 => x"7e",
          4641 => x"81",
          4642 => x"82",
          4643 => x"82",
          4644 => x"70",
          4645 => x"29",
          4646 => x"05",
          4647 => x"82",
          4648 => x"5a",
          4649 => x"74",
          4650 => x"38",
          4651 => x"08",
          4652 => x"70",
          4653 => x"ff",
          4654 => x"74",
          4655 => x"29",
          4656 => x"05",
          4657 => x"82",
          4658 => x"56",
          4659 => x"75",
          4660 => x"82",
          4661 => x"70",
          4662 => x"98",
          4663 => x"a4",
          4664 => x"56",
          4665 => x"25",
          4666 => x"82",
          4667 => x"52",
          4668 => x"a1",
          4669 => x"81",
          4670 => x"81",
          4671 => x"70",
          4672 => x"ed",
          4673 => x"51",
          4674 => x"24",
          4675 => x"ee",
          4676 => x"34",
          4677 => x"1b",
          4678 => x"a8",
          4679 => x"82",
          4680 => x"f3",
          4681 => x"fd",
          4682 => x"a8",
          4683 => x"ff",
          4684 => x"73",
          4685 => x"c6",
          4686 => x"a4",
          4687 => x"54",
          4688 => x"a4",
          4689 => x"54",
          4690 => x"a8",
          4691 => x"c8",
          4692 => x"51",
          4693 => x"3f",
          4694 => x"33",
          4695 => x"70",
          4696 => x"ed",
          4697 => x"51",
          4698 => x"74",
          4699 => x"74",
          4700 => x"14",
          4701 => x"82",
          4702 => x"52",
          4703 => x"ff",
          4704 => x"74",
          4705 => x"29",
          4706 => x"05",
          4707 => x"82",
          4708 => x"58",
          4709 => x"75",
          4710 => x"82",
          4711 => x"52",
          4712 => x"a0",
          4713 => x"ed",
          4714 => x"98",
          4715 => x"2c",
          4716 => x"33",
          4717 => x"57",
          4718 => x"fa",
          4719 => x"f1",
          4720 => x"88",
          4721 => x"ea",
          4722 => x"80",
          4723 => x"80",
          4724 => x"98",
          4725 => x"a4",
          4726 => x"55",
          4727 => x"de",
          4728 => x"39",
          4729 => x"33",
          4730 => x"80",
          4731 => x"f1",
          4732 => x"8a",
          4733 => x"ba",
          4734 => x"a4",
          4735 => x"f6",
          4736 => x"d5",
          4737 => x"ff",
          4738 => x"96",
          4739 => x"a4",
          4740 => x"80",
          4741 => x"81",
          4742 => x"79",
          4743 => x"3f",
          4744 => x"7a",
          4745 => x"82",
          4746 => x"80",
          4747 => x"a4",
          4748 => x"d5",
          4749 => x"3d",
          4750 => x"ed",
          4751 => x"73",
          4752 => x"ba",
          4753 => x"c8",
          4754 => x"51",
          4755 => x"3f",
          4756 => x"33",
          4757 => x"73",
          4758 => x"34",
          4759 => x"06",
          4760 => x"82",
          4761 => x"82",
          4762 => x"55",
          4763 => x"2e",
          4764 => x"ff",
          4765 => x"82",
          4766 => x"74",
          4767 => x"98",
          4768 => x"ff",
          4769 => x"55",
          4770 => x"ad",
          4771 => x"54",
          4772 => x"74",
          4773 => x"c8",
          4774 => x"33",
          4775 => x"92",
          4776 => x"80",
          4777 => x"80",
          4778 => x"98",
          4779 => x"a4",
          4780 => x"55",
          4781 => x"d5",
          4782 => x"c8",
          4783 => x"51",
          4784 => x"3f",
          4785 => x"33",
          4786 => x"70",
          4787 => x"ed",
          4788 => x"51",
          4789 => x"74",
          4790 => x"38",
          4791 => x"08",
          4792 => x"ff",
          4793 => x"74",
          4794 => x"29",
          4795 => x"05",
          4796 => x"82",
          4797 => x"58",
          4798 => x"75",
          4799 => x"f7",
          4800 => x"ed",
          4801 => x"81",
          4802 => x"ed",
          4803 => x"56",
          4804 => x"27",
          4805 => x"82",
          4806 => x"52",
          4807 => x"73",
          4808 => x"34",
          4809 => x"33",
          4810 => x"9d",
          4811 => x"ed",
          4812 => x"81",
          4813 => x"ed",
          4814 => x"56",
          4815 => x"26",
          4816 => x"ba",
          4817 => x"a8",
          4818 => x"82",
          4819 => x"ee",
          4820 => x"0b",
          4821 => x"34",
          4822 => x"ed",
          4823 => x"9e",
          4824 => x"38",
          4825 => x"08",
          4826 => x"2e",
          4827 => x"51",
          4828 => x"3f",
          4829 => x"08",
          4830 => x"34",
          4831 => x"08",
          4832 => x"81",
          4833 => x"52",
          4834 => x"a6",
          4835 => x"5b",
          4836 => x"7a",
          4837 => x"d4",
          4838 => x"11",
          4839 => x"74",
          4840 => x"38",
          4841 => x"a4",
          4842 => x"d5",
          4843 => x"ed",
          4844 => x"d5",
          4845 => x"ff",
          4846 => x"53",
          4847 => x"51",
          4848 => x"3f",
          4849 => x"80",
          4850 => x"08",
          4851 => x"2e",
          4852 => x"74",
          4853 => x"ad",
          4854 => x"7a",
          4855 => x"81",
          4856 => x"82",
          4857 => x"55",
          4858 => x"a4",
          4859 => x"ff",
          4860 => x"82",
          4861 => x"82",
          4862 => x"82",
          4863 => x"81",
          4864 => x"05",
          4865 => x"79",
          4866 => x"d9",
          4867 => x"39",
          4868 => x"82",
          4869 => x"70",
          4870 => x"74",
          4871 => x"38",
          4872 => x"a3",
          4873 => x"d5",
          4874 => x"ed",
          4875 => x"d5",
          4876 => x"ff",
          4877 => x"53",
          4878 => x"51",
          4879 => x"3f",
          4880 => x"73",
          4881 => x"5b",
          4882 => x"82",
          4883 => x"74",
          4884 => x"ed",
          4885 => x"ed",
          4886 => x"79",
          4887 => x"3f",
          4888 => x"82",
          4889 => x"70",
          4890 => x"82",
          4891 => x"59",
          4892 => x"77",
          4893 => x"38",
          4894 => x"08",
          4895 => x"54",
          4896 => x"a8",
          4897 => x"70",
          4898 => x"ff",
          4899 => x"f4",
          4900 => x"ed",
          4901 => x"73",
          4902 => x"e2",
          4903 => x"c8",
          4904 => x"51",
          4905 => x"3f",
          4906 => x"33",
          4907 => x"73",
          4908 => x"34",
          4909 => x"f9",
          4910 => x"fa",
          4911 => x"d5",
          4912 => x"80",
          4913 => x"d0",
          4914 => x"80",
          4915 => x"84",
          4916 => x"ff",
          4917 => x"82",
          4918 => x"54",
          4919 => x"74",
          4920 => x"76",
          4921 => x"82",
          4922 => x"54",
          4923 => x"34",
          4924 => x"34",
          4925 => x"08",
          4926 => x"15",
          4927 => x"15",
          4928 => x"d4",
          4929 => x"d0",
          4930 => x"fe",
          4931 => x"70",
          4932 => x"06",
          4933 => x"58",
          4934 => x"74",
          4935 => x"73",
          4936 => x"82",
          4937 => x"70",
          4938 => x"d5",
          4939 => x"f8",
          4940 => x"55",
          4941 => x"34",
          4942 => x"34",
          4943 => x"04",
          4944 => x"73",
          4945 => x"84",
          4946 => x"38",
          4947 => x"2a",
          4948 => x"83",
          4949 => x"51",
          4950 => x"82",
          4951 => x"83",
          4952 => x"f9",
          4953 => x"a6",
          4954 => x"84",
          4955 => x"22",
          4956 => x"d5",
          4957 => x"83",
          4958 => x"74",
          4959 => x"11",
          4960 => x"12",
          4961 => x"2b",
          4962 => x"05",
          4963 => x"71",
          4964 => x"06",
          4965 => x"2a",
          4966 => x"59",
          4967 => x"57",
          4968 => x"71",
          4969 => x"81",
          4970 => x"d5",
          4971 => x"75",
          4972 => x"54",
          4973 => x"34",
          4974 => x"34",
          4975 => x"08",
          4976 => x"33",
          4977 => x"71",
          4978 => x"70",
          4979 => x"ff",
          4980 => x"52",
          4981 => x"05",
          4982 => x"ff",
          4983 => x"2a",
          4984 => x"71",
          4985 => x"72",
          4986 => x"53",
          4987 => x"34",
          4988 => x"08",
          4989 => x"76",
          4990 => x"17",
          4991 => x"0d",
          4992 => x"0d",
          4993 => x"08",
          4994 => x"9e",
          4995 => x"83",
          4996 => x"86",
          4997 => x"12",
          4998 => x"2b",
          4999 => x"07",
          5000 => x"52",
          5001 => x"05",
          5002 => x"85",
          5003 => x"88",
          5004 => x"88",
          5005 => x"56",
          5006 => x"13",
          5007 => x"13",
          5008 => x"d4",
          5009 => x"84",
          5010 => x"12",
          5011 => x"2b",
          5012 => x"07",
          5013 => x"52",
          5014 => x"12",
          5015 => x"33",
          5016 => x"07",
          5017 => x"54",
          5018 => x"70",
          5019 => x"73",
          5020 => x"82",
          5021 => x"13",
          5022 => x"12",
          5023 => x"2b",
          5024 => x"ff",
          5025 => x"88",
          5026 => x"53",
          5027 => x"73",
          5028 => x"14",
          5029 => x"0d",
          5030 => x"0d",
          5031 => x"22",
          5032 => x"08",
          5033 => x"71",
          5034 => x"81",
          5035 => x"88",
          5036 => x"88",
          5037 => x"33",
          5038 => x"71",
          5039 => x"90",
          5040 => x"5f",
          5041 => x"5a",
          5042 => x"54",
          5043 => x"80",
          5044 => x"51",
          5045 => x"82",
          5046 => x"70",
          5047 => x"81",
          5048 => x"8b",
          5049 => x"2b",
          5050 => x"70",
          5051 => x"33",
          5052 => x"07",
          5053 => x"8f",
          5054 => x"51",
          5055 => x"53",
          5056 => x"72",
          5057 => x"2a",
          5058 => x"82",
          5059 => x"83",
          5060 => x"d5",
          5061 => x"16",
          5062 => x"12",
          5063 => x"2b",
          5064 => x"07",
          5065 => x"55",
          5066 => x"33",
          5067 => x"71",
          5068 => x"70",
          5069 => x"06",
          5070 => x"57",
          5071 => x"52",
          5072 => x"71",
          5073 => x"88",
          5074 => x"fb",
          5075 => x"d5",
          5076 => x"84",
          5077 => x"22",
          5078 => x"72",
          5079 => x"33",
          5080 => x"71",
          5081 => x"83",
          5082 => x"5b",
          5083 => x"52",
          5084 => x"33",
          5085 => x"71",
          5086 => x"02",
          5087 => x"05",
          5088 => x"70",
          5089 => x"51",
          5090 => x"71",
          5091 => x"81",
          5092 => x"d5",
          5093 => x"15",
          5094 => x"12",
          5095 => x"2b",
          5096 => x"07",
          5097 => x"52",
          5098 => x"12",
          5099 => x"33",
          5100 => x"07",
          5101 => x"54",
          5102 => x"70",
          5103 => x"72",
          5104 => x"82",
          5105 => x"14",
          5106 => x"83",
          5107 => x"88",
          5108 => x"d5",
          5109 => x"54",
          5110 => x"04",
          5111 => x"7b",
          5112 => x"08",
          5113 => x"70",
          5114 => x"06",
          5115 => x"53",
          5116 => x"82",
          5117 => x"76",
          5118 => x"11",
          5119 => x"83",
          5120 => x"8b",
          5121 => x"2b",
          5122 => x"70",
          5123 => x"33",
          5124 => x"71",
          5125 => x"53",
          5126 => x"53",
          5127 => x"59",
          5128 => x"25",
          5129 => x"80",
          5130 => x"51",
          5131 => x"81",
          5132 => x"14",
          5133 => x"33",
          5134 => x"71",
          5135 => x"76",
          5136 => x"2a",
          5137 => x"58",
          5138 => x"14",
          5139 => x"ff",
          5140 => x"87",
          5141 => x"d5",
          5142 => x"19",
          5143 => x"85",
          5144 => x"88",
          5145 => x"88",
          5146 => x"5b",
          5147 => x"84",
          5148 => x"85",
          5149 => x"d5",
          5150 => x"53",
          5151 => x"14",
          5152 => x"87",
          5153 => x"d5",
          5154 => x"76",
          5155 => x"75",
          5156 => x"82",
          5157 => x"18",
          5158 => x"12",
          5159 => x"2b",
          5160 => x"80",
          5161 => x"88",
          5162 => x"55",
          5163 => x"74",
          5164 => x"15",
          5165 => x"0d",
          5166 => x"0d",
          5167 => x"d5",
          5168 => x"38",
          5169 => x"71",
          5170 => x"38",
          5171 => x"8c",
          5172 => x"0d",
          5173 => x"0d",
          5174 => x"58",
          5175 => x"82",
          5176 => x"83",
          5177 => x"82",
          5178 => x"84",
          5179 => x"12",
          5180 => x"2b",
          5181 => x"59",
          5182 => x"81",
          5183 => x"75",
          5184 => x"cb",
          5185 => x"29",
          5186 => x"81",
          5187 => x"88",
          5188 => x"81",
          5189 => x"79",
          5190 => x"ff",
          5191 => x"7f",
          5192 => x"51",
          5193 => x"77",
          5194 => x"38",
          5195 => x"85",
          5196 => x"5a",
          5197 => x"33",
          5198 => x"71",
          5199 => x"57",
          5200 => x"38",
          5201 => x"ff",
          5202 => x"7a",
          5203 => x"80",
          5204 => x"82",
          5205 => x"11",
          5206 => x"12",
          5207 => x"2b",
          5208 => x"ff",
          5209 => x"52",
          5210 => x"55",
          5211 => x"83",
          5212 => x"80",
          5213 => x"26",
          5214 => x"74",
          5215 => x"2e",
          5216 => x"77",
          5217 => x"81",
          5218 => x"75",
          5219 => x"3f",
          5220 => x"82",
          5221 => x"79",
          5222 => x"f7",
          5223 => x"d5",
          5224 => x"1c",
          5225 => x"87",
          5226 => x"8b",
          5227 => x"2b",
          5228 => x"5e",
          5229 => x"7a",
          5230 => x"ff",
          5231 => x"88",
          5232 => x"56",
          5233 => x"15",
          5234 => x"ff",
          5235 => x"85",
          5236 => x"d5",
          5237 => x"83",
          5238 => x"72",
          5239 => x"33",
          5240 => x"71",
          5241 => x"70",
          5242 => x"5b",
          5243 => x"56",
          5244 => x"19",
          5245 => x"19",
          5246 => x"d4",
          5247 => x"84",
          5248 => x"12",
          5249 => x"2b",
          5250 => x"07",
          5251 => x"55",
          5252 => x"78",
          5253 => x"76",
          5254 => x"82",
          5255 => x"70",
          5256 => x"84",
          5257 => x"12",
          5258 => x"2b",
          5259 => x"2a",
          5260 => x"52",
          5261 => x"84",
          5262 => x"85",
          5263 => x"d5",
          5264 => x"84",
          5265 => x"82",
          5266 => x"8d",
          5267 => x"fe",
          5268 => x"52",
          5269 => x"08",
          5270 => x"db",
          5271 => x"71",
          5272 => x"38",
          5273 => x"ed",
          5274 => x"e4",
          5275 => x"82",
          5276 => x"84",
          5277 => x"ee",
          5278 => x"66",
          5279 => x"70",
          5280 => x"d5",
          5281 => x"2e",
          5282 => x"84",
          5283 => x"3f",
          5284 => x"7e",
          5285 => x"3f",
          5286 => x"08",
          5287 => x"39",
          5288 => x"7b",
          5289 => x"3f",
          5290 => x"ba",
          5291 => x"f5",
          5292 => x"d5",
          5293 => x"ff",
          5294 => x"d5",
          5295 => x"71",
          5296 => x"70",
          5297 => x"06",
          5298 => x"73",
          5299 => x"81",
          5300 => x"88",
          5301 => x"75",
          5302 => x"ff",
          5303 => x"88",
          5304 => x"73",
          5305 => x"70",
          5306 => x"33",
          5307 => x"07",
          5308 => x"53",
          5309 => x"48",
          5310 => x"54",
          5311 => x"56",
          5312 => x"80",
          5313 => x"76",
          5314 => x"06",
          5315 => x"83",
          5316 => x"42",
          5317 => x"33",
          5318 => x"71",
          5319 => x"70",
          5320 => x"70",
          5321 => x"33",
          5322 => x"71",
          5323 => x"53",
          5324 => x"56",
          5325 => x"25",
          5326 => x"75",
          5327 => x"ff",
          5328 => x"54",
          5329 => x"81",
          5330 => x"18",
          5331 => x"2e",
          5332 => x"8f",
          5333 => x"f6",
          5334 => x"83",
          5335 => x"58",
          5336 => x"7f",
          5337 => x"74",
          5338 => x"78",
          5339 => x"3f",
          5340 => x"7f",
          5341 => x"75",
          5342 => x"38",
          5343 => x"11",
          5344 => x"33",
          5345 => x"07",
          5346 => x"f4",
          5347 => x"52",
          5348 => x"b7",
          5349 => x"e4",
          5350 => x"ff",
          5351 => x"7c",
          5352 => x"2b",
          5353 => x"08",
          5354 => x"53",
          5355 => x"91",
          5356 => x"d5",
          5357 => x"84",
          5358 => x"ff",
          5359 => x"5c",
          5360 => x"60",
          5361 => x"74",
          5362 => x"38",
          5363 => x"c9",
          5364 => x"d4",
          5365 => x"11",
          5366 => x"33",
          5367 => x"07",
          5368 => x"f4",
          5369 => x"52",
          5370 => x"df",
          5371 => x"e4",
          5372 => x"ff",
          5373 => x"7c",
          5374 => x"2b",
          5375 => x"08",
          5376 => x"53",
          5377 => x"91",
          5378 => x"d5",
          5379 => x"84",
          5380 => x"05",
          5381 => x"73",
          5382 => x"06",
          5383 => x"7b",
          5384 => x"f9",
          5385 => x"d5",
          5386 => x"82",
          5387 => x"80",
          5388 => x"7d",
          5389 => x"82",
          5390 => x"51",
          5391 => x"3f",
          5392 => x"98",
          5393 => x"7a",
          5394 => x"38",
          5395 => x"52",
          5396 => x"8f",
          5397 => x"83",
          5398 => x"d4",
          5399 => x"05",
          5400 => x"3f",
          5401 => x"82",
          5402 => x"94",
          5403 => x"fc",
          5404 => x"77",
          5405 => x"54",
          5406 => x"82",
          5407 => x"55",
          5408 => x"08",
          5409 => x"38",
          5410 => x"52",
          5411 => x"08",
          5412 => x"fd",
          5413 => x"d5",
          5414 => x"3d",
          5415 => x"3d",
          5416 => x"05",
          5417 => x"52",
          5418 => x"87",
          5419 => x"e0",
          5420 => x"71",
          5421 => x"0c",
          5422 => x"04",
          5423 => x"02",
          5424 => x"02",
          5425 => x"05",
          5426 => x"83",
          5427 => x"26",
          5428 => x"72",
          5429 => x"c0",
          5430 => x"53",
          5431 => x"74",
          5432 => x"38",
          5433 => x"73",
          5434 => x"c0",
          5435 => x"51",
          5436 => x"85",
          5437 => x"98",
          5438 => x"52",
          5439 => x"82",
          5440 => x"70",
          5441 => x"38",
          5442 => x"8c",
          5443 => x"ec",
          5444 => x"fc",
          5445 => x"52",
          5446 => x"87",
          5447 => x"08",
          5448 => x"2e",
          5449 => x"82",
          5450 => x"34",
          5451 => x"13",
          5452 => x"82",
          5453 => x"86",
          5454 => x"f3",
          5455 => x"62",
          5456 => x"05",
          5457 => x"57",
          5458 => x"83",
          5459 => x"fe",
          5460 => x"d5",
          5461 => x"06",
          5462 => x"71",
          5463 => x"71",
          5464 => x"2b",
          5465 => x"80",
          5466 => x"92",
          5467 => x"c0",
          5468 => x"41",
          5469 => x"5a",
          5470 => x"87",
          5471 => x"0c",
          5472 => x"84",
          5473 => x"08",
          5474 => x"70",
          5475 => x"53",
          5476 => x"2e",
          5477 => x"08",
          5478 => x"70",
          5479 => x"34",
          5480 => x"80",
          5481 => x"53",
          5482 => x"2e",
          5483 => x"53",
          5484 => x"26",
          5485 => x"80",
          5486 => x"87",
          5487 => x"08",
          5488 => x"38",
          5489 => x"8c",
          5490 => x"80",
          5491 => x"78",
          5492 => x"99",
          5493 => x"0c",
          5494 => x"8c",
          5495 => x"08",
          5496 => x"51",
          5497 => x"38",
          5498 => x"8d",
          5499 => x"17",
          5500 => x"81",
          5501 => x"53",
          5502 => x"2e",
          5503 => x"fc",
          5504 => x"52",
          5505 => x"7d",
          5506 => x"ed",
          5507 => x"80",
          5508 => x"71",
          5509 => x"38",
          5510 => x"53",
          5511 => x"e4",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"02",
          5515 => x"05",
          5516 => x"58",
          5517 => x"80",
          5518 => x"fc",
          5519 => x"d5",
          5520 => x"06",
          5521 => x"71",
          5522 => x"81",
          5523 => x"38",
          5524 => x"2b",
          5525 => x"80",
          5526 => x"92",
          5527 => x"c0",
          5528 => x"40",
          5529 => x"5a",
          5530 => x"c0",
          5531 => x"76",
          5532 => x"76",
          5533 => x"75",
          5534 => x"2a",
          5535 => x"51",
          5536 => x"80",
          5537 => x"7a",
          5538 => x"5c",
          5539 => x"81",
          5540 => x"81",
          5541 => x"06",
          5542 => x"80",
          5543 => x"87",
          5544 => x"08",
          5545 => x"38",
          5546 => x"8c",
          5547 => x"80",
          5548 => x"77",
          5549 => x"99",
          5550 => x"0c",
          5551 => x"8c",
          5552 => x"08",
          5553 => x"51",
          5554 => x"38",
          5555 => x"8d",
          5556 => x"70",
          5557 => x"84",
          5558 => x"5b",
          5559 => x"2e",
          5560 => x"fc",
          5561 => x"52",
          5562 => x"7d",
          5563 => x"f8",
          5564 => x"80",
          5565 => x"71",
          5566 => x"38",
          5567 => x"53",
          5568 => x"e4",
          5569 => x"0d",
          5570 => x"0d",
          5571 => x"05",
          5572 => x"02",
          5573 => x"05",
          5574 => x"54",
          5575 => x"fe",
          5576 => x"e4",
          5577 => x"53",
          5578 => x"80",
          5579 => x"0b",
          5580 => x"8c",
          5581 => x"71",
          5582 => x"dc",
          5583 => x"24",
          5584 => x"84",
          5585 => x"92",
          5586 => x"54",
          5587 => x"8d",
          5588 => x"39",
          5589 => x"80",
          5590 => x"cb",
          5591 => x"70",
          5592 => x"81",
          5593 => x"52",
          5594 => x"8a",
          5595 => x"98",
          5596 => x"71",
          5597 => x"c0",
          5598 => x"52",
          5599 => x"81",
          5600 => x"c0",
          5601 => x"53",
          5602 => x"82",
          5603 => x"71",
          5604 => x"39",
          5605 => x"39",
          5606 => x"77",
          5607 => x"81",
          5608 => x"72",
          5609 => x"84",
          5610 => x"73",
          5611 => x"0c",
          5612 => x"04",
          5613 => x"74",
          5614 => x"71",
          5615 => x"2b",
          5616 => x"e4",
          5617 => x"84",
          5618 => x"fd",
          5619 => x"83",
          5620 => x"12",
          5621 => x"2b",
          5622 => x"07",
          5623 => x"70",
          5624 => x"2b",
          5625 => x"07",
          5626 => x"0c",
          5627 => x"56",
          5628 => x"3d",
          5629 => x"3d",
          5630 => x"84",
          5631 => x"22",
          5632 => x"72",
          5633 => x"54",
          5634 => x"2a",
          5635 => x"34",
          5636 => x"04",
          5637 => x"73",
          5638 => x"70",
          5639 => x"05",
          5640 => x"88",
          5641 => x"72",
          5642 => x"54",
          5643 => x"2a",
          5644 => x"70",
          5645 => x"34",
          5646 => x"51",
          5647 => x"83",
          5648 => x"fe",
          5649 => x"75",
          5650 => x"51",
          5651 => x"92",
          5652 => x"81",
          5653 => x"73",
          5654 => x"55",
          5655 => x"51",
          5656 => x"3d",
          5657 => x"3d",
          5658 => x"76",
          5659 => x"72",
          5660 => x"05",
          5661 => x"11",
          5662 => x"38",
          5663 => x"04",
          5664 => x"78",
          5665 => x"56",
          5666 => x"81",
          5667 => x"74",
          5668 => x"56",
          5669 => x"31",
          5670 => x"52",
          5671 => x"80",
          5672 => x"71",
          5673 => x"38",
          5674 => x"e4",
          5675 => x"0d",
          5676 => x"0d",
          5677 => x"51",
          5678 => x"73",
          5679 => x"81",
          5680 => x"33",
          5681 => x"38",
          5682 => x"d5",
          5683 => x"3d",
          5684 => x"0b",
          5685 => x"0c",
          5686 => x"0d",
          5687 => x"70",
          5688 => x"52",
          5689 => x"55",
          5690 => x"3f",
          5691 => x"d5",
          5692 => x"38",
          5693 => x"98",
          5694 => x"52",
          5695 => x"f9",
          5696 => x"d5",
          5697 => x"ff",
          5698 => x"72",
          5699 => x"38",
          5700 => x"72",
          5701 => x"d5",
          5702 => x"3d",
          5703 => x"3d",
          5704 => x"80",
          5705 => x"33",
          5706 => x"7a",
          5707 => x"38",
          5708 => x"16",
          5709 => x"16",
          5710 => x"17",
          5711 => x"f9",
          5712 => x"d5",
          5713 => x"2e",
          5714 => x"b7",
          5715 => x"e4",
          5716 => x"34",
          5717 => x"70",
          5718 => x"31",
          5719 => x"59",
          5720 => x"77",
          5721 => x"82",
          5722 => x"74",
          5723 => x"81",
          5724 => x"81",
          5725 => x"53",
          5726 => x"16",
          5727 => x"a5",
          5728 => x"81",
          5729 => x"d5",
          5730 => x"3d",
          5731 => x"3d",
          5732 => x"56",
          5733 => x"74",
          5734 => x"2e",
          5735 => x"51",
          5736 => x"82",
          5737 => x"57",
          5738 => x"08",
          5739 => x"54",
          5740 => x"16",
          5741 => x"33",
          5742 => x"3f",
          5743 => x"08",
          5744 => x"38",
          5745 => x"57",
          5746 => x"0c",
          5747 => x"e4",
          5748 => x"0d",
          5749 => x"0d",
          5750 => x"57",
          5751 => x"82",
          5752 => x"58",
          5753 => x"08",
          5754 => x"76",
          5755 => x"83",
          5756 => x"06",
          5757 => x"84",
          5758 => x"78",
          5759 => x"81",
          5760 => x"38",
          5761 => x"82",
          5762 => x"52",
          5763 => x"52",
          5764 => x"3f",
          5765 => x"52",
          5766 => x"51",
          5767 => x"84",
          5768 => x"d2",
          5769 => x"fb",
          5770 => x"8a",
          5771 => x"52",
          5772 => x"51",
          5773 => x"94",
          5774 => x"84",
          5775 => x"fb",
          5776 => x"17",
          5777 => x"a4",
          5778 => x"c8",
          5779 => x"08",
          5780 => x"b4",
          5781 => x"55",
          5782 => x"81",
          5783 => x"f7",
          5784 => x"84",
          5785 => x"53",
          5786 => x"17",
          5787 => x"99",
          5788 => x"e4",
          5789 => x"83",
          5790 => x"77",
          5791 => x"0c",
          5792 => x"04",
          5793 => x"77",
          5794 => x"12",
          5795 => x"55",
          5796 => x"56",
          5797 => x"8d",
          5798 => x"22",
          5799 => x"b0",
          5800 => x"57",
          5801 => x"d5",
          5802 => x"3d",
          5803 => x"3d",
          5804 => x"70",
          5805 => x"57",
          5806 => x"81",
          5807 => x"9c",
          5808 => x"81",
          5809 => x"74",
          5810 => x"72",
          5811 => x"f5",
          5812 => x"24",
          5813 => x"81",
          5814 => x"81",
          5815 => x"83",
          5816 => x"38",
          5817 => x"76",
          5818 => x"70",
          5819 => x"16",
          5820 => x"74",
          5821 => x"96",
          5822 => x"e4",
          5823 => x"38",
          5824 => x"06",
          5825 => x"33",
          5826 => x"89",
          5827 => x"08",
          5828 => x"54",
          5829 => x"fc",
          5830 => x"d5",
          5831 => x"fe",
          5832 => x"ff",
          5833 => x"11",
          5834 => x"2b",
          5835 => x"81",
          5836 => x"2a",
          5837 => x"51",
          5838 => x"e2",
          5839 => x"ff",
          5840 => x"da",
          5841 => x"2a",
          5842 => x"05",
          5843 => x"fc",
          5844 => x"d5",
          5845 => x"c6",
          5846 => x"83",
          5847 => x"05",
          5848 => x"f8",
          5849 => x"d5",
          5850 => x"ff",
          5851 => x"ae",
          5852 => x"2a",
          5853 => x"05",
          5854 => x"fc",
          5855 => x"d5",
          5856 => x"38",
          5857 => x"83",
          5858 => x"05",
          5859 => x"f8",
          5860 => x"d5",
          5861 => x"0a",
          5862 => x"39",
          5863 => x"82",
          5864 => x"89",
          5865 => x"f8",
          5866 => x"7c",
          5867 => x"56",
          5868 => x"77",
          5869 => x"38",
          5870 => x"08",
          5871 => x"38",
          5872 => x"72",
          5873 => x"9d",
          5874 => x"24",
          5875 => x"81",
          5876 => x"82",
          5877 => x"83",
          5878 => x"38",
          5879 => x"76",
          5880 => x"70",
          5881 => x"18",
          5882 => x"76",
          5883 => x"9e",
          5884 => x"e4",
          5885 => x"d5",
          5886 => x"d9",
          5887 => x"ff",
          5888 => x"05",
          5889 => x"81",
          5890 => x"54",
          5891 => x"80",
          5892 => x"77",
          5893 => x"f0",
          5894 => x"8f",
          5895 => x"51",
          5896 => x"34",
          5897 => x"17",
          5898 => x"2a",
          5899 => x"05",
          5900 => x"fa",
          5901 => x"d5",
          5902 => x"82",
          5903 => x"81",
          5904 => x"83",
          5905 => x"b8",
          5906 => x"2a",
          5907 => x"8f",
          5908 => x"2a",
          5909 => x"f0",
          5910 => x"06",
          5911 => x"72",
          5912 => x"ec",
          5913 => x"2a",
          5914 => x"05",
          5915 => x"fa",
          5916 => x"d5",
          5917 => x"82",
          5918 => x"80",
          5919 => x"83",
          5920 => x"52",
          5921 => x"fe",
          5922 => x"b8",
          5923 => x"e6",
          5924 => x"76",
          5925 => x"17",
          5926 => x"75",
          5927 => x"3f",
          5928 => x"08",
          5929 => x"e4",
          5930 => x"77",
          5931 => x"77",
          5932 => x"fc",
          5933 => x"b8",
          5934 => x"51",
          5935 => x"8b",
          5936 => x"e4",
          5937 => x"06",
          5938 => x"72",
          5939 => x"3f",
          5940 => x"17",
          5941 => x"d5",
          5942 => x"3d",
          5943 => x"3d",
          5944 => x"7e",
          5945 => x"56",
          5946 => x"75",
          5947 => x"74",
          5948 => x"27",
          5949 => x"80",
          5950 => x"ff",
          5951 => x"75",
          5952 => x"3f",
          5953 => x"08",
          5954 => x"e4",
          5955 => x"38",
          5956 => x"54",
          5957 => x"81",
          5958 => x"39",
          5959 => x"08",
          5960 => x"39",
          5961 => x"51",
          5962 => x"82",
          5963 => x"58",
          5964 => x"08",
          5965 => x"c7",
          5966 => x"e4",
          5967 => x"d2",
          5968 => x"e4",
          5969 => x"cf",
          5970 => x"74",
          5971 => x"fc",
          5972 => x"d5",
          5973 => x"38",
          5974 => x"fe",
          5975 => x"08",
          5976 => x"74",
          5977 => x"38",
          5978 => x"17",
          5979 => x"33",
          5980 => x"73",
          5981 => x"77",
          5982 => x"26",
          5983 => x"80",
          5984 => x"d5",
          5985 => x"3d",
          5986 => x"3d",
          5987 => x"71",
          5988 => x"5b",
          5989 => x"90",
          5990 => x"77",
          5991 => x"38",
          5992 => x"78",
          5993 => x"81",
          5994 => x"79",
          5995 => x"f9",
          5996 => x"55",
          5997 => x"e4",
          5998 => x"e0",
          5999 => x"e4",
          6000 => x"d5",
          6001 => x"2e",
          6002 => x"9c",
          6003 => x"d5",
          6004 => x"82",
          6005 => x"58",
          6006 => x"70",
          6007 => x"80",
          6008 => x"38",
          6009 => x"09",
          6010 => x"e2",
          6011 => x"56",
          6012 => x"76",
          6013 => x"82",
          6014 => x"7a",
          6015 => x"3f",
          6016 => x"d5",
          6017 => x"2e",
          6018 => x"86",
          6019 => x"e4",
          6020 => x"d5",
          6021 => x"70",
          6022 => x"07",
          6023 => x"7c",
          6024 => x"e4",
          6025 => x"51",
          6026 => x"81",
          6027 => x"d5",
          6028 => x"2e",
          6029 => x"17",
          6030 => x"74",
          6031 => x"73",
          6032 => x"27",
          6033 => x"58",
          6034 => x"80",
          6035 => x"56",
          6036 => x"9c",
          6037 => x"26",
          6038 => x"56",
          6039 => x"81",
          6040 => x"52",
          6041 => x"c6",
          6042 => x"e4",
          6043 => x"b8",
          6044 => x"82",
          6045 => x"81",
          6046 => x"06",
          6047 => x"d5",
          6048 => x"82",
          6049 => x"09",
          6050 => x"72",
          6051 => x"70",
          6052 => x"51",
          6053 => x"80",
          6054 => x"78",
          6055 => x"06",
          6056 => x"73",
          6057 => x"39",
          6058 => x"52",
          6059 => x"f7",
          6060 => x"e4",
          6061 => x"e4",
          6062 => x"82",
          6063 => x"07",
          6064 => x"55",
          6065 => x"2e",
          6066 => x"80",
          6067 => x"75",
          6068 => x"76",
          6069 => x"3f",
          6070 => x"08",
          6071 => x"38",
          6072 => x"0c",
          6073 => x"fe",
          6074 => x"08",
          6075 => x"74",
          6076 => x"ff",
          6077 => x"0c",
          6078 => x"81",
          6079 => x"84",
          6080 => x"39",
          6081 => x"81",
          6082 => x"8c",
          6083 => x"8c",
          6084 => x"e4",
          6085 => x"39",
          6086 => x"55",
          6087 => x"e4",
          6088 => x"0d",
          6089 => x"0d",
          6090 => x"55",
          6091 => x"82",
          6092 => x"58",
          6093 => x"d5",
          6094 => x"d8",
          6095 => x"74",
          6096 => x"3f",
          6097 => x"08",
          6098 => x"08",
          6099 => x"59",
          6100 => x"77",
          6101 => x"70",
          6102 => x"8a",
          6103 => x"84",
          6104 => x"56",
          6105 => x"58",
          6106 => x"97",
          6107 => x"75",
          6108 => x"52",
          6109 => x"51",
          6110 => x"82",
          6111 => x"80",
          6112 => x"8a",
          6113 => x"32",
          6114 => x"72",
          6115 => x"2a",
          6116 => x"56",
          6117 => x"e4",
          6118 => x"0d",
          6119 => x"0d",
          6120 => x"08",
          6121 => x"74",
          6122 => x"26",
          6123 => x"74",
          6124 => x"72",
          6125 => x"74",
          6126 => x"88",
          6127 => x"73",
          6128 => x"33",
          6129 => x"27",
          6130 => x"16",
          6131 => x"9b",
          6132 => x"2a",
          6133 => x"88",
          6134 => x"58",
          6135 => x"80",
          6136 => x"16",
          6137 => x"0c",
          6138 => x"8a",
          6139 => x"89",
          6140 => x"72",
          6141 => x"38",
          6142 => x"51",
          6143 => x"82",
          6144 => x"54",
          6145 => x"08",
          6146 => x"38",
          6147 => x"d5",
          6148 => x"8b",
          6149 => x"08",
          6150 => x"08",
          6151 => x"82",
          6152 => x"74",
          6153 => x"cb",
          6154 => x"75",
          6155 => x"3f",
          6156 => x"08",
          6157 => x"73",
          6158 => x"98",
          6159 => x"82",
          6160 => x"2e",
          6161 => x"39",
          6162 => x"39",
          6163 => x"13",
          6164 => x"74",
          6165 => x"16",
          6166 => x"18",
          6167 => x"77",
          6168 => x"0c",
          6169 => x"04",
          6170 => x"7a",
          6171 => x"12",
          6172 => x"59",
          6173 => x"80",
          6174 => x"86",
          6175 => x"98",
          6176 => x"14",
          6177 => x"55",
          6178 => x"81",
          6179 => x"83",
          6180 => x"77",
          6181 => x"81",
          6182 => x"0c",
          6183 => x"55",
          6184 => x"76",
          6185 => x"17",
          6186 => x"74",
          6187 => x"9b",
          6188 => x"39",
          6189 => x"ff",
          6190 => x"2a",
          6191 => x"81",
          6192 => x"52",
          6193 => x"e6",
          6194 => x"e4",
          6195 => x"55",
          6196 => x"d5",
          6197 => x"80",
          6198 => x"55",
          6199 => x"08",
          6200 => x"f4",
          6201 => x"08",
          6202 => x"08",
          6203 => x"38",
          6204 => x"77",
          6205 => x"84",
          6206 => x"39",
          6207 => x"52",
          6208 => x"86",
          6209 => x"e4",
          6210 => x"55",
          6211 => x"08",
          6212 => x"c4",
          6213 => x"82",
          6214 => x"81",
          6215 => x"81",
          6216 => x"e4",
          6217 => x"b0",
          6218 => x"e4",
          6219 => x"51",
          6220 => x"82",
          6221 => x"a0",
          6222 => x"15",
          6223 => x"75",
          6224 => x"3f",
          6225 => x"08",
          6226 => x"76",
          6227 => x"77",
          6228 => x"9c",
          6229 => x"55",
          6230 => x"e4",
          6231 => x"0d",
          6232 => x"0d",
          6233 => x"08",
          6234 => x"80",
          6235 => x"fc",
          6236 => x"d5",
          6237 => x"82",
          6238 => x"80",
          6239 => x"d5",
          6240 => x"98",
          6241 => x"78",
          6242 => x"3f",
          6243 => x"08",
          6244 => x"e4",
          6245 => x"38",
          6246 => x"08",
          6247 => x"70",
          6248 => x"58",
          6249 => x"2e",
          6250 => x"83",
          6251 => x"82",
          6252 => x"55",
          6253 => x"81",
          6254 => x"07",
          6255 => x"2e",
          6256 => x"16",
          6257 => x"2e",
          6258 => x"88",
          6259 => x"82",
          6260 => x"56",
          6261 => x"51",
          6262 => x"82",
          6263 => x"54",
          6264 => x"08",
          6265 => x"9b",
          6266 => x"2e",
          6267 => x"83",
          6268 => x"73",
          6269 => x"0c",
          6270 => x"04",
          6271 => x"76",
          6272 => x"54",
          6273 => x"82",
          6274 => x"83",
          6275 => x"76",
          6276 => x"53",
          6277 => x"2e",
          6278 => x"90",
          6279 => x"51",
          6280 => x"82",
          6281 => x"90",
          6282 => x"53",
          6283 => x"e4",
          6284 => x"0d",
          6285 => x"0d",
          6286 => x"83",
          6287 => x"54",
          6288 => x"55",
          6289 => x"3f",
          6290 => x"51",
          6291 => x"2e",
          6292 => x"8b",
          6293 => x"2a",
          6294 => x"51",
          6295 => x"86",
          6296 => x"fd",
          6297 => x"54",
          6298 => x"53",
          6299 => x"71",
          6300 => x"05",
          6301 => x"05",
          6302 => x"05",
          6303 => x"06",
          6304 => x"51",
          6305 => x"e4",
          6306 => x"d5",
          6307 => x"3d",
          6308 => x"3d",
          6309 => x"40",
          6310 => x"08",
          6311 => x"ff",
          6312 => x"98",
          6313 => x"2e",
          6314 => x"98",
          6315 => x"7d",
          6316 => x"3f",
          6317 => x"08",
          6318 => x"e4",
          6319 => x"38",
          6320 => x"70",
          6321 => x"73",
          6322 => x"5b",
          6323 => x"8b",
          6324 => x"06",
          6325 => x"06",
          6326 => x"86",
          6327 => x"d5",
          6328 => x"73",
          6329 => x"09",
          6330 => x"38",
          6331 => x"d5",
          6332 => x"73",
          6333 => x"81",
          6334 => x"81",
          6335 => x"07",
          6336 => x"38",
          6337 => x"08",
          6338 => x"54",
          6339 => x"2e",
          6340 => x"83",
          6341 => x"75",
          6342 => x"38",
          6343 => x"81",
          6344 => x"8f",
          6345 => x"06",
          6346 => x"73",
          6347 => x"81",
          6348 => x"72",
          6349 => x"38",
          6350 => x"74",
          6351 => x"70",
          6352 => x"ac",
          6353 => x"5d",
          6354 => x"2e",
          6355 => x"81",
          6356 => x"15",
          6357 => x"73",
          6358 => x"06",
          6359 => x"8c",
          6360 => x"16",
          6361 => x"cc",
          6362 => x"e4",
          6363 => x"ff",
          6364 => x"80",
          6365 => x"33",
          6366 => x"06",
          6367 => x"05",
          6368 => x"7b",
          6369 => x"c7",
          6370 => x"75",
          6371 => x"a4",
          6372 => x"e4",
          6373 => x"ff",
          6374 => x"80",
          6375 => x"73",
          6376 => x"80",
          6377 => x"10",
          6378 => x"53",
          6379 => x"81",
          6380 => x"39",
          6381 => x"ff",
          6382 => x"06",
          6383 => x"17",
          6384 => x"27",
          6385 => x"33",
          6386 => x"70",
          6387 => x"54",
          6388 => x"2e",
          6389 => x"81",
          6390 => x"38",
          6391 => x"53",
          6392 => x"ff",
          6393 => x"ff",
          6394 => x"84",
          6395 => x"53",
          6396 => x"39",
          6397 => x"74",
          6398 => x"3f",
          6399 => x"08",
          6400 => x"53",
          6401 => x"a7",
          6402 => x"ac",
          6403 => x"39",
          6404 => x"51",
          6405 => x"82",
          6406 => x"5b",
          6407 => x"08",
          6408 => x"19",
          6409 => x"38",
          6410 => x"0b",
          6411 => x"7a",
          6412 => x"0c",
          6413 => x"04",
          6414 => x"60",
          6415 => x"59",
          6416 => x"51",
          6417 => x"82",
          6418 => x"58",
          6419 => x"08",
          6420 => x"81",
          6421 => x"5c",
          6422 => x"1a",
          6423 => x"08",
          6424 => x"ea",
          6425 => x"d5",
          6426 => x"82",
          6427 => x"83",
          6428 => x"19",
          6429 => x"57",
          6430 => x"38",
          6431 => x"f6",
          6432 => x"33",
          6433 => x"81",
          6434 => x"54",
          6435 => x"34",
          6436 => x"2e",
          6437 => x"74",
          6438 => x"81",
          6439 => x"74",
          6440 => x"38",
          6441 => x"38",
          6442 => x"09",
          6443 => x"f7",
          6444 => x"33",
          6445 => x"70",
          6446 => x"55",
          6447 => x"a1",
          6448 => x"2a",
          6449 => x"51",
          6450 => x"2e",
          6451 => x"17",
          6452 => x"bf",
          6453 => x"1c",
          6454 => x"0c",
          6455 => x"75",
          6456 => x"81",
          6457 => x"38",
          6458 => x"56",
          6459 => x"09",
          6460 => x"ac",
          6461 => x"08",
          6462 => x"5d",
          6463 => x"82",
          6464 => x"83",
          6465 => x"55",
          6466 => x"38",
          6467 => x"bf",
          6468 => x"f3",
          6469 => x"81",
          6470 => x"82",
          6471 => x"33",
          6472 => x"e5",
          6473 => x"d5",
          6474 => x"ff",
          6475 => x"79",
          6476 => x"38",
          6477 => x"26",
          6478 => x"75",
          6479 => x"a0",
          6480 => x"e4",
          6481 => x"1e",
          6482 => x"55",
          6483 => x"55",
          6484 => x"3f",
          6485 => x"e4",
          6486 => x"81",
          6487 => x"38",
          6488 => x"39",
          6489 => x"ff",
          6490 => x"06",
          6491 => x"1b",
          6492 => x"27",
          6493 => x"76",
          6494 => x"2a",
          6495 => x"51",
          6496 => x"80",
          6497 => x"73",
          6498 => x"38",
          6499 => x"70",
          6500 => x"73",
          6501 => x"1c",
          6502 => x"06",
          6503 => x"39",
          6504 => x"73",
          6505 => x"7b",
          6506 => x"51",
          6507 => x"82",
          6508 => x"81",
          6509 => x"73",
          6510 => x"38",
          6511 => x"81",
          6512 => x"95",
          6513 => x"a0",
          6514 => x"19",
          6515 => x"b0",
          6516 => x"e4",
          6517 => x"9e",
          6518 => x"5c",
          6519 => x"1a",
          6520 => x"78",
          6521 => x"3f",
          6522 => x"08",
          6523 => x"e4",
          6524 => x"fc",
          6525 => x"82",
          6526 => x"90",
          6527 => x"ee",
          6528 => x"70",
          6529 => x"33",
          6530 => x"56",
          6531 => x"55",
          6532 => x"38",
          6533 => x"08",
          6534 => x"56",
          6535 => x"2e",
          6536 => x"1d",
          6537 => x"70",
          6538 => x"5d",
          6539 => x"53",
          6540 => x"53",
          6541 => x"53",
          6542 => x"87",
          6543 => x"cb",
          6544 => x"06",
          6545 => x"2e",
          6546 => x"80",
          6547 => x"1b",
          6548 => x"8c",
          6549 => x"56",
          6550 => x"7d",
          6551 => x"e3",
          6552 => x"7b",
          6553 => x"38",
          6554 => x"22",
          6555 => x"ff",
          6556 => x"73",
          6557 => x"38",
          6558 => x"ff",
          6559 => x"59",
          6560 => x"74",
          6561 => x"10",
          6562 => x"2a",
          6563 => x"70",
          6564 => x"56",
          6565 => x"80",
          6566 => x"75",
          6567 => x"32",
          6568 => x"57",
          6569 => x"db",
          6570 => x"75",
          6571 => x"84",
          6572 => x"57",
          6573 => x"07",
          6574 => x"b9",
          6575 => x"38",
          6576 => x"73",
          6577 => x"16",
          6578 => x"84",
          6579 => x"56",
          6580 => x"94",
          6581 => x"17",
          6582 => x"74",
          6583 => x"27",
          6584 => x"33",
          6585 => x"2e",
          6586 => x"19",
          6587 => x"54",
          6588 => x"82",
          6589 => x"80",
          6590 => x"ff",
          6591 => x"74",
          6592 => x"81",
          6593 => x"15",
          6594 => x"27",
          6595 => x"19",
          6596 => x"54",
          6597 => x"3d",
          6598 => x"05",
          6599 => x"81",
          6600 => x"a0",
          6601 => x"26",
          6602 => x"17",
          6603 => x"33",
          6604 => x"75",
          6605 => x"75",
          6606 => x"79",
          6607 => x"3f",
          6608 => x"08",
          6609 => x"1b",
          6610 => x"7b",
          6611 => x"38",
          6612 => x"80",
          6613 => x"f0",
          6614 => x"e4",
          6615 => x"d5",
          6616 => x"2e",
          6617 => x"82",
          6618 => x"80",
          6619 => x"ab",
          6620 => x"80",
          6621 => x"70",
          6622 => x"81",
          6623 => x"5e",
          6624 => x"80",
          6625 => x"8d",
          6626 => x"51",
          6627 => x"3f",
          6628 => x"08",
          6629 => x"52",
          6630 => x"c5",
          6631 => x"e4",
          6632 => x"d5",
          6633 => x"9e",
          6634 => x"59",
          6635 => x"81",
          6636 => x"85",
          6637 => x"08",
          6638 => x"54",
          6639 => x"dd",
          6640 => x"e4",
          6641 => x"d5",
          6642 => x"fa",
          6643 => x"51",
          6644 => x"82",
          6645 => x"81",
          6646 => x"98",
          6647 => x"7b",
          6648 => x"3f",
          6649 => x"08",
          6650 => x"e4",
          6651 => x"38",
          6652 => x"9c",
          6653 => x"81",
          6654 => x"57",
          6655 => x"17",
          6656 => x"8b",
          6657 => x"d5",
          6658 => x"17",
          6659 => x"e4",
          6660 => x"16",
          6661 => x"3f",
          6662 => x"f3",
          6663 => x"55",
          6664 => x"ff",
          6665 => x"74",
          6666 => x"22",
          6667 => x"51",
          6668 => x"82",
          6669 => x"33",
          6670 => x"df",
          6671 => x"85",
          6672 => x"ff",
          6673 => x"57",
          6674 => x"d4",
          6675 => x"ff",
          6676 => x"38",
          6677 => x"70",
          6678 => x"73",
          6679 => x"80",
          6680 => x"77",
          6681 => x"0b",
          6682 => x"80",
          6683 => x"ef",
          6684 => x"d5",
          6685 => x"82",
          6686 => x"80",
          6687 => x"19",
          6688 => x"d7",
          6689 => x"08",
          6690 => x"e2",
          6691 => x"d5",
          6692 => x"82",
          6693 => x"ae",
          6694 => x"82",
          6695 => x"52",
          6696 => x"51",
          6697 => x"8b",
          6698 => x"52",
          6699 => x"51",
          6700 => x"9c",
          6701 => x"1b",
          6702 => x"55",
          6703 => x"16",
          6704 => x"83",
          6705 => x"55",
          6706 => x"e4",
          6707 => x"0d",
          6708 => x"0d",
          6709 => x"90",
          6710 => x"13",
          6711 => x"57",
          6712 => x"2e",
          6713 => x"52",
          6714 => x"b1",
          6715 => x"e4",
          6716 => x"d5",
          6717 => x"c9",
          6718 => x"08",
          6719 => x"e1",
          6720 => x"d5",
          6721 => x"82",
          6722 => x"ab",
          6723 => x"08",
          6724 => x"34",
          6725 => x"17",
          6726 => x"08",
          6727 => x"38",
          6728 => x"08",
          6729 => x"ee",
          6730 => x"d5",
          6731 => x"82",
          6732 => x"80",
          6733 => x"73",
          6734 => x"81",
          6735 => x"82",
          6736 => x"d5",
          6737 => x"3d",
          6738 => x"3d",
          6739 => x"71",
          6740 => x"5c",
          6741 => x"19",
          6742 => x"08",
          6743 => x"e2",
          6744 => x"08",
          6745 => x"bb",
          6746 => x"71",
          6747 => x"08",
          6748 => x"57",
          6749 => x"72",
          6750 => x"9d",
          6751 => x"14",
          6752 => x"1b",
          6753 => x"7a",
          6754 => x"d0",
          6755 => x"83",
          6756 => x"51",
          6757 => x"ff",
          6758 => x"74",
          6759 => x"39",
          6760 => x"11",
          6761 => x"31",
          6762 => x"83",
          6763 => x"90",
          6764 => x"51",
          6765 => x"3f",
          6766 => x"08",
          6767 => x"06",
          6768 => x"75",
          6769 => x"81",
          6770 => x"38",
          6771 => x"53",
          6772 => x"74",
          6773 => x"82",
          6774 => x"74",
          6775 => x"70",
          6776 => x"25",
          6777 => x"07",
          6778 => x"73",
          6779 => x"38",
          6780 => x"39",
          6781 => x"81",
          6782 => x"57",
          6783 => x"1d",
          6784 => x"11",
          6785 => x"54",
          6786 => x"f1",
          6787 => x"70",
          6788 => x"30",
          6789 => x"51",
          6790 => x"94",
          6791 => x"0b",
          6792 => x"80",
          6793 => x"58",
          6794 => x"1c",
          6795 => x"33",
          6796 => x"56",
          6797 => x"2e",
          6798 => x"85",
          6799 => x"06",
          6800 => x"e5",
          6801 => x"32",
          6802 => x"72",
          6803 => x"51",
          6804 => x"8b",
          6805 => x"72",
          6806 => x"38",
          6807 => x"81",
          6808 => x"81",
          6809 => x"76",
          6810 => x"58",
          6811 => x"57",
          6812 => x"ff",
          6813 => x"17",
          6814 => x"80",
          6815 => x"34",
          6816 => x"53",
          6817 => x"38",
          6818 => x"bf",
          6819 => x"34",
          6820 => x"e1",
          6821 => x"89",
          6822 => x"5a",
          6823 => x"2e",
          6824 => x"96",
          6825 => x"55",
          6826 => x"ff",
          6827 => x"55",
          6828 => x"aa",
          6829 => x"08",
          6830 => x"51",
          6831 => x"27",
          6832 => x"84",
          6833 => x"39",
          6834 => x"53",
          6835 => x"53",
          6836 => x"8a",
          6837 => x"70",
          6838 => x"06",
          6839 => x"76",
          6840 => x"58",
          6841 => x"81",
          6842 => x"71",
          6843 => x"55",
          6844 => x"b5",
          6845 => x"94",
          6846 => x"0b",
          6847 => x"9c",
          6848 => x"11",
          6849 => x"72",
          6850 => x"89",
          6851 => x"1c",
          6852 => x"13",
          6853 => x"34",
          6854 => x"9c",
          6855 => x"d9",
          6856 => x"d5",
          6857 => x"0c",
          6858 => x"d9",
          6859 => x"d5",
          6860 => x"19",
          6861 => x"51",
          6862 => x"82",
          6863 => x"84",
          6864 => x"3d",
          6865 => x"3d",
          6866 => x"08",
          6867 => x"64",
          6868 => x"55",
          6869 => x"2e",
          6870 => x"55",
          6871 => x"2e",
          6872 => x"80",
          6873 => x"7f",
          6874 => x"88",
          6875 => x"39",
          6876 => x"80",
          6877 => x"56",
          6878 => x"af",
          6879 => x"06",
          6880 => x"56",
          6881 => x"32",
          6882 => x"80",
          6883 => x"51",
          6884 => x"dc",
          6885 => x"1f",
          6886 => x"33",
          6887 => x"9f",
          6888 => x"ff",
          6889 => x"1f",
          6890 => x"7d",
          6891 => x"3f",
          6892 => x"08",
          6893 => x"39",
          6894 => x"08",
          6895 => x"5b",
          6896 => x"92",
          6897 => x"51",
          6898 => x"82",
          6899 => x"ff",
          6900 => x"38",
          6901 => x"0b",
          6902 => x"08",
          6903 => x"78",
          6904 => x"d5",
          6905 => x"2a",
          6906 => x"75",
          6907 => x"59",
          6908 => x"08",
          6909 => x"06",
          6910 => x"70",
          6911 => x"27",
          6912 => x"07",
          6913 => x"56",
          6914 => x"75",
          6915 => x"ae",
          6916 => x"ff",
          6917 => x"75",
          6918 => x"80",
          6919 => x"3f",
          6920 => x"08",
          6921 => x"78",
          6922 => x"81",
          6923 => x"10",
          6924 => x"74",
          6925 => x"59",
          6926 => x"81",
          6927 => x"61",
          6928 => x"56",
          6929 => x"2e",
          6930 => x"83",
          6931 => x"73",
          6932 => x"70",
          6933 => x"25",
          6934 => x"51",
          6935 => x"38",
          6936 => x"76",
          6937 => x"57",
          6938 => x"09",
          6939 => x"38",
          6940 => x"73",
          6941 => x"38",
          6942 => x"78",
          6943 => x"81",
          6944 => x"38",
          6945 => x"54",
          6946 => x"09",
          6947 => x"c1",
          6948 => x"54",
          6949 => x"09",
          6950 => x"38",
          6951 => x"54",
          6952 => x"80",
          6953 => x"56",
          6954 => x"78",
          6955 => x"38",
          6956 => x"75",
          6957 => x"57",
          6958 => x"58",
          6959 => x"e9",
          6960 => x"07",
          6961 => x"1f",
          6962 => x"39",
          6963 => x"a8",
          6964 => x"1a",
          6965 => x"74",
          6966 => x"71",
          6967 => x"70",
          6968 => x"2a",
          6969 => x"58",
          6970 => x"ae",
          6971 => x"73",
          6972 => x"19",
          6973 => x"38",
          6974 => x"11",
          6975 => x"74",
          6976 => x"38",
          6977 => x"90",
          6978 => x"07",
          6979 => x"39",
          6980 => x"70",
          6981 => x"06",
          6982 => x"73",
          6983 => x"81",
          6984 => x"81",
          6985 => x"1b",
          6986 => x"55",
          6987 => x"2e",
          6988 => x"8f",
          6989 => x"ff",
          6990 => x"73",
          6991 => x"81",
          6992 => x"76",
          6993 => x"78",
          6994 => x"38",
          6995 => x"05",
          6996 => x"54",
          6997 => x"9d",
          6998 => x"1a",
          6999 => x"ff",
          7000 => x"80",
          7001 => x"fe",
          7002 => x"55",
          7003 => x"2e",
          7004 => x"eb",
          7005 => x"a0",
          7006 => x"51",
          7007 => x"80",
          7008 => x"88",
          7009 => x"1a",
          7010 => x"1f",
          7011 => x"75",
          7012 => x"94",
          7013 => x"2e",
          7014 => x"ae",
          7015 => x"70",
          7016 => x"51",
          7017 => x"2e",
          7018 => x"80",
          7019 => x"76",
          7020 => x"d1",
          7021 => x"73",
          7022 => x"26",
          7023 => x"5b",
          7024 => x"70",
          7025 => x"07",
          7026 => x"7e",
          7027 => x"55",
          7028 => x"2e",
          7029 => x"8b",
          7030 => x"38",
          7031 => x"8b",
          7032 => x"07",
          7033 => x"26",
          7034 => x"78",
          7035 => x"8b",
          7036 => x"81",
          7037 => x"5f",
          7038 => x"80",
          7039 => x"af",
          7040 => x"07",
          7041 => x"52",
          7042 => x"ce",
          7043 => x"d5",
          7044 => x"ff",
          7045 => x"87",
          7046 => x"06",
          7047 => x"73",
          7048 => x"38",
          7049 => x"06",
          7050 => x"11",
          7051 => x"81",
          7052 => x"a4",
          7053 => x"54",
          7054 => x"8a",
          7055 => x"07",
          7056 => x"fe",
          7057 => x"18",
          7058 => x"88",
          7059 => x"73",
          7060 => x"18",
          7061 => x"39",
          7062 => x"92",
          7063 => x"82",
          7064 => x"d4",
          7065 => x"d5",
          7066 => x"2e",
          7067 => x"df",
          7068 => x"58",
          7069 => x"ff",
          7070 => x"73",
          7071 => x"38",
          7072 => x"5c",
          7073 => x"54",
          7074 => x"8e",
          7075 => x"07",
          7076 => x"83",
          7077 => x"58",
          7078 => x"18",
          7079 => x"75",
          7080 => x"18",
          7081 => x"39",
          7082 => x"54",
          7083 => x"2e",
          7084 => x"86",
          7085 => x"a0",
          7086 => x"88",
          7087 => x"06",
          7088 => x"82",
          7089 => x"06",
          7090 => x"06",
          7091 => x"2e",
          7092 => x"83",
          7093 => x"83",
          7094 => x"06",
          7095 => x"82",
          7096 => x"81",
          7097 => x"06",
          7098 => x"9f",
          7099 => x"06",
          7100 => x"2e",
          7101 => x"90",
          7102 => x"82",
          7103 => x"06",
          7104 => x"80",
          7105 => x"76",
          7106 => x"76",
          7107 => x"7d",
          7108 => x"3f",
          7109 => x"08",
          7110 => x"56",
          7111 => x"e4",
          7112 => x"be",
          7113 => x"e4",
          7114 => x"09",
          7115 => x"e8",
          7116 => x"2a",
          7117 => x"76",
          7118 => x"51",
          7119 => x"2e",
          7120 => x"81",
          7121 => x"80",
          7122 => x"38",
          7123 => x"ab",
          7124 => x"56",
          7125 => x"74",
          7126 => x"73",
          7127 => x"56",
          7128 => x"82",
          7129 => x"06",
          7130 => x"ac",
          7131 => x"33",
          7132 => x"70",
          7133 => x"55",
          7134 => x"2e",
          7135 => x"1e",
          7136 => x"06",
          7137 => x"05",
          7138 => x"e4",
          7139 => x"d5",
          7140 => x"1f",
          7141 => x"39",
          7142 => x"e4",
          7143 => x"0d",
          7144 => x"0d",
          7145 => x"7b",
          7146 => x"73",
          7147 => x"55",
          7148 => x"2e",
          7149 => x"75",
          7150 => x"57",
          7151 => x"26",
          7152 => x"ba",
          7153 => x"70",
          7154 => x"ba",
          7155 => x"06",
          7156 => x"73",
          7157 => x"70",
          7158 => x"51",
          7159 => x"89",
          7160 => x"82",
          7161 => x"ff",
          7162 => x"56",
          7163 => x"2e",
          7164 => x"80",
          7165 => x"d4",
          7166 => x"08",
          7167 => x"76",
          7168 => x"58",
          7169 => x"81",
          7170 => x"ff",
          7171 => x"53",
          7172 => x"26",
          7173 => x"13",
          7174 => x"06",
          7175 => x"9f",
          7176 => x"99",
          7177 => x"e0",
          7178 => x"ff",
          7179 => x"72",
          7180 => x"2a",
          7181 => x"72",
          7182 => x"06",
          7183 => x"ff",
          7184 => x"30",
          7185 => x"70",
          7186 => x"07",
          7187 => x"9f",
          7188 => x"54",
          7189 => x"80",
          7190 => x"81",
          7191 => x"59",
          7192 => x"25",
          7193 => x"8b",
          7194 => x"24",
          7195 => x"76",
          7196 => x"78",
          7197 => x"82",
          7198 => x"51",
          7199 => x"e4",
          7200 => x"0d",
          7201 => x"0d",
          7202 => x"0b",
          7203 => x"ff",
          7204 => x"0c",
          7205 => x"51",
          7206 => x"84",
          7207 => x"e4",
          7208 => x"38",
          7209 => x"51",
          7210 => x"82",
          7211 => x"83",
          7212 => x"54",
          7213 => x"82",
          7214 => x"09",
          7215 => x"e3",
          7216 => x"b8",
          7217 => x"57",
          7218 => x"2e",
          7219 => x"83",
          7220 => x"74",
          7221 => x"70",
          7222 => x"25",
          7223 => x"51",
          7224 => x"38",
          7225 => x"2e",
          7226 => x"b5",
          7227 => x"82",
          7228 => x"80",
          7229 => x"cf",
          7230 => x"d5",
          7231 => x"82",
          7232 => x"80",
          7233 => x"85",
          7234 => x"98",
          7235 => x"16",
          7236 => x"3f",
          7237 => x"08",
          7238 => x"e4",
          7239 => x"83",
          7240 => x"74",
          7241 => x"0c",
          7242 => x"04",
          7243 => x"61",
          7244 => x"80",
          7245 => x"58",
          7246 => x"0c",
          7247 => x"e1",
          7248 => x"e4",
          7249 => x"56",
          7250 => x"d5",
          7251 => x"87",
          7252 => x"d5",
          7253 => x"29",
          7254 => x"05",
          7255 => x"53",
          7256 => x"80",
          7257 => x"38",
          7258 => x"76",
          7259 => x"74",
          7260 => x"72",
          7261 => x"38",
          7262 => x"51",
          7263 => x"82",
          7264 => x"81",
          7265 => x"81",
          7266 => x"72",
          7267 => x"80",
          7268 => x"38",
          7269 => x"70",
          7270 => x"53",
          7271 => x"86",
          7272 => x"f2",
          7273 => x"34",
          7274 => x"82",
          7275 => x"33",
          7276 => x"81",
          7277 => x"33",
          7278 => x"3f",
          7279 => x"08",
          7280 => x"70",
          7281 => x"55",
          7282 => x"86",
          7283 => x"80",
          7284 => x"74",
          7285 => x"81",
          7286 => x"8a",
          7287 => x"b8",
          7288 => x"53",
          7289 => x"fd",
          7290 => x"d5",
          7291 => x"ff",
          7292 => x"82",
          7293 => x"76",
          7294 => x"9c",
          7295 => x"d9",
          7296 => x"72",
          7297 => x"90",
          7298 => x"74",
          7299 => x"56",
          7300 => x"33",
          7301 => x"72",
          7302 => x"38",
          7303 => x"51",
          7304 => x"82",
          7305 => x"57",
          7306 => x"84",
          7307 => x"ff",
          7308 => x"56",
          7309 => x"25",
          7310 => x"18",
          7311 => x"11",
          7312 => x"70",
          7313 => x"71",
          7314 => x"71",
          7315 => x"f0",
          7316 => x"51",
          7317 => x"74",
          7318 => x"57",
          7319 => x"90",
          7320 => x"73",
          7321 => x"3f",
          7322 => x"08",
          7323 => x"57",
          7324 => x"d5",
          7325 => x"54",
          7326 => x"2e",
          7327 => x"83",
          7328 => x"81",
          7329 => x"38",
          7330 => x"8c",
          7331 => x"84",
          7332 => x"83",
          7333 => x"38",
          7334 => x"84",
          7335 => x"38",
          7336 => x"81",
          7337 => x"38",
          7338 => x"51",
          7339 => x"82",
          7340 => x"83",
          7341 => x"53",
          7342 => x"2e",
          7343 => x"84",
          7344 => x"ce",
          7345 => x"ec",
          7346 => x"e4",
          7347 => x"ff",
          7348 => x"8d",
          7349 => x"14",
          7350 => x"3f",
          7351 => x"08",
          7352 => x"15",
          7353 => x"14",
          7354 => x"34",
          7355 => x"33",
          7356 => x"81",
          7357 => x"54",
          7358 => x"72",
          7359 => x"98",
          7360 => x"ff",
          7361 => x"29",
          7362 => x"33",
          7363 => x"72",
          7364 => x"72",
          7365 => x"38",
          7366 => x"06",
          7367 => x"2e",
          7368 => x"56",
          7369 => x"80",
          7370 => x"c9",
          7371 => x"d5",
          7372 => x"82",
          7373 => x"88",
          7374 => x"8f",
          7375 => x"56",
          7376 => x"38",
          7377 => x"51",
          7378 => x"82",
          7379 => x"83",
          7380 => x"55",
          7381 => x"80",
          7382 => x"c8",
          7383 => x"d5",
          7384 => x"80",
          7385 => x"c8",
          7386 => x"d5",
          7387 => x"ff",
          7388 => x"8d",
          7389 => x"2e",
          7390 => x"88",
          7391 => x"14",
          7392 => x"05",
          7393 => x"75",
          7394 => x"38",
          7395 => x"52",
          7396 => x"51",
          7397 => x"3f",
          7398 => x"08",
          7399 => x"e4",
          7400 => x"82",
          7401 => x"d5",
          7402 => x"ff",
          7403 => x"26",
          7404 => x"57",
          7405 => x"f5",
          7406 => x"82",
          7407 => x"f5",
          7408 => x"81",
          7409 => x"8d",
          7410 => x"2e",
          7411 => x"82",
          7412 => x"16",
          7413 => x"16",
          7414 => x"70",
          7415 => x"7a",
          7416 => x"0c",
          7417 => x"83",
          7418 => x"06",
          7419 => x"e2",
          7420 => x"c0",
          7421 => x"e4",
          7422 => x"ff",
          7423 => x"56",
          7424 => x"38",
          7425 => x"38",
          7426 => x"51",
          7427 => x"82",
          7428 => x"ac",
          7429 => x"82",
          7430 => x"39",
          7431 => x"80",
          7432 => x"38",
          7433 => x"15",
          7434 => x"53",
          7435 => x"8d",
          7436 => x"15",
          7437 => x"76",
          7438 => x"51",
          7439 => x"13",
          7440 => x"8d",
          7441 => x"15",
          7442 => x"cc",
          7443 => x"94",
          7444 => x"0b",
          7445 => x"ff",
          7446 => x"15",
          7447 => x"2e",
          7448 => x"81",
          7449 => x"e8",
          7450 => x"c8",
          7451 => x"e4",
          7452 => x"ff",
          7453 => x"81",
          7454 => x"06",
          7455 => x"81",
          7456 => x"51",
          7457 => x"82",
          7458 => x"80",
          7459 => x"d5",
          7460 => x"15",
          7461 => x"14",
          7462 => x"3f",
          7463 => x"08",
          7464 => x"06",
          7465 => x"d4",
          7466 => x"81",
          7467 => x"38",
          7468 => x"c6",
          7469 => x"d5",
          7470 => x"8b",
          7471 => x"2e",
          7472 => x"b3",
          7473 => x"14",
          7474 => x"3f",
          7475 => x"08",
          7476 => x"e4",
          7477 => x"81",
          7478 => x"84",
          7479 => x"c5",
          7480 => x"d5",
          7481 => x"15",
          7482 => x"14",
          7483 => x"3f",
          7484 => x"08",
          7485 => x"76",
          7486 => x"ed",
          7487 => x"05",
          7488 => x"ed",
          7489 => x"86",
          7490 => x"ed",
          7491 => x"15",
          7492 => x"98",
          7493 => x"56",
          7494 => x"e4",
          7495 => x"0d",
          7496 => x"0d",
          7497 => x"55",
          7498 => x"ba",
          7499 => x"53",
          7500 => x"b2",
          7501 => x"52",
          7502 => x"aa",
          7503 => x"22",
          7504 => x"57",
          7505 => x"2e",
          7506 => x"9a",
          7507 => x"33",
          7508 => x"ca",
          7509 => x"e4",
          7510 => x"52",
          7511 => x"71",
          7512 => x"55",
          7513 => x"53",
          7514 => x"0c",
          7515 => x"d5",
          7516 => x"3d",
          7517 => x"3d",
          7518 => x"05",
          7519 => x"89",
          7520 => x"52",
          7521 => x"3f",
          7522 => x"0b",
          7523 => x"08",
          7524 => x"82",
          7525 => x"84",
          7526 => x"ac",
          7527 => x"55",
          7528 => x"2e",
          7529 => x"74",
          7530 => x"73",
          7531 => x"38",
          7532 => x"78",
          7533 => x"54",
          7534 => x"92",
          7535 => x"89",
          7536 => x"84",
          7537 => x"e4",
          7538 => x"e4",
          7539 => x"82",
          7540 => x"88",
          7541 => x"ea",
          7542 => x"02",
          7543 => x"eb",
          7544 => x"59",
          7545 => x"80",
          7546 => x"38",
          7547 => x"70",
          7548 => x"cc",
          7549 => x"3d",
          7550 => x"58",
          7551 => x"82",
          7552 => x"55",
          7553 => x"08",
          7554 => x"7a",
          7555 => x"8c",
          7556 => x"56",
          7557 => x"82",
          7558 => x"55",
          7559 => x"08",
          7560 => x"80",
          7561 => x"70",
          7562 => x"57",
          7563 => x"83",
          7564 => x"77",
          7565 => x"73",
          7566 => x"ab",
          7567 => x"2e",
          7568 => x"84",
          7569 => x"06",
          7570 => x"51",
          7571 => x"82",
          7572 => x"55",
          7573 => x"b2",
          7574 => x"06",
          7575 => x"b8",
          7576 => x"2a",
          7577 => x"51",
          7578 => x"2e",
          7579 => x"55",
          7580 => x"77",
          7581 => x"74",
          7582 => x"77",
          7583 => x"81",
          7584 => x"73",
          7585 => x"af",
          7586 => x"7a",
          7587 => x"3f",
          7588 => x"08",
          7589 => x"b2",
          7590 => x"8e",
          7591 => x"f4",
          7592 => x"a0",
          7593 => x"34",
          7594 => x"52",
          7595 => x"85",
          7596 => x"62",
          7597 => x"c2",
          7598 => x"54",
          7599 => x"15",
          7600 => x"2e",
          7601 => x"7a",
          7602 => x"51",
          7603 => x"75",
          7604 => x"d0",
          7605 => x"86",
          7606 => x"e4",
          7607 => x"d5",
          7608 => x"ca",
          7609 => x"74",
          7610 => x"02",
          7611 => x"70",
          7612 => x"81",
          7613 => x"56",
          7614 => x"86",
          7615 => x"82",
          7616 => x"81",
          7617 => x"06",
          7618 => x"80",
          7619 => x"75",
          7620 => x"73",
          7621 => x"38",
          7622 => x"92",
          7623 => x"7a",
          7624 => x"3f",
          7625 => x"08",
          7626 => x"90",
          7627 => x"55",
          7628 => x"08",
          7629 => x"77",
          7630 => x"81",
          7631 => x"73",
          7632 => x"38",
          7633 => x"07",
          7634 => x"11",
          7635 => x"0c",
          7636 => x"0c",
          7637 => x"52",
          7638 => x"3f",
          7639 => x"08",
          7640 => x"08",
          7641 => x"63",
          7642 => x"5a",
          7643 => x"82",
          7644 => x"82",
          7645 => x"8c",
          7646 => x"7a",
          7647 => x"17",
          7648 => x"23",
          7649 => x"34",
          7650 => x"1a",
          7651 => x"9c",
          7652 => x"0b",
          7653 => x"77",
          7654 => x"81",
          7655 => x"73",
          7656 => x"8d",
          7657 => x"e4",
          7658 => x"81",
          7659 => x"d5",
          7660 => x"1a",
          7661 => x"22",
          7662 => x"7b",
          7663 => x"a8",
          7664 => x"78",
          7665 => x"3f",
          7666 => x"08",
          7667 => x"e4",
          7668 => x"83",
          7669 => x"82",
          7670 => x"ff",
          7671 => x"06",
          7672 => x"55",
          7673 => x"56",
          7674 => x"76",
          7675 => x"51",
          7676 => x"27",
          7677 => x"70",
          7678 => x"5a",
          7679 => x"76",
          7680 => x"74",
          7681 => x"83",
          7682 => x"73",
          7683 => x"38",
          7684 => x"51",
          7685 => x"82",
          7686 => x"85",
          7687 => x"8e",
          7688 => x"2a",
          7689 => x"08",
          7690 => x"0c",
          7691 => x"79",
          7692 => x"73",
          7693 => x"0c",
          7694 => x"04",
          7695 => x"60",
          7696 => x"40",
          7697 => x"80",
          7698 => x"3d",
          7699 => x"78",
          7700 => x"3f",
          7701 => x"08",
          7702 => x"e4",
          7703 => x"91",
          7704 => x"74",
          7705 => x"38",
          7706 => x"c7",
          7707 => x"33",
          7708 => x"87",
          7709 => x"2e",
          7710 => x"95",
          7711 => x"91",
          7712 => x"56",
          7713 => x"81",
          7714 => x"34",
          7715 => x"a3",
          7716 => x"08",
          7717 => x"31",
          7718 => x"27",
          7719 => x"5c",
          7720 => x"82",
          7721 => x"19",
          7722 => x"ff",
          7723 => x"74",
          7724 => x"7e",
          7725 => x"ff",
          7726 => x"2a",
          7727 => x"79",
          7728 => x"87",
          7729 => x"08",
          7730 => x"98",
          7731 => x"78",
          7732 => x"3f",
          7733 => x"08",
          7734 => x"27",
          7735 => x"74",
          7736 => x"a3",
          7737 => x"1a",
          7738 => x"08",
          7739 => x"c3",
          7740 => x"d5",
          7741 => x"2e",
          7742 => x"82",
          7743 => x"1a",
          7744 => x"59",
          7745 => x"2e",
          7746 => x"77",
          7747 => x"11",
          7748 => x"55",
          7749 => x"85",
          7750 => x"31",
          7751 => x"76",
          7752 => x"81",
          7753 => x"ff",
          7754 => x"82",
          7755 => x"fe",
          7756 => x"83",
          7757 => x"56",
          7758 => x"a0",
          7759 => x"08",
          7760 => x"74",
          7761 => x"38",
          7762 => x"b8",
          7763 => x"16",
          7764 => x"89",
          7765 => x"51",
          7766 => x"3f",
          7767 => x"56",
          7768 => x"9c",
          7769 => x"19",
          7770 => x"06",
          7771 => x"31",
          7772 => x"76",
          7773 => x"7b",
          7774 => x"08",
          7775 => x"c0",
          7776 => x"d5",
          7777 => x"ff",
          7778 => x"94",
          7779 => x"ff",
          7780 => x"05",
          7781 => x"ff",
          7782 => x"7b",
          7783 => x"08",
          7784 => x"76",
          7785 => x"08",
          7786 => x"0c",
          7787 => x"f0",
          7788 => x"75",
          7789 => x"0c",
          7790 => x"04",
          7791 => x"60",
          7792 => x"40",
          7793 => x"80",
          7794 => x"3d",
          7795 => x"77",
          7796 => x"3f",
          7797 => x"08",
          7798 => x"e4",
          7799 => x"91",
          7800 => x"74",
          7801 => x"38",
          7802 => x"bf",
          7803 => x"33",
          7804 => x"70",
          7805 => x"56",
          7806 => x"74",
          7807 => x"ab",
          7808 => x"82",
          7809 => x"34",
          7810 => x"9f",
          7811 => x"91",
          7812 => x"56",
          7813 => x"94",
          7814 => x"11",
          7815 => x"76",
          7816 => x"75",
          7817 => x"80",
          7818 => x"38",
          7819 => x"70",
          7820 => x"56",
          7821 => x"82",
          7822 => x"11",
          7823 => x"77",
          7824 => x"5c",
          7825 => x"38",
          7826 => x"88",
          7827 => x"74",
          7828 => x"52",
          7829 => x"18",
          7830 => x"51",
          7831 => x"82",
          7832 => x"55",
          7833 => x"08",
          7834 => x"b2",
          7835 => x"2e",
          7836 => x"74",
          7837 => x"95",
          7838 => x"19",
          7839 => x"08",
          7840 => x"88",
          7841 => x"55",
          7842 => x"9c",
          7843 => x"09",
          7844 => x"38",
          7845 => x"bd",
          7846 => x"d5",
          7847 => x"ed",
          7848 => x"08",
          7849 => x"ff",
          7850 => x"82",
          7851 => x"80",
          7852 => x"38",
          7853 => x"08",
          7854 => x"2a",
          7855 => x"80",
          7856 => x"38",
          7857 => x"8a",
          7858 => x"5b",
          7859 => x"27",
          7860 => x"7b",
          7861 => x"54",
          7862 => x"52",
          7863 => x"51",
          7864 => x"3f",
          7865 => x"08",
          7866 => x"7e",
          7867 => x"78",
          7868 => x"74",
          7869 => x"38",
          7870 => x"b4",
          7871 => x"31",
          7872 => x"05",
          7873 => x"51",
          7874 => x"3f",
          7875 => x"0b",
          7876 => x"78",
          7877 => x"80",
          7878 => x"18",
          7879 => x"08",
          7880 => x"7e",
          7881 => x"f6",
          7882 => x"e4",
          7883 => x"38",
          7884 => x"12",
          7885 => x"9c",
          7886 => x"18",
          7887 => x"06",
          7888 => x"31",
          7889 => x"76",
          7890 => x"7b",
          7891 => x"08",
          7892 => x"ff",
          7893 => x"82",
          7894 => x"fd",
          7895 => x"53",
          7896 => x"18",
          7897 => x"06",
          7898 => x"51",
          7899 => x"3f",
          7900 => x"0b",
          7901 => x"7b",
          7902 => x"08",
          7903 => x"76",
          7904 => x"08",
          7905 => x"1c",
          7906 => x"08",
          7907 => x"5c",
          7908 => x"83",
          7909 => x"74",
          7910 => x"fd",
          7911 => x"18",
          7912 => x"07",
          7913 => x"19",
          7914 => x"75",
          7915 => x"0c",
          7916 => x"04",
          7917 => x"7a",
          7918 => x"05",
          7919 => x"56",
          7920 => x"82",
          7921 => x"57",
          7922 => x"08",
          7923 => x"90",
          7924 => x"86",
          7925 => x"06",
          7926 => x"73",
          7927 => x"ee",
          7928 => x"08",
          7929 => x"ff",
          7930 => x"82",
          7931 => x"57",
          7932 => x"08",
          7933 => x"a4",
          7934 => x"11",
          7935 => x"55",
          7936 => x"16",
          7937 => x"08",
          7938 => x"75",
          7939 => x"a5",
          7940 => x"08",
          7941 => x"51",
          7942 => x"3f",
          7943 => x"0a",
          7944 => x"51",
          7945 => x"3f",
          7946 => x"15",
          7947 => x"c6",
          7948 => x"81",
          7949 => x"34",
          7950 => x"bb",
          7951 => x"d5",
          7952 => x"17",
          7953 => x"06",
          7954 => x"90",
          7955 => x"82",
          7956 => x"8a",
          7957 => x"fc",
          7958 => x"70",
          7959 => x"d4",
          7960 => x"e4",
          7961 => x"d5",
          7962 => x"38",
          7963 => x"05",
          7964 => x"f1",
          7965 => x"d5",
          7966 => x"82",
          7967 => x"87",
          7968 => x"e4",
          7969 => x"72",
          7970 => x"0c",
          7971 => x"04",
          7972 => x"84",
          7973 => x"89",
          7974 => x"80",
          7975 => x"e4",
          7976 => x"38",
          7977 => x"08",
          7978 => x"34",
          7979 => x"82",
          7980 => x"83",
          7981 => x"ee",
          7982 => x"53",
          7983 => x"05",
          7984 => x"51",
          7985 => x"82",
          7986 => x"55",
          7987 => x"08",
          7988 => x"76",
          7989 => x"94",
          7990 => x"51",
          7991 => x"82",
          7992 => x"55",
          7993 => x"08",
          7994 => x"80",
          7995 => x"70",
          7996 => x"56",
          7997 => x"89",
          7998 => x"98",
          7999 => x"b2",
          8000 => x"05",
          8001 => x"2a",
          8002 => x"51",
          8003 => x"80",
          8004 => x"76",
          8005 => x"52",
          8006 => x"3f",
          8007 => x"08",
          8008 => x"8e",
          8009 => x"e4",
          8010 => x"09",
          8011 => x"38",
          8012 => x"82",
          8013 => x"94",
          8014 => x"ff",
          8015 => x"80",
          8016 => x"80",
          8017 => x"5b",
          8018 => x"34",
          8019 => x"df",
          8020 => x"05",
          8021 => x"3d",
          8022 => x"3f",
          8023 => x"08",
          8024 => x"e4",
          8025 => x"38",
          8026 => x"3d",
          8027 => x"98",
          8028 => x"d8",
          8029 => x"58",
          8030 => x"08",
          8031 => x"2e",
          8032 => x"a0",
          8033 => x"3d",
          8034 => x"c4",
          8035 => x"d5",
          8036 => x"82",
          8037 => x"82",
          8038 => x"d9",
          8039 => x"7b",
          8040 => x"ea",
          8041 => x"e4",
          8042 => x"d5",
          8043 => x"d8",
          8044 => x"3d",
          8045 => x"51",
          8046 => x"82",
          8047 => x"80",
          8048 => x"76",
          8049 => x"c3",
          8050 => x"d5",
          8051 => x"82",
          8052 => x"82",
          8053 => x"52",
          8054 => x"b6",
          8055 => x"e4",
          8056 => x"d5",
          8057 => x"38",
          8058 => x"08",
          8059 => x"c8",
          8060 => x"82",
          8061 => x"2e",
          8062 => x"52",
          8063 => x"e8",
          8064 => x"e4",
          8065 => x"d5",
          8066 => x"2e",
          8067 => x"84",
          8068 => x"06",
          8069 => x"57",
          8070 => x"76",
          8071 => x"80",
          8072 => x"b8",
          8073 => x"51",
          8074 => x"76",
          8075 => x"11",
          8076 => x"51",
          8077 => x"73",
          8078 => x"38",
          8079 => x"05",
          8080 => x"81",
          8081 => x"56",
          8082 => x"f5",
          8083 => x"54",
          8084 => x"81",
          8085 => x"80",
          8086 => x"78",
          8087 => x"55",
          8088 => x"e1",
          8089 => x"ff",
          8090 => x"58",
          8091 => x"74",
          8092 => x"75",
          8093 => x"18",
          8094 => x"08",
          8095 => x"af",
          8096 => x"f4",
          8097 => x"2e",
          8098 => x"8d",
          8099 => x"80",
          8100 => x"11",
          8101 => x"74",
          8102 => x"82",
          8103 => x"70",
          8104 => x"c7",
          8105 => x"08",
          8106 => x"5c",
          8107 => x"73",
          8108 => x"38",
          8109 => x"1a",
          8110 => x"55",
          8111 => x"38",
          8112 => x"73",
          8113 => x"38",
          8114 => x"76",
          8115 => x"74",
          8116 => x"33",
          8117 => x"05",
          8118 => x"15",
          8119 => x"ba",
          8120 => x"05",
          8121 => x"ff",
          8122 => x"06",
          8123 => x"57",
          8124 => x"e0",
          8125 => x"81",
          8126 => x"73",
          8127 => x"81",
          8128 => x"7a",
          8129 => x"38",
          8130 => x"76",
          8131 => x"0c",
          8132 => x"0d",
          8133 => x"0d",
          8134 => x"3d",
          8135 => x"71",
          8136 => x"eb",
          8137 => x"d5",
          8138 => x"82",
          8139 => x"82",
          8140 => x"15",
          8141 => x"82",
          8142 => x"15",
          8143 => x"76",
          8144 => x"90",
          8145 => x"81",
          8146 => x"06",
          8147 => x"72",
          8148 => x"56",
          8149 => x"54",
          8150 => x"17",
          8151 => x"78",
          8152 => x"38",
          8153 => x"22",
          8154 => x"59",
          8155 => x"78",
          8156 => x"76",
          8157 => x"51",
          8158 => x"3f",
          8159 => x"08",
          8160 => x"54",
          8161 => x"53",
          8162 => x"3f",
          8163 => x"08",
          8164 => x"38",
          8165 => x"75",
          8166 => x"18",
          8167 => x"31",
          8168 => x"57",
          8169 => x"b2",
          8170 => x"08",
          8171 => x"38",
          8172 => x"51",
          8173 => x"3f",
          8174 => x"08",
          8175 => x"e4",
          8176 => x"81",
          8177 => x"d5",
          8178 => x"2e",
          8179 => x"82",
          8180 => x"88",
          8181 => x"98",
          8182 => x"80",
          8183 => x"38",
          8184 => x"80",
          8185 => x"77",
          8186 => x"08",
          8187 => x"0c",
          8188 => x"70",
          8189 => x"81",
          8190 => x"5a",
          8191 => x"2e",
          8192 => x"52",
          8193 => x"bb",
          8194 => x"d5",
          8195 => x"82",
          8196 => x"95",
          8197 => x"e4",
          8198 => x"39",
          8199 => x"51",
          8200 => x"3f",
          8201 => x"08",
          8202 => x"2e",
          8203 => x"74",
          8204 => x"79",
          8205 => x"14",
          8206 => x"38",
          8207 => x"0c",
          8208 => x"94",
          8209 => x"94",
          8210 => x"83",
          8211 => x"72",
          8212 => x"38",
          8213 => x"51",
          8214 => x"3f",
          8215 => x"08",
          8216 => x"0b",
          8217 => x"82",
          8218 => x"39",
          8219 => x"16",
          8220 => x"bb",
          8221 => x"2a",
          8222 => x"08",
          8223 => x"15",
          8224 => x"15",
          8225 => x"90",
          8226 => x"16",
          8227 => x"33",
          8228 => x"53",
          8229 => x"34",
          8230 => x"06",
          8231 => x"2e",
          8232 => x"9c",
          8233 => x"85",
          8234 => x"16",
          8235 => x"72",
          8236 => x"0c",
          8237 => x"04",
          8238 => x"79",
          8239 => x"75",
          8240 => x"8b",
          8241 => x"89",
          8242 => x"52",
          8243 => x"05",
          8244 => x"3f",
          8245 => x"08",
          8246 => x"e4",
          8247 => x"38",
          8248 => x"7a",
          8249 => x"d4",
          8250 => x"d5",
          8251 => x"82",
          8252 => x"80",
          8253 => x"16",
          8254 => x"2b",
          8255 => x"74",
          8256 => x"86",
          8257 => x"84",
          8258 => x"06",
          8259 => x"73",
          8260 => x"38",
          8261 => x"52",
          8262 => x"e0",
          8263 => x"e4",
          8264 => x"0c",
          8265 => x"14",
          8266 => x"23",
          8267 => x"51",
          8268 => x"3f",
          8269 => x"08",
          8270 => x"2e",
          8271 => x"85",
          8272 => x"86",
          8273 => x"2e",
          8274 => x"76",
          8275 => x"73",
          8276 => x"0c",
          8277 => x"04",
          8278 => x"76",
          8279 => x"05",
          8280 => x"53",
          8281 => x"82",
          8282 => x"87",
          8283 => x"e4",
          8284 => x"86",
          8285 => x"fb",
          8286 => x"79",
          8287 => x"05",
          8288 => x"56",
          8289 => x"3f",
          8290 => x"08",
          8291 => x"e4",
          8292 => x"38",
          8293 => x"82",
          8294 => x"52",
          8295 => x"bb",
          8296 => x"d5",
          8297 => x"80",
          8298 => x"d5",
          8299 => x"73",
          8300 => x"3f",
          8301 => x"08",
          8302 => x"e4",
          8303 => x"09",
          8304 => x"38",
          8305 => x"39",
          8306 => x"08",
          8307 => x"52",
          8308 => x"f6",
          8309 => x"73",
          8310 => x"8c",
          8311 => x"e4",
          8312 => x"70",
          8313 => x"07",
          8314 => x"82",
          8315 => x"06",
          8316 => x"54",
          8317 => x"e4",
          8318 => x"0d",
          8319 => x"0d",
          8320 => x"53",
          8321 => x"53",
          8322 => x"56",
          8323 => x"82",
          8324 => x"55",
          8325 => x"08",
          8326 => x"52",
          8327 => x"a6",
          8328 => x"e4",
          8329 => x"d5",
          8330 => x"38",
          8331 => x"05",
          8332 => x"2b",
          8333 => x"80",
          8334 => x"86",
          8335 => x"76",
          8336 => x"38",
          8337 => x"51",
          8338 => x"74",
          8339 => x"0c",
          8340 => x"04",
          8341 => x"63",
          8342 => x"80",
          8343 => x"ec",
          8344 => x"3d",
          8345 => x"3f",
          8346 => x"08",
          8347 => x"e4",
          8348 => x"38",
          8349 => x"73",
          8350 => x"08",
          8351 => x"13",
          8352 => x"58",
          8353 => x"26",
          8354 => x"7c",
          8355 => x"39",
          8356 => x"ce",
          8357 => x"81",
          8358 => x"d5",
          8359 => x"33",
          8360 => x"81",
          8361 => x"06",
          8362 => x"82",
          8363 => x"76",
          8364 => x"f0",
          8365 => x"af",
          8366 => x"d5",
          8367 => x"2e",
          8368 => x"d5",
          8369 => x"2e",
          8370 => x"d5",
          8371 => x"70",
          8372 => x"08",
          8373 => x"7a",
          8374 => x"7f",
          8375 => x"54",
          8376 => x"77",
          8377 => x"80",
          8378 => x"15",
          8379 => x"e4",
          8380 => x"75",
          8381 => x"52",
          8382 => x"52",
          8383 => x"8e",
          8384 => x"e4",
          8385 => x"d5",
          8386 => x"d6",
          8387 => x"33",
          8388 => x"1a",
          8389 => x"54",
          8390 => x"09",
          8391 => x"38",
          8392 => x"ff",
          8393 => x"82",
          8394 => x"83",
          8395 => x"70",
          8396 => x"25",
          8397 => x"59",
          8398 => x"9b",
          8399 => x"51",
          8400 => x"3f",
          8401 => x"08",
          8402 => x"70",
          8403 => x"25",
          8404 => x"59",
          8405 => x"75",
          8406 => x"7a",
          8407 => x"ff",
          8408 => x"7c",
          8409 => x"94",
          8410 => x"11",
          8411 => x"56",
          8412 => x"15",
          8413 => x"d5",
          8414 => x"3d",
          8415 => x"3d",
          8416 => x"3d",
          8417 => x"70",
          8418 => x"95",
          8419 => x"e4",
          8420 => x"d5",
          8421 => x"aa",
          8422 => x"33",
          8423 => x"a2",
          8424 => x"33",
          8425 => x"70",
          8426 => x"55",
          8427 => x"73",
          8428 => x"90",
          8429 => x"08",
          8430 => x"18",
          8431 => x"82",
          8432 => x"38",
          8433 => x"08",
          8434 => x"08",
          8435 => x"ff",
          8436 => x"82",
          8437 => x"74",
          8438 => x"56",
          8439 => x"98",
          8440 => x"76",
          8441 => x"c6",
          8442 => x"e4",
          8443 => x"09",
          8444 => x"38",
          8445 => x"d5",
          8446 => x"2e",
          8447 => x"85",
          8448 => x"a4",
          8449 => x"38",
          8450 => x"d5",
          8451 => x"15",
          8452 => x"38",
          8453 => x"53",
          8454 => x"08",
          8455 => x"ff",
          8456 => x"82",
          8457 => x"56",
          8458 => x"8c",
          8459 => x"17",
          8460 => x"07",
          8461 => x"18",
          8462 => x"2e",
          8463 => x"91",
          8464 => x"55",
          8465 => x"e4",
          8466 => x"0d",
          8467 => x"0d",
          8468 => x"3d",
          8469 => x"52",
          8470 => x"d9",
          8471 => x"d5",
          8472 => x"82",
          8473 => x"81",
          8474 => x"46",
          8475 => x"52",
          8476 => x"52",
          8477 => x"3f",
          8478 => x"08",
          8479 => x"e4",
          8480 => x"38",
          8481 => x"05",
          8482 => x"2a",
          8483 => x"51",
          8484 => x"55",
          8485 => x"38",
          8486 => x"54",
          8487 => x"81",
          8488 => x"80",
          8489 => x"70",
          8490 => x"54",
          8491 => x"81",
          8492 => x"52",
          8493 => x"ba",
          8494 => x"d5",
          8495 => x"84",
          8496 => x"06",
          8497 => x"73",
          8498 => x"d6",
          8499 => x"82",
          8500 => x"98",
          8501 => x"81",
          8502 => x"5a",
          8503 => x"08",
          8504 => x"8a",
          8505 => x"54",
          8506 => x"3f",
          8507 => x"08",
          8508 => x"e4",
          8509 => x"38",
          8510 => x"08",
          8511 => x"ff",
          8512 => x"82",
          8513 => x"55",
          8514 => x"08",
          8515 => x"55",
          8516 => x"82",
          8517 => x"84",
          8518 => x"82",
          8519 => x"80",
          8520 => x"51",
          8521 => x"82",
          8522 => x"82",
          8523 => x"30",
          8524 => x"e4",
          8525 => x"25",
          8526 => x"75",
          8527 => x"38",
          8528 => x"90",
          8529 => x"75",
          8530 => x"ff",
          8531 => x"82",
          8532 => x"55",
          8533 => x"78",
          8534 => x"f9",
          8535 => x"e4",
          8536 => x"82",
          8537 => x"a2",
          8538 => x"e8",
          8539 => x"53",
          8540 => x"bc",
          8541 => x"3d",
          8542 => x"3f",
          8543 => x"08",
          8544 => x"e4",
          8545 => x"38",
          8546 => x"52",
          8547 => x"52",
          8548 => x"3f",
          8549 => x"08",
          8550 => x"e4",
          8551 => x"88",
          8552 => x"39",
          8553 => x"08",
          8554 => x"81",
          8555 => x"38",
          8556 => x"05",
          8557 => x"2a",
          8558 => x"55",
          8559 => x"81",
          8560 => x"5a",
          8561 => x"3d",
          8562 => x"ff",
          8563 => x"82",
          8564 => x"75",
          8565 => x"d5",
          8566 => x"38",
          8567 => x"d5",
          8568 => x"2e",
          8569 => x"83",
          8570 => x"82",
          8571 => x"ff",
          8572 => x"06",
          8573 => x"54",
          8574 => x"73",
          8575 => x"82",
          8576 => x"52",
          8577 => x"b2",
          8578 => x"d5",
          8579 => x"82",
          8580 => x"81",
          8581 => x"53",
          8582 => x"19",
          8583 => x"c6",
          8584 => x"ae",
          8585 => x"34",
          8586 => x"0b",
          8587 => x"34",
          8588 => x"0a",
          8589 => x"19",
          8590 => x"d8",
          8591 => x"78",
          8592 => x"51",
          8593 => x"3f",
          8594 => x"b8",
          8595 => x"d8",
          8596 => x"a3",
          8597 => x"54",
          8598 => x"d9",
          8599 => x"53",
          8600 => x"11",
          8601 => x"b7",
          8602 => x"54",
          8603 => x"15",
          8604 => x"ff",
          8605 => x"82",
          8606 => x"54",
          8607 => x"08",
          8608 => x"88",
          8609 => x"64",
          8610 => x"ff",
          8611 => x"75",
          8612 => x"78",
          8613 => x"9d",
          8614 => x"90",
          8615 => x"34",
          8616 => x"0b",
          8617 => x"78",
          8618 => x"a9",
          8619 => x"e4",
          8620 => x"39",
          8621 => x"52",
          8622 => x"ac",
          8623 => x"82",
          8624 => x"9a",
          8625 => x"d8",
          8626 => x"3d",
          8627 => x"d1",
          8628 => x"53",
          8629 => x"fc",
          8630 => x"3d",
          8631 => x"3f",
          8632 => x"08",
          8633 => x"e4",
          8634 => x"38",
          8635 => x"3d",
          8636 => x"3d",
          8637 => x"c8",
          8638 => x"d5",
          8639 => x"82",
          8640 => x"82",
          8641 => x"81",
          8642 => x"81",
          8643 => x"86",
          8644 => x"af",
          8645 => x"a5",
          8646 => x"aa",
          8647 => x"05",
          8648 => x"9f",
          8649 => x"77",
          8650 => x"70",
          8651 => x"a2",
          8652 => x"3d",
          8653 => x"51",
          8654 => x"82",
          8655 => x"55",
          8656 => x"08",
          8657 => x"a1",
          8658 => x"09",
          8659 => x"38",
          8660 => x"08",
          8661 => x"88",
          8662 => x"39",
          8663 => x"08",
          8664 => x"81",
          8665 => x"38",
          8666 => x"bd",
          8667 => x"d5",
          8668 => x"82",
          8669 => x"81",
          8670 => x"56",
          8671 => x"3d",
          8672 => x"52",
          8673 => x"ff",
          8674 => x"02",
          8675 => x"8b",
          8676 => x"16",
          8677 => x"2a",
          8678 => x"51",
          8679 => x"89",
          8680 => x"07",
          8681 => x"17",
          8682 => x"81",
          8683 => x"34",
          8684 => x"70",
          8685 => x"81",
          8686 => x"55",
          8687 => x"80",
          8688 => x"64",
          8689 => x"38",
          8690 => x"51",
          8691 => x"3f",
          8692 => x"08",
          8693 => x"ff",
          8694 => x"82",
          8695 => x"e4",
          8696 => x"80",
          8697 => x"d5",
          8698 => x"78",
          8699 => x"9e",
          8700 => x"e4",
          8701 => x"d8",
          8702 => x"55",
          8703 => x"08",
          8704 => x"81",
          8705 => x"73",
          8706 => x"81",
          8707 => x"63",
          8708 => x"76",
          8709 => x"9d",
          8710 => x"81",
          8711 => x"34",
          8712 => x"d5",
          8713 => x"38",
          8714 => x"a5",
          8715 => x"e4",
          8716 => x"d5",
          8717 => x"38",
          8718 => x"a3",
          8719 => x"d5",
          8720 => x"74",
          8721 => x"0c",
          8722 => x"04",
          8723 => x"02",
          8724 => x"33",
          8725 => x"80",
          8726 => x"57",
          8727 => x"96",
          8728 => x"52",
          8729 => x"d1",
          8730 => x"d5",
          8731 => x"82",
          8732 => x"80",
          8733 => x"5a",
          8734 => x"3d",
          8735 => x"c5",
          8736 => x"d5",
          8737 => x"82",
          8738 => x"b8",
          8739 => x"cf",
          8740 => x"a0",
          8741 => x"55",
          8742 => x"75",
          8743 => x"71",
          8744 => x"33",
          8745 => x"74",
          8746 => x"57",
          8747 => x"8b",
          8748 => x"54",
          8749 => x"15",
          8750 => x"ff",
          8751 => x"82",
          8752 => x"55",
          8753 => x"e4",
          8754 => x"0d",
          8755 => x"0d",
          8756 => x"53",
          8757 => x"05",
          8758 => x"51",
          8759 => x"82",
          8760 => x"55",
          8761 => x"08",
          8762 => x"76",
          8763 => x"94",
          8764 => x"51",
          8765 => x"82",
          8766 => x"55",
          8767 => x"08",
          8768 => x"80",
          8769 => x"81",
          8770 => x"86",
          8771 => x"38",
          8772 => x"86",
          8773 => x"90",
          8774 => x"54",
          8775 => x"ff",
          8776 => x"76",
          8777 => x"83",
          8778 => x"51",
          8779 => x"3f",
          8780 => x"08",
          8781 => x"d5",
          8782 => x"3d",
          8783 => x"3d",
          8784 => x"5c",
          8785 => x"99",
          8786 => x"52",
          8787 => x"cf",
          8788 => x"d5",
          8789 => x"d5",
          8790 => x"70",
          8791 => x"08",
          8792 => x"51",
          8793 => x"80",
          8794 => x"38",
          8795 => x"06",
          8796 => x"80",
          8797 => x"38",
          8798 => x"5f",
          8799 => x"3d",
          8800 => x"ff",
          8801 => x"82",
          8802 => x"57",
          8803 => x"08",
          8804 => x"74",
          8805 => x"ff",
          8806 => x"82",
          8807 => x"57",
          8808 => x"08",
          8809 => x"d5",
          8810 => x"d5",
          8811 => x"5b",
          8812 => x"18",
          8813 => x"18",
          8814 => x"74",
          8815 => x"81",
          8816 => x"78",
          8817 => x"8b",
          8818 => x"54",
          8819 => x"75",
          8820 => x"38",
          8821 => x"1b",
          8822 => x"55",
          8823 => x"2e",
          8824 => x"39",
          8825 => x"09",
          8826 => x"38",
          8827 => x"80",
          8828 => x"70",
          8829 => x"25",
          8830 => x"80",
          8831 => x"38",
          8832 => x"bc",
          8833 => x"11",
          8834 => x"ff",
          8835 => x"82",
          8836 => x"57",
          8837 => x"08",
          8838 => x"70",
          8839 => x"80",
          8840 => x"83",
          8841 => x"80",
          8842 => x"84",
          8843 => x"a7",
          8844 => x"b8",
          8845 => x"9b",
          8846 => x"d5",
          8847 => x"0c",
          8848 => x"e4",
          8849 => x"0d",
          8850 => x"0d",
          8851 => x"3d",
          8852 => x"52",
          8853 => x"cd",
          8854 => x"d5",
          8855 => x"d5",
          8856 => x"54",
          8857 => x"08",
          8858 => x"8b",
          8859 => x"8a",
          8860 => x"58",
          8861 => x"3f",
          8862 => x"33",
          8863 => x"9f",
          8864 => x"86",
          8865 => x"9d",
          8866 => x"9c",
          8867 => x"d5",
          8868 => x"ff",
          8869 => x"c4",
          8870 => x"e4",
          8871 => x"c0",
          8872 => x"52",
          8873 => x"08",
          8874 => x"3f",
          8875 => x"08",
          8876 => x"06",
          8877 => x"2e",
          8878 => x"52",
          8879 => x"51",
          8880 => x"3f",
          8881 => x"08",
          8882 => x"ff",
          8883 => x"38",
          8884 => x"88",
          8885 => x"8a",
          8886 => x"38",
          8887 => x"e7",
          8888 => x"75",
          8889 => x"74",
          8890 => x"73",
          8891 => x"05",
          8892 => x"16",
          8893 => x"70",
          8894 => x"34",
          8895 => x"70",
          8896 => x"56",
          8897 => x"fe",
          8898 => x"3d",
          8899 => x"55",
          8900 => x"2e",
          8901 => x"75",
          8902 => x"38",
          8903 => x"55",
          8904 => x"33",
          8905 => x"a0",
          8906 => x"06",
          8907 => x"16",
          8908 => x"38",
          8909 => x"42",
          8910 => x"3d",
          8911 => x"ff",
          8912 => x"82",
          8913 => x"54",
          8914 => x"08",
          8915 => x"81",
          8916 => x"ff",
          8917 => x"82",
          8918 => x"54",
          8919 => x"08",
          8920 => x"80",
          8921 => x"54",
          8922 => x"80",
          8923 => x"d5",
          8924 => x"2e",
          8925 => x"80",
          8926 => x"54",
          8927 => x"80",
          8928 => x"52",
          8929 => x"ab",
          8930 => x"d5",
          8931 => x"82",
          8932 => x"b1",
          8933 => x"82",
          8934 => x"52",
          8935 => x"99",
          8936 => x"54",
          8937 => x"15",
          8938 => x"77",
          8939 => x"ff",
          8940 => x"78",
          8941 => x"83",
          8942 => x"51",
          8943 => x"3f",
          8944 => x"08",
          8945 => x"74",
          8946 => x"0c",
          8947 => x"04",
          8948 => x"60",
          8949 => x"05",
          8950 => x"33",
          8951 => x"05",
          8952 => x"40",
          8953 => x"b9",
          8954 => x"e4",
          8955 => x"d5",
          8956 => x"bd",
          8957 => x"33",
          8958 => x"b5",
          8959 => x"2e",
          8960 => x"1a",
          8961 => x"90",
          8962 => x"33",
          8963 => x"70",
          8964 => x"55",
          8965 => x"38",
          8966 => x"97",
          8967 => x"82",
          8968 => x"58",
          8969 => x"7e",
          8970 => x"70",
          8971 => x"55",
          8972 => x"56",
          8973 => x"f6",
          8974 => x"7d",
          8975 => x"70",
          8976 => x"2a",
          8977 => x"08",
          8978 => x"08",
          8979 => x"5d",
          8980 => x"77",
          8981 => x"9c",
          8982 => x"26",
          8983 => x"57",
          8984 => x"59",
          8985 => x"52",
          8986 => x"9c",
          8987 => x"15",
          8988 => x"9c",
          8989 => x"26",
          8990 => x"55",
          8991 => x"08",
          8992 => x"99",
          8993 => x"e4",
          8994 => x"ff",
          8995 => x"d5",
          8996 => x"38",
          8997 => x"75",
          8998 => x"81",
          8999 => x"93",
          9000 => x"80",
          9001 => x"2e",
          9002 => x"ff",
          9003 => x"58",
          9004 => x"7d",
          9005 => x"38",
          9006 => x"55",
          9007 => x"b4",
          9008 => x"56",
          9009 => x"09",
          9010 => x"38",
          9011 => x"53",
          9012 => x"51",
          9013 => x"3f",
          9014 => x"08",
          9015 => x"e4",
          9016 => x"38",
          9017 => x"ff",
          9018 => x"5c",
          9019 => x"84",
          9020 => x"5c",
          9021 => x"12",
          9022 => x"80",
          9023 => x"78",
          9024 => x"7c",
          9025 => x"90",
          9026 => x"c0",
          9027 => x"90",
          9028 => x"15",
          9029 => x"94",
          9030 => x"54",
          9031 => x"91",
          9032 => x"31",
          9033 => x"84",
          9034 => x"07",
          9035 => x"16",
          9036 => x"73",
          9037 => x"0c",
          9038 => x"04",
          9039 => x"6c",
          9040 => x"05",
          9041 => x"33",
          9042 => x"45",
          9043 => x"d1",
          9044 => x"80",
          9045 => x"e4",
          9046 => x"a0",
          9047 => x"e4",
          9048 => x"82",
          9049 => x"70",
          9050 => x"74",
          9051 => x"38",
          9052 => x"82",
          9053 => x"82",
          9054 => x"05",
          9055 => x"11",
          9056 => x"d9",
          9057 => x"41",
          9058 => x"7f",
          9059 => x"ac",
          9060 => x"e4",
          9061 => x"06",
          9062 => x"56",
          9063 => x"74",
          9064 => x"76",
          9065 => x"81",
          9066 => x"8a",
          9067 => x"cc",
          9068 => x"fc",
          9069 => x"52",
          9070 => x"92",
          9071 => x"d5",
          9072 => x"38",
          9073 => x"80",
          9074 => x"74",
          9075 => x"26",
          9076 => x"15",
          9077 => x"74",
          9078 => x"38",
          9079 => x"80",
          9080 => x"84",
          9081 => x"92",
          9082 => x"80",
          9083 => x"38",
          9084 => x"06",
          9085 => x"2e",
          9086 => x"56",
          9087 => x"78",
          9088 => x"89",
          9089 => x"2b",
          9090 => x"43",
          9091 => x"38",
          9092 => x"30",
          9093 => x"77",
          9094 => x"91",
          9095 => x"dc",
          9096 => x"2e",
          9097 => x"81",
          9098 => x"7a",
          9099 => x"ff",
          9100 => x"81",
          9101 => x"e4",
          9102 => x"38",
          9103 => x"51",
          9104 => x"3f",
          9105 => x"08",
          9106 => x"06",
          9107 => x"74",
          9108 => x"2e",
          9109 => x"8b",
          9110 => x"90",
          9111 => x"b2",
          9112 => x"57",
          9113 => x"8b",
          9114 => x"b6",
          9115 => x"92",
          9116 => x"d5",
          9117 => x"ba",
          9118 => x"ff",
          9119 => x"82",
          9120 => x"48",
          9121 => x"3d",
          9122 => x"81",
          9123 => x"ff",
          9124 => x"81",
          9125 => x"e4",
          9126 => x"38",
          9127 => x"70",
          9128 => x"d5",
          9129 => x"51",
          9130 => x"38",
          9131 => x"55",
          9132 => x"75",
          9133 => x"38",
          9134 => x"48",
          9135 => x"ff",
          9136 => x"b8",
          9137 => x"78",
          9138 => x"8a",
          9139 => x"81",
          9140 => x"06",
          9141 => x"80",
          9142 => x"62",
          9143 => x"74",
          9144 => x"8d",
          9145 => x"06",
          9146 => x"2e",
          9147 => x"62",
          9148 => x"93",
          9149 => x"74",
          9150 => x"80",
          9151 => x"7d",
          9152 => x"81",
          9153 => x"38",
          9154 => x"67",
          9155 => x"81",
          9156 => x"98",
          9157 => x"74",
          9158 => x"38",
          9159 => x"98",
          9160 => x"98",
          9161 => x"82",
          9162 => x"57",
          9163 => x"80",
          9164 => x"76",
          9165 => x"38",
          9166 => x"51",
          9167 => x"3f",
          9168 => x"08",
          9169 => x"87",
          9170 => x"2a",
          9171 => x"5c",
          9172 => x"d5",
          9173 => x"80",
          9174 => x"46",
          9175 => x"0a",
          9176 => x"ec",
          9177 => x"39",
          9178 => x"67",
          9179 => x"81",
          9180 => x"88",
          9181 => x"74",
          9182 => x"38",
          9183 => x"98",
          9184 => x"88",
          9185 => x"82",
          9186 => x"57",
          9187 => x"80",
          9188 => x"76",
          9189 => x"38",
          9190 => x"51",
          9191 => x"3f",
          9192 => x"08",
          9193 => x"57",
          9194 => x"08",
          9195 => x"96",
          9196 => x"82",
          9197 => x"10",
          9198 => x"08",
          9199 => x"72",
          9200 => x"59",
          9201 => x"ff",
          9202 => x"5d",
          9203 => x"46",
          9204 => x"11",
          9205 => x"70",
          9206 => x"71",
          9207 => x"06",
          9208 => x"52",
          9209 => x"41",
          9210 => x"09",
          9211 => x"38",
          9212 => x"18",
          9213 => x"39",
          9214 => x"79",
          9215 => x"70",
          9216 => x"58",
          9217 => x"76",
          9218 => x"38",
          9219 => x"7d",
          9220 => x"70",
          9221 => x"55",
          9222 => x"3f",
          9223 => x"08",
          9224 => x"2e",
          9225 => x"9b",
          9226 => x"e4",
          9227 => x"f5",
          9228 => x"38",
          9229 => x"38",
          9230 => x"59",
          9231 => x"38",
          9232 => x"7d",
          9233 => x"81",
          9234 => x"38",
          9235 => x"0b",
          9236 => x"08",
          9237 => x"78",
          9238 => x"1a",
          9239 => x"c0",
          9240 => x"74",
          9241 => x"39",
          9242 => x"55",
          9243 => x"8f",
          9244 => x"fd",
          9245 => x"d5",
          9246 => x"f5",
          9247 => x"78",
          9248 => x"79",
          9249 => x"80",
          9250 => x"f1",
          9251 => x"39",
          9252 => x"81",
          9253 => x"06",
          9254 => x"55",
          9255 => x"27",
          9256 => x"81",
          9257 => x"56",
          9258 => x"38",
          9259 => x"80",
          9260 => x"ff",
          9261 => x"8b",
          9262 => x"a0",
          9263 => x"ff",
          9264 => x"84",
          9265 => x"1b",
          9266 => x"aa",
          9267 => x"1c",
          9268 => x"ff",
          9269 => x"8e",
          9270 => x"8e",
          9271 => x"0b",
          9272 => x"7d",
          9273 => x"30",
          9274 => x"84",
          9275 => x"51",
          9276 => x"51",
          9277 => x"3f",
          9278 => x"83",
          9279 => x"90",
          9280 => x"ff",
          9281 => x"93",
          9282 => x"8d",
          9283 => x"39",
          9284 => x"1b",
          9285 => x"fc",
          9286 => x"95",
          9287 => x"52",
          9288 => x"ff",
          9289 => x"81",
          9290 => x"1b",
          9291 => x"c6",
          9292 => x"9c",
          9293 => x"8d",
          9294 => x"83",
          9295 => x"06",
          9296 => x"82",
          9297 => x"52",
          9298 => x"51",
          9299 => x"3f",
          9300 => x"1b",
          9301 => x"bc",
          9302 => x"ac",
          9303 => x"8d",
          9304 => x"52",
          9305 => x"ff",
          9306 => x"86",
          9307 => x"51",
          9308 => x"3f",
          9309 => x"80",
          9310 => x"a9",
          9311 => x"1c",
          9312 => x"82",
          9313 => x"80",
          9314 => x"ae",
          9315 => x"b2",
          9316 => x"1b",
          9317 => x"fc",
          9318 => x"ff",
          9319 => x"96",
          9320 => x"8c",
          9321 => x"80",
          9322 => x"34",
          9323 => x"1c",
          9324 => x"82",
          9325 => x"ab",
          9326 => x"8d",
          9327 => x"d4",
          9328 => x"fe",
          9329 => x"59",
          9330 => x"3f",
          9331 => x"53",
          9332 => x"51",
          9333 => x"3f",
          9334 => x"d5",
          9335 => x"9c",
          9336 => x"2e",
          9337 => x"80",
          9338 => x"54",
          9339 => x"7a",
          9340 => x"ff",
          9341 => x"84",
          9342 => x"52",
          9343 => x"8c",
          9344 => x"8b",
          9345 => x"52",
          9346 => x"8c",
          9347 => x"8a",
          9348 => x"52",
          9349 => x"51",
          9350 => x"3f",
          9351 => x"83",
          9352 => x"ff",
          9353 => x"82",
          9354 => x"1b",
          9355 => x"e4",
          9356 => x"d5",
          9357 => x"ff",
          9358 => x"75",
          9359 => x"53",
          9360 => x"51",
          9361 => x"3f",
          9362 => x"1f",
          9363 => x"7f",
          9364 => x"d1",
          9365 => x"80",
          9366 => x"ff",
          9367 => x"60",
          9368 => x"7d",
          9369 => x"81",
          9370 => x"f8",
          9371 => x"ff",
          9372 => x"ff",
          9373 => x"51",
          9374 => x"3f",
          9375 => x"88",
          9376 => x"39",
          9377 => x"f8",
          9378 => x"2e",
          9379 => x"55",
          9380 => x"51",
          9381 => x"3f",
          9382 => x"57",
          9383 => x"83",
          9384 => x"76",
          9385 => x"7a",
          9386 => x"ff",
          9387 => x"82",
          9388 => x"82",
          9389 => x"80",
          9390 => x"e4",
          9391 => x"51",
          9392 => x"3f",
          9393 => x"78",
          9394 => x"74",
          9395 => x"18",
          9396 => x"2e",
          9397 => x"79",
          9398 => x"2e",
          9399 => x"55",
          9400 => x"62",
          9401 => x"74",
          9402 => x"75",
          9403 => x"7f",
          9404 => x"b1",
          9405 => x"e4",
          9406 => x"38",
          9407 => x"78",
          9408 => x"74",
          9409 => x"57",
          9410 => x"93",
          9411 => x"67",
          9412 => x"26",
          9413 => x"57",
          9414 => x"83",
          9415 => x"64",
          9416 => x"38",
          9417 => x"53",
          9418 => x"51",
          9419 => x"3f",
          9420 => x"d5",
          9421 => x"c4",
          9422 => x"29",
          9423 => x"83",
          9424 => x"75",
          9425 => x"e4",
          9426 => x"52",
          9427 => x"85",
          9428 => x"81",
          9429 => x"2a",
          9430 => x"77",
          9431 => x"84",
          9432 => x"52",
          9433 => x"89",
          9434 => x"d4",
          9435 => x"51",
          9436 => x"3f",
          9437 => x"55",
          9438 => x"81",
          9439 => x"34",
          9440 => x"16",
          9441 => x"16",
          9442 => x"16",
          9443 => x"56",
          9444 => x"52",
          9445 => x"a1",
          9446 => x"0b",
          9447 => x"82",
          9448 => x"82",
          9449 => x"56",
          9450 => x"34",
          9451 => x"08",
          9452 => x"7e",
          9453 => x"1b",
          9454 => x"d8",
          9455 => x"83",
          9456 => x"ff",
          9457 => x"81",
          9458 => x"7a",
          9459 => x"ff",
          9460 => x"81",
          9461 => x"e4",
          9462 => x"80",
          9463 => x"7f",
          9464 => x"a5",
          9465 => x"82",
          9466 => x"90",
          9467 => x"8e",
          9468 => x"81",
          9469 => x"82",
          9470 => x"56",
          9471 => x"e4",
          9472 => x"0d",
          9473 => x"0d",
          9474 => x"59",
          9475 => x"ff",
          9476 => x"57",
          9477 => x"b4",
          9478 => x"f8",
          9479 => x"81",
          9480 => x"52",
          9481 => x"94",
          9482 => x"2e",
          9483 => x"9c",
          9484 => x"33",
          9485 => x"2e",
          9486 => x"76",
          9487 => x"58",
          9488 => x"57",
          9489 => x"09",
          9490 => x"38",
          9491 => x"78",
          9492 => x"38",
          9493 => x"82",
          9494 => x"8d",
          9495 => x"f7",
          9496 => x"02",
          9497 => x"05",
          9498 => x"77",
          9499 => x"81",
          9500 => x"8d",
          9501 => x"e7",
          9502 => x"08",
          9503 => x"24",
          9504 => x"17",
          9505 => x"8c",
          9506 => x"77",
          9507 => x"16",
          9508 => x"25",
          9509 => x"3d",
          9510 => x"75",
          9511 => x"52",
          9512 => x"ca",
          9513 => x"76",
          9514 => x"70",
          9515 => x"2a",
          9516 => x"51",
          9517 => x"84",
          9518 => x"19",
          9519 => x"8b",
          9520 => x"f9",
          9521 => x"84",
          9522 => x"56",
          9523 => x"a7",
          9524 => x"fc",
          9525 => x"53",
          9526 => x"75",
          9527 => x"dc",
          9528 => x"e4",
          9529 => x"84",
          9530 => x"2e",
          9531 => x"87",
          9532 => x"08",
          9533 => x"ff",
          9534 => x"d5",
          9535 => x"3d",
          9536 => x"3d",
          9537 => x"80",
          9538 => x"52",
          9539 => x"86",
          9540 => x"74",
          9541 => x"0d",
          9542 => x"0d",
          9543 => x"05",
          9544 => x"86",
          9545 => x"54",
          9546 => x"73",
          9547 => x"fe",
          9548 => x"51",
          9549 => x"98",
          9550 => x"fd",
          9551 => x"02",
          9552 => x"05",
          9553 => x"80",
          9554 => x"ff",
          9555 => x"72",
          9556 => x"06",
          9557 => x"39",
          9558 => x"73",
          9559 => x"83",
          9560 => x"81",
          9561 => x"70",
          9562 => x"38",
          9563 => x"22",
          9564 => x"2e",
          9565 => x"12",
          9566 => x"ff",
          9567 => x"71",
          9568 => x"8d",
          9569 => x"82",
          9570 => x"70",
          9571 => x"e1",
          9572 => x"12",
          9573 => x"06",
          9574 => x"82",
          9575 => x"85",
          9576 => x"fe",
          9577 => x"92",
          9578 => x"84",
          9579 => x"22",
          9580 => x"53",
          9581 => x"26",
          9582 => x"53",
          9583 => x"83",
          9584 => x"81",
          9585 => x"70",
          9586 => x"8b",
          9587 => x"82",
          9588 => x"70",
          9589 => x"72",
          9590 => x"0c",
          9591 => x"04",
          9592 => x"77",
          9593 => x"ff",
          9594 => x"a7",
          9595 => x"ff",
          9596 => x"cb",
          9597 => x"9f",
          9598 => x"85",
          9599 => x"9c",
          9600 => x"82",
          9601 => x"70",
          9602 => x"25",
          9603 => x"07",
          9604 => x"70",
          9605 => x"75",
          9606 => x"57",
          9607 => x"2a",
          9608 => x"06",
          9609 => x"52",
          9610 => x"71",
          9611 => x"38",
          9612 => x"80",
          9613 => x"84",
          9614 => x"e8",
          9615 => x"08",
          9616 => x"31",
          9617 => x"70",
          9618 => x"51",
          9619 => x"71",
          9620 => x"06",
          9621 => x"51",
          9622 => x"f0",
          9623 => x"39",
          9624 => x"9a",
          9625 => x"51",
          9626 => x"12",
          9627 => x"88",
          9628 => x"39",
          9629 => x"51",
          9630 => x"a0",
          9631 => x"83",
          9632 => x"52",
          9633 => x"fe",
          9634 => x"10",
          9635 => x"f1",
          9636 => x"70",
          9637 => x"0c",
          9638 => x"04",
          9639 => x"ff",
          9640 => x"ff",
          9641 => x"ff",
          9642 => x"00",
          9643 => x"51",
          9644 => x"d5",
          9645 => x"dc",
          9646 => x"e3",
          9647 => x"ea",
          9648 => x"f1",
          9649 => x"f8",
          9650 => x"ff",
          9651 => x"06",
          9652 => x"0d",
          9653 => x"14",
          9654 => x"1b",
          9655 => x"21",
          9656 => x"27",
          9657 => x"2d",
          9658 => x"33",
          9659 => x"39",
          9660 => x"3f",
          9661 => x"45",
          9662 => x"4b",
          9663 => x"33",
          9664 => x"39",
          9665 => x"3f",
          9666 => x"45",
          9667 => x"4b",
          9668 => x"29",
          9669 => x"29",
          9670 => x"3a",
          9671 => x"92",
          9672 => x"11",
          9673 => x"fe",
          9674 => x"02",
          9675 => x"63",
          9676 => x"45",
          9677 => x"db",
          9678 => x"61",
          9679 => x"e4",
          9680 => x"fe",
          9681 => x"3a",
          9682 => x"63",
          9683 => x"02",
          9684 => x"fe",
          9685 => x"fe",
          9686 => x"61",
          9687 => x"db",
          9688 => x"63",
          9689 => x"92",
          9690 => x"41",
          9691 => x"4f",
          9692 => x"5b",
          9693 => x"60",
          9694 => x"65",
          9695 => x"6a",
          9696 => x"6f",
          9697 => x"74",
          9698 => x"7a",
          9699 => x"31",
          9700 => x"1a",
          9701 => x"1a",
          9702 => x"60",
          9703 => x"1a",
          9704 => x"1a",
          9705 => x"1a",
          9706 => x"1a",
          9707 => x"1a",
          9708 => x"1a",
          9709 => x"1a",
          9710 => x"1d",
          9711 => x"1a",
          9712 => x"48",
          9713 => x"78",
          9714 => x"1a",
          9715 => x"1a",
          9716 => x"1a",
          9717 => x"1a",
          9718 => x"1a",
          9719 => x"1a",
          9720 => x"1a",
          9721 => x"1a",
          9722 => x"1a",
          9723 => x"1a",
          9724 => x"1a",
          9725 => x"1a",
          9726 => x"1a",
          9727 => x"1a",
          9728 => x"1a",
          9729 => x"1a",
          9730 => x"1a",
          9731 => x"1a",
          9732 => x"1a",
          9733 => x"1a",
          9734 => x"1a",
          9735 => x"1a",
          9736 => x"1a",
          9737 => x"1a",
          9738 => x"1a",
          9739 => x"1a",
          9740 => x"1a",
          9741 => x"1a",
          9742 => x"1a",
          9743 => x"1a",
          9744 => x"1a",
          9745 => x"1a",
          9746 => x"1a",
          9747 => x"1a",
          9748 => x"1a",
          9749 => x"1a",
          9750 => x"a8",
          9751 => x"1a",
          9752 => x"1a",
          9753 => x"1a",
          9754 => x"1a",
          9755 => x"16",
          9756 => x"1a",
          9757 => x"1a",
          9758 => x"1a",
          9759 => x"1a",
          9760 => x"1a",
          9761 => x"1a",
          9762 => x"1a",
          9763 => x"1a",
          9764 => x"1a",
          9765 => x"1a",
          9766 => x"d8",
          9767 => x"3f",
          9768 => x"af",
          9769 => x"af",
          9770 => x"af",
          9771 => x"1a",
          9772 => x"3f",
          9773 => x"1a",
          9774 => x"1a",
          9775 => x"98",
          9776 => x"1a",
          9777 => x"1a",
          9778 => x"ec",
          9779 => x"f7",
          9780 => x"1a",
          9781 => x"1a",
          9782 => x"11",
          9783 => x"1a",
          9784 => x"1f",
          9785 => x"1a",
          9786 => x"1a",
          9787 => x"16",
          9788 => x"69",
          9789 => x"00",
          9790 => x"63",
          9791 => x"00",
          9792 => x"69",
          9793 => x"00",
          9794 => x"61",
          9795 => x"00",
          9796 => x"65",
          9797 => x"00",
          9798 => x"65",
          9799 => x"00",
          9800 => x"70",
          9801 => x"00",
          9802 => x"66",
          9803 => x"00",
          9804 => x"6d",
          9805 => x"00",
          9806 => x"00",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"00",
          9811 => x"00",
          9812 => x"00",
          9813 => x"6c",
          9814 => x"00",
          9815 => x"00",
          9816 => x"74",
          9817 => x"00",
          9818 => x"65",
          9819 => x"00",
          9820 => x"6f",
          9821 => x"00",
          9822 => x"74",
          9823 => x"00",
          9824 => x"73",
          9825 => x"00",
          9826 => x"73",
          9827 => x"00",
          9828 => x"6f",
          9829 => x"00",
          9830 => x"00",
          9831 => x"6b",
          9832 => x"72",
          9833 => x"00",
          9834 => x"65",
          9835 => x"6c",
          9836 => x"72",
          9837 => x"00",
          9838 => x"6b",
          9839 => x"74",
          9840 => x"61",
          9841 => x"00",
          9842 => x"66",
          9843 => x"20",
          9844 => x"6e",
          9845 => x"00",
          9846 => x"70",
          9847 => x"20",
          9848 => x"6e",
          9849 => x"00",
          9850 => x"61",
          9851 => x"20",
          9852 => x"65",
          9853 => x"65",
          9854 => x"00",
          9855 => x"65",
          9856 => x"64",
          9857 => x"65",
          9858 => x"00",
          9859 => x"65",
          9860 => x"72",
          9861 => x"79",
          9862 => x"69",
          9863 => x"2e",
          9864 => x"00",
          9865 => x"65",
          9866 => x"6e",
          9867 => x"20",
          9868 => x"61",
          9869 => x"2e",
          9870 => x"00",
          9871 => x"69",
          9872 => x"72",
          9873 => x"20",
          9874 => x"74",
          9875 => x"65",
          9876 => x"00",
          9877 => x"76",
          9878 => x"75",
          9879 => x"72",
          9880 => x"20",
          9881 => x"61",
          9882 => x"2e",
          9883 => x"00",
          9884 => x"6b",
          9885 => x"74",
          9886 => x"61",
          9887 => x"64",
          9888 => x"00",
          9889 => x"63",
          9890 => x"61",
          9891 => x"6c",
          9892 => x"69",
          9893 => x"79",
          9894 => x"6d",
          9895 => x"75",
          9896 => x"6f",
          9897 => x"69",
          9898 => x"00",
          9899 => x"6d",
          9900 => x"61",
          9901 => x"74",
          9902 => x"00",
          9903 => x"65",
          9904 => x"2c",
          9905 => x"65",
          9906 => x"69",
          9907 => x"63",
          9908 => x"65",
          9909 => x"64",
          9910 => x"00",
          9911 => x"65",
          9912 => x"20",
          9913 => x"6b",
          9914 => x"00",
          9915 => x"75",
          9916 => x"63",
          9917 => x"74",
          9918 => x"6d",
          9919 => x"2e",
          9920 => x"00",
          9921 => x"20",
          9922 => x"79",
          9923 => x"65",
          9924 => x"69",
          9925 => x"2e",
          9926 => x"00",
          9927 => x"61",
          9928 => x"65",
          9929 => x"69",
          9930 => x"72",
          9931 => x"74",
          9932 => x"00",
          9933 => x"63",
          9934 => x"2e",
          9935 => x"00",
          9936 => x"6e",
          9937 => x"20",
          9938 => x"6f",
          9939 => x"00",
          9940 => x"75",
          9941 => x"74",
          9942 => x"25",
          9943 => x"74",
          9944 => x"75",
          9945 => x"74",
          9946 => x"73",
          9947 => x"0a",
          9948 => x"00",
          9949 => x"64",
          9950 => x"00",
          9951 => x"6c",
          9952 => x"00",
          9953 => x"00",
          9954 => x"58",
          9955 => x"00",
          9956 => x"20",
          9957 => x"20",
          9958 => x"00",
          9959 => x"58",
          9960 => x"00",
          9961 => x"00",
          9962 => x"00",
          9963 => x"00",
          9964 => x"00",
          9965 => x"20",
          9966 => x"28",
          9967 => x"00",
          9968 => x"31",
          9969 => x"30",
          9970 => x"00",
          9971 => x"31",
          9972 => x"00",
          9973 => x"55",
          9974 => x"65",
          9975 => x"30",
          9976 => x"20",
          9977 => x"25",
          9978 => x"2a",
          9979 => x"00",
          9980 => x"20",
          9981 => x"65",
          9982 => x"70",
          9983 => x"61",
          9984 => x"65",
          9985 => x"00",
          9986 => x"65",
          9987 => x"6e",
          9988 => x"72",
          9989 => x"00",
          9990 => x"20",
          9991 => x"65",
          9992 => x"70",
          9993 => x"00",
          9994 => x"54",
          9995 => x"44",
          9996 => x"74",
          9997 => x"75",
          9998 => x"00",
          9999 => x"54",
         10000 => x"52",
         10001 => x"74",
         10002 => x"75",
         10003 => x"00",
         10004 => x"54",
         10005 => x"58",
         10006 => x"74",
         10007 => x"75",
         10008 => x"00",
         10009 => x"54",
         10010 => x"58",
         10011 => x"74",
         10012 => x"75",
         10013 => x"00",
         10014 => x"54",
         10015 => x"58",
         10016 => x"74",
         10017 => x"75",
         10018 => x"00",
         10019 => x"54",
         10020 => x"58",
         10021 => x"74",
         10022 => x"75",
         10023 => x"00",
         10024 => x"74",
         10025 => x"20",
         10026 => x"74",
         10027 => x"72",
         10028 => x"00",
         10029 => x"62",
         10030 => x"67",
         10031 => x"6d",
         10032 => x"2e",
         10033 => x"00",
         10034 => x"6f",
         10035 => x"63",
         10036 => x"74",
         10037 => x"00",
         10038 => x"5f",
         10039 => x"2e",
         10040 => x"00",
         10041 => x"00",
         10042 => x"6c",
         10043 => x"74",
         10044 => x"6e",
         10045 => x"61",
         10046 => x"65",
         10047 => x"20",
         10048 => x"64",
         10049 => x"20",
         10050 => x"61",
         10051 => x"69",
         10052 => x"20",
         10053 => x"75",
         10054 => x"79",
         10055 => x"00",
         10056 => x"00",
         10057 => x"61",
         10058 => x"67",
         10059 => x"2e",
         10060 => x"00",
         10061 => x"79",
         10062 => x"2e",
         10063 => x"00",
         10064 => x"70",
         10065 => x"6e",
         10066 => x"2e",
         10067 => x"00",
         10068 => x"6c",
         10069 => x"30",
         10070 => x"2d",
         10071 => x"38",
         10072 => x"25",
         10073 => x"29",
         10074 => x"00",
         10075 => x"70",
         10076 => x"6d",
         10077 => x"00",
         10078 => x"6d",
         10079 => x"74",
         10080 => x"00",
         10081 => x"6c",
         10082 => x"30",
         10083 => x"00",
         10084 => x"00",
         10085 => x"6c",
         10086 => x"30",
         10087 => x"00",
         10088 => x"6c",
         10089 => x"30",
         10090 => x"2d",
         10091 => x"00",
         10092 => x"63",
         10093 => x"6e",
         10094 => x"6f",
         10095 => x"40",
         10096 => x"38",
         10097 => x"2e",
         10098 => x"00",
         10099 => x"6c",
         10100 => x"20",
         10101 => x"65",
         10102 => x"25",
         10103 => x"78",
         10104 => x"2e",
         10105 => x"00",
         10106 => x"6c",
         10107 => x"74",
         10108 => x"65",
         10109 => x"6f",
         10110 => x"28",
         10111 => x"2e",
         10112 => x"00",
         10113 => x"74",
         10114 => x"69",
         10115 => x"61",
         10116 => x"69",
         10117 => x"69",
         10118 => x"2e",
         10119 => x"00",
         10120 => x"64",
         10121 => x"62",
         10122 => x"69",
         10123 => x"2e",
         10124 => x"00",
         10125 => x"00",
         10126 => x"00",
         10127 => x"5c",
         10128 => x"25",
         10129 => x"73",
         10130 => x"00",
         10131 => x"5c",
         10132 => x"25",
         10133 => x"00",
         10134 => x"5c",
         10135 => x"00",
         10136 => x"20",
         10137 => x"6d",
         10138 => x"2e",
         10139 => x"00",
         10140 => x"6f",
         10141 => x"65",
         10142 => x"75",
         10143 => x"64",
         10144 => x"61",
         10145 => x"74",
         10146 => x"6f",
         10147 => x"73",
         10148 => x"6d",
         10149 => x"64",
         10150 => x"00",
         10151 => x"6e",
         10152 => x"2e",
         10153 => x"00",
         10154 => x"62",
         10155 => x"67",
         10156 => x"74",
         10157 => x"75",
         10158 => x"2e",
         10159 => x"00",
         10160 => x"25",
         10161 => x"64",
         10162 => x"3a",
         10163 => x"25",
         10164 => x"64",
         10165 => x"00",
         10166 => x"20",
         10167 => x"66",
         10168 => x"72",
         10169 => x"6f",
         10170 => x"00",
         10171 => x"72",
         10172 => x"53",
         10173 => x"63",
         10174 => x"69",
         10175 => x"00",
         10176 => x"65",
         10177 => x"65",
         10178 => x"6d",
         10179 => x"6d",
         10180 => x"65",
         10181 => x"00",
         10182 => x"20",
         10183 => x"53",
         10184 => x"4d",
         10185 => x"25",
         10186 => x"3a",
         10187 => x"58",
         10188 => x"00",
         10189 => x"20",
         10190 => x"41",
         10191 => x"20",
         10192 => x"25",
         10193 => x"3a",
         10194 => x"58",
         10195 => x"00",
         10196 => x"20",
         10197 => x"4e",
         10198 => x"41",
         10199 => x"25",
         10200 => x"3a",
         10201 => x"58",
         10202 => x"00",
         10203 => x"20",
         10204 => x"4d",
         10205 => x"20",
         10206 => x"25",
         10207 => x"3a",
         10208 => x"58",
         10209 => x"00",
         10210 => x"20",
         10211 => x"20",
         10212 => x"20",
         10213 => x"25",
         10214 => x"3a",
         10215 => x"58",
         10216 => x"00",
         10217 => x"20",
         10218 => x"43",
         10219 => x"20",
         10220 => x"44",
         10221 => x"63",
         10222 => x"3d",
         10223 => x"64",
         10224 => x"00",
         10225 => x"20",
         10226 => x"45",
         10227 => x"20",
         10228 => x"54",
         10229 => x"72",
         10230 => x"3d",
         10231 => x"64",
         10232 => x"00",
         10233 => x"20",
         10234 => x"52",
         10235 => x"52",
         10236 => x"43",
         10237 => x"6e",
         10238 => x"3d",
         10239 => x"64",
         10240 => x"00",
         10241 => x"20",
         10242 => x"48",
         10243 => x"45",
         10244 => x"53",
         10245 => x"00",
         10246 => x"20",
         10247 => x"49",
         10248 => x"00",
         10249 => x"20",
         10250 => x"54",
         10251 => x"00",
         10252 => x"20",
         10253 => x"00",
         10254 => x"20",
         10255 => x"00",
         10256 => x"72",
         10257 => x"65",
         10258 => x"00",
         10259 => x"20",
         10260 => x"20",
         10261 => x"65",
         10262 => x"65",
         10263 => x"72",
         10264 => x"64",
         10265 => x"73",
         10266 => x"25",
         10267 => x"0a",
         10268 => x"00",
         10269 => x"20",
         10270 => x"20",
         10271 => x"6f",
         10272 => x"53",
         10273 => x"74",
         10274 => x"64",
         10275 => x"73",
         10276 => x"25",
         10277 => x"0a",
         10278 => x"00",
         10279 => x"20",
         10280 => x"63",
         10281 => x"74",
         10282 => x"20",
         10283 => x"72",
         10284 => x"20",
         10285 => x"20",
         10286 => x"25",
         10287 => x"0a",
         10288 => x"00",
         10289 => x"63",
         10290 => x"00",
         10291 => x"20",
         10292 => x"20",
         10293 => x"20",
         10294 => x"20",
         10295 => x"20",
         10296 => x"20",
         10297 => x"20",
         10298 => x"25",
         10299 => x"0a",
         10300 => x"00",
         10301 => x"20",
         10302 => x"74",
         10303 => x"43",
         10304 => x"6b",
         10305 => x"65",
         10306 => x"20",
         10307 => x"20",
         10308 => x"25",
         10309 => x"30",
         10310 => x"48",
         10311 => x"00",
         10312 => x"20",
         10313 => x"41",
         10314 => x"6c",
         10315 => x"20",
         10316 => x"71",
         10317 => x"20",
         10318 => x"20",
         10319 => x"25",
         10320 => x"30",
         10321 => x"48",
         10322 => x"00",
         10323 => x"20",
         10324 => x"68",
         10325 => x"65",
         10326 => x"52",
         10327 => x"43",
         10328 => x"6b",
         10329 => x"65",
         10330 => x"25",
         10331 => x"30",
         10332 => x"48",
         10333 => x"00",
         10334 => x"6c",
         10335 => x"00",
         10336 => x"69",
         10337 => x"00",
         10338 => x"78",
         10339 => x"00",
         10340 => x"00",
         10341 => x"6d",
         10342 => x"00",
         10343 => x"6e",
         10344 => x"00",
         10345 => x"00",
         10346 => x"00",
         10347 => x"02",
         10348 => x"fc",
         10349 => x"00",
         10350 => x"03",
         10351 => x"f8",
         10352 => x"00",
         10353 => x"04",
         10354 => x"f4",
         10355 => x"00",
         10356 => x"05",
         10357 => x"f0",
         10358 => x"00",
         10359 => x"06",
         10360 => x"ec",
         10361 => x"00",
         10362 => x"07",
         10363 => x"e8",
         10364 => x"00",
         10365 => x"01",
         10366 => x"e4",
         10367 => x"00",
         10368 => x"08",
         10369 => x"e0",
         10370 => x"00",
         10371 => x"0b",
         10372 => x"dc",
         10373 => x"00",
         10374 => x"09",
         10375 => x"d8",
         10376 => x"00",
         10377 => x"0a",
         10378 => x"d4",
         10379 => x"00",
         10380 => x"0d",
         10381 => x"d0",
         10382 => x"00",
         10383 => x"0c",
         10384 => x"cc",
         10385 => x"00",
         10386 => x"0e",
         10387 => x"c8",
         10388 => x"00",
         10389 => x"0f",
         10390 => x"c4",
         10391 => x"00",
         10392 => x"0f",
         10393 => x"c0",
         10394 => x"00",
         10395 => x"10",
         10396 => x"bc",
         10397 => x"00",
         10398 => x"11",
         10399 => x"b8",
         10400 => x"00",
         10401 => x"12",
         10402 => x"b4",
         10403 => x"00",
         10404 => x"13",
         10405 => x"b0",
         10406 => x"00",
         10407 => x"14",
         10408 => x"ac",
         10409 => x"00",
         10410 => x"15",
         10411 => x"00",
         10412 => x"00",
         10413 => x"00",
         10414 => x"00",
         10415 => x"7e",
         10416 => x"7e",
         10417 => x"7e",
         10418 => x"00",
         10419 => x"7e",
         10420 => x"7e",
         10421 => x"7e",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"00",
         10430 => x"00",
         10431 => x"00",
         10432 => x"00",
         10433 => x"74",
         10434 => x"00",
         10435 => x"74",
         10436 => x"00",
         10437 => x"00",
         10438 => x"6c",
         10439 => x"25",
         10440 => x"00",
         10441 => x"6c",
         10442 => x"74",
         10443 => x"65",
         10444 => x"20",
         10445 => x"20",
         10446 => x"74",
         10447 => x"20",
         10448 => x"65",
         10449 => x"20",
         10450 => x"2e",
         10451 => x"00",
         10452 => x"6e",
         10453 => x"6f",
         10454 => x"2f",
         10455 => x"61",
         10456 => x"68",
         10457 => x"6f",
         10458 => x"66",
         10459 => x"2c",
         10460 => x"73",
         10461 => x"69",
         10462 => x"00",
         10463 => x"00",
         10464 => x"3c",
         10465 => x"7f",
         10466 => x"00",
         10467 => x"3d",
         10468 => x"00",
         10469 => x"00",
         10470 => x"33",
         10471 => x"00",
         10472 => x"4d",
         10473 => x"53",
         10474 => x"00",
         10475 => x"4e",
         10476 => x"20",
         10477 => x"46",
         10478 => x"32",
         10479 => x"00",
         10480 => x"4e",
         10481 => x"20",
         10482 => x"46",
         10483 => x"20",
         10484 => x"00",
         10485 => x"7c",
         10486 => x"00",
         10487 => x"00",
         10488 => x"00",
         10489 => x"07",
         10490 => x"12",
         10491 => x"1c",
         10492 => x"00",
         10493 => x"41",
         10494 => x"80",
         10495 => x"49",
         10496 => x"8f",
         10497 => x"4f",
         10498 => x"55",
         10499 => x"9b",
         10500 => x"9f",
         10501 => x"55",
         10502 => x"a7",
         10503 => x"ab",
         10504 => x"af",
         10505 => x"b3",
         10506 => x"b7",
         10507 => x"bb",
         10508 => x"bf",
         10509 => x"c3",
         10510 => x"c7",
         10511 => x"cb",
         10512 => x"cf",
         10513 => x"d3",
         10514 => x"d7",
         10515 => x"db",
         10516 => x"df",
         10517 => x"e3",
         10518 => x"e7",
         10519 => x"eb",
         10520 => x"ef",
         10521 => x"f3",
         10522 => x"f7",
         10523 => x"fb",
         10524 => x"ff",
         10525 => x"3b",
         10526 => x"2f",
         10527 => x"3a",
         10528 => x"7c",
         10529 => x"00",
         10530 => x"04",
         10531 => x"40",
         10532 => x"00",
         10533 => x"00",
         10534 => x"02",
         10535 => x"08",
         10536 => x"20",
         10537 => x"00",
         10538 => x"fc",
         10539 => x"e2",
         10540 => x"e0",
         10541 => x"e7",
         10542 => x"eb",
         10543 => x"ef",
         10544 => x"ec",
         10545 => x"c5",
         10546 => x"e6",
         10547 => x"f4",
         10548 => x"f2",
         10549 => x"f9",
         10550 => x"d6",
         10551 => x"a2",
         10552 => x"a5",
         10553 => x"92",
         10554 => x"ed",
         10555 => x"fa",
         10556 => x"d1",
         10557 => x"ba",
         10558 => x"10",
         10559 => x"bd",
         10560 => x"a1",
         10561 => x"bb",
         10562 => x"92",
         10563 => x"02",
         10564 => x"61",
         10565 => x"56",
         10566 => x"63",
         10567 => x"57",
         10568 => x"5c",
         10569 => x"10",
         10570 => x"34",
         10571 => x"1c",
         10572 => x"3c",
         10573 => x"5f",
         10574 => x"54",
         10575 => x"66",
         10576 => x"50",
         10577 => x"67",
         10578 => x"64",
         10579 => x"59",
         10580 => x"52",
         10581 => x"6b",
         10582 => x"18",
         10583 => x"88",
         10584 => x"8c",
         10585 => x"80",
         10586 => x"df",
         10587 => x"c0",
         10588 => x"c3",
         10589 => x"c4",
         10590 => x"98",
         10591 => x"b4",
         10592 => x"c6",
         10593 => x"29",
         10594 => x"b1",
         10595 => x"64",
         10596 => x"21",
         10597 => x"48",
         10598 => x"19",
         10599 => x"1a",
         10600 => x"b2",
         10601 => x"a0",
         10602 => x"1a",
         10603 => x"17",
         10604 => x"07",
         10605 => x"01",
         10606 => x"00",
         10607 => x"32",
         10608 => x"39",
         10609 => x"4a",
         10610 => x"79",
         10611 => x"80",
         10612 => x"43",
         10613 => x"82",
         10614 => x"84",
         10615 => x"86",
         10616 => x"87",
         10617 => x"8a",
         10618 => x"8b",
         10619 => x"8e",
         10620 => x"90",
         10621 => x"91",
         10622 => x"94",
         10623 => x"96",
         10624 => x"98",
         10625 => x"3d",
         10626 => x"9c",
         10627 => x"20",
         10628 => x"a0",
         10629 => x"a2",
         10630 => x"a4",
         10631 => x"a6",
         10632 => x"a7",
         10633 => x"aa",
         10634 => x"ac",
         10635 => x"ae",
         10636 => x"af",
         10637 => x"b2",
         10638 => x"b3",
         10639 => x"b5",
         10640 => x"b8",
         10641 => x"ba",
         10642 => x"bc",
         10643 => x"be",
         10644 => x"c0",
         10645 => x"c2",
         10646 => x"c4",
         10647 => x"c4",
         10648 => x"c8",
         10649 => x"ca",
         10650 => x"ca",
         10651 => x"10",
         10652 => x"01",
         10653 => x"de",
         10654 => x"f3",
         10655 => x"f1",
         10656 => x"f4",
         10657 => x"28",
         10658 => x"12",
         10659 => x"09",
         10660 => x"3b",
         10661 => x"3d",
         10662 => x"3f",
         10663 => x"41",
         10664 => x"46",
         10665 => x"53",
         10666 => x"81",
         10667 => x"55",
         10668 => x"8a",
         10669 => x"8f",
         10670 => x"90",
         10671 => x"5d",
         10672 => x"5f",
         10673 => x"61",
         10674 => x"94",
         10675 => x"65",
         10676 => x"67",
         10677 => x"96",
         10678 => x"62",
         10679 => x"6d",
         10680 => x"9c",
         10681 => x"71",
         10682 => x"73",
         10683 => x"9f",
         10684 => x"77",
         10685 => x"79",
         10686 => x"7b",
         10687 => x"64",
         10688 => x"7f",
         10689 => x"81",
         10690 => x"a9",
         10691 => x"85",
         10692 => x"87",
         10693 => x"44",
         10694 => x"b2",
         10695 => x"8d",
         10696 => x"8f",
         10697 => x"91",
         10698 => x"7b",
         10699 => x"fd",
         10700 => x"ff",
         10701 => x"04",
         10702 => x"88",
         10703 => x"8a",
         10704 => x"11",
         10705 => x"02",
         10706 => x"a3",
         10707 => x"08",
         10708 => x"03",
         10709 => x"8e",
         10710 => x"d8",
         10711 => x"f2",
         10712 => x"f9",
         10713 => x"f4",
         10714 => x"f6",
         10715 => x"f7",
         10716 => x"fa",
         10717 => x"30",
         10718 => x"50",
         10719 => x"60",
         10720 => x"8a",
         10721 => x"c1",
         10722 => x"cf",
         10723 => x"c0",
         10724 => x"44",
         10725 => x"26",
         10726 => x"00",
         10727 => x"01",
         10728 => x"00",
         10729 => x"a0",
         10730 => x"00",
         10731 => x"10",
         10732 => x"20",
         10733 => x"30",
         10734 => x"40",
         10735 => x"51",
         10736 => x"59",
         10737 => x"5b",
         10738 => x"5d",
         10739 => x"5f",
         10740 => x"08",
         10741 => x"0e",
         10742 => x"bb",
         10743 => x"c9",
         10744 => x"cb",
         10745 => x"db",
         10746 => x"f9",
         10747 => x"eb",
         10748 => x"fb",
         10749 => x"08",
         10750 => x"08",
         10751 => x"08",
         10752 => x"04",
         10753 => x"b9",
         10754 => x"bc",
         10755 => x"01",
         10756 => x"d0",
         10757 => x"e0",
         10758 => x"e5",
         10759 => x"ec",
         10760 => x"01",
         10761 => x"4e",
         10762 => x"32",
         10763 => x"10",
         10764 => x"01",
         10765 => x"d0",
         10766 => x"30",
         10767 => x"60",
         10768 => x"67",
         10769 => x"75",
         10770 => x"80",
         10771 => x"00",
         10772 => x"41",
         10773 => x"00",
         10774 => x"00",
         10775 => x"f0",
         10776 => x"00",
         10777 => x"00",
         10778 => x"00",
         10779 => x"f8",
         10780 => x"00",
         10781 => x"00",
         10782 => x"00",
         10783 => x"00",
         10784 => x"00",
         10785 => x"00",
         10786 => x"00",
         10787 => x"08",
         10788 => x"00",
         10789 => x"00",
         10790 => x"00",
         10791 => x"10",
         10792 => x"00",
         10793 => x"00",
         10794 => x"00",
         10795 => x"18",
         10796 => x"00",
         10797 => x"00",
         10798 => x"00",
         10799 => x"20",
         10800 => x"00",
         10801 => x"00",
         10802 => x"00",
         10803 => x"28",
         10804 => x"00",
         10805 => x"00",
         10806 => x"00",
         10807 => x"30",
         10808 => x"00",
         10809 => x"00",
         10810 => x"00",
         10811 => x"38",
         10812 => x"00",
         10813 => x"00",
         10814 => x"00",
         10815 => x"3c",
         10816 => x"00",
         10817 => x"00",
         10818 => x"00",
         10819 => x"40",
         10820 => x"00",
         10821 => x"00",
         10822 => x"00",
         10823 => x"44",
         10824 => x"00",
         10825 => x"00",
         10826 => x"00",
         10827 => x"48",
         10828 => x"00",
         10829 => x"00",
         10830 => x"00",
         10831 => x"4c",
         10832 => x"00",
         10833 => x"00",
         10834 => x"00",
         10835 => x"50",
         10836 => x"00",
         10837 => x"00",
         10838 => x"00",
         10839 => x"54",
         10840 => x"00",
         10841 => x"00",
         10842 => x"00",
         10843 => x"5c",
         10844 => x"00",
         10845 => x"00",
         10846 => x"00",
         10847 => x"60",
         10848 => x"00",
         10849 => x"00",
         10850 => x"00",
         10851 => x"68",
         10852 => x"00",
         10853 => x"00",
         10854 => x"00",
         10855 => x"70",
         10856 => x"00",
         10857 => x"00",
         10858 => x"00",
         10859 => x"78",
         10860 => x"00",
         10861 => x"00",
         10862 => x"00",
         10863 => x"80",
         10864 => x"00",
         10865 => x"00",
         10866 => x"00",
         10867 => x"88",
         10868 => x"00",
         10869 => x"00",
         10870 => x"00",
         10871 => x"90",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"98",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"ff",
         10882 => x"00",
         10883 => x"ff",
         10884 => x"00",
         10885 => x"ff",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"ff",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"01",
         10899 => x"01",
         10900 => x"01",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"04",
         10927 => x"00",
         10928 => x"0c",
         10929 => x"00",
         10930 => x"14",
         10931 => x"00",
         10932 => x"00",
         10933 => x"00",
         10934 => x"02",
         10935 => x"04",
         10936 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"b9",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a4",
           270 => x"0b",
           271 => x"0b",
           272 => x"c2",
           273 => x"0b",
           274 => x"0b",
           275 => x"e0",
           276 => x"0b",
           277 => x"0b",
           278 => x"80",
           279 => x"0b",
           280 => x"0b",
           281 => x"9e",
           282 => x"0b",
           283 => x"0b",
           284 => x"bd",
           285 => x"0b",
           286 => x"0b",
           287 => x"dd",
           288 => x"0b",
           289 => x"0b",
           290 => x"fd",
           291 => x"0b",
           292 => x"0b",
           293 => x"9d",
           294 => x"0b",
           295 => x"0b",
           296 => x"bd",
           297 => x"0b",
           298 => x"0b",
           299 => x"dd",
           300 => x"0b",
           301 => x"0b",
           302 => x"fd",
           303 => x"0b",
           304 => x"0b",
           305 => x"9d",
           306 => x"0b",
           307 => x"0b",
           308 => x"bd",
           309 => x"0b",
           310 => x"0b",
           311 => x"dd",
           312 => x"0b",
           313 => x"0b",
           314 => x"fd",
           315 => x"0b",
           316 => x"0b",
           317 => x"9d",
           318 => x"0b",
           319 => x"0b",
           320 => x"bd",
           321 => x"0b",
           322 => x"0b",
           323 => x"dd",
           324 => x"0b",
           325 => x"0b",
           326 => x"fd",
           327 => x"0b",
           328 => x"0b",
           329 => x"9d",
           330 => x"0b",
           331 => x"0b",
           332 => x"bd",
           333 => x"0b",
           334 => x"0b",
           335 => x"dd",
           336 => x"0b",
           337 => x"0b",
           338 => x"fd",
           339 => x"0b",
           340 => x"0b",
           341 => x"9d",
           342 => x"0b",
           343 => x"0b",
           344 => x"bd",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"d5",
           386 => x"f6",
           387 => x"d5",
           388 => x"80",
           389 => x"d5",
           390 => x"b2",
           391 => x"f0",
           392 => x"90",
           393 => x"f0",
           394 => x"2d",
           395 => x"08",
           396 => x"04",
           397 => x"0c",
           398 => x"82",
           399 => x"84",
           400 => x"82",
           401 => x"94",
           402 => x"d5",
           403 => x"80",
           404 => x"d5",
           405 => x"c2",
           406 => x"f0",
           407 => x"90",
           408 => x"f0",
           409 => x"f7",
           410 => x"f0",
           411 => x"90",
           412 => x"f0",
           413 => x"a6",
           414 => x"f0",
           415 => x"90",
           416 => x"f0",
           417 => x"2d",
           418 => x"08",
           419 => x"04",
           420 => x"0c",
           421 => x"82",
           422 => x"84",
           423 => x"82",
           424 => x"97",
           425 => x"d5",
           426 => x"80",
           427 => x"d5",
           428 => x"f9",
           429 => x"d5",
           430 => x"80",
           431 => x"d5",
           432 => x"fa",
           433 => x"d5",
           434 => x"80",
           435 => x"d5",
           436 => x"f2",
           437 => x"d5",
           438 => x"80",
           439 => x"d5",
           440 => x"f3",
           441 => x"d5",
           442 => x"80",
           443 => x"d5",
           444 => x"f5",
           445 => x"d5",
           446 => x"80",
           447 => x"d5",
           448 => x"eb",
           449 => x"d5",
           450 => x"80",
           451 => x"d5",
           452 => x"f8",
           453 => x"d5",
           454 => x"80",
           455 => x"d5",
           456 => x"f0",
           457 => x"d5",
           458 => x"80",
           459 => x"d5",
           460 => x"f3",
           461 => x"d5",
           462 => x"80",
           463 => x"d5",
           464 => x"fe",
           465 => x"d5",
           466 => x"80",
           467 => x"d5",
           468 => x"86",
           469 => x"d5",
           470 => x"80",
           471 => x"d5",
           472 => x"f7",
           473 => x"d5",
           474 => x"80",
           475 => x"d5",
           476 => x"81",
           477 => x"d5",
           478 => x"80",
           479 => x"d5",
           480 => x"82",
           481 => x"d5",
           482 => x"80",
           483 => x"d5",
           484 => x"82",
           485 => x"d5",
           486 => x"80",
           487 => x"d5",
           488 => x"8a",
           489 => x"d5",
           490 => x"80",
           491 => x"d5",
           492 => x"88",
           493 => x"d5",
           494 => x"80",
           495 => x"d5",
           496 => x"8d",
           497 => x"d5",
           498 => x"80",
           499 => x"d5",
           500 => x"83",
           501 => x"d5",
           502 => x"80",
           503 => x"d5",
           504 => x"90",
           505 => x"d5",
           506 => x"80",
           507 => x"d5",
           508 => x"91",
           509 => x"d5",
           510 => x"80",
           511 => x"d5",
           512 => x"f9",
           513 => x"d5",
           514 => x"80",
           515 => x"d5",
           516 => x"f9",
           517 => x"d5",
           518 => x"80",
           519 => x"d5",
           520 => x"fa",
           521 => x"d5",
           522 => x"80",
           523 => x"d5",
           524 => x"84",
           525 => x"d5",
           526 => x"80",
           527 => x"d5",
           528 => x"92",
           529 => x"d5",
           530 => x"80",
           531 => x"d5",
           532 => x"94",
           533 => x"d5",
           534 => x"80",
           535 => x"d5",
           536 => x"97",
           537 => x"d5",
           538 => x"80",
           539 => x"d5",
           540 => x"ea",
           541 => x"d5",
           542 => x"80",
           543 => x"d5",
           544 => x"9a",
           545 => x"d5",
           546 => x"80",
           547 => x"d5",
           548 => x"aa",
           549 => x"d5",
           550 => x"80",
           551 => x"d5",
           552 => x"a8",
           553 => x"d5",
           554 => x"80",
           555 => x"d5",
           556 => x"aa",
           557 => x"d5",
           558 => x"80",
           559 => x"d5",
           560 => x"ac",
           561 => x"d5",
           562 => x"80",
           563 => x"d5",
           564 => x"ae",
           565 => x"d5",
           566 => x"80",
           567 => x"d5",
           568 => x"f2",
           569 => x"d5",
           570 => x"80",
           571 => x"d5",
           572 => x"f3",
           573 => x"d5",
           574 => x"80",
           575 => x"d5",
           576 => x"f7",
           577 => x"d5",
           578 => x"80",
           579 => x"d5",
           580 => x"d7",
           581 => x"d5",
           582 => x"80",
           583 => x"d5",
           584 => x"a4",
           585 => x"d5",
           586 => x"80",
           587 => x"d5",
           588 => x"a4",
           589 => x"d5",
           590 => x"80",
           591 => x"d5",
           592 => x"a8",
           593 => x"d5",
           594 => x"80",
           595 => x"d5",
           596 => x"a1",
           597 => x"d5",
           598 => x"80",
           599 => x"04",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"04",
           609 => x"81",
           610 => x"83",
           611 => x"05",
           612 => x"10",
           613 => x"72",
           614 => x"51",
           615 => x"72",
           616 => x"06",
           617 => x"72",
           618 => x"10",
           619 => x"10",
           620 => x"ed",
           621 => x"53",
           622 => x"d5",
           623 => x"f1",
           624 => x"38",
           625 => x"84",
           626 => x"0b",
           627 => x"bc",
           628 => x"51",
           629 => x"04",
           630 => x"f0",
           631 => x"d5",
           632 => x"3d",
           633 => x"f0",
           634 => x"70",
           635 => x"08",
           636 => x"82",
           637 => x"fc",
           638 => x"82",
           639 => x"88",
           640 => x"82",
           641 => x"52",
           642 => x"3f",
           643 => x"08",
           644 => x"f0",
           645 => x"0c",
           646 => x"08",
           647 => x"70",
           648 => x"0c",
           649 => x"3d",
           650 => x"f0",
           651 => x"d5",
           652 => x"82",
           653 => x"fb",
           654 => x"d5",
           655 => x"05",
           656 => x"33",
           657 => x"70",
           658 => x"51",
           659 => x"8f",
           660 => x"82",
           661 => x"8c",
           662 => x"83",
           663 => x"80",
           664 => x"f0",
           665 => x"0c",
           666 => x"82",
           667 => x"8c",
           668 => x"05",
           669 => x"08",
           670 => x"80",
           671 => x"f0",
           672 => x"0c",
           673 => x"08",
           674 => x"82",
           675 => x"fc",
           676 => x"d5",
           677 => x"05",
           678 => x"80",
           679 => x"0b",
           680 => x"08",
           681 => x"25",
           682 => x"82",
           683 => x"90",
           684 => x"a0",
           685 => x"d5",
           686 => x"82",
           687 => x"f8",
           688 => x"82",
           689 => x"f8",
           690 => x"2e",
           691 => x"8d",
           692 => x"82",
           693 => x"f4",
           694 => x"d2",
           695 => x"f0",
           696 => x"08",
           697 => x"08",
           698 => x"53",
           699 => x"34",
           700 => x"08",
           701 => x"ff",
           702 => x"f0",
           703 => x"0c",
           704 => x"08",
           705 => x"81",
           706 => x"f0",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"80",
           711 => x"d5",
           712 => x"05",
           713 => x"d5",
           714 => x"05",
           715 => x"d5",
           716 => x"05",
           717 => x"e4",
           718 => x"0d",
           719 => x"0c",
           720 => x"f0",
           721 => x"d5",
           722 => x"3d",
           723 => x"82",
           724 => x"e5",
           725 => x"d5",
           726 => x"05",
           727 => x"f0",
           728 => x"0c",
           729 => x"82",
           730 => x"e8",
           731 => x"d5",
           732 => x"05",
           733 => x"f0",
           734 => x"0c",
           735 => x"08",
           736 => x"54",
           737 => x"08",
           738 => x"53",
           739 => x"08",
           740 => x"53",
           741 => x"8d",
           742 => x"e4",
           743 => x"d5",
           744 => x"05",
           745 => x"f0",
           746 => x"08",
           747 => x"08",
           748 => x"05",
           749 => x"74",
           750 => x"f0",
           751 => x"08",
           752 => x"e4",
           753 => x"3d",
           754 => x"f0",
           755 => x"d5",
           756 => x"82",
           757 => x"fb",
           758 => x"d5",
           759 => x"05",
           760 => x"f0",
           761 => x"0c",
           762 => x"08",
           763 => x"54",
           764 => x"08",
           765 => x"53",
           766 => x"08",
           767 => x"52",
           768 => x"82",
           769 => x"70",
           770 => x"08",
           771 => x"82",
           772 => x"f8",
           773 => x"82",
           774 => x"51",
           775 => x"0d",
           776 => x"0c",
           777 => x"f0",
           778 => x"d5",
           779 => x"3d",
           780 => x"82",
           781 => x"e4",
           782 => x"d5",
           783 => x"05",
           784 => x"0b",
           785 => x"82",
           786 => x"88",
           787 => x"11",
           788 => x"2a",
           789 => x"70",
           790 => x"51",
           791 => x"72",
           792 => x"38",
           793 => x"d5",
           794 => x"05",
           795 => x"39",
           796 => x"08",
           797 => x"53",
           798 => x"72",
           799 => x"08",
           800 => x"72",
           801 => x"53",
           802 => x"95",
           803 => x"d5",
           804 => x"05",
           805 => x"82",
           806 => x"8c",
           807 => x"d5",
           808 => x"05",
           809 => x"06",
           810 => x"80",
           811 => x"38",
           812 => x"08",
           813 => x"53",
           814 => x"81",
           815 => x"d5",
           816 => x"05",
           817 => x"b9",
           818 => x"38",
           819 => x"08",
           820 => x"53",
           821 => x"09",
           822 => x"c5",
           823 => x"f0",
           824 => x"33",
           825 => x"70",
           826 => x"51",
           827 => x"38",
           828 => x"08",
           829 => x"70",
           830 => x"81",
           831 => x"06",
           832 => x"53",
           833 => x"99",
           834 => x"f0",
           835 => x"22",
           836 => x"07",
           837 => x"82",
           838 => x"e4",
           839 => x"d0",
           840 => x"f0",
           841 => x"33",
           842 => x"70",
           843 => x"70",
           844 => x"11",
           845 => x"51",
           846 => x"55",
           847 => x"d5",
           848 => x"05",
           849 => x"f0",
           850 => x"33",
           851 => x"f0",
           852 => x"33",
           853 => x"11",
           854 => x"72",
           855 => x"08",
           856 => x"82",
           857 => x"e8",
           858 => x"98",
           859 => x"2c",
           860 => x"72",
           861 => x"38",
           862 => x"82",
           863 => x"e8",
           864 => x"d5",
           865 => x"05",
           866 => x"2a",
           867 => x"51",
           868 => x"fd",
           869 => x"d5",
           870 => x"05",
           871 => x"2b",
           872 => x"70",
           873 => x"88",
           874 => x"51",
           875 => x"82",
           876 => x"ec",
           877 => x"b8",
           878 => x"f0",
           879 => x"22",
           880 => x"70",
           881 => x"51",
           882 => x"2e",
           883 => x"d5",
           884 => x"05",
           885 => x"2b",
           886 => x"51",
           887 => x"8a",
           888 => x"82",
           889 => x"e8",
           890 => x"d5",
           891 => x"05",
           892 => x"82",
           893 => x"c4",
           894 => x"82",
           895 => x"c4",
           896 => x"d8",
           897 => x"38",
           898 => x"08",
           899 => x"70",
           900 => x"af",
           901 => x"08",
           902 => x"53",
           903 => x"d5",
           904 => x"05",
           905 => x"07",
           906 => x"82",
           907 => x"e4",
           908 => x"d5",
           909 => x"05",
           910 => x"07",
           911 => x"82",
           912 => x"e4",
           913 => x"a8",
           914 => x"f0",
           915 => x"22",
           916 => x"07",
           917 => x"82",
           918 => x"e4",
           919 => x"90",
           920 => x"f0",
           921 => x"22",
           922 => x"07",
           923 => x"82",
           924 => x"e4",
           925 => x"f8",
           926 => x"f0",
           927 => x"22",
           928 => x"51",
           929 => x"d5",
           930 => x"05",
           931 => x"82",
           932 => x"e8",
           933 => x"d8",
           934 => x"f0",
           935 => x"22",
           936 => x"51",
           937 => x"d5",
           938 => x"05",
           939 => x"39",
           940 => x"d5",
           941 => x"05",
           942 => x"f0",
           943 => x"22",
           944 => x"53",
           945 => x"f0",
           946 => x"23",
           947 => x"82",
           948 => x"f8",
           949 => x"a8",
           950 => x"f0",
           951 => x"08",
           952 => x"08",
           953 => x"84",
           954 => x"f0",
           955 => x"0c",
           956 => x"53",
           957 => x"f0",
           958 => x"34",
           959 => x"08",
           960 => x"ff",
           961 => x"72",
           962 => x"08",
           963 => x"8c",
           964 => x"d5",
           965 => x"05",
           966 => x"f0",
           967 => x"08",
           968 => x"d5",
           969 => x"05",
           970 => x"82",
           971 => x"fc",
           972 => x"d5",
           973 => x"05",
           974 => x"2a",
           975 => x"51",
           976 => x"72",
           977 => x"38",
           978 => x"08",
           979 => x"70",
           980 => x"72",
           981 => x"82",
           982 => x"fc",
           983 => x"53",
           984 => x"82",
           985 => x"53",
           986 => x"f0",
           987 => x"23",
           988 => x"d5",
           989 => x"05",
           990 => x"8a",
           991 => x"e4",
           992 => x"82",
           993 => x"f4",
           994 => x"d5",
           995 => x"05",
           996 => x"d5",
           997 => x"05",
           998 => x"31",
           999 => x"82",
          1000 => x"ec",
          1001 => x"d8",
          1002 => x"f0",
          1003 => x"08",
          1004 => x"08",
          1005 => x"84",
          1006 => x"f0",
          1007 => x"0c",
          1008 => x"d5",
          1009 => x"05",
          1010 => x"f0",
          1011 => x"22",
          1012 => x"70",
          1013 => x"51",
          1014 => x"80",
          1015 => x"82",
          1016 => x"e8",
          1017 => x"98",
          1018 => x"98",
          1019 => x"d5",
          1020 => x"05",
          1021 => x"a2",
          1022 => x"d5",
          1023 => x"72",
          1024 => x"08",
          1025 => x"99",
          1026 => x"f0",
          1027 => x"08",
          1028 => x"3f",
          1029 => x"08",
          1030 => x"d5",
          1031 => x"05",
          1032 => x"f0",
          1033 => x"22",
          1034 => x"f0",
          1035 => x"22",
          1036 => x"54",
          1037 => x"d5",
          1038 => x"05",
          1039 => x"39",
          1040 => x"08",
          1041 => x"70",
          1042 => x"81",
          1043 => x"53",
          1044 => x"a4",
          1045 => x"f0",
          1046 => x"08",
          1047 => x"08",
          1048 => x"84",
          1049 => x"f0",
          1050 => x"0c",
          1051 => x"d5",
          1052 => x"05",
          1053 => x"39",
          1054 => x"08",
          1055 => x"82",
          1056 => x"90",
          1057 => x"05",
          1058 => x"08",
          1059 => x"70",
          1060 => x"f0",
          1061 => x"0c",
          1062 => x"f0",
          1063 => x"08",
          1064 => x"08",
          1065 => x"82",
          1066 => x"fc",
          1067 => x"25",
          1068 => x"d5",
          1069 => x"05",
          1070 => x"07",
          1071 => x"82",
          1072 => x"e4",
          1073 => x"d5",
          1074 => x"05",
          1075 => x"d5",
          1076 => x"05",
          1077 => x"f0",
          1078 => x"22",
          1079 => x"06",
          1080 => x"82",
          1081 => x"e4",
          1082 => x"af",
          1083 => x"82",
          1084 => x"f4",
          1085 => x"39",
          1086 => x"08",
          1087 => x"70",
          1088 => x"51",
          1089 => x"d5",
          1090 => x"05",
          1091 => x"0b",
          1092 => x"08",
          1093 => x"90",
          1094 => x"f0",
          1095 => x"23",
          1096 => x"08",
          1097 => x"70",
          1098 => x"81",
          1099 => x"53",
          1100 => x"a4",
          1101 => x"f0",
          1102 => x"08",
          1103 => x"08",
          1104 => x"84",
          1105 => x"f0",
          1106 => x"0c",
          1107 => x"d5",
          1108 => x"05",
          1109 => x"39",
          1110 => x"08",
          1111 => x"82",
          1112 => x"90",
          1113 => x"05",
          1114 => x"08",
          1115 => x"70",
          1116 => x"f0",
          1117 => x"0c",
          1118 => x"f0",
          1119 => x"08",
          1120 => x"08",
          1121 => x"82",
          1122 => x"e4",
          1123 => x"cf",
          1124 => x"72",
          1125 => x"08",
          1126 => x"82",
          1127 => x"82",
          1128 => x"f0",
          1129 => x"d5",
          1130 => x"05",
          1131 => x"f0",
          1132 => x"22",
          1133 => x"08",
          1134 => x"71",
          1135 => x"56",
          1136 => x"9e",
          1137 => x"e4",
          1138 => x"75",
          1139 => x"f0",
          1140 => x"08",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"33",
          1145 => x"73",
          1146 => x"82",
          1147 => x"f0",
          1148 => x"72",
          1149 => x"d5",
          1150 => x"05",
          1151 => x"df",
          1152 => x"53",
          1153 => x"f0",
          1154 => x"34",
          1155 => x"d5",
          1156 => x"05",
          1157 => x"33",
          1158 => x"53",
          1159 => x"f0",
          1160 => x"34",
          1161 => x"08",
          1162 => x"53",
          1163 => x"08",
          1164 => x"73",
          1165 => x"f0",
          1166 => x"08",
          1167 => x"d5",
          1168 => x"05",
          1169 => x"f0",
          1170 => x"22",
          1171 => x"d5",
          1172 => x"05",
          1173 => x"a3",
          1174 => x"d5",
          1175 => x"82",
          1176 => x"fc",
          1177 => x"82",
          1178 => x"fc",
          1179 => x"2e",
          1180 => x"b2",
          1181 => x"f0",
          1182 => x"08",
          1183 => x"54",
          1184 => x"74",
          1185 => x"51",
          1186 => x"d5",
          1187 => x"05",
          1188 => x"f0",
          1189 => x"22",
          1190 => x"51",
          1191 => x"2e",
          1192 => x"d5",
          1193 => x"05",
          1194 => x"51",
          1195 => x"d5",
          1196 => x"05",
          1197 => x"f0",
          1198 => x"22",
          1199 => x"70",
          1200 => x"51",
          1201 => x"2e",
          1202 => x"82",
          1203 => x"ec",
          1204 => x"90",
          1205 => x"f0",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"90",
          1209 => x"f0",
          1210 => x"0c",
          1211 => x"08",
          1212 => x"51",
          1213 => x"2e",
          1214 => x"95",
          1215 => x"f0",
          1216 => x"08",
          1217 => x"72",
          1218 => x"08",
          1219 => x"93",
          1220 => x"f0",
          1221 => x"08",
          1222 => x"72",
          1223 => x"08",
          1224 => x"82",
          1225 => x"c8",
          1226 => x"d5",
          1227 => x"05",
          1228 => x"f0",
          1229 => x"22",
          1230 => x"70",
          1231 => x"51",
          1232 => x"2e",
          1233 => x"82",
          1234 => x"e8",
          1235 => x"98",
          1236 => x"2c",
          1237 => x"08",
          1238 => x"57",
          1239 => x"72",
          1240 => x"38",
          1241 => x"08",
          1242 => x"70",
          1243 => x"53",
          1244 => x"f0",
          1245 => x"23",
          1246 => x"d5",
          1247 => x"05",
          1248 => x"d5",
          1249 => x"05",
          1250 => x"31",
          1251 => x"82",
          1252 => x"e8",
          1253 => x"d5",
          1254 => x"05",
          1255 => x"2a",
          1256 => x"51",
          1257 => x"80",
          1258 => x"82",
          1259 => x"e8",
          1260 => x"88",
          1261 => x"2b",
          1262 => x"70",
          1263 => x"51",
          1264 => x"72",
          1265 => x"f0",
          1266 => x"22",
          1267 => x"51",
          1268 => x"d5",
          1269 => x"05",
          1270 => x"82",
          1271 => x"fc",
          1272 => x"88",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"51",
          1276 => x"72",
          1277 => x"f0",
          1278 => x"22",
          1279 => x"51",
          1280 => x"d5",
          1281 => x"05",
          1282 => x"f0",
          1283 => x"22",
          1284 => x"06",
          1285 => x"b0",
          1286 => x"f0",
          1287 => x"22",
          1288 => x"54",
          1289 => x"f0",
          1290 => x"23",
          1291 => x"70",
          1292 => x"53",
          1293 => x"90",
          1294 => x"f0",
          1295 => x"08",
          1296 => x"8a",
          1297 => x"39",
          1298 => x"08",
          1299 => x"70",
          1300 => x"81",
          1301 => x"53",
          1302 => x"91",
          1303 => x"f0",
          1304 => x"08",
          1305 => x"8a",
          1306 => x"c7",
          1307 => x"f0",
          1308 => x"22",
          1309 => x"70",
          1310 => x"51",
          1311 => x"2e",
          1312 => x"d5",
          1313 => x"05",
          1314 => x"51",
          1315 => x"a3",
          1316 => x"f0",
          1317 => x"22",
          1318 => x"70",
          1319 => x"51",
          1320 => x"2e",
          1321 => x"d5",
          1322 => x"05",
          1323 => x"51",
          1324 => x"82",
          1325 => x"e4",
          1326 => x"86",
          1327 => x"06",
          1328 => x"72",
          1329 => x"38",
          1330 => x"08",
          1331 => x"52",
          1332 => x"df",
          1333 => x"f0",
          1334 => x"22",
          1335 => x"2e",
          1336 => x"94",
          1337 => x"f0",
          1338 => x"08",
          1339 => x"f0",
          1340 => x"33",
          1341 => x"3f",
          1342 => x"08",
          1343 => x"70",
          1344 => x"81",
          1345 => x"53",
          1346 => x"b0",
          1347 => x"f0",
          1348 => x"22",
          1349 => x"54",
          1350 => x"f0",
          1351 => x"23",
          1352 => x"70",
          1353 => x"53",
          1354 => x"90",
          1355 => x"f0",
          1356 => x"08",
          1357 => x"88",
          1358 => x"39",
          1359 => x"08",
          1360 => x"70",
          1361 => x"81",
          1362 => x"53",
          1363 => x"b0",
          1364 => x"f0",
          1365 => x"33",
          1366 => x"54",
          1367 => x"f0",
          1368 => x"34",
          1369 => x"70",
          1370 => x"53",
          1371 => x"90",
          1372 => x"f0",
          1373 => x"08",
          1374 => x"88",
          1375 => x"39",
          1376 => x"08",
          1377 => x"70",
          1378 => x"81",
          1379 => x"53",
          1380 => x"82",
          1381 => x"ec",
          1382 => x"11",
          1383 => x"82",
          1384 => x"ec",
          1385 => x"90",
          1386 => x"2c",
          1387 => x"73",
          1388 => x"82",
          1389 => x"88",
          1390 => x"a0",
          1391 => x"3f",
          1392 => x"d5",
          1393 => x"05",
          1394 => x"80",
          1395 => x"81",
          1396 => x"82",
          1397 => x"88",
          1398 => x"82",
          1399 => x"fc",
          1400 => x"87",
          1401 => x"ee",
          1402 => x"f0",
          1403 => x"33",
          1404 => x"f3",
          1405 => x"06",
          1406 => x"82",
          1407 => x"f4",
          1408 => x"11",
          1409 => x"82",
          1410 => x"f4",
          1411 => x"83",
          1412 => x"53",
          1413 => x"ff",
          1414 => x"38",
          1415 => x"08",
          1416 => x"52",
          1417 => x"08",
          1418 => x"70",
          1419 => x"d5",
          1420 => x"05",
          1421 => x"82",
          1422 => x"fc",
          1423 => x"86",
          1424 => x"b7",
          1425 => x"f0",
          1426 => x"33",
          1427 => x"d3",
          1428 => x"06",
          1429 => x"82",
          1430 => x"f4",
          1431 => x"11",
          1432 => x"82",
          1433 => x"f4",
          1434 => x"83",
          1435 => x"53",
          1436 => x"ff",
          1437 => x"38",
          1438 => x"08",
          1439 => x"52",
          1440 => x"08",
          1441 => x"70",
          1442 => x"86",
          1443 => x"d5",
          1444 => x"05",
          1445 => x"82",
          1446 => x"fc",
          1447 => x"b7",
          1448 => x"f0",
          1449 => x"08",
          1450 => x"2e",
          1451 => x"d5",
          1452 => x"05",
          1453 => x"d5",
          1454 => x"05",
          1455 => x"82",
          1456 => x"f0",
          1457 => x"d5",
          1458 => x"05",
          1459 => x"52",
          1460 => x"3f",
          1461 => x"d5",
          1462 => x"05",
          1463 => x"2a",
          1464 => x"51",
          1465 => x"80",
          1466 => x"38",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"72",
          1470 => x"08",
          1471 => x"73",
          1472 => x"90",
          1473 => x"80",
          1474 => x"38",
          1475 => x"08",
          1476 => x"52",
          1477 => x"9b",
          1478 => x"82",
          1479 => x"88",
          1480 => x"82",
          1481 => x"f8",
          1482 => x"85",
          1483 => x"0b",
          1484 => x"08",
          1485 => x"ea",
          1486 => x"d5",
          1487 => x"05",
          1488 => x"a5",
          1489 => x"06",
          1490 => x"0b",
          1491 => x"08",
          1492 => x"80",
          1493 => x"f0",
          1494 => x"23",
          1495 => x"d5",
          1496 => x"05",
          1497 => x"82",
          1498 => x"f4",
          1499 => x"80",
          1500 => x"f0",
          1501 => x"08",
          1502 => x"f0",
          1503 => x"33",
          1504 => x"3f",
          1505 => x"82",
          1506 => x"88",
          1507 => x"11",
          1508 => x"d5",
          1509 => x"05",
          1510 => x"82",
          1511 => x"e0",
          1512 => x"d5",
          1513 => x"3d",
          1514 => x"f0",
          1515 => x"d5",
          1516 => x"82",
          1517 => x"fd",
          1518 => x"f1",
          1519 => x"82",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"88",
          1523 => x"e4",
          1524 => x"d5",
          1525 => x"82",
          1526 => x"54",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"f0",
          1531 => x"0d",
          1532 => x"d5",
          1533 => x"05",
          1534 => x"c8",
          1535 => x"33",
          1536 => x"70",
          1537 => x"81",
          1538 => x"51",
          1539 => x"80",
          1540 => x"ff",
          1541 => x"f0",
          1542 => x"0c",
          1543 => x"82",
          1544 => x"88",
          1545 => x"72",
          1546 => x"f0",
          1547 => x"08",
          1548 => x"d5",
          1549 => x"05",
          1550 => x"82",
          1551 => x"fc",
          1552 => x"81",
          1553 => x"72",
          1554 => x"38",
          1555 => x"08",
          1556 => x"08",
          1557 => x"f0",
          1558 => x"33",
          1559 => x"08",
          1560 => x"2d",
          1561 => x"08",
          1562 => x"2e",
          1563 => x"ff",
          1564 => x"f0",
          1565 => x"0c",
          1566 => x"82",
          1567 => x"82",
          1568 => x"53",
          1569 => x"90",
          1570 => x"72",
          1571 => x"e4",
          1572 => x"80",
          1573 => x"ff",
          1574 => x"f0",
          1575 => x"0c",
          1576 => x"08",
          1577 => x"70",
          1578 => x"08",
          1579 => x"53",
          1580 => x"08",
          1581 => x"82",
          1582 => x"87",
          1583 => x"d5",
          1584 => x"82",
          1585 => x"02",
          1586 => x"0c",
          1587 => x"80",
          1588 => x"f0",
          1589 => x"0c",
          1590 => x"08",
          1591 => x"85",
          1592 => x"81",
          1593 => x"32",
          1594 => x"51",
          1595 => x"53",
          1596 => x"8d",
          1597 => x"82",
          1598 => x"f4",
          1599 => x"f3",
          1600 => x"f0",
          1601 => x"08",
          1602 => x"82",
          1603 => x"88",
          1604 => x"05",
          1605 => x"08",
          1606 => x"53",
          1607 => x"f0",
          1608 => x"34",
          1609 => x"06",
          1610 => x"2e",
          1611 => x"d5",
          1612 => x"05",
          1613 => x"f0",
          1614 => x"08",
          1615 => x"f0",
          1616 => x"33",
          1617 => x"08",
          1618 => x"2d",
          1619 => x"08",
          1620 => x"2e",
          1621 => x"ff",
          1622 => x"f0",
          1623 => x"0c",
          1624 => x"82",
          1625 => x"f8",
          1626 => x"82",
          1627 => x"f4",
          1628 => x"82",
          1629 => x"f4",
          1630 => x"d5",
          1631 => x"3d",
          1632 => x"f0",
          1633 => x"d5",
          1634 => x"82",
          1635 => x"fe",
          1636 => x"f1",
          1637 => x"82",
          1638 => x"88",
          1639 => x"93",
          1640 => x"e4",
          1641 => x"d5",
          1642 => x"84",
          1643 => x"d5",
          1644 => x"82",
          1645 => x"02",
          1646 => x"0c",
          1647 => x"82",
          1648 => x"8c",
          1649 => x"11",
          1650 => x"2a",
          1651 => x"70",
          1652 => x"51",
          1653 => x"72",
          1654 => x"38",
          1655 => x"d5",
          1656 => x"05",
          1657 => x"39",
          1658 => x"08",
          1659 => x"85",
          1660 => x"82",
          1661 => x"06",
          1662 => x"53",
          1663 => x"80",
          1664 => x"d5",
          1665 => x"05",
          1666 => x"f0",
          1667 => x"08",
          1668 => x"14",
          1669 => x"08",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"08",
          1673 => x"f0",
          1674 => x"08",
          1675 => x"54",
          1676 => x"73",
          1677 => x"74",
          1678 => x"f0",
          1679 => x"08",
          1680 => x"81",
          1681 => x"0c",
          1682 => x"08",
          1683 => x"70",
          1684 => x"08",
          1685 => x"51",
          1686 => x"39",
          1687 => x"08",
          1688 => x"82",
          1689 => x"8c",
          1690 => x"82",
          1691 => x"88",
          1692 => x"81",
          1693 => x"90",
          1694 => x"54",
          1695 => x"82",
          1696 => x"53",
          1697 => x"82",
          1698 => x"8c",
          1699 => x"11",
          1700 => x"8c",
          1701 => x"d5",
          1702 => x"05",
          1703 => x"d5",
          1704 => x"05",
          1705 => x"8a",
          1706 => x"82",
          1707 => x"fc",
          1708 => x"d5",
          1709 => x"05",
          1710 => x"e4",
          1711 => x"0d",
          1712 => x"0c",
          1713 => x"f0",
          1714 => x"d5",
          1715 => x"3d",
          1716 => x"f0",
          1717 => x"08",
          1718 => x"70",
          1719 => x"81",
          1720 => x"51",
          1721 => x"2e",
          1722 => x"0b",
          1723 => x"08",
          1724 => x"83",
          1725 => x"d5",
          1726 => x"05",
          1727 => x"33",
          1728 => x"70",
          1729 => x"51",
          1730 => x"80",
          1731 => x"38",
          1732 => x"08",
          1733 => x"82",
          1734 => x"88",
          1735 => x"53",
          1736 => x"70",
          1737 => x"51",
          1738 => x"14",
          1739 => x"f0",
          1740 => x"08",
          1741 => x"81",
          1742 => x"0c",
          1743 => x"08",
          1744 => x"84",
          1745 => x"82",
          1746 => x"f8",
          1747 => x"51",
          1748 => x"39",
          1749 => x"08",
          1750 => x"85",
          1751 => x"82",
          1752 => x"06",
          1753 => x"52",
          1754 => x"80",
          1755 => x"d5",
          1756 => x"05",
          1757 => x"70",
          1758 => x"f0",
          1759 => x"0c",
          1760 => x"d5",
          1761 => x"05",
          1762 => x"82",
          1763 => x"88",
          1764 => x"d5",
          1765 => x"05",
          1766 => x"85",
          1767 => x"a0",
          1768 => x"71",
          1769 => x"ff",
          1770 => x"f0",
          1771 => x"0c",
          1772 => x"82",
          1773 => x"88",
          1774 => x"08",
          1775 => x"0c",
          1776 => x"39",
          1777 => x"08",
          1778 => x"82",
          1779 => x"88",
          1780 => x"94",
          1781 => x"52",
          1782 => x"d5",
          1783 => x"82",
          1784 => x"fc",
          1785 => x"82",
          1786 => x"fc",
          1787 => x"25",
          1788 => x"82",
          1789 => x"88",
          1790 => x"d5",
          1791 => x"05",
          1792 => x"f0",
          1793 => x"08",
          1794 => x"82",
          1795 => x"f0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"2e",
          1799 => x"95",
          1800 => x"f0",
          1801 => x"08",
          1802 => x"71",
          1803 => x"08",
          1804 => x"93",
          1805 => x"f0",
          1806 => x"08",
          1807 => x"71",
          1808 => x"08",
          1809 => x"82",
          1810 => x"f4",
          1811 => x"82",
          1812 => x"ec",
          1813 => x"13",
          1814 => x"82",
          1815 => x"f8",
          1816 => x"39",
          1817 => x"08",
          1818 => x"8c",
          1819 => x"05",
          1820 => x"82",
          1821 => x"fc",
          1822 => x"81",
          1823 => x"82",
          1824 => x"f8",
          1825 => x"51",
          1826 => x"f0",
          1827 => x"08",
          1828 => x"0c",
          1829 => x"82",
          1830 => x"04",
          1831 => x"08",
          1832 => x"f0",
          1833 => x"0d",
          1834 => x"08",
          1835 => x"82",
          1836 => x"fc",
          1837 => x"d5",
          1838 => x"05",
          1839 => x"f0",
          1840 => x"0c",
          1841 => x"08",
          1842 => x"80",
          1843 => x"38",
          1844 => x"08",
          1845 => x"82",
          1846 => x"fc",
          1847 => x"81",
          1848 => x"d5",
          1849 => x"05",
          1850 => x"f0",
          1851 => x"08",
          1852 => x"d5",
          1853 => x"05",
          1854 => x"81",
          1855 => x"d5",
          1856 => x"05",
          1857 => x"f0",
          1858 => x"08",
          1859 => x"f0",
          1860 => x"0c",
          1861 => x"08",
          1862 => x"82",
          1863 => x"90",
          1864 => x"82",
          1865 => x"f8",
          1866 => x"d5",
          1867 => x"05",
          1868 => x"82",
          1869 => x"90",
          1870 => x"d5",
          1871 => x"05",
          1872 => x"82",
          1873 => x"90",
          1874 => x"d5",
          1875 => x"05",
          1876 => x"81",
          1877 => x"d5",
          1878 => x"05",
          1879 => x"82",
          1880 => x"fc",
          1881 => x"d5",
          1882 => x"05",
          1883 => x"82",
          1884 => x"f8",
          1885 => x"d5",
          1886 => x"05",
          1887 => x"f0",
          1888 => x"08",
          1889 => x"33",
          1890 => x"ae",
          1891 => x"f0",
          1892 => x"08",
          1893 => x"d5",
          1894 => x"05",
          1895 => x"f0",
          1896 => x"08",
          1897 => x"d5",
          1898 => x"05",
          1899 => x"f0",
          1900 => x"08",
          1901 => x"38",
          1902 => x"08",
          1903 => x"51",
          1904 => x"d5",
          1905 => x"05",
          1906 => x"82",
          1907 => x"f8",
          1908 => x"d5",
          1909 => x"05",
          1910 => x"71",
          1911 => x"d5",
          1912 => x"05",
          1913 => x"82",
          1914 => x"fc",
          1915 => x"ad",
          1916 => x"f0",
          1917 => x"08",
          1918 => x"e4",
          1919 => x"3d",
          1920 => x"f0",
          1921 => x"d5",
          1922 => x"82",
          1923 => x"fe",
          1924 => x"d5",
          1925 => x"05",
          1926 => x"f0",
          1927 => x"0c",
          1928 => x"08",
          1929 => x"52",
          1930 => x"d5",
          1931 => x"05",
          1932 => x"82",
          1933 => x"fc",
          1934 => x"81",
          1935 => x"51",
          1936 => x"83",
          1937 => x"82",
          1938 => x"fc",
          1939 => x"05",
          1940 => x"08",
          1941 => x"82",
          1942 => x"fc",
          1943 => x"d5",
          1944 => x"05",
          1945 => x"82",
          1946 => x"51",
          1947 => x"82",
          1948 => x"04",
          1949 => x"08",
          1950 => x"f0",
          1951 => x"0d",
          1952 => x"08",
          1953 => x"82",
          1954 => x"fc",
          1955 => x"d5",
          1956 => x"05",
          1957 => x"33",
          1958 => x"08",
          1959 => x"81",
          1960 => x"f0",
          1961 => x"0c",
          1962 => x"08",
          1963 => x"53",
          1964 => x"34",
          1965 => x"08",
          1966 => x"81",
          1967 => x"f0",
          1968 => x"0c",
          1969 => x"06",
          1970 => x"2e",
          1971 => x"be",
          1972 => x"f0",
          1973 => x"08",
          1974 => x"e4",
          1975 => x"3d",
          1976 => x"f0",
          1977 => x"d5",
          1978 => x"82",
          1979 => x"fd",
          1980 => x"d5",
          1981 => x"05",
          1982 => x"f0",
          1983 => x"0c",
          1984 => x"08",
          1985 => x"82",
          1986 => x"f8",
          1987 => x"d5",
          1988 => x"05",
          1989 => x"80",
          1990 => x"d5",
          1991 => x"05",
          1992 => x"82",
          1993 => x"90",
          1994 => x"d5",
          1995 => x"05",
          1996 => x"82",
          1997 => x"90",
          1998 => x"d5",
          1999 => x"05",
          2000 => x"ba",
          2001 => x"f0",
          2002 => x"08",
          2003 => x"82",
          2004 => x"f8",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"fc",
          2009 => x"52",
          2010 => x"82",
          2011 => x"fc",
          2012 => x"05",
          2013 => x"08",
          2014 => x"ff",
          2015 => x"d5",
          2016 => x"05",
          2017 => x"d5",
          2018 => x"85",
          2019 => x"d5",
          2020 => x"82",
          2021 => x"02",
          2022 => x"0c",
          2023 => x"82",
          2024 => x"90",
          2025 => x"2e",
          2026 => x"82",
          2027 => x"8c",
          2028 => x"71",
          2029 => x"f0",
          2030 => x"08",
          2031 => x"d5",
          2032 => x"05",
          2033 => x"f0",
          2034 => x"08",
          2035 => x"81",
          2036 => x"54",
          2037 => x"71",
          2038 => x"80",
          2039 => x"d5",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"f0",
          2045 => x"0c",
          2046 => x"06",
          2047 => x"8d",
          2048 => x"82",
          2049 => x"fc",
          2050 => x"9b",
          2051 => x"f0",
          2052 => x"08",
          2053 => x"d5",
          2054 => x"05",
          2055 => x"f0",
          2056 => x"08",
          2057 => x"38",
          2058 => x"82",
          2059 => x"90",
          2060 => x"2e",
          2061 => x"82",
          2062 => x"88",
          2063 => x"33",
          2064 => x"8d",
          2065 => x"82",
          2066 => x"fc",
          2067 => x"d7",
          2068 => x"f0",
          2069 => x"08",
          2070 => x"d5",
          2071 => x"05",
          2072 => x"f0",
          2073 => x"08",
          2074 => x"52",
          2075 => x"81",
          2076 => x"f0",
          2077 => x"0c",
          2078 => x"d5",
          2079 => x"05",
          2080 => x"82",
          2081 => x"8c",
          2082 => x"33",
          2083 => x"70",
          2084 => x"08",
          2085 => x"53",
          2086 => x"53",
          2087 => x"0b",
          2088 => x"08",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"d5",
          2092 => x"3d",
          2093 => x"f0",
          2094 => x"d5",
          2095 => x"82",
          2096 => x"fa",
          2097 => x"d5",
          2098 => x"05",
          2099 => x"d5",
          2100 => x"05",
          2101 => x"8d",
          2102 => x"e4",
          2103 => x"d5",
          2104 => x"05",
          2105 => x"f0",
          2106 => x"08",
          2107 => x"53",
          2108 => x"e2",
          2109 => x"d5",
          2110 => x"82",
          2111 => x"fc",
          2112 => x"82",
          2113 => x"fc",
          2114 => x"38",
          2115 => x"d5",
          2116 => x"05",
          2117 => x"82",
          2118 => x"fc",
          2119 => x"d5",
          2120 => x"05",
          2121 => x"80",
          2122 => x"d5",
          2123 => x"05",
          2124 => x"d5",
          2125 => x"05",
          2126 => x"d5",
          2127 => x"05",
          2128 => x"a2",
          2129 => x"e4",
          2130 => x"d5",
          2131 => x"05",
          2132 => x"d5",
          2133 => x"05",
          2134 => x"e4",
          2135 => x"0d",
          2136 => x"0c",
          2137 => x"f0",
          2138 => x"d5",
          2139 => x"3d",
          2140 => x"f0",
          2141 => x"08",
          2142 => x"08",
          2143 => x"82",
          2144 => x"8c",
          2145 => x"38",
          2146 => x"d5",
          2147 => x"05",
          2148 => x"39",
          2149 => x"08",
          2150 => x"52",
          2151 => x"d5",
          2152 => x"05",
          2153 => x"82",
          2154 => x"f8",
          2155 => x"81",
          2156 => x"51",
          2157 => x"9f",
          2158 => x"f0",
          2159 => x"08",
          2160 => x"d5",
          2161 => x"05",
          2162 => x"f0",
          2163 => x"08",
          2164 => x"38",
          2165 => x"82",
          2166 => x"f8",
          2167 => x"05",
          2168 => x"08",
          2169 => x"82",
          2170 => x"f8",
          2171 => x"d5",
          2172 => x"05",
          2173 => x"82",
          2174 => x"fc",
          2175 => x"82",
          2176 => x"fc",
          2177 => x"d5",
          2178 => x"3d",
          2179 => x"f0",
          2180 => x"d5",
          2181 => x"82",
          2182 => x"fe",
          2183 => x"d5",
          2184 => x"05",
          2185 => x"f0",
          2186 => x"0c",
          2187 => x"08",
          2188 => x"80",
          2189 => x"38",
          2190 => x"08",
          2191 => x"81",
          2192 => x"f0",
          2193 => x"0c",
          2194 => x"08",
          2195 => x"ff",
          2196 => x"f0",
          2197 => x"0c",
          2198 => x"08",
          2199 => x"80",
          2200 => x"82",
          2201 => x"8c",
          2202 => x"70",
          2203 => x"08",
          2204 => x"52",
          2205 => x"34",
          2206 => x"08",
          2207 => x"81",
          2208 => x"f0",
          2209 => x"0c",
          2210 => x"82",
          2211 => x"88",
          2212 => x"82",
          2213 => x"51",
          2214 => x"82",
          2215 => x"04",
          2216 => x"08",
          2217 => x"f0",
          2218 => x"0d",
          2219 => x"d5",
          2220 => x"05",
          2221 => x"f0",
          2222 => x"08",
          2223 => x"38",
          2224 => x"08",
          2225 => x"30",
          2226 => x"08",
          2227 => x"80",
          2228 => x"f0",
          2229 => x"0c",
          2230 => x"08",
          2231 => x"8a",
          2232 => x"82",
          2233 => x"f4",
          2234 => x"d5",
          2235 => x"05",
          2236 => x"f0",
          2237 => x"0c",
          2238 => x"08",
          2239 => x"80",
          2240 => x"82",
          2241 => x"8c",
          2242 => x"82",
          2243 => x"8c",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"fc",
          2248 => x"38",
          2249 => x"d5",
          2250 => x"05",
          2251 => x"f0",
          2252 => x"08",
          2253 => x"08",
          2254 => x"80",
          2255 => x"f0",
          2256 => x"08",
          2257 => x"f0",
          2258 => x"08",
          2259 => x"3f",
          2260 => x"08",
          2261 => x"f0",
          2262 => x"0c",
          2263 => x"f0",
          2264 => x"08",
          2265 => x"38",
          2266 => x"08",
          2267 => x"30",
          2268 => x"08",
          2269 => x"82",
          2270 => x"f8",
          2271 => x"82",
          2272 => x"54",
          2273 => x"82",
          2274 => x"04",
          2275 => x"08",
          2276 => x"f0",
          2277 => x"0d",
          2278 => x"d5",
          2279 => x"05",
          2280 => x"f0",
          2281 => x"08",
          2282 => x"38",
          2283 => x"08",
          2284 => x"30",
          2285 => x"08",
          2286 => x"81",
          2287 => x"f0",
          2288 => x"0c",
          2289 => x"08",
          2290 => x"80",
          2291 => x"82",
          2292 => x"8c",
          2293 => x"82",
          2294 => x"8c",
          2295 => x"53",
          2296 => x"08",
          2297 => x"52",
          2298 => x"08",
          2299 => x"51",
          2300 => x"82",
          2301 => x"70",
          2302 => x"08",
          2303 => x"54",
          2304 => x"08",
          2305 => x"80",
          2306 => x"82",
          2307 => x"f8",
          2308 => x"82",
          2309 => x"f8",
          2310 => x"d5",
          2311 => x"05",
          2312 => x"d5",
          2313 => x"87",
          2314 => x"d5",
          2315 => x"82",
          2316 => x"02",
          2317 => x"0c",
          2318 => x"80",
          2319 => x"f0",
          2320 => x"08",
          2321 => x"f0",
          2322 => x"08",
          2323 => x"3f",
          2324 => x"08",
          2325 => x"e4",
          2326 => x"3d",
          2327 => x"f0",
          2328 => x"d5",
          2329 => x"82",
          2330 => x"fd",
          2331 => x"53",
          2332 => x"08",
          2333 => x"52",
          2334 => x"08",
          2335 => x"51",
          2336 => x"d5",
          2337 => x"82",
          2338 => x"54",
          2339 => x"82",
          2340 => x"04",
          2341 => x"08",
          2342 => x"f0",
          2343 => x"0d",
          2344 => x"d5",
          2345 => x"05",
          2346 => x"82",
          2347 => x"f8",
          2348 => x"d5",
          2349 => x"05",
          2350 => x"f0",
          2351 => x"08",
          2352 => x"82",
          2353 => x"fc",
          2354 => x"2e",
          2355 => x"0b",
          2356 => x"08",
          2357 => x"24",
          2358 => x"d5",
          2359 => x"05",
          2360 => x"d5",
          2361 => x"05",
          2362 => x"f0",
          2363 => x"08",
          2364 => x"f0",
          2365 => x"0c",
          2366 => x"82",
          2367 => x"fc",
          2368 => x"2e",
          2369 => x"82",
          2370 => x"8c",
          2371 => x"d5",
          2372 => x"05",
          2373 => x"38",
          2374 => x"08",
          2375 => x"82",
          2376 => x"8c",
          2377 => x"82",
          2378 => x"88",
          2379 => x"d5",
          2380 => x"05",
          2381 => x"f0",
          2382 => x"08",
          2383 => x"f0",
          2384 => x"0c",
          2385 => x"08",
          2386 => x"81",
          2387 => x"f0",
          2388 => x"0c",
          2389 => x"08",
          2390 => x"81",
          2391 => x"f0",
          2392 => x"0c",
          2393 => x"82",
          2394 => x"90",
          2395 => x"2e",
          2396 => x"d5",
          2397 => x"05",
          2398 => x"d5",
          2399 => x"05",
          2400 => x"39",
          2401 => x"08",
          2402 => x"70",
          2403 => x"08",
          2404 => x"51",
          2405 => x"08",
          2406 => x"82",
          2407 => x"85",
          2408 => x"d5",
          2409 => x"82",
          2410 => x"02",
          2411 => x"0c",
          2412 => x"80",
          2413 => x"f0",
          2414 => x"34",
          2415 => x"08",
          2416 => x"53",
          2417 => x"82",
          2418 => x"88",
          2419 => x"08",
          2420 => x"33",
          2421 => x"d5",
          2422 => x"05",
          2423 => x"ff",
          2424 => x"a0",
          2425 => x"06",
          2426 => x"d5",
          2427 => x"05",
          2428 => x"81",
          2429 => x"53",
          2430 => x"d5",
          2431 => x"05",
          2432 => x"ad",
          2433 => x"06",
          2434 => x"0b",
          2435 => x"08",
          2436 => x"82",
          2437 => x"88",
          2438 => x"08",
          2439 => x"0c",
          2440 => x"53",
          2441 => x"d5",
          2442 => x"05",
          2443 => x"f0",
          2444 => x"33",
          2445 => x"2e",
          2446 => x"81",
          2447 => x"d5",
          2448 => x"05",
          2449 => x"81",
          2450 => x"70",
          2451 => x"72",
          2452 => x"f0",
          2453 => x"34",
          2454 => x"08",
          2455 => x"82",
          2456 => x"e8",
          2457 => x"d5",
          2458 => x"05",
          2459 => x"2e",
          2460 => x"d5",
          2461 => x"05",
          2462 => x"2e",
          2463 => x"cd",
          2464 => x"82",
          2465 => x"f4",
          2466 => x"d5",
          2467 => x"05",
          2468 => x"81",
          2469 => x"70",
          2470 => x"72",
          2471 => x"f0",
          2472 => x"34",
          2473 => x"82",
          2474 => x"f0",
          2475 => x"34",
          2476 => x"08",
          2477 => x"70",
          2478 => x"71",
          2479 => x"51",
          2480 => x"82",
          2481 => x"f8",
          2482 => x"fe",
          2483 => x"f0",
          2484 => x"33",
          2485 => x"26",
          2486 => x"0b",
          2487 => x"08",
          2488 => x"83",
          2489 => x"d5",
          2490 => x"05",
          2491 => x"73",
          2492 => x"82",
          2493 => x"f8",
          2494 => x"72",
          2495 => x"38",
          2496 => x"0b",
          2497 => x"08",
          2498 => x"82",
          2499 => x"0b",
          2500 => x"08",
          2501 => x"b2",
          2502 => x"f0",
          2503 => x"33",
          2504 => x"27",
          2505 => x"d5",
          2506 => x"05",
          2507 => x"b9",
          2508 => x"8d",
          2509 => x"82",
          2510 => x"ec",
          2511 => x"a5",
          2512 => x"82",
          2513 => x"f4",
          2514 => x"0b",
          2515 => x"08",
          2516 => x"82",
          2517 => x"f8",
          2518 => x"a0",
          2519 => x"cf",
          2520 => x"f0",
          2521 => x"33",
          2522 => x"73",
          2523 => x"82",
          2524 => x"f8",
          2525 => x"11",
          2526 => x"82",
          2527 => x"f8",
          2528 => x"d5",
          2529 => x"05",
          2530 => x"51",
          2531 => x"d5",
          2532 => x"05",
          2533 => x"f0",
          2534 => x"33",
          2535 => x"27",
          2536 => x"d5",
          2537 => x"05",
          2538 => x"51",
          2539 => x"d5",
          2540 => x"05",
          2541 => x"f0",
          2542 => x"33",
          2543 => x"26",
          2544 => x"0b",
          2545 => x"08",
          2546 => x"81",
          2547 => x"d5",
          2548 => x"05",
          2549 => x"f0",
          2550 => x"33",
          2551 => x"74",
          2552 => x"80",
          2553 => x"f0",
          2554 => x"0c",
          2555 => x"82",
          2556 => x"f4",
          2557 => x"82",
          2558 => x"fc",
          2559 => x"82",
          2560 => x"f8",
          2561 => x"12",
          2562 => x"08",
          2563 => x"82",
          2564 => x"88",
          2565 => x"08",
          2566 => x"0c",
          2567 => x"51",
          2568 => x"72",
          2569 => x"f0",
          2570 => x"34",
          2571 => x"82",
          2572 => x"f0",
          2573 => x"72",
          2574 => x"38",
          2575 => x"08",
          2576 => x"30",
          2577 => x"08",
          2578 => x"82",
          2579 => x"8c",
          2580 => x"d5",
          2581 => x"05",
          2582 => x"53",
          2583 => x"d5",
          2584 => x"05",
          2585 => x"f0",
          2586 => x"08",
          2587 => x"0c",
          2588 => x"82",
          2589 => x"04",
          2590 => x"08",
          2591 => x"f0",
          2592 => x"0d",
          2593 => x"d5",
          2594 => x"05",
          2595 => x"f0",
          2596 => x"08",
          2597 => x"0c",
          2598 => x"08",
          2599 => x"70",
          2600 => x"72",
          2601 => x"82",
          2602 => x"f8",
          2603 => x"81",
          2604 => x"72",
          2605 => x"81",
          2606 => x"82",
          2607 => x"88",
          2608 => x"08",
          2609 => x"0c",
          2610 => x"82",
          2611 => x"f8",
          2612 => x"72",
          2613 => x"81",
          2614 => x"81",
          2615 => x"f0",
          2616 => x"34",
          2617 => x"08",
          2618 => x"70",
          2619 => x"71",
          2620 => x"51",
          2621 => x"82",
          2622 => x"f8",
          2623 => x"d5",
          2624 => x"05",
          2625 => x"b0",
          2626 => x"06",
          2627 => x"82",
          2628 => x"88",
          2629 => x"08",
          2630 => x"0c",
          2631 => x"53",
          2632 => x"d5",
          2633 => x"05",
          2634 => x"f0",
          2635 => x"33",
          2636 => x"08",
          2637 => x"82",
          2638 => x"e8",
          2639 => x"e2",
          2640 => x"82",
          2641 => x"e8",
          2642 => x"f8",
          2643 => x"80",
          2644 => x"0b",
          2645 => x"08",
          2646 => x"82",
          2647 => x"88",
          2648 => x"08",
          2649 => x"0c",
          2650 => x"53",
          2651 => x"d5",
          2652 => x"05",
          2653 => x"39",
          2654 => x"d5",
          2655 => x"05",
          2656 => x"f0",
          2657 => x"08",
          2658 => x"05",
          2659 => x"08",
          2660 => x"33",
          2661 => x"08",
          2662 => x"80",
          2663 => x"d5",
          2664 => x"05",
          2665 => x"a0",
          2666 => x"81",
          2667 => x"f0",
          2668 => x"0c",
          2669 => x"82",
          2670 => x"f8",
          2671 => x"af",
          2672 => x"38",
          2673 => x"08",
          2674 => x"53",
          2675 => x"83",
          2676 => x"80",
          2677 => x"f0",
          2678 => x"0c",
          2679 => x"88",
          2680 => x"f0",
          2681 => x"34",
          2682 => x"d5",
          2683 => x"05",
          2684 => x"73",
          2685 => x"82",
          2686 => x"f8",
          2687 => x"72",
          2688 => x"38",
          2689 => x"0b",
          2690 => x"08",
          2691 => x"82",
          2692 => x"0b",
          2693 => x"08",
          2694 => x"80",
          2695 => x"f0",
          2696 => x"0c",
          2697 => x"08",
          2698 => x"53",
          2699 => x"81",
          2700 => x"d5",
          2701 => x"05",
          2702 => x"e0",
          2703 => x"38",
          2704 => x"08",
          2705 => x"e0",
          2706 => x"72",
          2707 => x"08",
          2708 => x"82",
          2709 => x"f8",
          2710 => x"11",
          2711 => x"82",
          2712 => x"f8",
          2713 => x"d5",
          2714 => x"05",
          2715 => x"73",
          2716 => x"82",
          2717 => x"f8",
          2718 => x"11",
          2719 => x"82",
          2720 => x"f8",
          2721 => x"d5",
          2722 => x"05",
          2723 => x"89",
          2724 => x"80",
          2725 => x"f0",
          2726 => x"0c",
          2727 => x"82",
          2728 => x"f8",
          2729 => x"d5",
          2730 => x"05",
          2731 => x"72",
          2732 => x"38",
          2733 => x"d5",
          2734 => x"05",
          2735 => x"39",
          2736 => x"08",
          2737 => x"70",
          2738 => x"08",
          2739 => x"29",
          2740 => x"08",
          2741 => x"70",
          2742 => x"f0",
          2743 => x"0c",
          2744 => x"08",
          2745 => x"70",
          2746 => x"71",
          2747 => x"51",
          2748 => x"53",
          2749 => x"d5",
          2750 => x"05",
          2751 => x"39",
          2752 => x"08",
          2753 => x"53",
          2754 => x"90",
          2755 => x"f0",
          2756 => x"08",
          2757 => x"f0",
          2758 => x"0c",
          2759 => x"08",
          2760 => x"82",
          2761 => x"fc",
          2762 => x"0c",
          2763 => x"82",
          2764 => x"ec",
          2765 => x"d5",
          2766 => x"05",
          2767 => x"e4",
          2768 => x"0d",
          2769 => x"0c",
          2770 => x"0d",
          2771 => x"70",
          2772 => x"74",
          2773 => x"df",
          2774 => x"77",
          2775 => x"85",
          2776 => x"80",
          2777 => x"33",
          2778 => x"2e",
          2779 => x"86",
          2780 => x"55",
          2781 => x"57",
          2782 => x"82",
          2783 => x"70",
          2784 => x"e5",
          2785 => x"d5",
          2786 => x"d5",
          2787 => x"75",
          2788 => x"52",
          2789 => x"3f",
          2790 => x"08",
          2791 => x"16",
          2792 => x"81",
          2793 => x"38",
          2794 => x"81",
          2795 => x"54",
          2796 => x"c4",
          2797 => x"73",
          2798 => x"0c",
          2799 => x"04",
          2800 => x"73",
          2801 => x"26",
          2802 => x"71",
          2803 => x"ad",
          2804 => x"71",
          2805 => x"b3",
          2806 => x"80",
          2807 => x"a8",
          2808 => x"39",
          2809 => x"51",
          2810 => x"82",
          2811 => x"80",
          2812 => x"b3",
          2813 => x"e4",
          2814 => x"e8",
          2815 => x"39",
          2816 => x"51",
          2817 => x"82",
          2818 => x"80",
          2819 => x"b4",
          2820 => x"c8",
          2821 => x"bc",
          2822 => x"39",
          2823 => x"51",
          2824 => x"b4",
          2825 => x"39",
          2826 => x"51",
          2827 => x"b5",
          2828 => x"39",
          2829 => x"51",
          2830 => x"b5",
          2831 => x"39",
          2832 => x"51",
          2833 => x"b6",
          2834 => x"39",
          2835 => x"51",
          2836 => x"b6",
          2837 => x"39",
          2838 => x"51",
          2839 => x"83",
          2840 => x"fb",
          2841 => x"79",
          2842 => x"87",
          2843 => x"38",
          2844 => x"87",
          2845 => x"90",
          2846 => x"52",
          2847 => x"af",
          2848 => x"e4",
          2849 => x"51",
          2850 => x"82",
          2851 => x"54",
          2852 => x"52",
          2853 => x"51",
          2854 => x"3f",
          2855 => x"04",
          2856 => x"66",
          2857 => x"80",
          2858 => x"5b",
          2859 => x"78",
          2860 => x"07",
          2861 => x"57",
          2862 => x"56",
          2863 => x"26",
          2864 => x"56",
          2865 => x"70",
          2866 => x"51",
          2867 => x"74",
          2868 => x"81",
          2869 => x"8c",
          2870 => x"56",
          2871 => x"3f",
          2872 => x"08",
          2873 => x"e4",
          2874 => x"82",
          2875 => x"87",
          2876 => x"0c",
          2877 => x"08",
          2878 => x"d4",
          2879 => x"80",
          2880 => x"75",
          2881 => x"b5",
          2882 => x"e4",
          2883 => x"d5",
          2884 => x"38",
          2885 => x"80",
          2886 => x"74",
          2887 => x"59",
          2888 => x"96",
          2889 => x"51",
          2890 => x"3f",
          2891 => x"78",
          2892 => x"7b",
          2893 => x"2a",
          2894 => x"57",
          2895 => x"80",
          2896 => x"82",
          2897 => x"87",
          2898 => x"08",
          2899 => x"fe",
          2900 => x"56",
          2901 => x"e4",
          2902 => x"0d",
          2903 => x"0d",
          2904 => x"05",
          2905 => x"58",
          2906 => x"80",
          2907 => x"7a",
          2908 => x"3f",
          2909 => x"08",
          2910 => x"80",
          2911 => x"76",
          2912 => x"38",
          2913 => x"f1",
          2914 => x"55",
          2915 => x"d5",
          2916 => x"52",
          2917 => x"2d",
          2918 => x"08",
          2919 => x"78",
          2920 => x"d5",
          2921 => x"3d",
          2922 => x"3d",
          2923 => x"63",
          2924 => x"80",
          2925 => x"73",
          2926 => x"41",
          2927 => x"5e",
          2928 => x"52",
          2929 => x"51",
          2930 => x"3f",
          2931 => x"51",
          2932 => x"3f",
          2933 => x"79",
          2934 => x"38",
          2935 => x"89",
          2936 => x"2e",
          2937 => x"c6",
          2938 => x"53",
          2939 => x"8e",
          2940 => x"52",
          2941 => x"51",
          2942 => x"3f",
          2943 => x"b7",
          2944 => x"b7",
          2945 => x"15",
          2946 => x"39",
          2947 => x"72",
          2948 => x"38",
          2949 => x"82",
          2950 => x"ff",
          2951 => x"89",
          2952 => x"90",
          2953 => x"b1",
          2954 => x"55",
          2955 => x"18",
          2956 => x"27",
          2957 => x"33",
          2958 => x"9c",
          2959 => x"99",
          2960 => x"82",
          2961 => x"ff",
          2962 => x"81",
          2963 => x"f1",
          2964 => x"a0",
          2965 => x"3f",
          2966 => x"82",
          2967 => x"ff",
          2968 => x"80",
          2969 => x"27",
          2970 => x"74",
          2971 => x"55",
          2972 => x"72",
          2973 => x"38",
          2974 => x"53",
          2975 => x"83",
          2976 => x"75",
          2977 => x"81",
          2978 => x"53",
          2979 => x"90",
          2980 => x"fe",
          2981 => x"82",
          2982 => x"52",
          2983 => x"39",
          2984 => x"08",
          2985 => x"d6",
          2986 => x"15",
          2987 => x"39",
          2988 => x"51",
          2989 => x"78",
          2990 => x"5c",
          2991 => x"3f",
          2992 => x"08",
          2993 => x"98",
          2994 => x"76",
          2995 => x"81",
          2996 => x"9c",
          2997 => x"d5",
          2998 => x"2b",
          2999 => x"70",
          3000 => x"30",
          3001 => x"70",
          3002 => x"07",
          3003 => x"06",
          3004 => x"59",
          3005 => x"80",
          3006 => x"38",
          3007 => x"09",
          3008 => x"38",
          3009 => x"39",
          3010 => x"72",
          3011 => x"b2",
          3012 => x"72",
          3013 => x"0c",
          3014 => x"04",
          3015 => x"02",
          3016 => x"82",
          3017 => x"82",
          3018 => x"55",
          3019 => x"3f",
          3020 => x"22",
          3021 => x"3f",
          3022 => x"54",
          3023 => x"53",
          3024 => x"33",
          3025 => x"d4",
          3026 => x"8d",
          3027 => x"2e",
          3028 => x"97",
          3029 => x"0d",
          3030 => x"0d",
          3031 => x"80",
          3032 => x"ff",
          3033 => x"98",
          3034 => x"b7",
          3035 => x"e2",
          3036 => x"98",
          3037 => x"81",
          3038 => x"06",
          3039 => x"80",
          3040 => x"81",
          3041 => x"3f",
          3042 => x"51",
          3043 => x"80",
          3044 => x"3f",
          3045 => x"70",
          3046 => x"52",
          3047 => x"92",
          3048 => x"98",
          3049 => x"b8",
          3050 => x"a6",
          3051 => x"98",
          3052 => x"83",
          3053 => x"06",
          3054 => x"80",
          3055 => x"81",
          3056 => x"3f",
          3057 => x"51",
          3058 => x"80",
          3059 => x"3f",
          3060 => x"70",
          3061 => x"52",
          3062 => x"92",
          3063 => x"97",
          3064 => x"b8",
          3065 => x"ea",
          3066 => x"97",
          3067 => x"85",
          3068 => x"06",
          3069 => x"80",
          3070 => x"81",
          3071 => x"3f",
          3072 => x"51",
          3073 => x"80",
          3074 => x"3f",
          3075 => x"70",
          3076 => x"52",
          3077 => x"92",
          3078 => x"97",
          3079 => x"b8",
          3080 => x"ae",
          3081 => x"97",
          3082 => x"87",
          3083 => x"06",
          3084 => x"80",
          3085 => x"81",
          3086 => x"3f",
          3087 => x"51",
          3088 => x"80",
          3089 => x"3f",
          3090 => x"70",
          3091 => x"52",
          3092 => x"92",
          3093 => x"96",
          3094 => x"b9",
          3095 => x"f2",
          3096 => x"96",
          3097 => x"83",
          3098 => x"0d",
          3099 => x"0d",
          3100 => x"05",
          3101 => x"70",
          3102 => x"80",
          3103 => x"e3",
          3104 => x"0b",
          3105 => x"33",
          3106 => x"38",
          3107 => x"b9",
          3108 => x"ec",
          3109 => x"8a",
          3110 => x"d5",
          3111 => x"70",
          3112 => x"08",
          3113 => x"82",
          3114 => x"51",
          3115 => x"0b",
          3116 => x"34",
          3117 => x"d0",
          3118 => x"73",
          3119 => x"81",
          3120 => x"82",
          3121 => x"74",
          3122 => x"81",
          3123 => x"82",
          3124 => x"80",
          3125 => x"82",
          3126 => x"51",
          3127 => x"91",
          3128 => x"f4",
          3129 => x"f0",
          3130 => x"0b",
          3131 => x"d8",
          3132 => x"82",
          3133 => x"54",
          3134 => x"09",
          3135 => x"38",
          3136 => x"53",
          3137 => x"51",
          3138 => x"80",
          3139 => x"e4",
          3140 => x"0d",
          3141 => x"0d",
          3142 => x"5e",
          3143 => x"ec",
          3144 => x"81",
          3145 => x"80",
          3146 => x"82",
          3147 => x"81",
          3148 => x"78",
          3149 => x"81",
          3150 => x"97",
          3151 => x"53",
          3152 => x"52",
          3153 => x"9e",
          3154 => x"78",
          3155 => x"90",
          3156 => x"a3",
          3157 => x"e4",
          3158 => x"88",
          3159 => x"e8",
          3160 => x"39",
          3161 => x"5e",
          3162 => x"51",
          3163 => x"3f",
          3164 => x"47",
          3165 => x"52",
          3166 => x"f1",
          3167 => x"ff",
          3168 => x"f3",
          3169 => x"d5",
          3170 => x"2b",
          3171 => x"51",
          3172 => x"c2",
          3173 => x"38",
          3174 => x"24",
          3175 => x"bd",
          3176 => x"38",
          3177 => x"90",
          3178 => x"2e",
          3179 => x"78",
          3180 => x"da",
          3181 => x"39",
          3182 => x"2e",
          3183 => x"78",
          3184 => x"85",
          3185 => x"bf",
          3186 => x"38",
          3187 => x"78",
          3188 => x"89",
          3189 => x"80",
          3190 => x"38",
          3191 => x"2e",
          3192 => x"78",
          3193 => x"89",
          3194 => x"a1",
          3195 => x"83",
          3196 => x"38",
          3197 => x"24",
          3198 => x"81",
          3199 => x"ed",
          3200 => x"39",
          3201 => x"2e",
          3202 => x"8a",
          3203 => x"3d",
          3204 => x"53",
          3205 => x"51",
          3206 => x"82",
          3207 => x"80",
          3208 => x"38",
          3209 => x"fc",
          3210 => x"84",
          3211 => x"c8",
          3212 => x"e4",
          3213 => x"fe",
          3214 => x"3d",
          3215 => x"53",
          3216 => x"51",
          3217 => x"82",
          3218 => x"86",
          3219 => x"e4",
          3220 => x"ba",
          3221 => x"af",
          3222 => x"64",
          3223 => x"7b",
          3224 => x"38",
          3225 => x"7a",
          3226 => x"5c",
          3227 => x"26",
          3228 => x"db",
          3229 => x"ff",
          3230 => x"ff",
          3231 => x"eb",
          3232 => x"d5",
          3233 => x"2e",
          3234 => x"b5",
          3235 => x"11",
          3236 => x"05",
          3237 => x"3f",
          3238 => x"08",
          3239 => x"c8",
          3240 => x"fe",
          3241 => x"ff",
          3242 => x"eb",
          3243 => x"d5",
          3244 => x"2e",
          3245 => x"82",
          3246 => x"ff",
          3247 => x"64",
          3248 => x"27",
          3249 => x"62",
          3250 => x"81",
          3251 => x"79",
          3252 => x"05",
          3253 => x"b5",
          3254 => x"11",
          3255 => x"05",
          3256 => x"3f",
          3257 => x"08",
          3258 => x"fc",
          3259 => x"fe",
          3260 => x"ff",
          3261 => x"ea",
          3262 => x"d5",
          3263 => x"2e",
          3264 => x"b5",
          3265 => x"11",
          3266 => x"05",
          3267 => x"3f",
          3268 => x"08",
          3269 => x"d0",
          3270 => x"c0",
          3271 => x"b9",
          3272 => x"79",
          3273 => x"38",
          3274 => x"7b",
          3275 => x"5b",
          3276 => x"92",
          3277 => x"7a",
          3278 => x"53",
          3279 => x"ba",
          3280 => x"ad",
          3281 => x"1a",
          3282 => x"44",
          3283 => x"8a",
          3284 => x"3f",
          3285 => x"b5",
          3286 => x"11",
          3287 => x"05",
          3288 => x"3f",
          3289 => x"08",
          3290 => x"82",
          3291 => x"59",
          3292 => x"89",
          3293 => x"80",
          3294 => x"cd",
          3295 => x"c9",
          3296 => x"80",
          3297 => x"82",
          3298 => x"45",
          3299 => x"d4",
          3300 => x"78",
          3301 => x"38",
          3302 => x"08",
          3303 => x"82",
          3304 => x"59",
          3305 => x"88",
          3306 => x"98",
          3307 => x"39",
          3308 => x"33",
          3309 => x"2e",
          3310 => x"d4",
          3311 => x"89",
          3312 => x"b0",
          3313 => x"05",
          3314 => x"fe",
          3315 => x"ff",
          3316 => x"e9",
          3317 => x"d5",
          3318 => x"de",
          3319 => x"c8",
          3320 => x"80",
          3321 => x"82",
          3322 => x"44",
          3323 => x"82",
          3324 => x"59",
          3325 => x"88",
          3326 => x"8c",
          3327 => x"39",
          3328 => x"33",
          3329 => x"2e",
          3330 => x"d4",
          3331 => x"aa",
          3332 => x"cb",
          3333 => x"80",
          3334 => x"82",
          3335 => x"44",
          3336 => x"d4",
          3337 => x"78",
          3338 => x"38",
          3339 => x"08",
          3340 => x"82",
          3341 => x"88",
          3342 => x"3d",
          3343 => x"53",
          3344 => x"51",
          3345 => x"82",
          3346 => x"80",
          3347 => x"80",
          3348 => x"7a",
          3349 => x"38",
          3350 => x"90",
          3351 => x"70",
          3352 => x"2a",
          3353 => x"51",
          3354 => x"78",
          3355 => x"38",
          3356 => x"83",
          3357 => x"82",
          3358 => x"c6",
          3359 => x"55",
          3360 => x"53",
          3361 => x"51",
          3362 => x"82",
          3363 => x"87",
          3364 => x"3d",
          3365 => x"53",
          3366 => x"51",
          3367 => x"82",
          3368 => x"80",
          3369 => x"38",
          3370 => x"fc",
          3371 => x"84",
          3372 => x"c4",
          3373 => x"e4",
          3374 => x"a4",
          3375 => x"02",
          3376 => x"33",
          3377 => x"81",
          3378 => x"3d",
          3379 => x"53",
          3380 => x"51",
          3381 => x"82",
          3382 => x"e1",
          3383 => x"39",
          3384 => x"54",
          3385 => x"84",
          3386 => x"ed",
          3387 => x"c4",
          3388 => x"f8",
          3389 => x"ff",
          3390 => x"79",
          3391 => x"59",
          3392 => x"f8",
          3393 => x"79",
          3394 => x"b5",
          3395 => x"11",
          3396 => x"05",
          3397 => x"3f",
          3398 => x"08",
          3399 => x"38",
          3400 => x"80",
          3401 => x"79",
          3402 => x"05",
          3403 => x"39",
          3404 => x"51",
          3405 => x"ff",
          3406 => x"3d",
          3407 => x"53",
          3408 => x"51",
          3409 => x"82",
          3410 => x"80",
          3411 => x"38",
          3412 => x"f0",
          3413 => x"84",
          3414 => x"cb",
          3415 => x"e4",
          3416 => x"a6",
          3417 => x"02",
          3418 => x"22",
          3419 => x"05",
          3420 => x"42",
          3421 => x"f0",
          3422 => x"84",
          3423 => x"a7",
          3424 => x"e4",
          3425 => x"f7",
          3426 => x"70",
          3427 => x"82",
          3428 => x"ff",
          3429 => x"82",
          3430 => x"53",
          3431 => x"79",
          3432 => x"8a",
          3433 => x"79",
          3434 => x"ae",
          3435 => x"38",
          3436 => x"87",
          3437 => x"05",
          3438 => x"b5",
          3439 => x"11",
          3440 => x"05",
          3441 => x"3f",
          3442 => x"08",
          3443 => x"38",
          3444 => x"80",
          3445 => x"79",
          3446 => x"5b",
          3447 => x"ff",
          3448 => x"bb",
          3449 => x"fc",
          3450 => x"39",
          3451 => x"f4",
          3452 => x"84",
          3453 => x"af",
          3454 => x"e4",
          3455 => x"f6",
          3456 => x"3d",
          3457 => x"53",
          3458 => x"51",
          3459 => x"82",
          3460 => x"80",
          3461 => x"61",
          3462 => x"59",
          3463 => x"42",
          3464 => x"f0",
          3465 => x"84",
          3466 => x"fb",
          3467 => x"e4",
          3468 => x"f6",
          3469 => x"70",
          3470 => x"82",
          3471 => x"ff",
          3472 => x"82",
          3473 => x"53",
          3474 => x"79",
          3475 => x"de",
          3476 => x"79",
          3477 => x"ae",
          3478 => x"38",
          3479 => x"9b",
          3480 => x"fe",
          3481 => x"ff",
          3482 => x"de",
          3483 => x"d5",
          3484 => x"2e",
          3485 => x"61",
          3486 => x"61",
          3487 => x"ff",
          3488 => x"bb",
          3489 => x"dc",
          3490 => x"39",
          3491 => x"80",
          3492 => x"84",
          3493 => x"e0",
          3494 => x"e4",
          3495 => x"f5",
          3496 => x"52",
          3497 => x"51",
          3498 => x"3f",
          3499 => x"04",
          3500 => x"80",
          3501 => x"84",
          3502 => x"bc",
          3503 => x"e4",
          3504 => x"f5",
          3505 => x"52",
          3506 => x"51",
          3507 => x"3f",
          3508 => x"2d",
          3509 => x"08",
          3510 => x"8c",
          3511 => x"e4",
          3512 => x"bb",
          3513 => x"a5",
          3514 => x"fc",
          3515 => x"84",
          3516 => x"3f",
          3517 => x"3f",
          3518 => x"82",
          3519 => x"c1",
          3520 => x"59",
          3521 => x"91",
          3522 => x"dc",
          3523 => x"33",
          3524 => x"2e",
          3525 => x"80",
          3526 => x"51",
          3527 => x"82",
          3528 => x"5d",
          3529 => x"08",
          3530 => x"92",
          3531 => x"e4",
          3532 => x"3d",
          3533 => x"51",
          3534 => x"82",
          3535 => x"60",
          3536 => x"5c",
          3537 => x"81",
          3538 => x"d5",
          3539 => x"cd",
          3540 => x"d5",
          3541 => x"26",
          3542 => x"81",
          3543 => x"2e",
          3544 => x"82",
          3545 => x"7a",
          3546 => x"38",
          3547 => x"7a",
          3548 => x"38",
          3549 => x"82",
          3550 => x"7b",
          3551 => x"b8",
          3552 => x"82",
          3553 => x"b5",
          3554 => x"05",
          3555 => x"b1",
          3556 => x"7b",
          3557 => x"ff",
          3558 => x"cd",
          3559 => x"39",
          3560 => x"bc",
          3561 => x"53",
          3562 => x"52",
          3563 => x"b0",
          3564 => x"a7",
          3565 => x"39",
          3566 => x"53",
          3567 => x"52",
          3568 => x"b0",
          3569 => x"a6",
          3570 => x"d4",
          3571 => x"d6",
          3572 => x"56",
          3573 => x"54",
          3574 => x"53",
          3575 => x"52",
          3576 => x"b0",
          3577 => x"f5",
          3578 => x"e4",
          3579 => x"e4",
          3580 => x"30",
          3581 => x"80",
          3582 => x"5b",
          3583 => x"7a",
          3584 => x"38",
          3585 => x"7a",
          3586 => x"80",
          3587 => x"81",
          3588 => x"ff",
          3589 => x"7a",
          3590 => x"7f",
          3591 => x"81",
          3592 => x"78",
          3593 => x"ff",
          3594 => x"06",
          3595 => x"bc",
          3596 => x"bf",
          3597 => x"51",
          3598 => x"f2",
          3599 => x"bc",
          3600 => x"bf",
          3601 => x"a0",
          3602 => x"0d",
          3603 => x"d6",
          3604 => x"c0",
          3605 => x"08",
          3606 => x"84",
          3607 => x"51",
          3608 => x"82",
          3609 => x"90",
          3610 => x"55",
          3611 => x"80",
          3612 => x"d7",
          3613 => x"82",
          3614 => x"07",
          3615 => x"c0",
          3616 => x"08",
          3617 => x"84",
          3618 => x"51",
          3619 => x"82",
          3620 => x"90",
          3621 => x"55",
          3622 => x"80",
          3623 => x"d7",
          3624 => x"82",
          3625 => x"07",
          3626 => x"80",
          3627 => x"c0",
          3628 => x"8c",
          3629 => x"87",
          3630 => x"0c",
          3631 => x"5a",
          3632 => x"5b",
          3633 => x"05",
          3634 => x"80",
          3635 => x"c4",
          3636 => x"70",
          3637 => x"70",
          3638 => x"f1",
          3639 => x"89",
          3640 => x"ff",
          3641 => x"9c",
          3642 => x"f8",
          3643 => x"a8",
          3644 => x"f0",
          3645 => x"d8",
          3646 => x"3f",
          3647 => x"9c",
          3648 => x"3f",
          3649 => x"3d",
          3650 => x"83",
          3651 => x"2b",
          3652 => x"3f",
          3653 => x"08",
          3654 => x"72",
          3655 => x"54",
          3656 => x"25",
          3657 => x"82",
          3658 => x"84",
          3659 => x"fc",
          3660 => x"70",
          3661 => x"80",
          3662 => x"72",
          3663 => x"8a",
          3664 => x"51",
          3665 => x"09",
          3666 => x"38",
          3667 => x"f1",
          3668 => x"51",
          3669 => x"09",
          3670 => x"38",
          3671 => x"81",
          3672 => x"73",
          3673 => x"81",
          3674 => x"84",
          3675 => x"52",
          3676 => x"52",
          3677 => x"2e",
          3678 => x"54",
          3679 => x"9d",
          3680 => x"38",
          3681 => x"12",
          3682 => x"33",
          3683 => x"a0",
          3684 => x"81",
          3685 => x"2e",
          3686 => x"ea",
          3687 => x"33",
          3688 => x"a0",
          3689 => x"06",
          3690 => x"54",
          3691 => x"70",
          3692 => x"25",
          3693 => x"51",
          3694 => x"2e",
          3695 => x"72",
          3696 => x"54",
          3697 => x"0c",
          3698 => x"82",
          3699 => x"86",
          3700 => x"fc",
          3701 => x"53",
          3702 => x"2e",
          3703 => x"3d",
          3704 => x"72",
          3705 => x"3f",
          3706 => x"08",
          3707 => x"53",
          3708 => x"53",
          3709 => x"e4",
          3710 => x"0d",
          3711 => x"0d",
          3712 => x"33",
          3713 => x"53",
          3714 => x"8b",
          3715 => x"38",
          3716 => x"ff",
          3717 => x"52",
          3718 => x"81",
          3719 => x"13",
          3720 => x"52",
          3721 => x"80",
          3722 => x"13",
          3723 => x"52",
          3724 => x"80",
          3725 => x"13",
          3726 => x"52",
          3727 => x"80",
          3728 => x"13",
          3729 => x"52",
          3730 => x"26",
          3731 => x"8a",
          3732 => x"87",
          3733 => x"e7",
          3734 => x"38",
          3735 => x"c0",
          3736 => x"72",
          3737 => x"98",
          3738 => x"13",
          3739 => x"98",
          3740 => x"13",
          3741 => x"98",
          3742 => x"13",
          3743 => x"98",
          3744 => x"13",
          3745 => x"98",
          3746 => x"13",
          3747 => x"98",
          3748 => x"87",
          3749 => x"0c",
          3750 => x"98",
          3751 => x"0b",
          3752 => x"9c",
          3753 => x"71",
          3754 => x"0c",
          3755 => x"04",
          3756 => x"7f",
          3757 => x"98",
          3758 => x"7d",
          3759 => x"98",
          3760 => x"7d",
          3761 => x"c0",
          3762 => x"5a",
          3763 => x"34",
          3764 => x"b4",
          3765 => x"83",
          3766 => x"c0",
          3767 => x"5a",
          3768 => x"34",
          3769 => x"ac",
          3770 => x"85",
          3771 => x"c0",
          3772 => x"5a",
          3773 => x"34",
          3774 => x"a4",
          3775 => x"88",
          3776 => x"c0",
          3777 => x"5a",
          3778 => x"23",
          3779 => x"79",
          3780 => x"06",
          3781 => x"ff",
          3782 => x"86",
          3783 => x"85",
          3784 => x"84",
          3785 => x"83",
          3786 => x"82",
          3787 => x"7d",
          3788 => x"06",
          3789 => x"c0",
          3790 => x"9d",
          3791 => x"0d",
          3792 => x"0d",
          3793 => x"33",
          3794 => x"33",
          3795 => x"06",
          3796 => x"87",
          3797 => x"51",
          3798 => x"86",
          3799 => x"94",
          3800 => x"08",
          3801 => x"70",
          3802 => x"54",
          3803 => x"2e",
          3804 => x"91",
          3805 => x"06",
          3806 => x"d7",
          3807 => x"32",
          3808 => x"51",
          3809 => x"2e",
          3810 => x"93",
          3811 => x"06",
          3812 => x"ff",
          3813 => x"81",
          3814 => x"87",
          3815 => x"52",
          3816 => x"86",
          3817 => x"94",
          3818 => x"72",
          3819 => x"d5",
          3820 => x"3d",
          3821 => x"3d",
          3822 => x"05",
          3823 => x"70",
          3824 => x"52",
          3825 => x"d3",
          3826 => x"3d",
          3827 => x"3d",
          3828 => x"05",
          3829 => x"8a",
          3830 => x"06",
          3831 => x"52",
          3832 => x"3f",
          3833 => x"33",
          3834 => x"06",
          3835 => x"c0",
          3836 => x"76",
          3837 => x"38",
          3838 => x"94",
          3839 => x"70",
          3840 => x"81",
          3841 => x"54",
          3842 => x"8c",
          3843 => x"2a",
          3844 => x"51",
          3845 => x"38",
          3846 => x"70",
          3847 => x"53",
          3848 => x"8d",
          3849 => x"2a",
          3850 => x"51",
          3851 => x"be",
          3852 => x"ff",
          3853 => x"c0",
          3854 => x"72",
          3855 => x"38",
          3856 => x"90",
          3857 => x"0c",
          3858 => x"d5",
          3859 => x"3d",
          3860 => x"3d",
          3861 => x"80",
          3862 => x"81",
          3863 => x"53",
          3864 => x"2e",
          3865 => x"71",
          3866 => x"81",
          3867 => x"fc",
          3868 => x"ff",
          3869 => x"55",
          3870 => x"94",
          3871 => x"80",
          3872 => x"87",
          3873 => x"51",
          3874 => x"96",
          3875 => x"06",
          3876 => x"70",
          3877 => x"38",
          3878 => x"70",
          3879 => x"51",
          3880 => x"72",
          3881 => x"81",
          3882 => x"70",
          3883 => x"38",
          3884 => x"70",
          3885 => x"51",
          3886 => x"38",
          3887 => x"06",
          3888 => x"94",
          3889 => x"80",
          3890 => x"87",
          3891 => x"52",
          3892 => x"81",
          3893 => x"70",
          3894 => x"53",
          3895 => x"ff",
          3896 => x"82",
          3897 => x"89",
          3898 => x"fe",
          3899 => x"d3",
          3900 => x"81",
          3901 => x"52",
          3902 => x"84",
          3903 => x"2e",
          3904 => x"c0",
          3905 => x"70",
          3906 => x"2a",
          3907 => x"51",
          3908 => x"80",
          3909 => x"71",
          3910 => x"51",
          3911 => x"80",
          3912 => x"2e",
          3913 => x"c0",
          3914 => x"71",
          3915 => x"ff",
          3916 => x"e4",
          3917 => x"3d",
          3918 => x"af",
          3919 => x"e4",
          3920 => x"06",
          3921 => x"0c",
          3922 => x"0d",
          3923 => x"33",
          3924 => x"06",
          3925 => x"c0",
          3926 => x"70",
          3927 => x"38",
          3928 => x"94",
          3929 => x"70",
          3930 => x"81",
          3931 => x"51",
          3932 => x"80",
          3933 => x"72",
          3934 => x"51",
          3935 => x"80",
          3936 => x"2e",
          3937 => x"c0",
          3938 => x"71",
          3939 => x"2b",
          3940 => x"51",
          3941 => x"82",
          3942 => x"84",
          3943 => x"ff",
          3944 => x"c0",
          3945 => x"70",
          3946 => x"06",
          3947 => x"80",
          3948 => x"38",
          3949 => x"a4",
          3950 => x"80",
          3951 => x"9e",
          3952 => x"d4",
          3953 => x"c0",
          3954 => x"82",
          3955 => x"87",
          3956 => x"08",
          3957 => x"0c",
          3958 => x"9c",
          3959 => x"90",
          3960 => x"9e",
          3961 => x"d4",
          3962 => x"c0",
          3963 => x"82",
          3964 => x"87",
          3965 => x"08",
          3966 => x"0c",
          3967 => x"b4",
          3968 => x"a0",
          3969 => x"9e",
          3970 => x"d4",
          3971 => x"c0",
          3972 => x"82",
          3973 => x"87",
          3974 => x"08",
          3975 => x"0c",
          3976 => x"c4",
          3977 => x"b0",
          3978 => x"9e",
          3979 => x"70",
          3980 => x"23",
          3981 => x"84",
          3982 => x"b8",
          3983 => x"9e",
          3984 => x"d4",
          3985 => x"c0",
          3986 => x"82",
          3987 => x"81",
          3988 => x"c4",
          3989 => x"87",
          3990 => x"08",
          3991 => x"0a",
          3992 => x"52",
          3993 => x"83",
          3994 => x"71",
          3995 => x"34",
          3996 => x"c0",
          3997 => x"70",
          3998 => x"06",
          3999 => x"70",
          4000 => x"38",
          4001 => x"82",
          4002 => x"80",
          4003 => x"9e",
          4004 => x"90",
          4005 => x"51",
          4006 => x"80",
          4007 => x"81",
          4008 => x"d4",
          4009 => x"0b",
          4010 => x"90",
          4011 => x"80",
          4012 => x"52",
          4013 => x"2e",
          4014 => x"52",
          4015 => x"c8",
          4016 => x"87",
          4017 => x"08",
          4018 => x"80",
          4019 => x"52",
          4020 => x"83",
          4021 => x"71",
          4022 => x"34",
          4023 => x"c0",
          4024 => x"70",
          4025 => x"06",
          4026 => x"70",
          4027 => x"38",
          4028 => x"82",
          4029 => x"80",
          4030 => x"9e",
          4031 => x"84",
          4032 => x"51",
          4033 => x"80",
          4034 => x"81",
          4035 => x"d4",
          4036 => x"0b",
          4037 => x"90",
          4038 => x"80",
          4039 => x"52",
          4040 => x"2e",
          4041 => x"52",
          4042 => x"cc",
          4043 => x"87",
          4044 => x"08",
          4045 => x"80",
          4046 => x"52",
          4047 => x"83",
          4048 => x"71",
          4049 => x"34",
          4050 => x"c0",
          4051 => x"70",
          4052 => x"06",
          4053 => x"70",
          4054 => x"38",
          4055 => x"82",
          4056 => x"80",
          4057 => x"9e",
          4058 => x"a0",
          4059 => x"52",
          4060 => x"2e",
          4061 => x"52",
          4062 => x"cf",
          4063 => x"9e",
          4064 => x"98",
          4065 => x"8a",
          4066 => x"51",
          4067 => x"d0",
          4068 => x"87",
          4069 => x"08",
          4070 => x"06",
          4071 => x"70",
          4072 => x"38",
          4073 => x"82",
          4074 => x"87",
          4075 => x"08",
          4076 => x"06",
          4077 => x"51",
          4078 => x"82",
          4079 => x"80",
          4080 => x"9e",
          4081 => x"88",
          4082 => x"52",
          4083 => x"83",
          4084 => x"71",
          4085 => x"34",
          4086 => x"90",
          4087 => x"06",
          4088 => x"82",
          4089 => x"83",
          4090 => x"fb",
          4091 => x"bd",
          4092 => x"93",
          4093 => x"d4",
          4094 => x"73",
          4095 => x"38",
          4096 => x"51",
          4097 => x"3f",
          4098 => x"51",
          4099 => x"3f",
          4100 => x"33",
          4101 => x"2e",
          4102 => x"d4",
          4103 => x"d4",
          4104 => x"54",
          4105 => x"98",
          4106 => x"ad",
          4107 => x"cb",
          4108 => x"80",
          4109 => x"82",
          4110 => x"82",
          4111 => x"11",
          4112 => x"be",
          4113 => x"93",
          4114 => x"d4",
          4115 => x"73",
          4116 => x"38",
          4117 => x"08",
          4118 => x"08",
          4119 => x"82",
          4120 => x"ff",
          4121 => x"82",
          4122 => x"54",
          4123 => x"94",
          4124 => x"88",
          4125 => x"8c",
          4126 => x"52",
          4127 => x"51",
          4128 => x"3f",
          4129 => x"33",
          4130 => x"2e",
          4131 => x"d4",
          4132 => x"d4",
          4133 => x"54",
          4134 => x"88",
          4135 => x"b9",
          4136 => x"cf",
          4137 => x"80",
          4138 => x"82",
          4139 => x"52",
          4140 => x"51",
          4141 => x"3f",
          4142 => x"33",
          4143 => x"2e",
          4144 => x"d4",
          4145 => x"82",
          4146 => x"ff",
          4147 => x"82",
          4148 => x"54",
          4149 => x"8e",
          4150 => x"d2",
          4151 => x"bf",
          4152 => x"91",
          4153 => x"d4",
          4154 => x"73",
          4155 => x"38",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"33",
          4159 => x"2e",
          4160 => x"c0",
          4161 => x"ad",
          4162 => x"d4",
          4163 => x"73",
          4164 => x"38",
          4165 => x"51",
          4166 => x"3f",
          4167 => x"33",
          4168 => x"2e",
          4169 => x"c0",
          4170 => x"ad",
          4171 => x"d4",
          4172 => x"73",
          4173 => x"38",
          4174 => x"51",
          4175 => x"3f",
          4176 => x"51",
          4177 => x"3f",
          4178 => x"08",
          4179 => x"cc",
          4180 => x"85",
          4181 => x"ac",
          4182 => x"c0",
          4183 => x"90",
          4184 => x"d4",
          4185 => x"82",
          4186 => x"ff",
          4187 => x"82",
          4188 => x"ff",
          4189 => x"82",
          4190 => x"52",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"08",
          4194 => x"c0",
          4195 => x"c5",
          4196 => x"d5",
          4197 => x"84",
          4198 => x"71",
          4199 => x"82",
          4200 => x"52",
          4201 => x"51",
          4202 => x"3f",
          4203 => x"33",
          4204 => x"2e",
          4205 => x"d4",
          4206 => x"bd",
          4207 => x"75",
          4208 => x"3f",
          4209 => x"08",
          4210 => x"29",
          4211 => x"54",
          4212 => x"e4",
          4213 => x"c2",
          4214 => x"8f",
          4215 => x"d4",
          4216 => x"73",
          4217 => x"38",
          4218 => x"08",
          4219 => x"c0",
          4220 => x"c4",
          4221 => x"d5",
          4222 => x"84",
          4223 => x"71",
          4224 => x"82",
          4225 => x"52",
          4226 => x"51",
          4227 => x"3f",
          4228 => x"ae",
          4229 => x"3d",
          4230 => x"3d",
          4231 => x"05",
          4232 => x"52",
          4233 => x"aa",
          4234 => x"29",
          4235 => x"05",
          4236 => x"04",
          4237 => x"51",
          4238 => x"c3",
          4239 => x"39",
          4240 => x"51",
          4241 => x"c3",
          4242 => x"39",
          4243 => x"51",
          4244 => x"c3",
          4245 => x"8f",
          4246 => x"3d",
          4247 => x"88",
          4248 => x"80",
          4249 => x"96",
          4250 => x"82",
          4251 => x"87",
          4252 => x"0c",
          4253 => x"0d",
          4254 => x"70",
          4255 => x"98",
          4256 => x"2c",
          4257 => x"70",
          4258 => x"53",
          4259 => x"51",
          4260 => x"c3",
          4261 => x"55",
          4262 => x"25",
          4263 => x"c3",
          4264 => x"12",
          4265 => x"97",
          4266 => x"33",
          4267 => x"70",
          4268 => x"81",
          4269 => x"81",
          4270 => x"d5",
          4271 => x"3d",
          4272 => x"3d",
          4273 => x"84",
          4274 => x"33",
          4275 => x"56",
          4276 => x"2e",
          4277 => x"f1",
          4278 => x"88",
          4279 => x"d3",
          4280 => x"c8",
          4281 => x"51",
          4282 => x"3f",
          4283 => x"08",
          4284 => x"ff",
          4285 => x"73",
          4286 => x"53",
          4287 => x"72",
          4288 => x"53",
          4289 => x"51",
          4290 => x"3f",
          4291 => x"87",
          4292 => x"f6",
          4293 => x"02",
          4294 => x"05",
          4295 => x"05",
          4296 => x"82",
          4297 => x"70",
          4298 => x"d4",
          4299 => x"08",
          4300 => x"5a",
          4301 => x"80",
          4302 => x"74",
          4303 => x"3f",
          4304 => x"33",
          4305 => x"82",
          4306 => x"81",
          4307 => x"58",
          4308 => x"fc",
          4309 => x"e4",
          4310 => x"82",
          4311 => x"70",
          4312 => x"d4",
          4313 => x"08",
          4314 => x"74",
          4315 => x"38",
          4316 => x"52",
          4317 => x"b6",
          4318 => x"d5",
          4319 => x"05",
          4320 => x"d5",
          4321 => x"81",
          4322 => x"93",
          4323 => x"38",
          4324 => x"d5",
          4325 => x"80",
          4326 => x"82",
          4327 => x"56",
          4328 => x"ac",
          4329 => x"ac",
          4330 => x"a4",
          4331 => x"fc",
          4332 => x"53",
          4333 => x"51",
          4334 => x"3f",
          4335 => x"08",
          4336 => x"81",
          4337 => x"82",
          4338 => x"51",
          4339 => x"3f",
          4340 => x"04",
          4341 => x"82",
          4342 => x"93",
          4343 => x"52",
          4344 => x"89",
          4345 => x"99",
          4346 => x"73",
          4347 => x"84",
          4348 => x"73",
          4349 => x"38",
          4350 => x"d5",
          4351 => x"d5",
          4352 => x"71",
          4353 => x"38",
          4354 => x"f0",
          4355 => x"d5",
          4356 => x"99",
          4357 => x"0b",
          4358 => x"0c",
          4359 => x"04",
          4360 => x"81",
          4361 => x"82",
          4362 => x"51",
          4363 => x"3f",
          4364 => x"08",
          4365 => x"82",
          4366 => x"53",
          4367 => x"88",
          4368 => x"56",
          4369 => x"3f",
          4370 => x"08",
          4371 => x"38",
          4372 => x"b3",
          4373 => x"d5",
          4374 => x"80",
          4375 => x"e4",
          4376 => x"38",
          4377 => x"08",
          4378 => x"17",
          4379 => x"74",
          4380 => x"76",
          4381 => x"82",
          4382 => x"57",
          4383 => x"3f",
          4384 => x"09",
          4385 => x"af",
          4386 => x"0d",
          4387 => x"0d",
          4388 => x"ad",
          4389 => x"5a",
          4390 => x"58",
          4391 => x"d5",
          4392 => x"80",
          4393 => x"82",
          4394 => x"81",
          4395 => x"0b",
          4396 => x"08",
          4397 => x"f8",
          4398 => x"70",
          4399 => x"9e",
          4400 => x"d5",
          4401 => x"2e",
          4402 => x"51",
          4403 => x"3f",
          4404 => x"08",
          4405 => x"55",
          4406 => x"d5",
          4407 => x"8e",
          4408 => x"e4",
          4409 => x"70",
          4410 => x"80",
          4411 => x"09",
          4412 => x"72",
          4413 => x"51",
          4414 => x"77",
          4415 => x"73",
          4416 => x"82",
          4417 => x"8c",
          4418 => x"51",
          4419 => x"3f",
          4420 => x"08",
          4421 => x"38",
          4422 => x"51",
          4423 => x"3f",
          4424 => x"09",
          4425 => x"38",
          4426 => x"51",
          4427 => x"3f",
          4428 => x"b1",
          4429 => x"3d",
          4430 => x"d5",
          4431 => x"34",
          4432 => x"82",
          4433 => x"a9",
          4434 => x"f6",
          4435 => x"7e",
          4436 => x"72",
          4437 => x"5a",
          4438 => x"2e",
          4439 => x"a2",
          4440 => x"78",
          4441 => x"76",
          4442 => x"81",
          4443 => x"70",
          4444 => x"58",
          4445 => x"2e",
          4446 => x"86",
          4447 => x"26",
          4448 => x"54",
          4449 => x"82",
          4450 => x"70",
          4451 => x"ff",
          4452 => x"82",
          4453 => x"53",
          4454 => x"08",
          4455 => x"f3",
          4456 => x"e4",
          4457 => x"38",
          4458 => x"55",
          4459 => x"88",
          4460 => x"2e",
          4461 => x"39",
          4462 => x"ac",
          4463 => x"5a",
          4464 => x"11",
          4465 => x"51",
          4466 => x"82",
          4467 => x"80",
          4468 => x"ff",
          4469 => x"52",
          4470 => x"b1",
          4471 => x"e4",
          4472 => x"06",
          4473 => x"38",
          4474 => x"39",
          4475 => x"81",
          4476 => x"54",
          4477 => x"ff",
          4478 => x"54",
          4479 => x"e4",
          4480 => x"0d",
          4481 => x"0d",
          4482 => x"b2",
          4483 => x"3d",
          4484 => x"5a",
          4485 => x"3d",
          4486 => x"b4",
          4487 => x"b0",
          4488 => x"73",
          4489 => x"73",
          4490 => x"33",
          4491 => x"83",
          4492 => x"76",
          4493 => x"bc",
          4494 => x"76",
          4495 => x"73",
          4496 => x"ad",
          4497 => x"98",
          4498 => x"d5",
          4499 => x"d5",
          4500 => x"d5",
          4501 => x"2e",
          4502 => x"93",
          4503 => x"82",
          4504 => x"51",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"38",
          4508 => x"51",
          4509 => x"3f",
          4510 => x"82",
          4511 => x"5b",
          4512 => x"08",
          4513 => x"52",
          4514 => x"52",
          4515 => x"f6",
          4516 => x"e4",
          4517 => x"d5",
          4518 => x"2e",
          4519 => x"80",
          4520 => x"d5",
          4521 => x"ff",
          4522 => x"82",
          4523 => x"55",
          4524 => x"d5",
          4525 => x"a9",
          4526 => x"e4",
          4527 => x"70",
          4528 => x"80",
          4529 => x"53",
          4530 => x"06",
          4531 => x"f8",
          4532 => x"1b",
          4533 => x"06",
          4534 => x"7b",
          4535 => x"80",
          4536 => x"2e",
          4537 => x"ff",
          4538 => x"39",
          4539 => x"ac",
          4540 => x"38",
          4541 => x"08",
          4542 => x"38",
          4543 => x"8f",
          4544 => x"c5",
          4545 => x"e4",
          4546 => x"70",
          4547 => x"59",
          4548 => x"ee",
          4549 => x"ff",
          4550 => x"a0",
          4551 => x"2b",
          4552 => x"82",
          4553 => x"70",
          4554 => x"97",
          4555 => x"2c",
          4556 => x"29",
          4557 => x"05",
          4558 => x"70",
          4559 => x"51",
          4560 => x"51",
          4561 => x"81",
          4562 => x"2e",
          4563 => x"77",
          4564 => x"38",
          4565 => x"0a",
          4566 => x"0a",
          4567 => x"2c",
          4568 => x"75",
          4569 => x"38",
          4570 => x"52",
          4571 => x"85",
          4572 => x"e4",
          4573 => x"06",
          4574 => x"2e",
          4575 => x"82",
          4576 => x"81",
          4577 => x"74",
          4578 => x"29",
          4579 => x"05",
          4580 => x"70",
          4581 => x"56",
          4582 => x"95",
          4583 => x"76",
          4584 => x"77",
          4585 => x"3f",
          4586 => x"08",
          4587 => x"54",
          4588 => x"d3",
          4589 => x"75",
          4590 => x"ca",
          4591 => x"55",
          4592 => x"a0",
          4593 => x"2b",
          4594 => x"82",
          4595 => x"70",
          4596 => x"98",
          4597 => x"11",
          4598 => x"82",
          4599 => x"33",
          4600 => x"51",
          4601 => x"55",
          4602 => x"09",
          4603 => x"92",
          4604 => x"ac",
          4605 => x"0c",
          4606 => x"ed",
          4607 => x"0b",
          4608 => x"34",
          4609 => x"82",
          4610 => x"75",
          4611 => x"34",
          4612 => x"34",
          4613 => x"7e",
          4614 => x"26",
          4615 => x"73",
          4616 => x"ae",
          4617 => x"73",
          4618 => x"ed",
          4619 => x"73",
          4620 => x"cb",
          4621 => x"a4",
          4622 => x"75",
          4623 => x"74",
          4624 => x"98",
          4625 => x"73",
          4626 => x"38",
          4627 => x"73",
          4628 => x"34",
          4629 => x"0a",
          4630 => x"0a",
          4631 => x"2c",
          4632 => x"33",
          4633 => x"df",
          4634 => x"a8",
          4635 => x"56",
          4636 => x"ed",
          4637 => x"1a",
          4638 => x"33",
          4639 => x"ed",
          4640 => x"73",
          4641 => x"38",
          4642 => x"73",
          4643 => x"34",
          4644 => x"33",
          4645 => x"0a",
          4646 => x"0a",
          4647 => x"2c",
          4648 => x"33",
          4649 => x"56",
          4650 => x"a8",
          4651 => x"c8",
          4652 => x"1a",
          4653 => x"54",
          4654 => x"3f",
          4655 => x"0a",
          4656 => x"0a",
          4657 => x"2c",
          4658 => x"33",
          4659 => x"73",
          4660 => x"38",
          4661 => x"33",
          4662 => x"70",
          4663 => x"ed",
          4664 => x"51",
          4665 => x"77",
          4666 => x"38",
          4667 => x"08",
          4668 => x"ff",
          4669 => x"74",
          4670 => x"29",
          4671 => x"05",
          4672 => x"82",
          4673 => x"56",
          4674 => x"75",
          4675 => x"fb",
          4676 => x"7a",
          4677 => x"81",
          4678 => x"ed",
          4679 => x"52",
          4680 => x"51",
          4681 => x"81",
          4682 => x"ed",
          4683 => x"81",
          4684 => x"55",
          4685 => x"fb",
          4686 => x"ed",
          4687 => x"05",
          4688 => x"ed",
          4689 => x"15",
          4690 => x"ed",
          4691 => x"f1",
          4692 => x"88",
          4693 => x"db",
          4694 => x"a8",
          4695 => x"2b",
          4696 => x"82",
          4697 => x"57",
          4698 => x"74",
          4699 => x"38",
          4700 => x"81",
          4701 => x"34",
          4702 => x"08",
          4703 => x"51",
          4704 => x"3f",
          4705 => x"0a",
          4706 => x"0a",
          4707 => x"2c",
          4708 => x"33",
          4709 => x"75",
          4710 => x"38",
          4711 => x"08",
          4712 => x"ff",
          4713 => x"82",
          4714 => x"70",
          4715 => x"98",
          4716 => x"a4",
          4717 => x"56",
          4718 => x"24",
          4719 => x"82",
          4720 => x"52",
          4721 => x"9f",
          4722 => x"81",
          4723 => x"81",
          4724 => x"70",
          4725 => x"ed",
          4726 => x"51",
          4727 => x"25",
          4728 => x"9b",
          4729 => x"a4",
          4730 => x"54",
          4731 => x"82",
          4732 => x"52",
          4733 => x"9f",
          4734 => x"ed",
          4735 => x"51",
          4736 => x"82",
          4737 => x"81",
          4738 => x"73",
          4739 => x"ed",
          4740 => x"73",
          4741 => x"38",
          4742 => x"52",
          4743 => x"f3",
          4744 => x"80",
          4745 => x"0b",
          4746 => x"34",
          4747 => x"ed",
          4748 => x"82",
          4749 => x"af",
          4750 => x"82",
          4751 => x"54",
          4752 => x"f9",
          4753 => x"f1",
          4754 => x"88",
          4755 => x"e3",
          4756 => x"a8",
          4757 => x"54",
          4758 => x"a8",
          4759 => x"ff",
          4760 => x"39",
          4761 => x"33",
          4762 => x"33",
          4763 => x"75",
          4764 => x"38",
          4765 => x"73",
          4766 => x"34",
          4767 => x"70",
          4768 => x"81",
          4769 => x"51",
          4770 => x"25",
          4771 => x"1a",
          4772 => x"33",
          4773 => x"f1",
          4774 => x"73",
          4775 => x"9e",
          4776 => x"81",
          4777 => x"81",
          4778 => x"70",
          4779 => x"ed",
          4780 => x"51",
          4781 => x"24",
          4782 => x"f1",
          4783 => x"a0",
          4784 => x"ef",
          4785 => x"a8",
          4786 => x"2b",
          4787 => x"82",
          4788 => x"57",
          4789 => x"74",
          4790 => x"a3",
          4791 => x"c8",
          4792 => x"51",
          4793 => x"3f",
          4794 => x"0a",
          4795 => x"0a",
          4796 => x"2c",
          4797 => x"33",
          4798 => x"75",
          4799 => x"38",
          4800 => x"82",
          4801 => x"70",
          4802 => x"82",
          4803 => x"59",
          4804 => x"77",
          4805 => x"38",
          4806 => x"08",
          4807 => x"54",
          4808 => x"a8",
          4809 => x"70",
          4810 => x"ff",
          4811 => x"82",
          4812 => x"70",
          4813 => x"82",
          4814 => x"58",
          4815 => x"75",
          4816 => x"f7",
          4817 => x"ed",
          4818 => x"52",
          4819 => x"51",
          4820 => x"80",
          4821 => x"a8",
          4822 => x"82",
          4823 => x"f7",
          4824 => x"b0",
          4825 => x"a8",
          4826 => x"80",
          4827 => x"74",
          4828 => x"92",
          4829 => x"e4",
          4830 => x"a4",
          4831 => x"e4",
          4832 => x"06",
          4833 => x"74",
          4834 => x"ff",
          4835 => x"93",
          4836 => x"39",
          4837 => x"82",
          4838 => x"fc",
          4839 => x"54",
          4840 => x"a7",
          4841 => x"ff",
          4842 => x"82",
          4843 => x"82",
          4844 => x"82",
          4845 => x"81",
          4846 => x"05",
          4847 => x"79",
          4848 => x"a2",
          4849 => x"54",
          4850 => x"73",
          4851 => x"80",
          4852 => x"38",
          4853 => x"a4",
          4854 => x"39",
          4855 => x"09",
          4856 => x"38",
          4857 => x"08",
          4858 => x"2e",
          4859 => x"51",
          4860 => x"3f",
          4861 => x"08",
          4862 => x"34",
          4863 => x"08",
          4864 => x"81",
          4865 => x"52",
          4866 => x"a5",
          4867 => x"c3",
          4868 => x"29",
          4869 => x"05",
          4870 => x"54",
          4871 => x"ab",
          4872 => x"ff",
          4873 => x"82",
          4874 => x"82",
          4875 => x"82",
          4876 => x"81",
          4877 => x"05",
          4878 => x"79",
          4879 => x"a6",
          4880 => x"54",
          4881 => x"06",
          4882 => x"74",
          4883 => x"34",
          4884 => x"82",
          4885 => x"82",
          4886 => x"52",
          4887 => x"e2",
          4888 => x"39",
          4889 => x"33",
          4890 => x"06",
          4891 => x"33",
          4892 => x"74",
          4893 => x"87",
          4894 => x"c8",
          4895 => x"14",
          4896 => x"ed",
          4897 => x"1a",
          4898 => x"54",
          4899 => x"3f",
          4900 => x"82",
          4901 => x"54",
          4902 => x"f4",
          4903 => x"f1",
          4904 => x"88",
          4905 => x"8b",
          4906 => x"a8",
          4907 => x"54",
          4908 => x"a8",
          4909 => x"39",
          4910 => x"84",
          4911 => x"82",
          4912 => x"a0",
          4913 => x"d5",
          4914 => x"80",
          4915 => x"52",
          4916 => x"51",
          4917 => x"3f",
          4918 => x"08",
          4919 => x"77",
          4920 => x"57",
          4921 => x"34",
          4922 => x"08",
          4923 => x"15",
          4924 => x"15",
          4925 => x"d4",
          4926 => x"86",
          4927 => x"87",
          4928 => x"d5",
          4929 => x"d5",
          4930 => x"05",
          4931 => x"07",
          4932 => x"ff",
          4933 => x"2a",
          4934 => x"56",
          4935 => x"34",
          4936 => x"34",
          4937 => x"22",
          4938 => x"82",
          4939 => x"05",
          4940 => x"55",
          4941 => x"15",
          4942 => x"15",
          4943 => x"0d",
          4944 => x"0d",
          4945 => x"51",
          4946 => x"8f",
          4947 => x"83",
          4948 => x"70",
          4949 => x"06",
          4950 => x"70",
          4951 => x"0c",
          4952 => x"04",
          4953 => x"02",
          4954 => x"02",
          4955 => x"05",
          4956 => x"82",
          4957 => x"71",
          4958 => x"11",
          4959 => x"73",
          4960 => x"81",
          4961 => x"88",
          4962 => x"a4",
          4963 => x"22",
          4964 => x"ff",
          4965 => x"88",
          4966 => x"52",
          4967 => x"5b",
          4968 => x"55",
          4969 => x"70",
          4970 => x"82",
          4971 => x"14",
          4972 => x"52",
          4973 => x"15",
          4974 => x"15",
          4975 => x"d4",
          4976 => x"70",
          4977 => x"33",
          4978 => x"07",
          4979 => x"8f",
          4980 => x"51",
          4981 => x"71",
          4982 => x"ff",
          4983 => x"88",
          4984 => x"51",
          4985 => x"34",
          4986 => x"06",
          4987 => x"12",
          4988 => x"d4",
          4989 => x"71",
          4990 => x"81",
          4991 => x"3d",
          4992 => x"3d",
          4993 => x"d4",
          4994 => x"05",
          4995 => x"70",
          4996 => x"11",
          4997 => x"87",
          4998 => x"8b",
          4999 => x"2b",
          5000 => x"59",
          5001 => x"72",
          5002 => x"33",
          5003 => x"71",
          5004 => x"70",
          5005 => x"56",
          5006 => x"84",
          5007 => x"85",
          5008 => x"d5",
          5009 => x"14",
          5010 => x"85",
          5011 => x"8b",
          5012 => x"2b",
          5013 => x"57",
          5014 => x"86",
          5015 => x"13",
          5016 => x"2b",
          5017 => x"2a",
          5018 => x"52",
          5019 => x"34",
          5020 => x"34",
          5021 => x"08",
          5022 => x"81",
          5023 => x"88",
          5024 => x"81",
          5025 => x"70",
          5026 => x"51",
          5027 => x"71",
          5028 => x"81",
          5029 => x"3d",
          5030 => x"3d",
          5031 => x"05",
          5032 => x"d4",
          5033 => x"2b",
          5034 => x"33",
          5035 => x"71",
          5036 => x"70",
          5037 => x"70",
          5038 => x"33",
          5039 => x"71",
          5040 => x"53",
          5041 => x"52",
          5042 => x"53",
          5043 => x"25",
          5044 => x"72",
          5045 => x"3f",
          5046 => x"08",
          5047 => x"33",
          5048 => x"71",
          5049 => x"83",
          5050 => x"11",
          5051 => x"12",
          5052 => x"2b",
          5053 => x"2b",
          5054 => x"06",
          5055 => x"51",
          5056 => x"53",
          5057 => x"88",
          5058 => x"72",
          5059 => x"73",
          5060 => x"82",
          5061 => x"70",
          5062 => x"81",
          5063 => x"8b",
          5064 => x"2b",
          5065 => x"57",
          5066 => x"70",
          5067 => x"33",
          5068 => x"07",
          5069 => x"ff",
          5070 => x"2a",
          5071 => x"58",
          5072 => x"34",
          5073 => x"34",
          5074 => x"04",
          5075 => x"82",
          5076 => x"02",
          5077 => x"05",
          5078 => x"2b",
          5079 => x"11",
          5080 => x"33",
          5081 => x"71",
          5082 => x"59",
          5083 => x"56",
          5084 => x"71",
          5085 => x"33",
          5086 => x"07",
          5087 => x"a2",
          5088 => x"07",
          5089 => x"53",
          5090 => x"53",
          5091 => x"70",
          5092 => x"82",
          5093 => x"70",
          5094 => x"81",
          5095 => x"8b",
          5096 => x"2b",
          5097 => x"57",
          5098 => x"82",
          5099 => x"13",
          5100 => x"2b",
          5101 => x"2a",
          5102 => x"52",
          5103 => x"34",
          5104 => x"34",
          5105 => x"08",
          5106 => x"33",
          5107 => x"71",
          5108 => x"82",
          5109 => x"52",
          5110 => x"0d",
          5111 => x"0d",
          5112 => x"d4",
          5113 => x"2a",
          5114 => x"ff",
          5115 => x"57",
          5116 => x"3f",
          5117 => x"08",
          5118 => x"71",
          5119 => x"33",
          5120 => x"71",
          5121 => x"83",
          5122 => x"11",
          5123 => x"12",
          5124 => x"2b",
          5125 => x"07",
          5126 => x"51",
          5127 => x"55",
          5128 => x"80",
          5129 => x"82",
          5130 => x"75",
          5131 => x"3f",
          5132 => x"84",
          5133 => x"15",
          5134 => x"2b",
          5135 => x"07",
          5136 => x"88",
          5137 => x"55",
          5138 => x"86",
          5139 => x"81",
          5140 => x"75",
          5141 => x"82",
          5142 => x"70",
          5143 => x"33",
          5144 => x"71",
          5145 => x"70",
          5146 => x"57",
          5147 => x"72",
          5148 => x"73",
          5149 => x"82",
          5150 => x"18",
          5151 => x"86",
          5152 => x"0b",
          5153 => x"82",
          5154 => x"53",
          5155 => x"34",
          5156 => x"34",
          5157 => x"08",
          5158 => x"81",
          5159 => x"88",
          5160 => x"82",
          5161 => x"70",
          5162 => x"51",
          5163 => x"74",
          5164 => x"81",
          5165 => x"3d",
          5166 => x"3d",
          5167 => x"82",
          5168 => x"84",
          5169 => x"3f",
          5170 => x"86",
          5171 => x"fe",
          5172 => x"3d",
          5173 => x"3d",
          5174 => x"52",
          5175 => x"3f",
          5176 => x"08",
          5177 => x"06",
          5178 => x"08",
          5179 => x"85",
          5180 => x"88",
          5181 => x"5f",
          5182 => x"5a",
          5183 => x"59",
          5184 => x"80",
          5185 => x"88",
          5186 => x"33",
          5187 => x"71",
          5188 => x"70",
          5189 => x"06",
          5190 => x"83",
          5191 => x"70",
          5192 => x"53",
          5193 => x"55",
          5194 => x"8a",
          5195 => x"2e",
          5196 => x"78",
          5197 => x"15",
          5198 => x"33",
          5199 => x"07",
          5200 => x"c2",
          5201 => x"ff",
          5202 => x"38",
          5203 => x"56",
          5204 => x"2b",
          5205 => x"08",
          5206 => x"81",
          5207 => x"88",
          5208 => x"81",
          5209 => x"51",
          5210 => x"5c",
          5211 => x"2e",
          5212 => x"55",
          5213 => x"78",
          5214 => x"38",
          5215 => x"80",
          5216 => x"38",
          5217 => x"09",
          5218 => x"38",
          5219 => x"f2",
          5220 => x"39",
          5221 => x"53",
          5222 => x"51",
          5223 => x"82",
          5224 => x"70",
          5225 => x"33",
          5226 => x"71",
          5227 => x"83",
          5228 => x"5a",
          5229 => x"05",
          5230 => x"83",
          5231 => x"70",
          5232 => x"59",
          5233 => x"84",
          5234 => x"81",
          5235 => x"76",
          5236 => x"82",
          5237 => x"75",
          5238 => x"11",
          5239 => x"11",
          5240 => x"33",
          5241 => x"07",
          5242 => x"53",
          5243 => x"5a",
          5244 => x"86",
          5245 => x"87",
          5246 => x"d5",
          5247 => x"1c",
          5248 => x"85",
          5249 => x"8b",
          5250 => x"2b",
          5251 => x"5a",
          5252 => x"54",
          5253 => x"34",
          5254 => x"34",
          5255 => x"08",
          5256 => x"1d",
          5257 => x"85",
          5258 => x"88",
          5259 => x"88",
          5260 => x"5f",
          5261 => x"73",
          5262 => x"75",
          5263 => x"82",
          5264 => x"1b",
          5265 => x"73",
          5266 => x"0c",
          5267 => x"04",
          5268 => x"74",
          5269 => x"d4",
          5270 => x"f4",
          5271 => x"53",
          5272 => x"8b",
          5273 => x"fc",
          5274 => x"d5",
          5275 => x"72",
          5276 => x"0c",
          5277 => x"04",
          5278 => x"64",
          5279 => x"80",
          5280 => x"82",
          5281 => x"60",
          5282 => x"06",
          5283 => x"a8",
          5284 => x"38",
          5285 => x"b8",
          5286 => x"e4",
          5287 => x"c7",
          5288 => x"38",
          5289 => x"92",
          5290 => x"83",
          5291 => x"51",
          5292 => x"82",
          5293 => x"83",
          5294 => x"82",
          5295 => x"7d",
          5296 => x"2a",
          5297 => x"ff",
          5298 => x"2b",
          5299 => x"33",
          5300 => x"71",
          5301 => x"70",
          5302 => x"83",
          5303 => x"70",
          5304 => x"05",
          5305 => x"1a",
          5306 => x"12",
          5307 => x"2b",
          5308 => x"2b",
          5309 => x"53",
          5310 => x"5c",
          5311 => x"5c",
          5312 => x"73",
          5313 => x"38",
          5314 => x"ff",
          5315 => x"70",
          5316 => x"06",
          5317 => x"16",
          5318 => x"33",
          5319 => x"07",
          5320 => x"1c",
          5321 => x"12",
          5322 => x"2b",
          5323 => x"07",
          5324 => x"52",
          5325 => x"80",
          5326 => x"78",
          5327 => x"83",
          5328 => x"41",
          5329 => x"27",
          5330 => x"60",
          5331 => x"7b",
          5332 => x"06",
          5333 => x"51",
          5334 => x"7a",
          5335 => x"06",
          5336 => x"39",
          5337 => x"7a",
          5338 => x"38",
          5339 => x"aa",
          5340 => x"39",
          5341 => x"7a",
          5342 => x"c8",
          5343 => x"82",
          5344 => x"12",
          5345 => x"2b",
          5346 => x"54",
          5347 => x"80",
          5348 => x"f7",
          5349 => x"d5",
          5350 => x"ff",
          5351 => x"54",
          5352 => x"83",
          5353 => x"d4",
          5354 => x"05",
          5355 => x"ff",
          5356 => x"82",
          5357 => x"14",
          5358 => x"83",
          5359 => x"59",
          5360 => x"39",
          5361 => x"7a",
          5362 => x"d4",
          5363 => x"f5",
          5364 => x"d5",
          5365 => x"82",
          5366 => x"12",
          5367 => x"2b",
          5368 => x"54",
          5369 => x"80",
          5370 => x"f6",
          5371 => x"d5",
          5372 => x"ff",
          5373 => x"54",
          5374 => x"83",
          5375 => x"d4",
          5376 => x"05",
          5377 => x"ff",
          5378 => x"82",
          5379 => x"14",
          5380 => x"62",
          5381 => x"5c",
          5382 => x"ff",
          5383 => x"39",
          5384 => x"54",
          5385 => x"82",
          5386 => x"5c",
          5387 => x"08",
          5388 => x"38",
          5389 => x"52",
          5390 => x"08",
          5391 => x"a6",
          5392 => x"f7",
          5393 => x"58",
          5394 => x"99",
          5395 => x"7a",
          5396 => x"f2",
          5397 => x"19",
          5398 => x"d5",
          5399 => x"84",
          5400 => x"f9",
          5401 => x"73",
          5402 => x"0c",
          5403 => x"04",
          5404 => x"77",
          5405 => x"52",
          5406 => x"3f",
          5407 => x"08",
          5408 => x"e4",
          5409 => x"8e",
          5410 => x"80",
          5411 => x"e4",
          5412 => x"9a",
          5413 => x"82",
          5414 => x"86",
          5415 => x"ff",
          5416 => x"8f",
          5417 => x"81",
          5418 => x"26",
          5419 => x"d5",
          5420 => x"52",
          5421 => x"e4",
          5422 => x"0d",
          5423 => x"0d",
          5424 => x"33",
          5425 => x"9f",
          5426 => x"53",
          5427 => x"81",
          5428 => x"38",
          5429 => x"87",
          5430 => x"11",
          5431 => x"54",
          5432 => x"84",
          5433 => x"54",
          5434 => x"87",
          5435 => x"11",
          5436 => x"0c",
          5437 => x"c0",
          5438 => x"70",
          5439 => x"70",
          5440 => x"51",
          5441 => x"8a",
          5442 => x"98",
          5443 => x"70",
          5444 => x"08",
          5445 => x"06",
          5446 => x"38",
          5447 => x"8c",
          5448 => x"80",
          5449 => x"71",
          5450 => x"14",
          5451 => x"e0",
          5452 => x"70",
          5453 => x"0c",
          5454 => x"04",
          5455 => x"60",
          5456 => x"8c",
          5457 => x"33",
          5458 => x"5b",
          5459 => x"5a",
          5460 => x"82",
          5461 => x"81",
          5462 => x"52",
          5463 => x"38",
          5464 => x"84",
          5465 => x"92",
          5466 => x"c0",
          5467 => x"87",
          5468 => x"13",
          5469 => x"57",
          5470 => x"0b",
          5471 => x"8c",
          5472 => x"0c",
          5473 => x"75",
          5474 => x"2a",
          5475 => x"51",
          5476 => x"80",
          5477 => x"7b",
          5478 => x"7b",
          5479 => x"5d",
          5480 => x"59",
          5481 => x"06",
          5482 => x"73",
          5483 => x"81",
          5484 => x"ff",
          5485 => x"72",
          5486 => x"38",
          5487 => x"8c",
          5488 => x"c3",
          5489 => x"98",
          5490 => x"71",
          5491 => x"38",
          5492 => x"2e",
          5493 => x"76",
          5494 => x"92",
          5495 => x"72",
          5496 => x"06",
          5497 => x"f7",
          5498 => x"5a",
          5499 => x"80",
          5500 => x"70",
          5501 => x"5a",
          5502 => x"80",
          5503 => x"73",
          5504 => x"06",
          5505 => x"38",
          5506 => x"fe",
          5507 => x"fc",
          5508 => x"52",
          5509 => x"83",
          5510 => x"71",
          5511 => x"d5",
          5512 => x"3d",
          5513 => x"3d",
          5514 => x"64",
          5515 => x"bf",
          5516 => x"40",
          5517 => x"59",
          5518 => x"58",
          5519 => x"82",
          5520 => x"81",
          5521 => x"52",
          5522 => x"09",
          5523 => x"b1",
          5524 => x"84",
          5525 => x"92",
          5526 => x"c0",
          5527 => x"87",
          5528 => x"13",
          5529 => x"56",
          5530 => x"87",
          5531 => x"0c",
          5532 => x"82",
          5533 => x"58",
          5534 => x"84",
          5535 => x"06",
          5536 => x"71",
          5537 => x"38",
          5538 => x"05",
          5539 => x"0c",
          5540 => x"73",
          5541 => x"81",
          5542 => x"71",
          5543 => x"38",
          5544 => x"8c",
          5545 => x"d0",
          5546 => x"98",
          5547 => x"71",
          5548 => x"38",
          5549 => x"2e",
          5550 => x"76",
          5551 => x"92",
          5552 => x"72",
          5553 => x"06",
          5554 => x"f7",
          5555 => x"59",
          5556 => x"1a",
          5557 => x"06",
          5558 => x"59",
          5559 => x"80",
          5560 => x"73",
          5561 => x"06",
          5562 => x"38",
          5563 => x"fe",
          5564 => x"fc",
          5565 => x"52",
          5566 => x"83",
          5567 => x"71",
          5568 => x"d5",
          5569 => x"3d",
          5570 => x"3d",
          5571 => x"84",
          5572 => x"33",
          5573 => x"a7",
          5574 => x"54",
          5575 => x"fa",
          5576 => x"d5",
          5577 => x"06",
          5578 => x"72",
          5579 => x"85",
          5580 => x"98",
          5581 => x"56",
          5582 => x"80",
          5583 => x"76",
          5584 => x"74",
          5585 => x"c0",
          5586 => x"54",
          5587 => x"2e",
          5588 => x"d4",
          5589 => x"2e",
          5590 => x"80",
          5591 => x"08",
          5592 => x"70",
          5593 => x"51",
          5594 => x"2e",
          5595 => x"c0",
          5596 => x"52",
          5597 => x"87",
          5598 => x"08",
          5599 => x"38",
          5600 => x"87",
          5601 => x"14",
          5602 => x"70",
          5603 => x"52",
          5604 => x"96",
          5605 => x"92",
          5606 => x"0a",
          5607 => x"39",
          5608 => x"0c",
          5609 => x"39",
          5610 => x"54",
          5611 => x"e4",
          5612 => x"0d",
          5613 => x"0d",
          5614 => x"33",
          5615 => x"88",
          5616 => x"d5",
          5617 => x"51",
          5618 => x"04",
          5619 => x"75",
          5620 => x"82",
          5621 => x"90",
          5622 => x"2b",
          5623 => x"33",
          5624 => x"88",
          5625 => x"71",
          5626 => x"e4",
          5627 => x"54",
          5628 => x"85",
          5629 => x"ff",
          5630 => x"02",
          5631 => x"05",
          5632 => x"70",
          5633 => x"05",
          5634 => x"88",
          5635 => x"72",
          5636 => x"0d",
          5637 => x"0d",
          5638 => x"52",
          5639 => x"81",
          5640 => x"70",
          5641 => x"70",
          5642 => x"05",
          5643 => x"88",
          5644 => x"72",
          5645 => x"54",
          5646 => x"2a",
          5647 => x"34",
          5648 => x"04",
          5649 => x"76",
          5650 => x"54",
          5651 => x"2e",
          5652 => x"70",
          5653 => x"33",
          5654 => x"05",
          5655 => x"11",
          5656 => x"84",
          5657 => x"fe",
          5658 => x"77",
          5659 => x"53",
          5660 => x"81",
          5661 => x"ff",
          5662 => x"f4",
          5663 => x"0d",
          5664 => x"0d",
          5665 => x"56",
          5666 => x"70",
          5667 => x"33",
          5668 => x"05",
          5669 => x"71",
          5670 => x"56",
          5671 => x"72",
          5672 => x"38",
          5673 => x"e2",
          5674 => x"d5",
          5675 => x"3d",
          5676 => x"3d",
          5677 => x"54",
          5678 => x"71",
          5679 => x"38",
          5680 => x"70",
          5681 => x"f3",
          5682 => x"82",
          5683 => x"84",
          5684 => x"80",
          5685 => x"e4",
          5686 => x"3d",
          5687 => x"08",
          5688 => x"05",
          5689 => x"54",
          5690 => x"e7",
          5691 => x"82",
          5692 => x"a2",
          5693 => x"2e",
          5694 => x"b5",
          5695 => x"80",
          5696 => x"82",
          5697 => x"83",
          5698 => x"53",
          5699 => x"86",
          5700 => x"0c",
          5701 => x"82",
          5702 => x"87",
          5703 => x"f7",
          5704 => x"56",
          5705 => x"17",
          5706 => x"74",
          5707 => x"d6",
          5708 => x"b4",
          5709 => x"b8",
          5710 => x"81",
          5711 => x"59",
          5712 => x"82",
          5713 => x"7a",
          5714 => x"06",
          5715 => x"d5",
          5716 => x"17",
          5717 => x"08",
          5718 => x"08",
          5719 => x"08",
          5720 => x"74",
          5721 => x"38",
          5722 => x"55",
          5723 => x"09",
          5724 => x"38",
          5725 => x"18",
          5726 => x"81",
          5727 => x"f9",
          5728 => x"39",
          5729 => x"82",
          5730 => x"8b",
          5731 => x"fa",
          5732 => x"7a",
          5733 => x"57",
          5734 => x"08",
          5735 => x"75",
          5736 => x"3f",
          5737 => x"08",
          5738 => x"e4",
          5739 => x"81",
          5740 => x"b8",
          5741 => x"16",
          5742 => x"80",
          5743 => x"e4",
          5744 => x"85",
          5745 => x"81",
          5746 => x"17",
          5747 => x"d5",
          5748 => x"3d",
          5749 => x"3d",
          5750 => x"52",
          5751 => x"3f",
          5752 => x"08",
          5753 => x"e4",
          5754 => x"38",
          5755 => x"74",
          5756 => x"81",
          5757 => x"38",
          5758 => x"59",
          5759 => x"09",
          5760 => x"e3",
          5761 => x"53",
          5762 => x"08",
          5763 => x"70",
          5764 => x"d3",
          5765 => x"d5",
          5766 => x"17",
          5767 => x"3f",
          5768 => x"a4",
          5769 => x"51",
          5770 => x"86",
          5771 => x"f2",
          5772 => x"17",
          5773 => x"3f",
          5774 => x"52",
          5775 => x"51",
          5776 => x"90",
          5777 => x"84",
          5778 => x"fb",
          5779 => x"17",
          5780 => x"70",
          5781 => x"79",
          5782 => x"52",
          5783 => x"51",
          5784 => x"77",
          5785 => x"80",
          5786 => x"81",
          5787 => x"f9",
          5788 => x"d5",
          5789 => x"2e",
          5790 => x"58",
          5791 => x"e4",
          5792 => x"0d",
          5793 => x"0d",
          5794 => x"9c",
          5795 => x"05",
          5796 => x"80",
          5797 => x"27",
          5798 => x"14",
          5799 => x"29",
          5800 => x"05",
          5801 => x"82",
          5802 => x"87",
          5803 => x"f9",
          5804 => x"7a",
          5805 => x"54",
          5806 => x"27",
          5807 => x"76",
          5808 => x"27",
          5809 => x"ff",
          5810 => x"58",
          5811 => x"80",
          5812 => x"82",
          5813 => x"72",
          5814 => x"38",
          5815 => x"72",
          5816 => x"8e",
          5817 => x"39",
          5818 => x"17",
          5819 => x"a8",
          5820 => x"53",
          5821 => x"fd",
          5822 => x"d5",
          5823 => x"9f",
          5824 => x"ff",
          5825 => x"11",
          5826 => x"70",
          5827 => x"18",
          5828 => x"76",
          5829 => x"53",
          5830 => x"82",
          5831 => x"80",
          5832 => x"83",
          5833 => x"b8",
          5834 => x"88",
          5835 => x"79",
          5836 => x"84",
          5837 => x"58",
          5838 => x"80",
          5839 => x"9f",
          5840 => x"80",
          5841 => x"88",
          5842 => x"08",
          5843 => x"51",
          5844 => x"82",
          5845 => x"80",
          5846 => x"10",
          5847 => x"74",
          5848 => x"51",
          5849 => x"82",
          5850 => x"83",
          5851 => x"58",
          5852 => x"87",
          5853 => x"08",
          5854 => x"51",
          5855 => x"82",
          5856 => x"9b",
          5857 => x"2b",
          5858 => x"74",
          5859 => x"51",
          5860 => x"82",
          5861 => x"f0",
          5862 => x"83",
          5863 => x"77",
          5864 => x"0c",
          5865 => x"04",
          5866 => x"7a",
          5867 => x"58",
          5868 => x"81",
          5869 => x"9e",
          5870 => x"17",
          5871 => x"96",
          5872 => x"53",
          5873 => x"81",
          5874 => x"79",
          5875 => x"72",
          5876 => x"38",
          5877 => x"72",
          5878 => x"b8",
          5879 => x"39",
          5880 => x"17",
          5881 => x"a8",
          5882 => x"53",
          5883 => x"fb",
          5884 => x"d5",
          5885 => x"82",
          5886 => x"81",
          5887 => x"83",
          5888 => x"b8",
          5889 => x"78",
          5890 => x"56",
          5891 => x"76",
          5892 => x"38",
          5893 => x"9f",
          5894 => x"33",
          5895 => x"07",
          5896 => x"74",
          5897 => x"83",
          5898 => x"89",
          5899 => x"08",
          5900 => x"51",
          5901 => x"82",
          5902 => x"59",
          5903 => x"08",
          5904 => x"74",
          5905 => x"16",
          5906 => x"84",
          5907 => x"76",
          5908 => x"88",
          5909 => x"81",
          5910 => x"8f",
          5911 => x"53",
          5912 => x"80",
          5913 => x"88",
          5914 => x"08",
          5915 => x"51",
          5916 => x"82",
          5917 => x"59",
          5918 => x"08",
          5919 => x"77",
          5920 => x"06",
          5921 => x"83",
          5922 => x"05",
          5923 => x"f6",
          5924 => x"39",
          5925 => x"a8",
          5926 => x"52",
          5927 => x"ef",
          5928 => x"e4",
          5929 => x"d5",
          5930 => x"38",
          5931 => x"06",
          5932 => x"83",
          5933 => x"18",
          5934 => x"54",
          5935 => x"f6",
          5936 => x"d5",
          5937 => x"0a",
          5938 => x"52",
          5939 => x"c5",
          5940 => x"83",
          5941 => x"82",
          5942 => x"8a",
          5943 => x"f8",
          5944 => x"7c",
          5945 => x"59",
          5946 => x"81",
          5947 => x"38",
          5948 => x"08",
          5949 => x"73",
          5950 => x"38",
          5951 => x"52",
          5952 => x"a4",
          5953 => x"e4",
          5954 => x"d5",
          5955 => x"f2",
          5956 => x"82",
          5957 => x"39",
          5958 => x"e6",
          5959 => x"e4",
          5960 => x"de",
          5961 => x"78",
          5962 => x"3f",
          5963 => x"08",
          5964 => x"e4",
          5965 => x"80",
          5966 => x"d5",
          5967 => x"2e",
          5968 => x"d5",
          5969 => x"2e",
          5970 => x"53",
          5971 => x"51",
          5972 => x"82",
          5973 => x"c5",
          5974 => x"08",
          5975 => x"18",
          5976 => x"57",
          5977 => x"90",
          5978 => x"94",
          5979 => x"16",
          5980 => x"54",
          5981 => x"34",
          5982 => x"78",
          5983 => x"38",
          5984 => x"82",
          5985 => x"8a",
          5986 => x"f6",
          5987 => x"7e",
          5988 => x"5b",
          5989 => x"38",
          5990 => x"58",
          5991 => x"88",
          5992 => x"08",
          5993 => x"38",
          5994 => x"39",
          5995 => x"51",
          5996 => x"81",
          5997 => x"d5",
          5998 => x"82",
          5999 => x"d5",
          6000 => x"82",
          6001 => x"ff",
          6002 => x"38",
          6003 => x"82",
          6004 => x"26",
          6005 => x"79",
          6006 => x"08",
          6007 => x"73",
          6008 => x"b9",
          6009 => x"2e",
          6010 => x"80",
          6011 => x"1a",
          6012 => x"08",
          6013 => x"38",
          6014 => x"52",
          6015 => x"af",
          6016 => x"82",
          6017 => x"81",
          6018 => x"06",
          6019 => x"d5",
          6020 => x"82",
          6021 => x"09",
          6022 => x"72",
          6023 => x"70",
          6024 => x"d5",
          6025 => x"51",
          6026 => x"73",
          6027 => x"82",
          6028 => x"80",
          6029 => x"90",
          6030 => x"81",
          6031 => x"38",
          6032 => x"08",
          6033 => x"73",
          6034 => x"75",
          6035 => x"77",
          6036 => x"56",
          6037 => x"76",
          6038 => x"82",
          6039 => x"26",
          6040 => x"75",
          6041 => x"f8",
          6042 => x"d5",
          6043 => x"2e",
          6044 => x"59",
          6045 => x"08",
          6046 => x"81",
          6047 => x"82",
          6048 => x"59",
          6049 => x"08",
          6050 => x"70",
          6051 => x"25",
          6052 => x"51",
          6053 => x"73",
          6054 => x"75",
          6055 => x"81",
          6056 => x"38",
          6057 => x"f5",
          6058 => x"75",
          6059 => x"f9",
          6060 => x"d5",
          6061 => x"d5",
          6062 => x"70",
          6063 => x"08",
          6064 => x"51",
          6065 => x"80",
          6066 => x"73",
          6067 => x"38",
          6068 => x"52",
          6069 => x"d0",
          6070 => x"e4",
          6071 => x"a5",
          6072 => x"18",
          6073 => x"08",
          6074 => x"18",
          6075 => x"74",
          6076 => x"38",
          6077 => x"18",
          6078 => x"33",
          6079 => x"73",
          6080 => x"97",
          6081 => x"74",
          6082 => x"38",
          6083 => x"55",
          6084 => x"d5",
          6085 => x"85",
          6086 => x"75",
          6087 => x"d5",
          6088 => x"3d",
          6089 => x"3d",
          6090 => x"52",
          6091 => x"3f",
          6092 => x"08",
          6093 => x"82",
          6094 => x"80",
          6095 => x"52",
          6096 => x"c1",
          6097 => x"e4",
          6098 => x"e4",
          6099 => x"0c",
          6100 => x"53",
          6101 => x"15",
          6102 => x"f2",
          6103 => x"56",
          6104 => x"16",
          6105 => x"22",
          6106 => x"27",
          6107 => x"54",
          6108 => x"76",
          6109 => x"33",
          6110 => x"3f",
          6111 => x"08",
          6112 => x"38",
          6113 => x"76",
          6114 => x"70",
          6115 => x"9f",
          6116 => x"56",
          6117 => x"d5",
          6118 => x"3d",
          6119 => x"3d",
          6120 => x"71",
          6121 => x"57",
          6122 => x"0a",
          6123 => x"38",
          6124 => x"53",
          6125 => x"38",
          6126 => x"0c",
          6127 => x"54",
          6128 => x"75",
          6129 => x"73",
          6130 => x"ac",
          6131 => x"73",
          6132 => x"85",
          6133 => x"0b",
          6134 => x"5a",
          6135 => x"27",
          6136 => x"ac",
          6137 => x"18",
          6138 => x"39",
          6139 => x"70",
          6140 => x"58",
          6141 => x"b2",
          6142 => x"76",
          6143 => x"3f",
          6144 => x"08",
          6145 => x"e4",
          6146 => x"bd",
          6147 => x"82",
          6148 => x"27",
          6149 => x"16",
          6150 => x"e4",
          6151 => x"38",
          6152 => x"39",
          6153 => x"55",
          6154 => x"52",
          6155 => x"d5",
          6156 => x"e4",
          6157 => x"0c",
          6158 => x"0c",
          6159 => x"53",
          6160 => x"80",
          6161 => x"85",
          6162 => x"94",
          6163 => x"2a",
          6164 => x"0c",
          6165 => x"06",
          6166 => x"9c",
          6167 => x"58",
          6168 => x"e4",
          6169 => x"0d",
          6170 => x"0d",
          6171 => x"90",
          6172 => x"05",
          6173 => x"f0",
          6174 => x"27",
          6175 => x"0b",
          6176 => x"98",
          6177 => x"84",
          6178 => x"2e",
          6179 => x"76",
          6180 => x"58",
          6181 => x"38",
          6182 => x"15",
          6183 => x"08",
          6184 => x"38",
          6185 => x"88",
          6186 => x"53",
          6187 => x"81",
          6188 => x"c0",
          6189 => x"22",
          6190 => x"89",
          6191 => x"72",
          6192 => x"74",
          6193 => x"f3",
          6194 => x"d5",
          6195 => x"82",
          6196 => x"82",
          6197 => x"27",
          6198 => x"81",
          6199 => x"e4",
          6200 => x"80",
          6201 => x"16",
          6202 => x"e4",
          6203 => x"ca",
          6204 => x"38",
          6205 => x"0c",
          6206 => x"dd",
          6207 => x"08",
          6208 => x"f9",
          6209 => x"d5",
          6210 => x"87",
          6211 => x"e4",
          6212 => x"80",
          6213 => x"55",
          6214 => x"08",
          6215 => x"38",
          6216 => x"d5",
          6217 => x"2e",
          6218 => x"d5",
          6219 => x"75",
          6220 => x"3f",
          6221 => x"08",
          6222 => x"94",
          6223 => x"52",
          6224 => x"c1",
          6225 => x"e4",
          6226 => x"0c",
          6227 => x"0c",
          6228 => x"05",
          6229 => x"80",
          6230 => x"d5",
          6231 => x"3d",
          6232 => x"3d",
          6233 => x"71",
          6234 => x"57",
          6235 => x"51",
          6236 => x"82",
          6237 => x"54",
          6238 => x"08",
          6239 => x"82",
          6240 => x"56",
          6241 => x"52",
          6242 => x"83",
          6243 => x"e4",
          6244 => x"d5",
          6245 => x"d2",
          6246 => x"e4",
          6247 => x"08",
          6248 => x"54",
          6249 => x"e5",
          6250 => x"06",
          6251 => x"58",
          6252 => x"08",
          6253 => x"38",
          6254 => x"75",
          6255 => x"80",
          6256 => x"81",
          6257 => x"7a",
          6258 => x"06",
          6259 => x"39",
          6260 => x"08",
          6261 => x"76",
          6262 => x"3f",
          6263 => x"08",
          6264 => x"e4",
          6265 => x"ff",
          6266 => x"84",
          6267 => x"06",
          6268 => x"54",
          6269 => x"e4",
          6270 => x"0d",
          6271 => x"0d",
          6272 => x"52",
          6273 => x"3f",
          6274 => x"08",
          6275 => x"06",
          6276 => x"51",
          6277 => x"83",
          6278 => x"06",
          6279 => x"14",
          6280 => x"3f",
          6281 => x"08",
          6282 => x"07",
          6283 => x"d5",
          6284 => x"3d",
          6285 => x"3d",
          6286 => x"70",
          6287 => x"06",
          6288 => x"53",
          6289 => x"af",
          6290 => x"33",
          6291 => x"83",
          6292 => x"06",
          6293 => x"90",
          6294 => x"15",
          6295 => x"3f",
          6296 => x"04",
          6297 => x"75",
          6298 => x"8b",
          6299 => x"2a",
          6300 => x"29",
          6301 => x"81",
          6302 => x"71",
          6303 => x"ff",
          6304 => x"56",
          6305 => x"72",
          6306 => x"82",
          6307 => x"85",
          6308 => x"f2",
          6309 => x"62",
          6310 => x"79",
          6311 => x"81",
          6312 => x"5d",
          6313 => x"80",
          6314 => x"38",
          6315 => x"52",
          6316 => x"db",
          6317 => x"e4",
          6318 => x"d5",
          6319 => x"eb",
          6320 => x"08",
          6321 => x"55",
          6322 => x"84",
          6323 => x"39",
          6324 => x"bf",
          6325 => x"ff",
          6326 => x"72",
          6327 => x"82",
          6328 => x"56",
          6329 => x"2e",
          6330 => x"83",
          6331 => x"82",
          6332 => x"53",
          6333 => x"09",
          6334 => x"38",
          6335 => x"73",
          6336 => x"99",
          6337 => x"e4",
          6338 => x"06",
          6339 => x"88",
          6340 => x"06",
          6341 => x"56",
          6342 => x"87",
          6343 => x"5c",
          6344 => x"76",
          6345 => x"81",
          6346 => x"38",
          6347 => x"70",
          6348 => x"53",
          6349 => x"92",
          6350 => x"33",
          6351 => x"06",
          6352 => x"08",
          6353 => x"56",
          6354 => x"7c",
          6355 => x"06",
          6356 => x"8d",
          6357 => x"7c",
          6358 => x"81",
          6359 => x"38",
          6360 => x"9a",
          6361 => x"e8",
          6362 => x"d5",
          6363 => x"ff",
          6364 => x"72",
          6365 => x"74",
          6366 => x"bf",
          6367 => x"f3",
          6368 => x"81",
          6369 => x"82",
          6370 => x"33",
          6371 => x"e8",
          6372 => x"d5",
          6373 => x"ff",
          6374 => x"77",
          6375 => x"38",
          6376 => x"26",
          6377 => x"73",
          6378 => x"59",
          6379 => x"23",
          6380 => x"8b",
          6381 => x"ff",
          6382 => x"81",
          6383 => x"81",
          6384 => x"77",
          6385 => x"74",
          6386 => x"2a",
          6387 => x"51",
          6388 => x"80",
          6389 => x"73",
          6390 => x"92",
          6391 => x"1a",
          6392 => x"23",
          6393 => x"81",
          6394 => x"53",
          6395 => x"ff",
          6396 => x"9d",
          6397 => x"38",
          6398 => x"e8",
          6399 => x"e4",
          6400 => x"06",
          6401 => x"2e",
          6402 => x"0b",
          6403 => x"a0",
          6404 => x"78",
          6405 => x"3f",
          6406 => x"08",
          6407 => x"e4",
          6408 => x"98",
          6409 => x"84",
          6410 => x"80",
          6411 => x"0c",
          6412 => x"e4",
          6413 => x"0d",
          6414 => x"0d",
          6415 => x"40",
          6416 => x"78",
          6417 => x"3f",
          6418 => x"08",
          6419 => x"e4",
          6420 => x"38",
          6421 => x"5f",
          6422 => x"ac",
          6423 => x"19",
          6424 => x"51",
          6425 => x"82",
          6426 => x"58",
          6427 => x"08",
          6428 => x"9c",
          6429 => x"33",
          6430 => x"86",
          6431 => x"82",
          6432 => x"17",
          6433 => x"70",
          6434 => x"56",
          6435 => x"1a",
          6436 => x"e5",
          6437 => x"38",
          6438 => x"70",
          6439 => x"54",
          6440 => x"8e",
          6441 => x"b2",
          6442 => x"2e",
          6443 => x"81",
          6444 => x"19",
          6445 => x"2a",
          6446 => x"51",
          6447 => x"82",
          6448 => x"86",
          6449 => x"06",
          6450 => x"80",
          6451 => x"8d",
          6452 => x"81",
          6453 => x"90",
          6454 => x"1d",
          6455 => x"5e",
          6456 => x"09",
          6457 => x"b9",
          6458 => x"33",
          6459 => x"2e",
          6460 => x"81",
          6461 => x"1f",
          6462 => x"52",
          6463 => x"3f",
          6464 => x"08",
          6465 => x"06",
          6466 => x"95",
          6467 => x"70",
          6468 => x"29",
          6469 => x"56",
          6470 => x"5a",
          6471 => x"1b",
          6472 => x"51",
          6473 => x"82",
          6474 => x"83",
          6475 => x"56",
          6476 => x"b1",
          6477 => x"fe",
          6478 => x"38",
          6479 => x"e1",
          6480 => x"d5",
          6481 => x"10",
          6482 => x"53",
          6483 => x"59",
          6484 => x"8d",
          6485 => x"d5",
          6486 => x"09",
          6487 => x"c1",
          6488 => x"8b",
          6489 => x"ff",
          6490 => x"81",
          6491 => x"81",
          6492 => x"7b",
          6493 => x"38",
          6494 => x"86",
          6495 => x"06",
          6496 => x"79",
          6497 => x"38",
          6498 => x"8b",
          6499 => x"1d",
          6500 => x"54",
          6501 => x"ff",
          6502 => x"ff",
          6503 => x"84",
          6504 => x"54",
          6505 => x"39",
          6506 => x"76",
          6507 => x"3f",
          6508 => x"08",
          6509 => x"54",
          6510 => x"bb",
          6511 => x"33",
          6512 => x"73",
          6513 => x"53",
          6514 => x"9c",
          6515 => x"e5",
          6516 => x"d5",
          6517 => x"2e",
          6518 => x"ff",
          6519 => x"ac",
          6520 => x"52",
          6521 => x"81",
          6522 => x"e4",
          6523 => x"d5",
          6524 => x"2e",
          6525 => x"77",
          6526 => x"0c",
          6527 => x"04",
          6528 => x"64",
          6529 => x"12",
          6530 => x"06",
          6531 => x"86",
          6532 => x"b5",
          6533 => x"1d",
          6534 => x"56",
          6535 => x"80",
          6536 => x"81",
          6537 => x"16",
          6538 => x"55",
          6539 => x"8c",
          6540 => x"70",
          6541 => x"70",
          6542 => x"e4",
          6543 => x"80",
          6544 => x"81",
          6545 => x"80",
          6546 => x"38",
          6547 => x"ab",
          6548 => x"5b",
          6549 => x"7b",
          6550 => x"53",
          6551 => x"51",
          6552 => x"85",
          6553 => x"c6",
          6554 => x"77",
          6555 => x"ff",
          6556 => x"55",
          6557 => x"b4",
          6558 => x"ff",
          6559 => x"19",
          6560 => x"57",
          6561 => x"76",
          6562 => x"81",
          6563 => x"2a",
          6564 => x"51",
          6565 => x"73",
          6566 => x"38",
          6567 => x"a1",
          6568 => x"17",
          6569 => x"25",
          6570 => x"39",
          6571 => x"02",
          6572 => x"05",
          6573 => x"b0",
          6574 => x"54",
          6575 => x"84",
          6576 => x"54",
          6577 => x"ff",
          6578 => x"76",
          6579 => x"58",
          6580 => x"38",
          6581 => x"05",
          6582 => x"fe",
          6583 => x"77",
          6584 => x"78",
          6585 => x"a0",
          6586 => x"74",
          6587 => x"52",
          6588 => x"3f",
          6589 => x"08",
          6590 => x"38",
          6591 => x"74",
          6592 => x"38",
          6593 => x"81",
          6594 => x"77",
          6595 => x"74",
          6596 => x"51",
          6597 => x"94",
          6598 => x"eb",
          6599 => x"15",
          6600 => x"58",
          6601 => x"87",
          6602 => x"81",
          6603 => x"70",
          6604 => x"57",
          6605 => x"87",
          6606 => x"38",
          6607 => x"f9",
          6608 => x"e4",
          6609 => x"81",
          6610 => x"e3",
          6611 => x"84",
          6612 => x"7a",
          6613 => x"82",
          6614 => x"d5",
          6615 => x"82",
          6616 => x"84",
          6617 => x"06",
          6618 => x"02",
          6619 => x"33",
          6620 => x"02",
          6621 => x"33",
          6622 => x"70",
          6623 => x"55",
          6624 => x"73",
          6625 => x"38",
          6626 => x"1d",
          6627 => x"9f",
          6628 => x"e4",
          6629 => x"78",
          6630 => x"f3",
          6631 => x"d5",
          6632 => x"82",
          6633 => x"82",
          6634 => x"19",
          6635 => x"2e",
          6636 => x"78",
          6637 => x"1b",
          6638 => x"53",
          6639 => x"ef",
          6640 => x"d5",
          6641 => x"82",
          6642 => x"81",
          6643 => x"1a",
          6644 => x"3f",
          6645 => x"08",
          6646 => x"5d",
          6647 => x"52",
          6648 => x"ab",
          6649 => x"e4",
          6650 => x"d5",
          6651 => x"d7",
          6652 => x"08",
          6653 => x"7a",
          6654 => x"5a",
          6655 => x"8d",
          6656 => x"0b",
          6657 => x"82",
          6658 => x"8c",
          6659 => x"d5",
          6660 => x"9a",
          6661 => x"df",
          6662 => x"29",
          6663 => x"55",
          6664 => x"ff",
          6665 => x"38",
          6666 => x"70",
          6667 => x"57",
          6668 => x"52",
          6669 => x"17",
          6670 => x"51",
          6671 => x"73",
          6672 => x"ff",
          6673 => x"17",
          6674 => x"27",
          6675 => x"83",
          6676 => x"8b",
          6677 => x"1b",
          6678 => x"54",
          6679 => x"77",
          6680 => x"58",
          6681 => x"81",
          6682 => x"34",
          6683 => x"51",
          6684 => x"82",
          6685 => x"57",
          6686 => x"08",
          6687 => x"ff",
          6688 => x"fe",
          6689 => x"1a",
          6690 => x"51",
          6691 => x"82",
          6692 => x"57",
          6693 => x"08",
          6694 => x"53",
          6695 => x"08",
          6696 => x"08",
          6697 => x"3f",
          6698 => x"1a",
          6699 => x"08",
          6700 => x"3f",
          6701 => x"ab",
          6702 => x"06",
          6703 => x"8c",
          6704 => x"0b",
          6705 => x"76",
          6706 => x"d5",
          6707 => x"3d",
          6708 => x"3d",
          6709 => x"08",
          6710 => x"ac",
          6711 => x"59",
          6712 => x"ff",
          6713 => x"72",
          6714 => x"ed",
          6715 => x"d5",
          6716 => x"82",
          6717 => x"80",
          6718 => x"15",
          6719 => x"51",
          6720 => x"82",
          6721 => x"54",
          6722 => x"08",
          6723 => x"15",
          6724 => x"73",
          6725 => x"83",
          6726 => x"15",
          6727 => x"a2",
          6728 => x"e4",
          6729 => x"51",
          6730 => x"82",
          6731 => x"54",
          6732 => x"08",
          6733 => x"38",
          6734 => x"09",
          6735 => x"38",
          6736 => x"82",
          6737 => x"88",
          6738 => x"f4",
          6739 => x"60",
          6740 => x"59",
          6741 => x"96",
          6742 => x"1c",
          6743 => x"83",
          6744 => x"1c",
          6745 => x"81",
          6746 => x"70",
          6747 => x"05",
          6748 => x"57",
          6749 => x"57",
          6750 => x"81",
          6751 => x"10",
          6752 => x"81",
          6753 => x"53",
          6754 => x"80",
          6755 => x"70",
          6756 => x"06",
          6757 => x"8f",
          6758 => x"38",
          6759 => x"df",
          6760 => x"96",
          6761 => x"79",
          6762 => x"54",
          6763 => x"7a",
          6764 => x"07",
          6765 => x"84",
          6766 => x"e4",
          6767 => x"ff",
          6768 => x"ff",
          6769 => x"38",
          6770 => x"a5",
          6771 => x"2a",
          6772 => x"34",
          6773 => x"34",
          6774 => x"39",
          6775 => x"30",
          6776 => x"80",
          6777 => x"25",
          6778 => x"54",
          6779 => x"85",
          6780 => x"9a",
          6781 => x"34",
          6782 => x"17",
          6783 => x"8c",
          6784 => x"10",
          6785 => x"51",
          6786 => x"fe",
          6787 => x"30",
          6788 => x"70",
          6789 => x"59",
          6790 => x"17",
          6791 => x"80",
          6792 => x"34",
          6793 => x"1a",
          6794 => x"9c",
          6795 => x"70",
          6796 => x"5b",
          6797 => x"a0",
          6798 => x"74",
          6799 => x"81",
          6800 => x"81",
          6801 => x"89",
          6802 => x"70",
          6803 => x"25",
          6804 => x"76",
          6805 => x"38",
          6806 => x"8b",
          6807 => x"70",
          6808 => x"34",
          6809 => x"74",
          6810 => x"05",
          6811 => x"17",
          6812 => x"27",
          6813 => x"77",
          6814 => x"53",
          6815 => x"14",
          6816 => x"33",
          6817 => x"87",
          6818 => x"38",
          6819 => x"19",
          6820 => x"80",
          6821 => x"73",
          6822 => x"55",
          6823 => x"80",
          6824 => x"38",
          6825 => x"19",
          6826 => x"33",
          6827 => x"54",
          6828 => x"26",
          6829 => x"1c",
          6830 => x"33",
          6831 => x"79",
          6832 => x"72",
          6833 => x"85",
          6834 => x"2a",
          6835 => x"06",
          6836 => x"2e",
          6837 => x"15",
          6838 => x"ff",
          6839 => x"74",
          6840 => x"05",
          6841 => x"19",
          6842 => x"19",
          6843 => x"59",
          6844 => x"ff",
          6845 => x"17",
          6846 => x"80",
          6847 => x"34",
          6848 => x"8c",
          6849 => x"53",
          6850 => x"72",
          6851 => x"9c",
          6852 => x"8b",
          6853 => x"19",
          6854 => x"08",
          6855 => x"53",
          6856 => x"82",
          6857 => x"78",
          6858 => x"51",
          6859 => x"82",
          6860 => x"86",
          6861 => x"13",
          6862 => x"3f",
          6863 => x"08",
          6864 => x"8e",
          6865 => x"f0",
          6866 => x"70",
          6867 => x"80",
          6868 => x"51",
          6869 => x"af",
          6870 => x"81",
          6871 => x"dc",
          6872 => x"74",
          6873 => x"38",
          6874 => x"08",
          6875 => x"aa",
          6876 => x"44",
          6877 => x"33",
          6878 => x"73",
          6879 => x"81",
          6880 => x"81",
          6881 => x"dc",
          6882 => x"70",
          6883 => x"07",
          6884 => x"73",
          6885 => x"88",
          6886 => x"70",
          6887 => x"73",
          6888 => x"38",
          6889 => x"ab",
          6890 => x"52",
          6891 => x"ee",
          6892 => x"e4",
          6893 => x"e1",
          6894 => x"7d",
          6895 => x"08",
          6896 => x"59",
          6897 => x"05",
          6898 => x"3f",
          6899 => x"08",
          6900 => x"b1",
          6901 => x"ff",
          6902 => x"e4",
          6903 => x"38",
          6904 => x"82",
          6905 => x"90",
          6906 => x"73",
          6907 => x"19",
          6908 => x"e4",
          6909 => x"ff",
          6910 => x"32",
          6911 => x"73",
          6912 => x"25",
          6913 => x"55",
          6914 => x"38",
          6915 => x"2e",
          6916 => x"80",
          6917 => x"38",
          6918 => x"c7",
          6919 => x"92",
          6920 => x"e4",
          6921 => x"38",
          6922 => x"26",
          6923 => x"78",
          6924 => x"75",
          6925 => x"19",
          6926 => x"39",
          6927 => x"80",
          6928 => x"56",
          6929 => x"af",
          6930 => x"06",
          6931 => x"57",
          6932 => x"32",
          6933 => x"80",
          6934 => x"51",
          6935 => x"dc",
          6936 => x"9f",
          6937 => x"2b",
          6938 => x"2e",
          6939 => x"8c",
          6940 => x"54",
          6941 => x"a5",
          6942 => x"39",
          6943 => x"09",
          6944 => x"c9",
          6945 => x"22",
          6946 => x"2e",
          6947 => x"80",
          6948 => x"22",
          6949 => x"2e",
          6950 => x"b6",
          6951 => x"1a",
          6952 => x"23",
          6953 => x"1f",
          6954 => x"54",
          6955 => x"83",
          6956 => x"73",
          6957 => x"05",
          6958 => x"18",
          6959 => x"27",
          6960 => x"a0",
          6961 => x"ab",
          6962 => x"c4",
          6963 => x"2e",
          6964 => x"10",
          6965 => x"55",
          6966 => x"16",
          6967 => x"32",
          6968 => x"9f",
          6969 => x"53",
          6970 => x"75",
          6971 => x"38",
          6972 => x"ff",
          6973 => x"e0",
          6974 => x"7a",
          6975 => x"80",
          6976 => x"8d",
          6977 => x"85",
          6978 => x"83",
          6979 => x"99",
          6980 => x"22",
          6981 => x"ff",
          6982 => x"5d",
          6983 => x"09",
          6984 => x"38",
          6985 => x"10",
          6986 => x"51",
          6987 => x"a0",
          6988 => x"7c",
          6989 => x"83",
          6990 => x"54",
          6991 => x"09",
          6992 => x"38",
          6993 => x"57",
          6994 => x"aa",
          6995 => x"fe",
          6996 => x"51",
          6997 => x"2e",
          6998 => x"10",
          6999 => x"55",
          7000 => x"78",
          7001 => x"38",
          7002 => x"22",
          7003 => x"ae",
          7004 => x"06",
          7005 => x"53",
          7006 => x"1e",
          7007 => x"3f",
          7008 => x"5c",
          7009 => x"10",
          7010 => x"81",
          7011 => x"54",
          7012 => x"82",
          7013 => x"a0",
          7014 => x"75",
          7015 => x"30",
          7016 => x"51",
          7017 => x"79",
          7018 => x"73",
          7019 => x"38",
          7020 => x"57",
          7021 => x"54",
          7022 => x"78",
          7023 => x"81",
          7024 => x"32",
          7025 => x"72",
          7026 => x"70",
          7027 => x"51",
          7028 => x"80",
          7029 => x"7e",
          7030 => x"ae",
          7031 => x"2e",
          7032 => x"83",
          7033 => x"79",
          7034 => x"38",
          7035 => x"58",
          7036 => x"2b",
          7037 => x"5d",
          7038 => x"39",
          7039 => x"27",
          7040 => x"82",
          7041 => x"b5",
          7042 => x"80",
          7043 => x"82",
          7044 => x"83",
          7045 => x"70",
          7046 => x"81",
          7047 => x"56",
          7048 => x"8c",
          7049 => x"ff",
          7050 => x"f4",
          7051 => x"54",
          7052 => x"27",
          7053 => x"1f",
          7054 => x"26",
          7055 => x"83",
          7056 => x"57",
          7057 => x"7d",
          7058 => x"76",
          7059 => x"55",
          7060 => x"81",
          7061 => x"c3",
          7062 => x"2e",
          7063 => x"52",
          7064 => x"51",
          7065 => x"82",
          7066 => x"80",
          7067 => x"80",
          7068 => x"07",
          7069 => x"39",
          7070 => x"54",
          7071 => x"85",
          7072 => x"07",
          7073 => x"16",
          7074 => x"26",
          7075 => x"81",
          7076 => x"70",
          7077 => x"06",
          7078 => x"7d",
          7079 => x"54",
          7080 => x"81",
          7081 => x"de",
          7082 => x"33",
          7083 => x"e5",
          7084 => x"06",
          7085 => x"0b",
          7086 => x"7e",
          7087 => x"81",
          7088 => x"7b",
          7089 => x"fc",
          7090 => x"8c",
          7091 => x"8c",
          7092 => x"7b",
          7093 => x"73",
          7094 => x"81",
          7095 => x"76",
          7096 => x"76",
          7097 => x"81",
          7098 => x"73",
          7099 => x"81",
          7100 => x"80",
          7101 => x"76",
          7102 => x"7b",
          7103 => x"81",
          7104 => x"73",
          7105 => x"38",
          7106 => x"57",
          7107 => x"34",
          7108 => x"a5",
          7109 => x"e4",
          7110 => x"33",
          7111 => x"d5",
          7112 => x"2e",
          7113 => x"d5",
          7114 => x"2e",
          7115 => x"80",
          7116 => x"85",
          7117 => x"06",
          7118 => x"57",
          7119 => x"80",
          7120 => x"74",
          7121 => x"73",
          7122 => x"ed",
          7123 => x"0b",
          7124 => x"80",
          7125 => x"39",
          7126 => x"54",
          7127 => x"85",
          7128 => x"74",
          7129 => x"81",
          7130 => x"73",
          7131 => x"1e",
          7132 => x"2a",
          7133 => x"51",
          7134 => x"80",
          7135 => x"90",
          7136 => x"ff",
          7137 => x"b8",
          7138 => x"51",
          7139 => x"82",
          7140 => x"88",
          7141 => x"a1",
          7142 => x"d5",
          7143 => x"3d",
          7144 => x"3d",
          7145 => x"ff",
          7146 => x"71",
          7147 => x"5c",
          7148 => x"80",
          7149 => x"38",
          7150 => x"05",
          7151 => x"9f",
          7152 => x"71",
          7153 => x"38",
          7154 => x"71",
          7155 => x"81",
          7156 => x"38",
          7157 => x"11",
          7158 => x"06",
          7159 => x"70",
          7160 => x"38",
          7161 => x"81",
          7162 => x"05",
          7163 => x"76",
          7164 => x"38",
          7165 => x"c7",
          7166 => x"77",
          7167 => x"57",
          7168 => x"05",
          7169 => x"70",
          7170 => x"33",
          7171 => x"53",
          7172 => x"99",
          7173 => x"e0",
          7174 => x"ff",
          7175 => x"ff",
          7176 => x"70",
          7177 => x"38",
          7178 => x"81",
          7179 => x"51",
          7180 => x"9f",
          7181 => x"72",
          7182 => x"81",
          7183 => x"70",
          7184 => x"72",
          7185 => x"32",
          7186 => x"72",
          7187 => x"73",
          7188 => x"53",
          7189 => x"70",
          7190 => x"38",
          7191 => x"19",
          7192 => x"75",
          7193 => x"38",
          7194 => x"83",
          7195 => x"74",
          7196 => x"59",
          7197 => x"39",
          7198 => x"33",
          7199 => x"d5",
          7200 => x"3d",
          7201 => x"3d",
          7202 => x"80",
          7203 => x"34",
          7204 => x"17",
          7205 => x"75",
          7206 => x"3f",
          7207 => x"d5",
          7208 => x"80",
          7209 => x"16",
          7210 => x"3f",
          7211 => x"08",
          7212 => x"06",
          7213 => x"73",
          7214 => x"2e",
          7215 => x"80",
          7216 => x"0b",
          7217 => x"56",
          7218 => x"e9",
          7219 => x"06",
          7220 => x"57",
          7221 => x"32",
          7222 => x"80",
          7223 => x"51",
          7224 => x"8a",
          7225 => x"e8",
          7226 => x"06",
          7227 => x"53",
          7228 => x"52",
          7229 => x"51",
          7230 => x"82",
          7231 => x"55",
          7232 => x"08",
          7233 => x"38",
          7234 => x"c7",
          7235 => x"8a",
          7236 => x"ed",
          7237 => x"e4",
          7238 => x"d5",
          7239 => x"2e",
          7240 => x"55",
          7241 => x"e4",
          7242 => x"0d",
          7243 => x"0d",
          7244 => x"05",
          7245 => x"33",
          7246 => x"75",
          7247 => x"fc",
          7248 => x"d5",
          7249 => x"8b",
          7250 => x"82",
          7251 => x"24",
          7252 => x"82",
          7253 => x"84",
          7254 => x"ac",
          7255 => x"55",
          7256 => x"73",
          7257 => x"b1",
          7258 => x"0c",
          7259 => x"06",
          7260 => x"57",
          7261 => x"ae",
          7262 => x"33",
          7263 => x"3f",
          7264 => x"08",
          7265 => x"70",
          7266 => x"55",
          7267 => x"76",
          7268 => x"83",
          7269 => x"2a",
          7270 => x"51",
          7271 => x"72",
          7272 => x"86",
          7273 => x"74",
          7274 => x"59",
          7275 => x"19",
          7276 => x"34",
          7277 => x"14",
          7278 => x"81",
          7279 => x"e4",
          7280 => x"06",
          7281 => x"54",
          7282 => x"72",
          7283 => x"76",
          7284 => x"38",
          7285 => x"70",
          7286 => x"53",
          7287 => x"86",
          7288 => x"70",
          7289 => x"5b",
          7290 => x"82",
          7291 => x"81",
          7292 => x"76",
          7293 => x"38",
          7294 => x"81",
          7295 => x"d5",
          7296 => x"53",
          7297 => x"81",
          7298 => x"3d",
          7299 => x"83",
          7300 => x"15",
          7301 => x"53",
          7302 => x"8d",
          7303 => x"15",
          7304 => x"3f",
          7305 => x"08",
          7306 => x"70",
          7307 => x"0c",
          7308 => x"16",
          7309 => x"80",
          7310 => x"77",
          7311 => x"d9",
          7312 => x"30",
          7313 => x"72",
          7314 => x"3d",
          7315 => x"05",
          7316 => x"53",
          7317 => x"59",
          7318 => x"83",
          7319 => x"2e",
          7320 => x"52",
          7321 => x"9e",
          7322 => x"e4",
          7323 => x"06",
          7324 => x"82",
          7325 => x"33",
          7326 => x"78",
          7327 => x"06",
          7328 => x"58",
          7329 => x"91",
          7330 => x"2e",
          7331 => x"16",
          7332 => x"56",
          7333 => x"c0",
          7334 => x"76",
          7335 => x"f9",
          7336 => x"76",
          7337 => x"f1",
          7338 => x"14",
          7339 => x"3f",
          7340 => x"08",
          7341 => x"06",
          7342 => x"80",
          7343 => x"06",
          7344 => x"80",
          7345 => x"c9",
          7346 => x"d5",
          7347 => x"ff",
          7348 => x"77",
          7349 => x"dc",
          7350 => x"f0",
          7351 => x"e4",
          7352 => x"a0",
          7353 => x"c8",
          7354 => x"15",
          7355 => x"14",
          7356 => x"70",
          7357 => x"51",
          7358 => x"56",
          7359 => x"84",
          7360 => x"81",
          7361 => x"71",
          7362 => x"16",
          7363 => x"53",
          7364 => x"23",
          7365 => x"8b",
          7366 => x"73",
          7367 => x"80",
          7368 => x"8d",
          7369 => x"39",
          7370 => x"51",
          7371 => x"82",
          7372 => x"53",
          7373 => x"08",
          7374 => x"72",
          7375 => x"8d",
          7376 => x"d5",
          7377 => x"14",
          7378 => x"3f",
          7379 => x"08",
          7380 => x"06",
          7381 => x"38",
          7382 => x"51",
          7383 => x"82",
          7384 => x"55",
          7385 => x"51",
          7386 => x"82",
          7387 => x"83",
          7388 => x"53",
          7389 => x"80",
          7390 => x"38",
          7391 => x"78",
          7392 => x"2a",
          7393 => x"78",
          7394 => x"8d",
          7395 => x"22",
          7396 => x"31",
          7397 => x"97",
          7398 => x"e4",
          7399 => x"d5",
          7400 => x"2e",
          7401 => x"82",
          7402 => x"80",
          7403 => x"f5",
          7404 => x"83",
          7405 => x"ff",
          7406 => x"38",
          7407 => x"9f",
          7408 => x"38",
          7409 => x"39",
          7410 => x"80",
          7411 => x"38",
          7412 => x"9c",
          7413 => x"a4",
          7414 => x"1c",
          7415 => x"0c",
          7416 => x"17",
          7417 => x"76",
          7418 => x"81",
          7419 => x"80",
          7420 => x"c7",
          7421 => x"d5",
          7422 => x"ff",
          7423 => x"8d",
          7424 => x"95",
          7425 => x"91",
          7426 => x"14",
          7427 => x"3f",
          7428 => x"08",
          7429 => x"74",
          7430 => x"a2",
          7431 => x"79",
          7432 => x"f5",
          7433 => x"ac",
          7434 => x"15",
          7435 => x"2e",
          7436 => x"10",
          7437 => x"2a",
          7438 => x"05",
          7439 => x"ff",
          7440 => x"53",
          7441 => x"a0",
          7442 => x"81",
          7443 => x"0b",
          7444 => x"ff",
          7445 => x"0c",
          7446 => x"84",
          7447 => x"83",
          7448 => x"06",
          7449 => x"80",
          7450 => x"c6",
          7451 => x"d5",
          7452 => x"ff",
          7453 => x"72",
          7454 => x"81",
          7455 => x"38",
          7456 => x"73",
          7457 => x"3f",
          7458 => x"08",
          7459 => x"82",
          7460 => x"84",
          7461 => x"b6",
          7462 => x"99",
          7463 => x"e4",
          7464 => x"ff",
          7465 => x"82",
          7466 => x"09",
          7467 => x"c8",
          7468 => x"51",
          7469 => x"82",
          7470 => x"84",
          7471 => x"d2",
          7472 => x"06",
          7473 => x"9c",
          7474 => x"80",
          7475 => x"e4",
          7476 => x"85",
          7477 => x"09",
          7478 => x"38",
          7479 => x"51",
          7480 => x"82",
          7481 => x"94",
          7482 => x"a4",
          7483 => x"dc",
          7484 => x"e4",
          7485 => x"0c",
          7486 => x"82",
          7487 => x"81",
          7488 => x"82",
          7489 => x"72",
          7490 => x"82",
          7491 => x"8c",
          7492 => x"0b",
          7493 => x"80",
          7494 => x"d5",
          7495 => x"3d",
          7496 => x"3d",
          7497 => x"89",
          7498 => x"2e",
          7499 => x"08",
          7500 => x"2e",
          7501 => x"33",
          7502 => x"2e",
          7503 => x"13",
          7504 => x"22",
          7505 => x"76",
          7506 => x"06",
          7507 => x"13",
          7508 => x"be",
          7509 => x"d5",
          7510 => x"06",
          7511 => x"38",
          7512 => x"54",
          7513 => x"80",
          7514 => x"71",
          7515 => x"82",
          7516 => x"87",
          7517 => x"fa",
          7518 => x"ab",
          7519 => x"58",
          7520 => x"05",
          7521 => x"9a",
          7522 => x"80",
          7523 => x"e4",
          7524 => x"38",
          7525 => x"08",
          7526 => x"ed",
          7527 => x"08",
          7528 => x"80",
          7529 => x"80",
          7530 => x"54",
          7531 => x"84",
          7532 => x"34",
          7533 => x"75",
          7534 => x"2e",
          7535 => x"53",
          7536 => x"53",
          7537 => x"f6",
          7538 => x"d5",
          7539 => x"73",
          7540 => x"0c",
          7541 => x"04",
          7542 => x"68",
          7543 => x"80",
          7544 => x"59",
          7545 => x"78",
          7546 => x"c8",
          7547 => x"06",
          7548 => x"3d",
          7549 => x"9a",
          7550 => x"52",
          7551 => x"3f",
          7552 => x"08",
          7553 => x"e4",
          7554 => x"38",
          7555 => x"52",
          7556 => x"52",
          7557 => x"3f",
          7558 => x"08",
          7559 => x"e4",
          7560 => x"02",
          7561 => x"33",
          7562 => x"55",
          7563 => x"25",
          7564 => x"55",
          7565 => x"54",
          7566 => x"81",
          7567 => x"80",
          7568 => x"74",
          7569 => x"81",
          7570 => x"75",
          7571 => x"3f",
          7572 => x"08",
          7573 => x"02",
          7574 => x"91",
          7575 => x"81",
          7576 => x"82",
          7577 => x"06",
          7578 => x"80",
          7579 => x"88",
          7580 => x"39",
          7581 => x"58",
          7582 => x"38",
          7583 => x"70",
          7584 => x"54",
          7585 => x"81",
          7586 => x"52",
          7587 => x"ed",
          7588 => x"e4",
          7589 => x"88",
          7590 => x"62",
          7591 => x"c2",
          7592 => x"54",
          7593 => x"15",
          7594 => x"62",
          7595 => x"d7",
          7596 => x"52",
          7597 => x"51",
          7598 => x"7a",
          7599 => x"83",
          7600 => x"80",
          7601 => x"38",
          7602 => x"08",
          7603 => x"53",
          7604 => x"3d",
          7605 => x"cc",
          7606 => x"d5",
          7607 => x"82",
          7608 => x"82",
          7609 => x"39",
          7610 => x"38",
          7611 => x"33",
          7612 => x"70",
          7613 => x"55",
          7614 => x"2e",
          7615 => x"55",
          7616 => x"77",
          7617 => x"81",
          7618 => x"73",
          7619 => x"38",
          7620 => x"54",
          7621 => x"a0",
          7622 => x"82",
          7623 => x"52",
          7624 => x"eb",
          7625 => x"e4",
          7626 => x"18",
          7627 => x"55",
          7628 => x"e4",
          7629 => x"38",
          7630 => x"70",
          7631 => x"54",
          7632 => x"86",
          7633 => x"c0",
          7634 => x"b4",
          7635 => x"1b",
          7636 => x"1b",
          7637 => x"70",
          7638 => x"a1",
          7639 => x"e4",
          7640 => x"e4",
          7641 => x"0c",
          7642 => x"52",
          7643 => x"3f",
          7644 => x"08",
          7645 => x"08",
          7646 => x"77",
          7647 => x"86",
          7648 => x"1a",
          7649 => x"1a",
          7650 => x"91",
          7651 => x"0b",
          7652 => x"80",
          7653 => x"0c",
          7654 => x"70",
          7655 => x"54",
          7656 => x"81",
          7657 => x"d5",
          7658 => x"2e",
          7659 => x"82",
          7660 => x"94",
          7661 => x"17",
          7662 => x"2b",
          7663 => x"57",
          7664 => x"52",
          7665 => x"e7",
          7666 => x"e4",
          7667 => x"d5",
          7668 => x"26",
          7669 => x"55",
          7670 => x"08",
          7671 => x"81",
          7672 => x"79",
          7673 => x"31",
          7674 => x"70",
          7675 => x"25",
          7676 => x"76",
          7677 => x"81",
          7678 => x"55",
          7679 => x"38",
          7680 => x"0c",
          7681 => x"75",
          7682 => x"54",
          7683 => x"a2",
          7684 => x"7a",
          7685 => x"3f",
          7686 => x"08",
          7687 => x"55",
          7688 => x"89",
          7689 => x"e4",
          7690 => x"1a",
          7691 => x"80",
          7692 => x"54",
          7693 => x"e4",
          7694 => x"0d",
          7695 => x"0d",
          7696 => x"64",
          7697 => x"59",
          7698 => x"90",
          7699 => x"52",
          7700 => x"ce",
          7701 => x"e4",
          7702 => x"d5",
          7703 => x"38",
          7704 => x"55",
          7705 => x"86",
          7706 => x"82",
          7707 => x"19",
          7708 => x"55",
          7709 => x"80",
          7710 => x"38",
          7711 => x"0b",
          7712 => x"82",
          7713 => x"39",
          7714 => x"1a",
          7715 => x"82",
          7716 => x"19",
          7717 => x"08",
          7718 => x"7c",
          7719 => x"74",
          7720 => x"2e",
          7721 => x"94",
          7722 => x"83",
          7723 => x"56",
          7724 => x"38",
          7725 => x"22",
          7726 => x"89",
          7727 => x"55",
          7728 => x"75",
          7729 => x"19",
          7730 => x"39",
          7731 => x"52",
          7732 => x"db",
          7733 => x"e4",
          7734 => x"75",
          7735 => x"38",
          7736 => x"ff",
          7737 => x"98",
          7738 => x"19",
          7739 => x"51",
          7740 => x"82",
          7741 => x"80",
          7742 => x"38",
          7743 => x"08",
          7744 => x"2a",
          7745 => x"80",
          7746 => x"38",
          7747 => x"8a",
          7748 => x"5c",
          7749 => x"27",
          7750 => x"7a",
          7751 => x"54",
          7752 => x"52",
          7753 => x"51",
          7754 => x"3f",
          7755 => x"08",
          7756 => x"7e",
          7757 => x"56",
          7758 => x"2e",
          7759 => x"16",
          7760 => x"55",
          7761 => x"95",
          7762 => x"53",
          7763 => x"b4",
          7764 => x"31",
          7765 => x"05",
          7766 => x"e8",
          7767 => x"2b",
          7768 => x"76",
          7769 => x"94",
          7770 => x"ff",
          7771 => x"71",
          7772 => x"7b",
          7773 => x"38",
          7774 => x"19",
          7775 => x"51",
          7776 => x"82",
          7777 => x"fd",
          7778 => x"53",
          7779 => x"83",
          7780 => x"b8",
          7781 => x"51",
          7782 => x"3f",
          7783 => x"7e",
          7784 => x"0c",
          7785 => x"1b",
          7786 => x"1c",
          7787 => x"fd",
          7788 => x"56",
          7789 => x"e4",
          7790 => x"0d",
          7791 => x"0d",
          7792 => x"64",
          7793 => x"58",
          7794 => x"90",
          7795 => x"52",
          7796 => x"ce",
          7797 => x"e4",
          7798 => x"d5",
          7799 => x"38",
          7800 => x"55",
          7801 => x"86",
          7802 => x"83",
          7803 => x"18",
          7804 => x"2a",
          7805 => x"51",
          7806 => x"56",
          7807 => x"83",
          7808 => x"39",
          7809 => x"19",
          7810 => x"83",
          7811 => x"0b",
          7812 => x"81",
          7813 => x"39",
          7814 => x"7c",
          7815 => x"74",
          7816 => x"38",
          7817 => x"7b",
          7818 => x"f3",
          7819 => x"08",
          7820 => x"06",
          7821 => x"82",
          7822 => x"8a",
          7823 => x"05",
          7824 => x"06",
          7825 => x"bf",
          7826 => x"38",
          7827 => x"55",
          7828 => x"7a",
          7829 => x"98",
          7830 => x"77",
          7831 => x"3f",
          7832 => x"08",
          7833 => x"e4",
          7834 => x"82",
          7835 => x"81",
          7836 => x"38",
          7837 => x"ff",
          7838 => x"98",
          7839 => x"18",
          7840 => x"74",
          7841 => x"7e",
          7842 => x"08",
          7843 => x"2e",
          7844 => x"8e",
          7845 => x"ff",
          7846 => x"82",
          7847 => x"fe",
          7848 => x"18",
          7849 => x"51",
          7850 => x"3f",
          7851 => x"08",
          7852 => x"d0",
          7853 => x"e4",
          7854 => x"89",
          7855 => x"78",
          7856 => x"d7",
          7857 => x"7f",
          7858 => x"58",
          7859 => x"75",
          7860 => x"75",
          7861 => x"78",
          7862 => x"7c",
          7863 => x"33",
          7864 => x"c2",
          7865 => x"e4",
          7866 => x"38",
          7867 => x"08",
          7868 => x"56",
          7869 => x"9c",
          7870 => x"53",
          7871 => x"77",
          7872 => x"7d",
          7873 => x"16",
          7874 => x"b8",
          7875 => x"80",
          7876 => x"34",
          7877 => x"56",
          7878 => x"8c",
          7879 => x"19",
          7880 => x"38",
          7881 => x"bb",
          7882 => x"d5",
          7883 => x"de",
          7884 => x"b4",
          7885 => x"76",
          7886 => x"94",
          7887 => x"ff",
          7888 => x"71",
          7889 => x"7b",
          7890 => x"38",
          7891 => x"18",
          7892 => x"51",
          7893 => x"3f",
          7894 => x"08",
          7895 => x"75",
          7896 => x"94",
          7897 => x"ff",
          7898 => x"05",
          7899 => x"d4",
          7900 => x"81",
          7901 => x"34",
          7902 => x"7e",
          7903 => x"0c",
          7904 => x"1a",
          7905 => x"94",
          7906 => x"1b",
          7907 => x"5e",
          7908 => x"27",
          7909 => x"55",
          7910 => x"0c",
          7911 => x"90",
          7912 => x"c0",
          7913 => x"90",
          7914 => x"56",
          7915 => x"e4",
          7916 => x"0d",
          7917 => x"0d",
          7918 => x"fc",
          7919 => x"52",
          7920 => x"3f",
          7921 => x"08",
          7922 => x"e4",
          7923 => x"38",
          7924 => x"70",
          7925 => x"81",
          7926 => x"55",
          7927 => x"80",
          7928 => x"16",
          7929 => x"51",
          7930 => x"3f",
          7931 => x"08",
          7932 => x"e4",
          7933 => x"38",
          7934 => x"8b",
          7935 => x"07",
          7936 => x"8b",
          7937 => x"16",
          7938 => x"52",
          7939 => x"cc",
          7940 => x"16",
          7941 => x"15",
          7942 => x"f9",
          7943 => x"b2",
          7944 => x"15",
          7945 => x"ed",
          7946 => x"92",
          7947 => x"b7",
          7948 => x"54",
          7949 => x"15",
          7950 => x"ff",
          7951 => x"82",
          7952 => x"90",
          7953 => x"bf",
          7954 => x"73",
          7955 => x"76",
          7956 => x"0c",
          7957 => x"04",
          7958 => x"76",
          7959 => x"fe",
          7960 => x"d5",
          7961 => x"82",
          7962 => x"9c",
          7963 => x"fc",
          7964 => x"51",
          7965 => x"82",
          7966 => x"53",
          7967 => x"08",
          7968 => x"d5",
          7969 => x"0c",
          7970 => x"e4",
          7971 => x"0d",
          7972 => x"0d",
          7973 => x"e6",
          7974 => x"52",
          7975 => x"d5",
          7976 => x"8b",
          7977 => x"e4",
          7978 => x"c0",
          7979 => x"71",
          7980 => x"0c",
          7981 => x"04",
          7982 => x"80",
          7983 => x"cc",
          7984 => x"3d",
          7985 => x"3f",
          7986 => x"08",
          7987 => x"e4",
          7988 => x"38",
          7989 => x"52",
          7990 => x"05",
          7991 => x"3f",
          7992 => x"08",
          7993 => x"e4",
          7994 => x"02",
          7995 => x"33",
          7996 => x"55",
          7997 => x"25",
          7998 => x"7a",
          7999 => x"54",
          8000 => x"a2",
          8001 => x"84",
          8002 => x"06",
          8003 => x"73",
          8004 => x"38",
          8005 => x"70",
          8006 => x"e1",
          8007 => x"e4",
          8008 => x"0c",
          8009 => x"d5",
          8010 => x"2e",
          8011 => x"83",
          8012 => x"74",
          8013 => x"0c",
          8014 => x"04",
          8015 => x"0d",
          8016 => x"08",
          8017 => x"08",
          8018 => x"7a",
          8019 => x"80",
          8020 => x"b4",
          8021 => x"e0",
          8022 => x"d1",
          8023 => x"e4",
          8024 => x"d5",
          8025 => x"a1",
          8026 => x"d4",
          8027 => x"7c",
          8028 => x"80",
          8029 => x"55",
          8030 => x"3d",
          8031 => x"80",
          8032 => x"38",
          8033 => x"d3",
          8034 => x"55",
          8035 => x"82",
          8036 => x"57",
          8037 => x"08",
          8038 => x"80",
          8039 => x"52",
          8040 => x"b7",
          8041 => x"d5",
          8042 => x"82",
          8043 => x"82",
          8044 => x"da",
          8045 => x"7b",
          8046 => x"3f",
          8047 => x"08",
          8048 => x"0c",
          8049 => x"51",
          8050 => x"82",
          8051 => x"57",
          8052 => x"08",
          8053 => x"80",
          8054 => x"c9",
          8055 => x"d5",
          8056 => x"82",
          8057 => x"a7",
          8058 => x"3d",
          8059 => x"51",
          8060 => x"73",
          8061 => x"08",
          8062 => x"76",
          8063 => x"c4",
          8064 => x"d5",
          8065 => x"82",
          8066 => x"80",
          8067 => x"76",
          8068 => x"81",
          8069 => x"82",
          8070 => x"39",
          8071 => x"38",
          8072 => x"fd",
          8073 => x"74",
          8074 => x"3f",
          8075 => x"78",
          8076 => x"33",
          8077 => x"56",
          8078 => x"92",
          8079 => x"c6",
          8080 => x"16",
          8081 => x"33",
          8082 => x"73",
          8083 => x"16",
          8084 => x"26",
          8085 => x"75",
          8086 => x"38",
          8087 => x"05",
          8088 => x"80",
          8089 => x"11",
          8090 => x"18",
          8091 => x"58",
          8092 => x"34",
          8093 => x"ff",
          8094 => x"3d",
          8095 => x"58",
          8096 => x"fd",
          8097 => x"7b",
          8098 => x"06",
          8099 => x"18",
          8100 => x"08",
          8101 => x"af",
          8102 => x"0b",
          8103 => x"33",
          8104 => x"82",
          8105 => x"70",
          8106 => x"52",
          8107 => x"56",
          8108 => x"8d",
          8109 => x"70",
          8110 => x"51",
          8111 => x"f5",
          8112 => x"54",
          8113 => x"a7",
          8114 => x"74",
          8115 => x"38",
          8116 => x"73",
          8117 => x"81",
          8118 => x"81",
          8119 => x"39",
          8120 => x"81",
          8121 => x"74",
          8122 => x"81",
          8123 => x"91",
          8124 => x"80",
          8125 => x"18",
          8126 => x"54",
          8127 => x"70",
          8128 => x"34",
          8129 => x"eb",
          8130 => x"34",
          8131 => x"e4",
          8132 => x"3d",
          8133 => x"3d",
          8134 => x"8d",
          8135 => x"54",
          8136 => x"55",
          8137 => x"82",
          8138 => x"53",
          8139 => x"08",
          8140 => x"91",
          8141 => x"72",
          8142 => x"8c",
          8143 => x"73",
          8144 => x"38",
          8145 => x"70",
          8146 => x"81",
          8147 => x"57",
          8148 => x"73",
          8149 => x"08",
          8150 => x"94",
          8151 => x"75",
          8152 => x"9b",
          8153 => x"11",
          8154 => x"2b",
          8155 => x"73",
          8156 => x"38",
          8157 => x"16",
          8158 => x"b3",
          8159 => x"e4",
          8160 => x"78",
          8161 => x"55",
          8162 => x"a3",
          8163 => x"e4",
          8164 => x"96",
          8165 => x"70",
          8166 => x"94",
          8167 => x"71",
          8168 => x"08",
          8169 => x"53",
          8170 => x"15",
          8171 => x"a7",
          8172 => x"74",
          8173 => x"d3",
          8174 => x"e4",
          8175 => x"d5",
          8176 => x"2e",
          8177 => x"82",
          8178 => x"ff",
          8179 => x"38",
          8180 => x"08",
          8181 => x"73",
          8182 => x"73",
          8183 => x"9f",
          8184 => x"27",
          8185 => x"75",
          8186 => x"16",
          8187 => x"17",
          8188 => x"33",
          8189 => x"70",
          8190 => x"55",
          8191 => x"80",
          8192 => x"73",
          8193 => x"ff",
          8194 => x"82",
          8195 => x"54",
          8196 => x"08",
          8197 => x"d5",
          8198 => x"a8",
          8199 => x"74",
          8200 => x"8b",
          8201 => x"e4",
          8202 => x"ff",
          8203 => x"81",
          8204 => x"38",
          8205 => x"9c",
          8206 => x"a7",
          8207 => x"16",
          8208 => x"39",
          8209 => x"16",
          8210 => x"75",
          8211 => x"53",
          8212 => x"ab",
          8213 => x"79",
          8214 => x"a9",
          8215 => x"e4",
          8216 => x"82",
          8217 => x"34",
          8218 => x"c4",
          8219 => x"91",
          8220 => x"53",
          8221 => x"89",
          8222 => x"e4",
          8223 => x"94",
          8224 => x"8c",
          8225 => x"27",
          8226 => x"8c",
          8227 => x"15",
          8228 => x"07",
          8229 => x"16",
          8230 => x"ff",
          8231 => x"80",
          8232 => x"77",
          8233 => x"2e",
          8234 => x"9c",
          8235 => x"53",
          8236 => x"e4",
          8237 => x"0d",
          8238 => x"0d",
          8239 => x"54",
          8240 => x"81",
          8241 => x"53",
          8242 => x"05",
          8243 => x"84",
          8244 => x"d9",
          8245 => x"e4",
          8246 => x"d5",
          8247 => x"eb",
          8248 => x"0c",
          8249 => x"51",
          8250 => x"82",
          8251 => x"55",
          8252 => x"08",
          8253 => x"ab",
          8254 => x"98",
          8255 => x"80",
          8256 => x"38",
          8257 => x"70",
          8258 => x"81",
          8259 => x"57",
          8260 => x"ae",
          8261 => x"08",
          8262 => x"c1",
          8263 => x"d5",
          8264 => x"17",
          8265 => x"86",
          8266 => x"17",
          8267 => x"75",
          8268 => x"ea",
          8269 => x"e4",
          8270 => x"84",
          8271 => x"06",
          8272 => x"55",
          8273 => x"80",
          8274 => x"80",
          8275 => x"54",
          8276 => x"e4",
          8277 => x"0d",
          8278 => x"0d",
          8279 => x"fc",
          8280 => x"52",
          8281 => x"3f",
          8282 => x"08",
          8283 => x"d5",
          8284 => x"0c",
          8285 => x"04",
          8286 => x"77",
          8287 => x"fc",
          8288 => x"53",
          8289 => x"9a",
          8290 => x"e4",
          8291 => x"d5",
          8292 => x"e1",
          8293 => x"38",
          8294 => x"08",
          8295 => x"ff",
          8296 => x"82",
          8297 => x"53",
          8298 => x"82",
          8299 => x"52",
          8300 => x"df",
          8301 => x"e4",
          8302 => x"d5",
          8303 => x"2e",
          8304 => x"85",
          8305 => x"87",
          8306 => x"e4",
          8307 => x"74",
          8308 => x"ce",
          8309 => x"52",
          8310 => x"bd",
          8311 => x"d5",
          8312 => x"32",
          8313 => x"72",
          8314 => x"70",
          8315 => x"08",
          8316 => x"54",
          8317 => x"d5",
          8318 => x"3d",
          8319 => x"3d",
          8320 => x"80",
          8321 => x"70",
          8322 => x"52",
          8323 => x"3f",
          8324 => x"08",
          8325 => x"e4",
          8326 => x"65",
          8327 => x"d2",
          8328 => x"d5",
          8329 => x"82",
          8330 => x"a0",
          8331 => x"cb",
          8332 => x"98",
          8333 => x"73",
          8334 => x"38",
          8335 => x"39",
          8336 => x"88",
          8337 => x"75",
          8338 => x"3f",
          8339 => x"e4",
          8340 => x"0d",
          8341 => x"0d",
          8342 => x"5c",
          8343 => x"3d",
          8344 => x"93",
          8345 => x"c5",
          8346 => x"e4",
          8347 => x"d5",
          8348 => x"82",
          8349 => x"0c",
          8350 => x"11",
          8351 => x"94",
          8352 => x"56",
          8353 => x"74",
          8354 => x"75",
          8355 => x"e6",
          8356 => x"81",
          8357 => x"5b",
          8358 => x"82",
          8359 => x"75",
          8360 => x"73",
          8361 => x"81",
          8362 => x"38",
          8363 => x"57",
          8364 => x"3d",
          8365 => x"ff",
          8366 => x"82",
          8367 => x"ff",
          8368 => x"82",
          8369 => x"81",
          8370 => x"82",
          8371 => x"30",
          8372 => x"e4",
          8373 => x"25",
          8374 => x"19",
          8375 => x"5a",
          8376 => x"08",
          8377 => x"38",
          8378 => x"a8",
          8379 => x"d5",
          8380 => x"58",
          8381 => x"77",
          8382 => x"7d",
          8383 => x"ad",
          8384 => x"d5",
          8385 => x"82",
          8386 => x"80",
          8387 => x"70",
          8388 => x"ff",
          8389 => x"56",
          8390 => x"2e",
          8391 => x"9e",
          8392 => x"51",
          8393 => x"3f",
          8394 => x"08",
          8395 => x"06",
          8396 => x"80",
          8397 => x"19",
          8398 => x"54",
          8399 => x"14",
          8400 => x"88",
          8401 => x"e4",
          8402 => x"06",
          8403 => x"80",
          8404 => x"19",
          8405 => x"54",
          8406 => x"06",
          8407 => x"79",
          8408 => x"78",
          8409 => x"79",
          8410 => x"84",
          8411 => x"07",
          8412 => x"84",
          8413 => x"82",
          8414 => x"92",
          8415 => x"f9",
          8416 => x"8a",
          8417 => x"53",
          8418 => x"e3",
          8419 => x"d5",
          8420 => x"82",
          8421 => x"81",
          8422 => x"17",
          8423 => x"81",
          8424 => x"17",
          8425 => x"2a",
          8426 => x"51",
          8427 => x"55",
          8428 => x"81",
          8429 => x"17",
          8430 => x"8c",
          8431 => x"81",
          8432 => x"9c",
          8433 => x"e4",
          8434 => x"17",
          8435 => x"51",
          8436 => x"3f",
          8437 => x"08",
          8438 => x"0c",
          8439 => x"39",
          8440 => x"52",
          8441 => x"ad",
          8442 => x"d5",
          8443 => x"2e",
          8444 => x"83",
          8445 => x"82",
          8446 => x"81",
          8447 => x"06",
          8448 => x"56",
          8449 => x"a1",
          8450 => x"82",
          8451 => x"9c",
          8452 => x"95",
          8453 => x"08",
          8454 => x"e4",
          8455 => x"51",
          8456 => x"3f",
          8457 => x"08",
          8458 => x"08",
          8459 => x"90",
          8460 => x"c0",
          8461 => x"90",
          8462 => x"80",
          8463 => x"75",
          8464 => x"75",
          8465 => x"d5",
          8466 => x"3d",
          8467 => x"3d",
          8468 => x"a2",
          8469 => x"05",
          8470 => x"51",
          8471 => x"82",
          8472 => x"55",
          8473 => x"08",
          8474 => x"78",
          8475 => x"08",
          8476 => x"70",
          8477 => x"cf",
          8478 => x"e4",
          8479 => x"d5",
          8480 => x"df",
          8481 => x"ff",
          8482 => x"85",
          8483 => x"06",
          8484 => x"86",
          8485 => x"cb",
          8486 => x"2b",
          8487 => x"24",
          8488 => x"02",
          8489 => x"33",
          8490 => x"58",
          8491 => x"76",
          8492 => x"6c",
          8493 => x"ff",
          8494 => x"82",
          8495 => x"74",
          8496 => x"81",
          8497 => x"56",
          8498 => x"80",
          8499 => x"54",
          8500 => x"08",
          8501 => x"2e",
          8502 => x"73",
          8503 => x"e4",
          8504 => x"52",
          8505 => x"52",
          8506 => x"b2",
          8507 => x"e4",
          8508 => x"d5",
          8509 => x"eb",
          8510 => x"e4",
          8511 => x"51",
          8512 => x"3f",
          8513 => x"08",
          8514 => x"e4",
          8515 => x"87",
          8516 => x"39",
          8517 => x"08",
          8518 => x"38",
          8519 => x"08",
          8520 => x"77",
          8521 => x"3f",
          8522 => x"08",
          8523 => x"08",
          8524 => x"d5",
          8525 => x"80",
          8526 => x"55",
          8527 => x"95",
          8528 => x"2e",
          8529 => x"53",
          8530 => x"51",
          8531 => x"3f",
          8532 => x"08",
          8533 => x"38",
          8534 => x"a8",
          8535 => x"d5",
          8536 => x"74",
          8537 => x"0c",
          8538 => x"04",
          8539 => x"82",
          8540 => x"ff",
          8541 => x"9b",
          8542 => x"b1",
          8543 => x"e4",
          8544 => x"d5",
          8545 => x"b7",
          8546 => x"6a",
          8547 => x"70",
          8548 => x"b3",
          8549 => x"e4",
          8550 => x"d5",
          8551 => x"38",
          8552 => x"9b",
          8553 => x"e4",
          8554 => x"09",
          8555 => x"8f",
          8556 => x"df",
          8557 => x"85",
          8558 => x"51",
          8559 => x"74",
          8560 => x"78",
          8561 => x"8a",
          8562 => x"57",
          8563 => x"3f",
          8564 => x"08",
          8565 => x"82",
          8566 => x"83",
          8567 => x"82",
          8568 => x"81",
          8569 => x"06",
          8570 => x"54",
          8571 => x"08",
          8572 => x"81",
          8573 => x"81",
          8574 => x"39",
          8575 => x"38",
          8576 => x"08",
          8577 => x"ff",
          8578 => x"82",
          8579 => x"54",
          8580 => x"08",
          8581 => x"8b",
          8582 => x"b8",
          8583 => x"a4",
          8584 => x"54",
          8585 => x"15",
          8586 => x"90",
          8587 => x"15",
          8588 => x"b2",
          8589 => x"ce",
          8590 => x"a3",
          8591 => x"53",
          8592 => x"53",
          8593 => x"ee",
          8594 => x"78",
          8595 => x"80",
          8596 => x"ff",
          8597 => x"78",
          8598 => x"80",
          8599 => x"7f",
          8600 => x"d8",
          8601 => x"ff",
          8602 => x"78",
          8603 => x"83",
          8604 => x"51",
          8605 => x"3f",
          8606 => x"08",
          8607 => x"e4",
          8608 => x"82",
          8609 => x"52",
          8610 => x"51",
          8611 => x"3f",
          8612 => x"52",
          8613 => x"b7",
          8614 => x"54",
          8615 => x"15",
          8616 => x"81",
          8617 => x"34",
          8618 => x"a6",
          8619 => x"d5",
          8620 => x"8b",
          8621 => x"75",
          8622 => x"ff",
          8623 => x"73",
          8624 => x"0c",
          8625 => x"04",
          8626 => x"ab",
          8627 => x"51",
          8628 => x"82",
          8629 => x"fe",
          8630 => x"ab",
          8631 => x"cd",
          8632 => x"e4",
          8633 => x"d5",
          8634 => x"d8",
          8635 => x"ab",
          8636 => x"9e",
          8637 => x"58",
          8638 => x"82",
          8639 => x"55",
          8640 => x"08",
          8641 => x"02",
          8642 => x"33",
          8643 => x"54",
          8644 => x"82",
          8645 => x"53",
          8646 => x"52",
          8647 => x"80",
          8648 => x"a2",
          8649 => x"53",
          8650 => x"3d",
          8651 => x"ff",
          8652 => x"ac",
          8653 => x"73",
          8654 => x"3f",
          8655 => x"08",
          8656 => x"e4",
          8657 => x"63",
          8658 => x"2e",
          8659 => x"88",
          8660 => x"3d",
          8661 => x"38",
          8662 => x"e8",
          8663 => x"e4",
          8664 => x"09",
          8665 => x"bb",
          8666 => x"ff",
          8667 => x"82",
          8668 => x"55",
          8669 => x"08",
          8670 => x"68",
          8671 => x"aa",
          8672 => x"05",
          8673 => x"51",
          8674 => x"3f",
          8675 => x"33",
          8676 => x"8b",
          8677 => x"84",
          8678 => x"06",
          8679 => x"73",
          8680 => x"a0",
          8681 => x"8b",
          8682 => x"54",
          8683 => x"15",
          8684 => x"33",
          8685 => x"70",
          8686 => x"55",
          8687 => x"2e",
          8688 => x"6f",
          8689 => x"e1",
          8690 => x"78",
          8691 => x"ad",
          8692 => x"e4",
          8693 => x"51",
          8694 => x"3f",
          8695 => x"d5",
          8696 => x"2e",
          8697 => x"82",
          8698 => x"52",
          8699 => x"a3",
          8700 => x"d5",
          8701 => x"80",
          8702 => x"58",
          8703 => x"e4",
          8704 => x"38",
          8705 => x"54",
          8706 => x"09",
          8707 => x"38",
          8708 => x"52",
          8709 => x"b4",
          8710 => x"54",
          8711 => x"15",
          8712 => x"82",
          8713 => x"9c",
          8714 => x"c1",
          8715 => x"d5",
          8716 => x"82",
          8717 => x"8c",
          8718 => x"ff",
          8719 => x"82",
          8720 => x"55",
          8721 => x"e4",
          8722 => x"0d",
          8723 => x"0d",
          8724 => x"05",
          8725 => x"05",
          8726 => x"33",
          8727 => x"53",
          8728 => x"05",
          8729 => x"51",
          8730 => x"82",
          8731 => x"55",
          8732 => x"08",
          8733 => x"78",
          8734 => x"96",
          8735 => x"51",
          8736 => x"82",
          8737 => x"55",
          8738 => x"08",
          8739 => x"80",
          8740 => x"81",
          8741 => x"86",
          8742 => x"38",
          8743 => x"61",
          8744 => x"12",
          8745 => x"7a",
          8746 => x"51",
          8747 => x"74",
          8748 => x"78",
          8749 => x"83",
          8750 => x"51",
          8751 => x"3f",
          8752 => x"08",
          8753 => x"d5",
          8754 => x"3d",
          8755 => x"3d",
          8756 => x"82",
          8757 => x"cc",
          8758 => x"3d",
          8759 => x"3f",
          8760 => x"08",
          8761 => x"e4",
          8762 => x"38",
          8763 => x"52",
          8764 => x"05",
          8765 => x"3f",
          8766 => x"08",
          8767 => x"e4",
          8768 => x"02",
          8769 => x"33",
          8770 => x"54",
          8771 => x"a6",
          8772 => x"22",
          8773 => x"71",
          8774 => x"53",
          8775 => x"51",
          8776 => x"3f",
          8777 => x"0b",
          8778 => x"76",
          8779 => x"a6",
          8780 => x"e4",
          8781 => x"82",
          8782 => x"94",
          8783 => x"e9",
          8784 => x"6c",
          8785 => x"53",
          8786 => x"05",
          8787 => x"51",
          8788 => x"82",
          8789 => x"82",
          8790 => x"30",
          8791 => x"e4",
          8792 => x"25",
          8793 => x"79",
          8794 => x"86",
          8795 => x"75",
          8796 => x"73",
          8797 => x"fa",
          8798 => x"80",
          8799 => x"8d",
          8800 => x"54",
          8801 => x"3f",
          8802 => x"08",
          8803 => x"e4",
          8804 => x"38",
          8805 => x"51",
          8806 => x"3f",
          8807 => x"08",
          8808 => x"e4",
          8809 => x"82",
          8810 => x"82",
          8811 => x"65",
          8812 => x"78",
          8813 => x"7b",
          8814 => x"55",
          8815 => x"34",
          8816 => x"8a",
          8817 => x"38",
          8818 => x"1a",
          8819 => x"34",
          8820 => x"9e",
          8821 => x"70",
          8822 => x"51",
          8823 => x"a0",
          8824 => x"8e",
          8825 => x"2e",
          8826 => x"86",
          8827 => x"34",
          8828 => x"30",
          8829 => x"80",
          8830 => x"7a",
          8831 => x"c1",
          8832 => x"2e",
          8833 => x"a4",
          8834 => x"51",
          8835 => x"3f",
          8836 => x"08",
          8837 => x"e4",
          8838 => x"7b",
          8839 => x"55",
          8840 => x"73",
          8841 => x"38",
          8842 => x"73",
          8843 => x"38",
          8844 => x"15",
          8845 => x"ff",
          8846 => x"82",
          8847 => x"7b",
          8848 => x"d5",
          8849 => x"3d",
          8850 => x"3d",
          8851 => x"9c",
          8852 => x"05",
          8853 => x"51",
          8854 => x"82",
          8855 => x"82",
          8856 => x"56",
          8857 => x"e4",
          8858 => x"38",
          8859 => x"52",
          8860 => x"52",
          8861 => x"ef",
          8862 => x"70",
          8863 => x"56",
          8864 => x"81",
          8865 => x"57",
          8866 => x"ff",
          8867 => x"82",
          8868 => x"83",
          8869 => x"80",
          8870 => x"d5",
          8871 => x"96",
          8872 => x"b5",
          8873 => x"e4",
          8874 => x"90",
          8875 => x"e4",
          8876 => x"ff",
          8877 => x"80",
          8878 => x"74",
          8879 => x"f4",
          8880 => x"ee",
          8881 => x"e4",
          8882 => x"81",
          8883 => x"88",
          8884 => x"26",
          8885 => x"39",
          8886 => x"86",
          8887 => x"81",
          8888 => x"ff",
          8889 => x"38",
          8890 => x"54",
          8891 => x"81",
          8892 => x"81",
          8893 => x"77",
          8894 => x"59",
          8895 => x"6d",
          8896 => x"55",
          8897 => x"26",
          8898 => x"8a",
          8899 => x"86",
          8900 => x"e5",
          8901 => x"38",
          8902 => x"99",
          8903 => x"05",
          8904 => x"70",
          8905 => x"73",
          8906 => x"81",
          8907 => x"ff",
          8908 => x"ed",
          8909 => x"80",
          8910 => x"90",
          8911 => x"55",
          8912 => x"3f",
          8913 => x"08",
          8914 => x"e4",
          8915 => x"38",
          8916 => x"51",
          8917 => x"3f",
          8918 => x"08",
          8919 => x"e4",
          8920 => x"75",
          8921 => x"66",
          8922 => x"34",
          8923 => x"82",
          8924 => x"84",
          8925 => x"06",
          8926 => x"80",
          8927 => x"2e",
          8928 => x"81",
          8929 => x"ff",
          8930 => x"82",
          8931 => x"54",
          8932 => x"08",
          8933 => x"53",
          8934 => x"08",
          8935 => x"ff",
          8936 => x"66",
          8937 => x"8b",
          8938 => x"53",
          8939 => x"51",
          8940 => x"3f",
          8941 => x"0b",
          8942 => x"78",
          8943 => x"96",
          8944 => x"e4",
          8945 => x"55",
          8946 => x"e4",
          8947 => x"0d",
          8948 => x"0d",
          8949 => x"88",
          8950 => x"05",
          8951 => x"fc",
          8952 => x"54",
          8953 => x"d2",
          8954 => x"d5",
          8955 => x"82",
          8956 => x"82",
          8957 => x"1a",
          8958 => x"82",
          8959 => x"80",
          8960 => x"8c",
          8961 => x"78",
          8962 => x"1a",
          8963 => x"2a",
          8964 => x"51",
          8965 => x"90",
          8966 => x"82",
          8967 => x"58",
          8968 => x"81",
          8969 => x"39",
          8970 => x"22",
          8971 => x"70",
          8972 => x"56",
          8973 => x"af",
          8974 => x"14",
          8975 => x"30",
          8976 => x"9f",
          8977 => x"e4",
          8978 => x"19",
          8979 => x"5a",
          8980 => x"81",
          8981 => x"38",
          8982 => x"77",
          8983 => x"82",
          8984 => x"56",
          8985 => x"74",
          8986 => x"ff",
          8987 => x"81",
          8988 => x"55",
          8989 => x"75",
          8990 => x"82",
          8991 => x"e4",
          8992 => x"ff",
          8993 => x"d5",
          8994 => x"2e",
          8995 => x"82",
          8996 => x"8e",
          8997 => x"56",
          8998 => x"09",
          8999 => x"38",
          9000 => x"59",
          9001 => x"77",
          9002 => x"06",
          9003 => x"87",
          9004 => x"39",
          9005 => x"ba",
          9006 => x"55",
          9007 => x"2e",
          9008 => x"15",
          9009 => x"2e",
          9010 => x"83",
          9011 => x"75",
          9012 => x"7e",
          9013 => x"d0",
          9014 => x"e4",
          9015 => x"d5",
          9016 => x"ce",
          9017 => x"16",
          9018 => x"56",
          9019 => x"38",
          9020 => x"19",
          9021 => x"90",
          9022 => x"7d",
          9023 => x"38",
          9024 => x"0c",
          9025 => x"0c",
          9026 => x"80",
          9027 => x"73",
          9028 => x"9c",
          9029 => x"05",
          9030 => x"57",
          9031 => x"26",
          9032 => x"7b",
          9033 => x"0c",
          9034 => x"81",
          9035 => x"84",
          9036 => x"54",
          9037 => x"e4",
          9038 => x"0d",
          9039 => x"0d",
          9040 => x"88",
          9041 => x"05",
          9042 => x"54",
          9043 => x"c4",
          9044 => x"56",
          9045 => x"d5",
          9046 => x"8d",
          9047 => x"d5",
          9048 => x"29",
          9049 => x"05",
          9050 => x"55",
          9051 => x"84",
          9052 => x"34",
          9053 => x"08",
          9054 => x"08",
          9055 => x"d8",
          9056 => x"d5",
          9057 => x"47",
          9058 => x"52",
          9059 => x"8e",
          9060 => x"d5",
          9061 => x"ff",
          9062 => x"06",
          9063 => x"56",
          9064 => x"38",
          9065 => x"70",
          9066 => x"55",
          9067 => x"8c",
          9068 => x"3d",
          9069 => x"83",
          9070 => x"ff",
          9071 => x"82",
          9072 => x"99",
          9073 => x"74",
          9074 => x"38",
          9075 => x"80",
          9076 => x"ff",
          9077 => x"55",
          9078 => x"83",
          9079 => x"78",
          9080 => x"38",
          9081 => x"26",
          9082 => x"81",
          9083 => x"8b",
          9084 => x"79",
          9085 => x"80",
          9086 => x"93",
          9087 => x"39",
          9088 => x"6f",
          9089 => x"89",
          9090 => x"49",
          9091 => x"83",
          9092 => x"61",
          9093 => x"25",
          9094 => x"55",
          9095 => x"8b",
          9096 => x"80",
          9097 => x"38",
          9098 => x"53",
          9099 => x"51",
          9100 => x"3f",
          9101 => x"d5",
          9102 => x"c1",
          9103 => x"1b",
          9104 => x"f1",
          9105 => x"e4",
          9106 => x"ff",
          9107 => x"56",
          9108 => x"d5",
          9109 => x"06",
          9110 => x"64",
          9111 => x"83",
          9112 => x"56",
          9113 => x"2e",
          9114 => x"83",
          9115 => x"ff",
          9116 => x"82",
          9117 => x"83",
          9118 => x"5f",
          9119 => x"3f",
          9120 => x"08",
          9121 => x"9a",
          9122 => x"53",
          9123 => x"51",
          9124 => x"3f",
          9125 => x"d5",
          9126 => x"e1",
          9127 => x"2a",
          9128 => x"82",
          9129 => x"41",
          9130 => x"83",
          9131 => x"67",
          9132 => x"7e",
          9133 => x"c5",
          9134 => x"31",
          9135 => x"80",
          9136 => x"8a",
          9137 => x"56",
          9138 => x"26",
          9139 => x"62",
          9140 => x"81",
          9141 => x"74",
          9142 => x"38",
          9143 => x"55",
          9144 => x"83",
          9145 => x"81",
          9146 => x"80",
          9147 => x"38",
          9148 => x"55",
          9149 => x"5e",
          9150 => x"8a",
          9151 => x"5a",
          9152 => x"09",
          9153 => x"e1",
          9154 => x"38",
          9155 => x"57",
          9156 => x"c9",
          9157 => x"5a",
          9158 => x"9d",
          9159 => x"26",
          9160 => x"c9",
          9161 => x"10",
          9162 => x"22",
          9163 => x"74",
          9164 => x"38",
          9165 => x"ee",
          9166 => x"67",
          9167 => x"ef",
          9168 => x"e4",
          9169 => x"84",
          9170 => x"89",
          9171 => x"a0",
          9172 => x"82",
          9173 => x"fc",
          9174 => x"56",
          9175 => x"f0",
          9176 => x"80",
          9177 => x"88",
          9178 => x"38",
          9179 => x"57",
          9180 => x"c9",
          9181 => x"5a",
          9182 => x"9d",
          9183 => x"26",
          9184 => x"c9",
          9185 => x"10",
          9186 => x"22",
          9187 => x"74",
          9188 => x"38",
          9189 => x"ee",
          9190 => x"67",
          9191 => x"8f",
          9192 => x"e4",
          9193 => x"05",
          9194 => x"e4",
          9195 => x"26",
          9196 => x"0b",
          9197 => x"08",
          9198 => x"e4",
          9199 => x"11",
          9200 => x"05",
          9201 => x"83",
          9202 => x"2a",
          9203 => x"a0",
          9204 => x"7d",
          9205 => x"6a",
          9206 => x"05",
          9207 => x"72",
          9208 => x"5c",
          9209 => x"59",
          9210 => x"2e",
          9211 => x"89",
          9212 => x"61",
          9213 => x"84",
          9214 => x"5d",
          9215 => x"18",
          9216 => x"69",
          9217 => x"74",
          9218 => x"e4",
          9219 => x"31",
          9220 => x"53",
          9221 => x"52",
          9222 => x"93",
          9223 => x"e4",
          9224 => x"83",
          9225 => x"06",
          9226 => x"d5",
          9227 => x"ff",
          9228 => x"dd",
          9229 => x"b8",
          9230 => x"2a",
          9231 => x"be",
          9232 => x"39",
          9233 => x"09",
          9234 => x"c5",
          9235 => x"f5",
          9236 => x"e4",
          9237 => x"38",
          9238 => x"79",
          9239 => x"80",
          9240 => x"38",
          9241 => x"96",
          9242 => x"06",
          9243 => x"2e",
          9244 => x"5e",
          9245 => x"82",
          9246 => x"9f",
          9247 => x"38",
          9248 => x"38",
          9249 => x"81",
          9250 => x"fc",
          9251 => x"e0",
          9252 => x"7d",
          9253 => x"81",
          9254 => x"7d",
          9255 => x"78",
          9256 => x"74",
          9257 => x"8e",
          9258 => x"d1",
          9259 => x"53",
          9260 => x"51",
          9261 => x"3f",
          9262 => x"c7",
          9263 => x"51",
          9264 => x"3f",
          9265 => x"8b",
          9266 => x"8e",
          9267 => x"8d",
          9268 => x"83",
          9269 => x"52",
          9270 => x"ff",
          9271 => x"81",
          9272 => x"34",
          9273 => x"70",
          9274 => x"2a",
          9275 => x"54",
          9276 => x"1b",
          9277 => x"ff",
          9278 => x"74",
          9279 => x"26",
          9280 => x"83",
          9281 => x"52",
          9282 => x"ff",
          9283 => x"8a",
          9284 => x"a0",
          9285 => x"8d",
          9286 => x"0b",
          9287 => x"bf",
          9288 => x"51",
          9289 => x"3f",
          9290 => x"9a",
          9291 => x"8d",
          9292 => x"52",
          9293 => x"ff",
          9294 => x"7d",
          9295 => x"81",
          9296 => x"38",
          9297 => x"0a",
          9298 => x"1b",
          9299 => x"c5",
          9300 => x"a4",
          9301 => x"8d",
          9302 => x"52",
          9303 => x"ff",
          9304 => x"81",
          9305 => x"51",
          9306 => x"3f",
          9307 => x"1b",
          9308 => x"83",
          9309 => x"0b",
          9310 => x"34",
          9311 => x"c2",
          9312 => x"53",
          9313 => x"52",
          9314 => x"51",
          9315 => x"88",
          9316 => x"a7",
          9317 => x"8c",
          9318 => x"83",
          9319 => x"52",
          9320 => x"ff",
          9321 => x"ff",
          9322 => x"1c",
          9323 => x"a6",
          9324 => x"53",
          9325 => x"52",
          9326 => x"ff",
          9327 => x"82",
          9328 => x"83",
          9329 => x"52",
          9330 => x"ab",
          9331 => x"7e",
          9332 => x"7f",
          9333 => x"ce",
          9334 => x"82",
          9335 => x"84",
          9336 => x"83",
          9337 => x"06",
          9338 => x"75",
          9339 => x"53",
          9340 => x"51",
          9341 => x"3f",
          9342 => x"80",
          9343 => x"ff",
          9344 => x"84",
          9345 => x"d2",
          9346 => x"ff",
          9347 => x"86",
          9348 => x"f2",
          9349 => x"1b",
          9350 => x"f9",
          9351 => x"52",
          9352 => x"51",
          9353 => x"3f",
          9354 => x"ec",
          9355 => x"8b",
          9356 => x"d4",
          9357 => x"51",
          9358 => x"3f",
          9359 => x"1f",
          9360 => x"7f",
          9361 => x"de",
          9362 => x"75",
          9363 => x"52",
          9364 => x"87",
          9365 => x"53",
          9366 => x"51",
          9367 => x"3f",
          9368 => x"58",
          9369 => x"09",
          9370 => x"38",
          9371 => x"51",
          9372 => x"3f",
          9373 => x"1b",
          9374 => x"99",
          9375 => x"52",
          9376 => x"91",
          9377 => x"ff",
          9378 => x"81",
          9379 => x"f8",
          9380 => x"7a",
          9381 => x"fd",
          9382 => x"61",
          9383 => x"26",
          9384 => x"57",
          9385 => x"53",
          9386 => x"51",
          9387 => x"3f",
          9388 => x"08",
          9389 => x"84",
          9390 => x"d5",
          9391 => x"7a",
          9392 => x"a3",
          9393 => x"75",
          9394 => x"56",
          9395 => x"81",
          9396 => x"80",
          9397 => x"38",
          9398 => x"83",
          9399 => x"65",
          9400 => x"74",
          9401 => x"38",
          9402 => x"54",
          9403 => x"52",
          9404 => x"86",
          9405 => x"d5",
          9406 => x"f8",
          9407 => x"75",
          9408 => x"56",
          9409 => x"8c",
          9410 => x"2e",
          9411 => x"57",
          9412 => x"ff",
          9413 => x"84",
          9414 => x"2e",
          9415 => x"57",
          9416 => x"b2",
          9417 => x"80",
          9418 => x"7f",
          9419 => x"8c",
          9420 => x"82",
          9421 => x"81",
          9422 => x"90",
          9423 => x"76",
          9424 => x"34",
          9425 => x"d5",
          9426 => x"7a",
          9427 => x"ff",
          9428 => x"81",
          9429 => x"83",
          9430 => x"58",
          9431 => x"38",
          9432 => x"77",
          9433 => x"ff",
          9434 => x"82",
          9435 => x"78",
          9436 => x"83",
          9437 => x"1b",
          9438 => x"34",
          9439 => x"16",
          9440 => x"82",
          9441 => x"83",
          9442 => x"84",
          9443 => x"1f",
          9444 => x"c1",
          9445 => x"fe",
          9446 => x"fe",
          9447 => x"34",
          9448 => x"08",
          9449 => x"07",
          9450 => x"16",
          9451 => x"e4",
          9452 => x"34",
          9453 => x"c6",
          9454 => x"88",
          9455 => x"52",
          9456 => x"51",
          9457 => x"3f",
          9458 => x"53",
          9459 => x"51",
          9460 => x"3f",
          9461 => x"d5",
          9462 => x"38",
          9463 => x"52",
          9464 => x"86",
          9465 => x"56",
          9466 => x"08",
          9467 => x"39",
          9468 => x"39",
          9469 => x"39",
          9470 => x"08",
          9471 => x"d5",
          9472 => x"3d",
          9473 => x"3d",
          9474 => x"5b",
          9475 => x"60",
          9476 => x"57",
          9477 => x"25",
          9478 => x"3d",
          9479 => x"55",
          9480 => x"15",
          9481 => x"c8",
          9482 => x"81",
          9483 => x"06",
          9484 => x"3d",
          9485 => x"8d",
          9486 => x"74",
          9487 => x"05",
          9488 => x"17",
          9489 => x"2e",
          9490 => x"c9",
          9491 => x"34",
          9492 => x"83",
          9493 => x"74",
          9494 => x"0c",
          9495 => x"04",
          9496 => x"7b",
          9497 => x"b3",
          9498 => x"57",
          9499 => x"09",
          9500 => x"38",
          9501 => x"51",
          9502 => x"17",
          9503 => x"76",
          9504 => x"88",
          9505 => x"17",
          9506 => x"59",
          9507 => x"81",
          9508 => x"76",
          9509 => x"8b",
          9510 => x"54",
          9511 => x"17",
          9512 => x"51",
          9513 => x"79",
          9514 => x"30",
          9515 => x"9f",
          9516 => x"53",
          9517 => x"75",
          9518 => x"81",
          9519 => x"0c",
          9520 => x"04",
          9521 => x"79",
          9522 => x"56",
          9523 => x"24",
          9524 => x"3d",
          9525 => x"74",
          9526 => x"52",
          9527 => x"c9",
          9528 => x"d5",
          9529 => x"38",
          9530 => x"78",
          9531 => x"06",
          9532 => x"16",
          9533 => x"39",
          9534 => x"82",
          9535 => x"89",
          9536 => x"fd",
          9537 => x"54",
          9538 => x"80",
          9539 => x"ff",
          9540 => x"76",
          9541 => x"3d",
          9542 => x"3d",
          9543 => x"e3",
          9544 => x"53",
          9545 => x"53",
          9546 => x"3f",
          9547 => x"51",
          9548 => x"72",
          9549 => x"3f",
          9550 => x"04",
          9551 => x"75",
          9552 => x"9a",
          9553 => x"53",
          9554 => x"80",
          9555 => x"38",
          9556 => x"ff",
          9557 => x"c3",
          9558 => x"ff",
          9559 => x"73",
          9560 => x"09",
          9561 => x"38",
          9562 => x"af",
          9563 => x"a8",
          9564 => x"71",
          9565 => x"81",
          9566 => x"ff",
          9567 => x"51",
          9568 => x"26",
          9569 => x"10",
          9570 => x"05",
          9571 => x"51",
          9572 => x"80",
          9573 => x"ff",
          9574 => x"71",
          9575 => x"0c",
          9576 => x"04",
          9577 => x"02",
          9578 => x"02",
          9579 => x"05",
          9580 => x"80",
          9581 => x"ff",
          9582 => x"70",
          9583 => x"71",
          9584 => x"09",
          9585 => x"38",
          9586 => x"26",
          9587 => x"10",
          9588 => x"05",
          9589 => x"51",
          9590 => x"e4",
          9591 => x"0d",
          9592 => x"0d",
          9593 => x"83",
          9594 => x"81",
          9595 => x"83",
          9596 => x"82",
          9597 => x"52",
          9598 => x"27",
          9599 => x"cf",
          9600 => x"70",
          9601 => x"22",
          9602 => x"80",
          9603 => x"26",
          9604 => x"55",
          9605 => x"38",
          9606 => x"05",
          9607 => x"88",
          9608 => x"ff",
          9609 => x"54",
          9610 => x"71",
          9611 => x"d7",
          9612 => x"26",
          9613 => x"73",
          9614 => x"ae",
          9615 => x"70",
          9616 => x"75",
          9617 => x"11",
          9618 => x"51",
          9619 => x"39",
          9620 => x"81",
          9621 => x"31",
          9622 => x"39",
          9623 => x"9f",
          9624 => x"51",
          9625 => x"12",
          9626 => x"e6",
          9627 => x"39",
          9628 => x"8b",
          9629 => x"12",
          9630 => x"c7",
          9631 => x"70",
          9632 => x"06",
          9633 => x"73",
          9634 => x"72",
          9635 => x"fe",
          9636 => x"51",
          9637 => x"e4",
          9638 => x"0d",
          9639 => x"ff",
          9640 => x"ff",
          9641 => x"00",
          9642 => x"ff",
          9643 => x"2c",
          9644 => x"2b",
          9645 => x"2b",
          9646 => x"2b",
          9647 => x"2b",
          9648 => x"2b",
          9649 => x"2b",
          9650 => x"2b",
          9651 => x"2c",
          9652 => x"2c",
          9653 => x"2c",
          9654 => x"2c",
          9655 => x"2c",
          9656 => x"2c",
          9657 => x"2c",
          9658 => x"2c",
          9659 => x"2c",
          9660 => x"2c",
          9661 => x"2c",
          9662 => x"2c",
          9663 => x"42",
          9664 => x"42",
          9665 => x"42",
          9666 => x"42",
          9667 => x"42",
          9668 => x"48",
          9669 => x"49",
          9670 => x"4a",
          9671 => x"4c",
          9672 => x"49",
          9673 => x"46",
          9674 => x"4b",
          9675 => x"4c",
          9676 => x"4b",
          9677 => x"4b",
          9678 => x"4b",
          9679 => x"49",
          9680 => x"46",
          9681 => x"4a",
          9682 => x"4a",
          9683 => x"4b",
          9684 => x"46",
          9685 => x"46",
          9686 => x"4b",
          9687 => x"4b",
          9688 => x"4c",
          9689 => x"4c",
          9690 => x"96",
          9691 => x"96",
          9692 => x"96",
          9693 => x"96",
          9694 => x"96",
          9695 => x"96",
          9696 => x"96",
          9697 => x"96",
          9698 => x"96",
          9699 => x"0e",
          9700 => x"17",
          9701 => x"17",
          9702 => x"0e",
          9703 => x"17",
          9704 => x"17",
          9705 => x"17",
          9706 => x"17",
          9707 => x"17",
          9708 => x"17",
          9709 => x"17",
          9710 => x"0e",
          9711 => x"17",
          9712 => x"0e",
          9713 => x"0e",
          9714 => x"17",
          9715 => x"17",
          9716 => x"17",
          9717 => x"17",
          9718 => x"17",
          9719 => x"17",
          9720 => x"17",
          9721 => x"17",
          9722 => x"17",
          9723 => x"17",
          9724 => x"17",
          9725 => x"17",
          9726 => x"17",
          9727 => x"17",
          9728 => x"17",
          9729 => x"17",
          9730 => x"17",
          9731 => x"17",
          9732 => x"17",
          9733 => x"17",
          9734 => x"17",
          9735 => x"17",
          9736 => x"17",
          9737 => x"17",
          9738 => x"17",
          9739 => x"17",
          9740 => x"17",
          9741 => x"17",
          9742 => x"17",
          9743 => x"17",
          9744 => x"17",
          9745 => x"17",
          9746 => x"17",
          9747 => x"17",
          9748 => x"17",
          9749 => x"17",
          9750 => x"0f",
          9751 => x"17",
          9752 => x"17",
          9753 => x"17",
          9754 => x"17",
          9755 => x"11",
          9756 => x"17",
          9757 => x"17",
          9758 => x"17",
          9759 => x"17",
          9760 => x"17",
          9761 => x"17",
          9762 => x"17",
          9763 => x"17",
          9764 => x"17",
          9765 => x"17",
          9766 => x"0e",
          9767 => x"10",
          9768 => x"0e",
          9769 => x"0e",
          9770 => x"0e",
          9771 => x"17",
          9772 => x"10",
          9773 => x"17",
          9774 => x"17",
          9775 => x"0e",
          9776 => x"17",
          9777 => x"17",
          9778 => x"10",
          9779 => x"10",
          9780 => x"17",
          9781 => x"17",
          9782 => x"0f",
          9783 => x"17",
          9784 => x"11",
          9785 => x"17",
          9786 => x"17",
          9787 => x"11",
          9788 => x"6e",
          9789 => x"00",
          9790 => x"6f",
          9791 => x"00",
          9792 => x"6e",
          9793 => x"00",
          9794 => x"6f",
          9795 => x"00",
          9796 => x"78",
          9797 => x"00",
          9798 => x"6c",
          9799 => x"00",
          9800 => x"6f",
          9801 => x"00",
          9802 => x"69",
          9803 => x"00",
          9804 => x"75",
          9805 => x"00",
          9806 => x"62",
          9807 => x"68",
          9808 => x"77",
          9809 => x"64",
          9810 => x"65",
          9811 => x"64",
          9812 => x"65",
          9813 => x"6c",
          9814 => x"00",
          9815 => x"70",
          9816 => x"73",
          9817 => x"74",
          9818 => x"73",
          9819 => x"00",
          9820 => x"66",
          9821 => x"00",
          9822 => x"73",
          9823 => x"00",
          9824 => x"61",
          9825 => x"00",
          9826 => x"61",
          9827 => x"00",
          9828 => x"6c",
          9829 => x"00",
          9830 => x"00",
          9831 => x"73",
          9832 => x"72",
          9833 => x"00",
          9834 => x"74",
          9835 => x"61",
          9836 => x"72",
          9837 => x"2e",
          9838 => x"73",
          9839 => x"6f",
          9840 => x"65",
          9841 => x"2e",
          9842 => x"20",
          9843 => x"65",
          9844 => x"75",
          9845 => x"00",
          9846 => x"20",
          9847 => x"68",
          9848 => x"75",
          9849 => x"00",
          9850 => x"76",
          9851 => x"64",
          9852 => x"6c",
          9853 => x"6d",
          9854 => x"00",
          9855 => x"63",
          9856 => x"20",
          9857 => x"69",
          9858 => x"00",
          9859 => x"6c",
          9860 => x"6c",
          9861 => x"64",
          9862 => x"78",
          9863 => x"73",
          9864 => x"00",
          9865 => x"6c",
          9866 => x"61",
          9867 => x"65",
          9868 => x"76",
          9869 => x"64",
          9870 => x"00",
          9871 => x"20",
          9872 => x"77",
          9873 => x"65",
          9874 => x"6f",
          9875 => x"74",
          9876 => x"00",
          9877 => x"69",
          9878 => x"6e",
          9879 => x"65",
          9880 => x"73",
          9881 => x"76",
          9882 => x"64",
          9883 => x"00",
          9884 => x"73",
          9885 => x"6f",
          9886 => x"6e",
          9887 => x"65",
          9888 => x"00",
          9889 => x"20",
          9890 => x"70",
          9891 => x"62",
          9892 => x"66",
          9893 => x"73",
          9894 => x"65",
          9895 => x"6f",
          9896 => x"20",
          9897 => x"64",
          9898 => x"2e",
          9899 => x"72",
          9900 => x"20",
          9901 => x"72",
          9902 => x"2e",
          9903 => x"6d",
          9904 => x"74",
          9905 => x"70",
          9906 => x"74",
          9907 => x"20",
          9908 => x"63",
          9909 => x"65",
          9910 => x"00",
          9911 => x"6c",
          9912 => x"73",
          9913 => x"63",
          9914 => x"2e",
          9915 => x"73",
          9916 => x"69",
          9917 => x"6e",
          9918 => x"65",
          9919 => x"79",
          9920 => x"00",
          9921 => x"6f",
          9922 => x"6e",
          9923 => x"70",
          9924 => x"66",
          9925 => x"73",
          9926 => x"00",
          9927 => x"72",
          9928 => x"74",
          9929 => x"20",
          9930 => x"6f",
          9931 => x"63",
          9932 => x"00",
          9933 => x"63",
          9934 => x"73",
          9935 => x"00",
          9936 => x"6b",
          9937 => x"6e",
          9938 => x"72",
          9939 => x"00",
          9940 => x"6c",
          9941 => x"79",
          9942 => x"20",
          9943 => x"61",
          9944 => x"6c",
          9945 => x"79",
          9946 => x"2f",
          9947 => x"2e",
          9948 => x"00",
          9949 => x"61",
          9950 => x"00",
          9951 => x"38",
          9952 => x"00",
          9953 => x"20",
          9954 => x"34",
          9955 => x"00",
          9956 => x"20",
          9957 => x"20",
          9958 => x"00",
          9959 => x"32",
          9960 => x"00",
          9961 => x"00",
          9962 => x"00",
          9963 => x"00",
          9964 => x"53",
          9965 => x"2a",
          9966 => x"20",
          9967 => x"00",
          9968 => x"2f",
          9969 => x"32",
          9970 => x"00",
          9971 => x"2e",
          9972 => x"00",
          9973 => x"50",
          9974 => x"72",
          9975 => x"25",
          9976 => x"29",
          9977 => x"20",
          9978 => x"2a",
          9979 => x"00",
          9980 => x"55",
          9981 => x"74",
          9982 => x"75",
          9983 => x"48",
          9984 => x"6c",
          9985 => x"00",
          9986 => x"6d",
          9987 => x"69",
          9988 => x"72",
          9989 => x"74",
          9990 => x"32",
          9991 => x"74",
          9992 => x"75",
          9993 => x"00",
          9994 => x"43",
          9995 => x"52",
          9996 => x"6e",
          9997 => x"72",
          9998 => x"00",
          9999 => x"43",
         10000 => x"57",
         10001 => x"6e",
         10002 => x"72",
         10003 => x"00",
         10004 => x"52",
         10005 => x"52",
         10006 => x"6e",
         10007 => x"72",
         10008 => x"00",
         10009 => x"52",
         10010 => x"54",
         10011 => x"6e",
         10012 => x"72",
         10013 => x"00",
         10014 => x"52",
         10015 => x"52",
         10016 => x"6e",
         10017 => x"72",
         10018 => x"00",
         10019 => x"52",
         10020 => x"54",
         10021 => x"6e",
         10022 => x"72",
         10023 => x"00",
         10024 => x"74",
         10025 => x"67",
         10026 => x"20",
         10027 => x"65",
         10028 => x"2e",
         10029 => x"61",
         10030 => x"6e",
         10031 => x"69",
         10032 => x"2e",
         10033 => x"00",
         10034 => x"74",
         10035 => x"65",
         10036 => x"61",
         10037 => x"00",
         10038 => x"53",
         10039 => x"75",
         10040 => x"74",
         10041 => x"00",
         10042 => x"69",
         10043 => x"20",
         10044 => x"69",
         10045 => x"69",
         10046 => x"73",
         10047 => x"64",
         10048 => x"72",
         10049 => x"2c",
         10050 => x"65",
         10051 => x"20",
         10052 => x"74",
         10053 => x"6e",
         10054 => x"6c",
         10055 => x"00",
         10056 => x"00",
         10057 => x"65",
         10058 => x"6e",
         10059 => x"2e",
         10060 => x"00",
         10061 => x"70",
         10062 => x"67",
         10063 => x"00",
         10064 => x"6d",
         10065 => x"69",
         10066 => x"2e",
         10067 => x"00",
         10068 => x"38",
         10069 => x"25",
         10070 => x"29",
         10071 => x"30",
         10072 => x"28",
         10073 => x"78",
         10074 => x"00",
         10075 => x"6d",
         10076 => x"65",
         10077 => x"79",
         10078 => x"6f",
         10079 => x"65",
         10080 => x"00",
         10081 => x"38",
         10082 => x"25",
         10083 => x"2d",
         10084 => x"3f",
         10085 => x"38",
         10086 => x"25",
         10087 => x"2d",
         10088 => x"38",
         10089 => x"25",
         10090 => x"58",
         10091 => x"00",
         10092 => x"65",
         10093 => x"69",
         10094 => x"63",
         10095 => x"20",
         10096 => x"30",
         10097 => x"20",
         10098 => x"0a",
         10099 => x"6c",
         10100 => x"67",
         10101 => x"64",
         10102 => x"20",
         10103 => x"6c",
         10104 => x"2e",
         10105 => x"00",
         10106 => x"6c",
         10107 => x"65",
         10108 => x"6e",
         10109 => x"63",
         10110 => x"20",
         10111 => x"29",
         10112 => x"00",
         10113 => x"73",
         10114 => x"74",
         10115 => x"20",
         10116 => x"6c",
         10117 => x"74",
         10118 => x"2e",
         10119 => x"00",
         10120 => x"6c",
         10121 => x"65",
         10122 => x"74",
         10123 => x"2e",
         10124 => x"00",
         10125 => x"55",
         10126 => x"6e",
         10127 => x"3a",
         10128 => x"5c",
         10129 => x"25",
         10130 => x"00",
         10131 => x"3a",
         10132 => x"5c",
         10133 => x"00",
         10134 => x"3a",
         10135 => x"00",
         10136 => x"64",
         10137 => x"6d",
         10138 => x"64",
         10139 => x"00",
         10140 => x"6d",
         10141 => x"20",
         10142 => x"61",
         10143 => x"65",
         10144 => x"63",
         10145 => x"6f",
         10146 => x"72",
         10147 => x"73",
         10148 => x"6f",
         10149 => x"6e",
         10150 => x"00",
         10151 => x"6e",
         10152 => x"67",
         10153 => x"00",
         10154 => x"61",
         10155 => x"6e",
         10156 => x"6e",
         10157 => x"72",
         10158 => x"73",
         10159 => x"00",
         10160 => x"2f",
         10161 => x"25",
         10162 => x"64",
         10163 => x"3a",
         10164 => x"25",
         10165 => x"0a",
         10166 => x"43",
         10167 => x"6e",
         10168 => x"75",
         10169 => x"69",
         10170 => x"00",
         10171 => x"66",
         10172 => x"20",
         10173 => x"20",
         10174 => x"66",
         10175 => x"00",
         10176 => x"44",
         10177 => x"63",
         10178 => x"69",
         10179 => x"65",
         10180 => x"74",
         10181 => x"00",
         10182 => x"20",
         10183 => x"20",
         10184 => x"41",
         10185 => x"28",
         10186 => x"58",
         10187 => x"38",
         10188 => x"0a",
         10189 => x"20",
         10190 => x"52",
         10191 => x"20",
         10192 => x"28",
         10193 => x"58",
         10194 => x"38",
         10195 => x"0a",
         10196 => x"20",
         10197 => x"53",
         10198 => x"52",
         10199 => x"28",
         10200 => x"58",
         10201 => x"38",
         10202 => x"0a",
         10203 => x"20",
         10204 => x"41",
         10205 => x"20",
         10206 => x"28",
         10207 => x"58",
         10208 => x"38",
         10209 => x"0a",
         10210 => x"20",
         10211 => x"4d",
         10212 => x"20",
         10213 => x"28",
         10214 => x"58",
         10215 => x"38",
         10216 => x"0a",
         10217 => x"20",
         10218 => x"20",
         10219 => x"44",
         10220 => x"28",
         10221 => x"69",
         10222 => x"20",
         10223 => x"32",
         10224 => x"0a",
         10225 => x"20",
         10226 => x"4d",
         10227 => x"20",
         10228 => x"28",
         10229 => x"65",
         10230 => x"20",
         10231 => x"32",
         10232 => x"0a",
         10233 => x"20",
         10234 => x"54",
         10235 => x"54",
         10236 => x"28",
         10237 => x"6e",
         10238 => x"73",
         10239 => x"32",
         10240 => x"0a",
         10241 => x"20",
         10242 => x"53",
         10243 => x"4e",
         10244 => x"55",
         10245 => x"00",
         10246 => x"20",
         10247 => x"20",
         10248 => x"00",
         10249 => x"20",
         10250 => x"43",
         10251 => x"00",
         10252 => x"20",
         10253 => x"32",
         10254 => x"20",
         10255 => x"49",
         10256 => x"64",
         10257 => x"73",
         10258 => x"00",
         10259 => x"20",
         10260 => x"55",
         10261 => x"73",
         10262 => x"56",
         10263 => x"6f",
         10264 => x"64",
         10265 => x"73",
         10266 => x"20",
         10267 => x"58",
         10268 => x"00",
         10269 => x"20",
         10270 => x"55",
         10271 => x"6d",
         10272 => x"20",
         10273 => x"72",
         10274 => x"64",
         10275 => x"73",
         10276 => x"20",
         10277 => x"58",
         10278 => x"00",
         10279 => x"20",
         10280 => x"61",
         10281 => x"53",
         10282 => x"74",
         10283 => x"64",
         10284 => x"73",
         10285 => x"20",
         10286 => x"20",
         10287 => x"58",
         10288 => x"00",
         10289 => x"73",
         10290 => x"00",
         10291 => x"20",
         10292 => x"55",
         10293 => x"20",
         10294 => x"20",
         10295 => x"20",
         10296 => x"20",
         10297 => x"20",
         10298 => x"20",
         10299 => x"58",
         10300 => x"00",
         10301 => x"20",
         10302 => x"73",
         10303 => x"20",
         10304 => x"63",
         10305 => x"72",
         10306 => x"20",
         10307 => x"20",
         10308 => x"20",
         10309 => x"25",
         10310 => x"4d",
         10311 => x"00",
         10312 => x"20",
         10313 => x"52",
         10314 => x"43",
         10315 => x"6b",
         10316 => x"65",
         10317 => x"20",
         10318 => x"20",
         10319 => x"20",
         10320 => x"25",
         10321 => x"4d",
         10322 => x"00",
         10323 => x"20",
         10324 => x"73",
         10325 => x"6e",
         10326 => x"44",
         10327 => x"20",
         10328 => x"63",
         10329 => x"72",
         10330 => x"20",
         10331 => x"25",
         10332 => x"4d",
         10333 => x"00",
         10334 => x"61",
         10335 => x"00",
         10336 => x"64",
         10337 => x"00",
         10338 => x"65",
         10339 => x"00",
         10340 => x"4f",
         10341 => x"4f",
         10342 => x"00",
         10343 => x"6b",
         10344 => x"6e",
         10345 => x"a3",
         10346 => x"00",
         10347 => x"00",
         10348 => x"a2",
         10349 => x"00",
         10350 => x"00",
         10351 => x"a2",
         10352 => x"00",
         10353 => x"00",
         10354 => x"a2",
         10355 => x"00",
         10356 => x"00",
         10357 => x"a2",
         10358 => x"00",
         10359 => x"00",
         10360 => x"a2",
         10361 => x"00",
         10362 => x"00",
         10363 => x"a2",
         10364 => x"00",
         10365 => x"00",
         10366 => x"a2",
         10367 => x"00",
         10368 => x"00",
         10369 => x"a2",
         10370 => x"00",
         10371 => x"00",
         10372 => x"a2",
         10373 => x"00",
         10374 => x"00",
         10375 => x"a2",
         10376 => x"00",
         10377 => x"00",
         10378 => x"a2",
         10379 => x"00",
         10380 => x"00",
         10381 => x"a2",
         10382 => x"00",
         10383 => x"00",
         10384 => x"a2",
         10385 => x"00",
         10386 => x"00",
         10387 => x"a2",
         10388 => x"00",
         10389 => x"00",
         10390 => x"a2",
         10391 => x"00",
         10392 => x"00",
         10393 => x"a2",
         10394 => x"00",
         10395 => x"00",
         10396 => x"a2",
         10397 => x"00",
         10398 => x"00",
         10399 => x"a2",
         10400 => x"00",
         10401 => x"00",
         10402 => x"a2",
         10403 => x"00",
         10404 => x"00",
         10405 => x"a2",
         10406 => x"00",
         10407 => x"00",
         10408 => x"a2",
         10409 => x"00",
         10410 => x"00",
         10411 => x"44",
         10412 => x"43",
         10413 => x"42",
         10414 => x"41",
         10415 => x"36",
         10416 => x"35",
         10417 => x"34",
         10418 => x"46",
         10419 => x"33",
         10420 => x"32",
         10421 => x"31",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"00",
         10430 => x"00",
         10431 => x"00",
         10432 => x"00",
         10433 => x"73",
         10434 => x"79",
         10435 => x"73",
         10436 => x"00",
         10437 => x"00",
         10438 => x"34",
         10439 => x"20",
         10440 => x"00",
         10441 => x"69",
         10442 => x"20",
         10443 => x"72",
         10444 => x"74",
         10445 => x"65",
         10446 => x"73",
         10447 => x"79",
         10448 => x"6c",
         10449 => x"6f",
         10450 => x"46",
         10451 => x"00",
         10452 => x"6e",
         10453 => x"20",
         10454 => x"6e",
         10455 => x"65",
         10456 => x"20",
         10457 => x"74",
         10458 => x"20",
         10459 => x"65",
         10460 => x"69",
         10461 => x"6c",
         10462 => x"2e",
         10463 => x"00",
         10464 => x"3a",
         10465 => x"7c",
         10466 => x"00",
         10467 => x"3b",
         10468 => x"00",
         10469 => x"54",
         10470 => x"54",
         10471 => x"00",
         10472 => x"90",
         10473 => x"4f",
         10474 => x"30",
         10475 => x"20",
         10476 => x"45",
         10477 => x"20",
         10478 => x"33",
         10479 => x"20",
         10480 => x"20",
         10481 => x"45",
         10482 => x"20",
         10483 => x"20",
         10484 => x"20",
         10485 => x"a3",
         10486 => x"00",
         10487 => x"00",
         10488 => x"00",
         10489 => x"05",
         10490 => x"10",
         10491 => x"18",
         10492 => x"00",
         10493 => x"45",
         10494 => x"8f",
         10495 => x"45",
         10496 => x"8e",
         10497 => x"92",
         10498 => x"55",
         10499 => x"9a",
         10500 => x"9e",
         10501 => x"4f",
         10502 => x"a6",
         10503 => x"aa",
         10504 => x"ae",
         10505 => x"b2",
         10506 => x"b6",
         10507 => x"ba",
         10508 => x"be",
         10509 => x"c2",
         10510 => x"c6",
         10511 => x"ca",
         10512 => x"ce",
         10513 => x"d2",
         10514 => x"d6",
         10515 => x"da",
         10516 => x"de",
         10517 => x"e2",
         10518 => x"e6",
         10519 => x"ea",
         10520 => x"ee",
         10521 => x"f2",
         10522 => x"f6",
         10523 => x"fa",
         10524 => x"fe",
         10525 => x"2c",
         10526 => x"5d",
         10527 => x"2a",
         10528 => x"3f",
         10529 => x"00",
         10530 => x"00",
         10531 => x"00",
         10532 => x"02",
         10533 => x"00",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"00",
         10538 => x"00",
         10539 => x"00",
         10540 => x"00",
         10541 => x"00",
         10542 => x"00",
         10543 => x"00",
         10544 => x"00",
         10545 => x"00",
         10546 => x"00",
         10547 => x"00",
         10548 => x"00",
         10549 => x"00",
         10550 => x"00",
         10551 => x"00",
         10552 => x"00",
         10553 => x"01",
         10554 => x"00",
         10555 => x"00",
         10556 => x"00",
         10557 => x"00",
         10558 => x"23",
         10559 => x"00",
         10560 => x"00",
         10561 => x"00",
         10562 => x"25",
         10563 => x"25",
         10564 => x"25",
         10565 => x"25",
         10566 => x"25",
         10567 => x"25",
         10568 => x"25",
         10569 => x"25",
         10570 => x"25",
         10571 => x"25",
         10572 => x"25",
         10573 => x"25",
         10574 => x"25",
         10575 => x"25",
         10576 => x"25",
         10577 => x"25",
         10578 => x"25",
         10579 => x"25",
         10580 => x"25",
         10581 => x"25",
         10582 => x"25",
         10583 => x"25",
         10584 => x"25",
         10585 => x"25",
         10586 => x"00",
         10587 => x"03",
         10588 => x"03",
         10589 => x"03",
         10590 => x"03",
         10591 => x"03",
         10592 => x"03",
         10593 => x"22",
         10594 => x"00",
         10595 => x"22",
         10596 => x"23",
         10597 => x"22",
         10598 => x"22",
         10599 => x"22",
         10600 => x"00",
         10601 => x"00",
         10602 => x"03",
         10603 => x"03",
         10604 => x"03",
         10605 => x"00",
         10606 => x"01",
         10607 => x"01",
         10608 => x"01",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"02",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"01",
         10622 => x"01",
         10623 => x"01",
         10624 => x"01",
         10625 => x"02",
         10626 => x"01",
         10627 => x"02",
         10628 => x"01",
         10629 => x"01",
         10630 => x"01",
         10631 => x"01",
         10632 => x"01",
         10633 => x"01",
         10634 => x"01",
         10635 => x"01",
         10636 => x"01",
         10637 => x"01",
         10638 => x"01",
         10639 => x"01",
         10640 => x"01",
         10641 => x"01",
         10642 => x"01",
         10643 => x"01",
         10644 => x"01",
         10645 => x"01",
         10646 => x"01",
         10647 => x"01",
         10648 => x"01",
         10649 => x"01",
         10650 => x"01",
         10651 => x"01",
         10652 => x"00",
         10653 => x"01",
         10654 => x"01",
         10655 => x"01",
         10656 => x"01",
         10657 => x"01",
         10658 => x"01",
         10659 => x"00",
         10660 => x"02",
         10661 => x"02",
         10662 => x"02",
         10663 => x"02",
         10664 => x"02",
         10665 => x"02",
         10666 => x"01",
         10667 => x"02",
         10668 => x"01",
         10669 => x"01",
         10670 => x"01",
         10671 => x"02",
         10672 => x"02",
         10673 => x"02",
         10674 => x"01",
         10675 => x"02",
         10676 => x"02",
         10677 => x"01",
         10678 => x"2c",
         10679 => x"02",
         10680 => x"01",
         10681 => x"02",
         10682 => x"02",
         10683 => x"01",
         10684 => x"02",
         10685 => x"02",
         10686 => x"02",
         10687 => x"2c",
         10688 => x"02",
         10689 => x"02",
         10690 => x"01",
         10691 => x"02",
         10692 => x"02",
         10693 => x"02",
         10694 => x"01",
         10695 => x"02",
         10696 => x"02",
         10697 => x"02",
         10698 => x"03",
         10699 => x"03",
         10700 => x"03",
         10701 => x"00",
         10702 => x"03",
         10703 => x"03",
         10704 => x"03",
         10705 => x"00",
         10706 => x"03",
         10707 => x"03",
         10708 => x"00",
         10709 => x"03",
         10710 => x"03",
         10711 => x"03",
         10712 => x"03",
         10713 => x"03",
         10714 => x"03",
         10715 => x"03",
         10716 => x"03",
         10717 => x"04",
         10718 => x"04",
         10719 => x"04",
         10720 => x"04",
         10721 => x"04",
         10722 => x"04",
         10723 => x"04",
         10724 => x"01",
         10725 => x"04",
         10726 => x"00",
         10727 => x"00",
         10728 => x"1e",
         10729 => x"1e",
         10730 => x"1f",
         10731 => x"1f",
         10732 => x"1f",
         10733 => x"1f",
         10734 => x"1f",
         10735 => x"1f",
         10736 => x"1f",
         10737 => x"1f",
         10738 => x"1f",
         10739 => x"1f",
         10740 => x"06",
         10741 => x"00",
         10742 => x"1f",
         10743 => x"1f",
         10744 => x"1f",
         10745 => x"1f",
         10746 => x"1f",
         10747 => x"1f",
         10748 => x"1f",
         10749 => x"06",
         10750 => x"06",
         10751 => x"06",
         10752 => x"00",
         10753 => x"1f",
         10754 => x"1f",
         10755 => x"00",
         10756 => x"1f",
         10757 => x"1f",
         10758 => x"1f",
         10759 => x"1f",
         10760 => x"00",
         10761 => x"21",
         10762 => x"21",
         10763 => x"02",
         10764 => x"00",
         10765 => x"24",
         10766 => x"2c",
         10767 => x"2c",
         10768 => x"2c",
         10769 => x"2c",
         10770 => x"2c",
         10771 => x"2d",
         10772 => x"ff",
         10773 => x"00",
         10774 => x"00",
         10775 => x"98",
         10776 => x"01",
         10777 => x"00",
         10778 => x"00",
         10779 => x"98",
         10780 => x"01",
         10781 => x"00",
         10782 => x"00",
         10783 => x"99",
         10784 => x"03",
         10785 => x"00",
         10786 => x"00",
         10787 => x"99",
         10788 => x"03",
         10789 => x"00",
         10790 => x"00",
         10791 => x"99",
         10792 => x"03",
         10793 => x"00",
         10794 => x"00",
         10795 => x"99",
         10796 => x"04",
         10797 => x"00",
         10798 => x"00",
         10799 => x"99",
         10800 => x"04",
         10801 => x"00",
         10802 => x"00",
         10803 => x"99",
         10804 => x"04",
         10805 => x"00",
         10806 => x"00",
         10807 => x"99",
         10808 => x"04",
         10809 => x"00",
         10810 => x"00",
         10811 => x"99",
         10812 => x"04",
         10813 => x"00",
         10814 => x"00",
         10815 => x"99",
         10816 => x"04",
         10817 => x"00",
         10818 => x"00",
         10819 => x"99",
         10820 => x"04",
         10821 => x"00",
         10822 => x"00",
         10823 => x"99",
         10824 => x"05",
         10825 => x"00",
         10826 => x"00",
         10827 => x"99",
         10828 => x"05",
         10829 => x"00",
         10830 => x"00",
         10831 => x"99",
         10832 => x"05",
         10833 => x"00",
         10834 => x"00",
         10835 => x"99",
         10836 => x"05",
         10837 => x"00",
         10838 => x"00",
         10839 => x"99",
         10840 => x"07",
         10841 => x"00",
         10842 => x"00",
         10843 => x"99",
         10844 => x"07",
         10845 => x"00",
         10846 => x"00",
         10847 => x"99",
         10848 => x"08",
         10849 => x"00",
         10850 => x"00",
         10851 => x"99",
         10852 => x"08",
         10853 => x"00",
         10854 => x"00",
         10855 => x"99",
         10856 => x"08",
         10857 => x"00",
         10858 => x"00",
         10859 => x"99",
         10860 => x"08",
         10861 => x"00",
         10862 => x"00",
         10863 => x"99",
         10864 => x"09",
         10865 => x"00",
         10866 => x"00",
         10867 => x"99",
         10868 => x"09",
         10869 => x"00",
         10870 => x"00",
         10871 => x"99",
         10872 => x"09",
         10873 => x"00",
         10874 => x"00",
         10875 => x"99",
         10876 => x"09",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"7f",
         10882 => x"00",
         10883 => x"7f",
         10884 => x"00",
         10885 => x"7f",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"ff",
         10890 => x"00",
         10891 => x"00",
         10892 => x"78",
         10893 => x"00",
         10894 => x"e1",
         10895 => x"e1",
         10896 => x"e1",
         10897 => x"00",
         10898 => x"01",
         10899 => x"01",
         10900 => x"10",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"a3",
         10927 => x"00",
         10928 => x"a3",
         10929 => x"00",
         10930 => x"a3",
         10931 => x"00",
         10932 => x"00",
         10933 => x"00",
         10934 => x"00",
         10935 => x"00",
         10936 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"85",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8d",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8e",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"8f",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"90",
           324 => x"0b",
           325 => x"04",
           326 => x"90",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"91",
           336 => x"0b",
           337 => x"04",
           338 => x"91",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"80",
           387 => x"82",
           388 => x"84",
           389 => x"82",
           390 => x"b3",
           391 => x"d5",
           392 => x"80",
           393 => x"d5",
           394 => x"e3",
           395 => x"f0",
           396 => x"90",
           397 => x"f0",
           398 => x"2d",
           399 => x"08",
           400 => x"04",
           401 => x"0c",
           402 => x"82",
           403 => x"84",
           404 => x"82",
           405 => x"b1",
           406 => x"d5",
           407 => x"80",
           408 => x"d5",
           409 => x"d0",
           410 => x"d5",
           411 => x"80",
           412 => x"d5",
           413 => x"cb",
           414 => x"d5",
           415 => x"80",
           416 => x"d5",
           417 => x"d8",
           418 => x"f0",
           419 => x"90",
           420 => x"f0",
           421 => x"2d",
           422 => x"08",
           423 => x"04",
           424 => x"0c",
           425 => x"82",
           426 => x"84",
           427 => x"82",
           428 => x"80",
           429 => x"82",
           430 => x"84",
           431 => x"82",
           432 => x"80",
           433 => x"82",
           434 => x"84",
           435 => x"82",
           436 => x"80",
           437 => x"82",
           438 => x"84",
           439 => x"82",
           440 => x"80",
           441 => x"82",
           442 => x"84",
           443 => x"82",
           444 => x"80",
           445 => x"82",
           446 => x"84",
           447 => x"82",
           448 => x"81",
           449 => x"82",
           450 => x"84",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"84",
           455 => x"82",
           456 => x"81",
           457 => x"82",
           458 => x"84",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"84",
           463 => x"82",
           464 => x"81",
           465 => x"82",
           466 => x"84",
           467 => x"82",
           468 => x"82",
           469 => x"82",
           470 => x"84",
           471 => x"82",
           472 => x"81",
           473 => x"82",
           474 => x"84",
           475 => x"82",
           476 => x"82",
           477 => x"82",
           478 => x"84",
           479 => x"82",
           480 => x"82",
           481 => x"82",
           482 => x"84",
           483 => x"82",
           484 => x"82",
           485 => x"82",
           486 => x"84",
           487 => x"82",
           488 => x"82",
           489 => x"82",
           490 => x"84",
           491 => x"82",
           492 => x"82",
           493 => x"82",
           494 => x"84",
           495 => x"82",
           496 => x"82",
           497 => x"82",
           498 => x"84",
           499 => x"82",
           500 => x"82",
           501 => x"82",
           502 => x"84",
           503 => x"82",
           504 => x"82",
           505 => x"82",
           506 => x"84",
           507 => x"82",
           508 => x"82",
           509 => x"82",
           510 => x"84",
           511 => x"82",
           512 => x"81",
           513 => x"82",
           514 => x"84",
           515 => x"82",
           516 => x"81",
           517 => x"82",
           518 => x"84",
           519 => x"82",
           520 => x"81",
           521 => x"82",
           522 => x"84",
           523 => x"82",
           524 => x"82",
           525 => x"82",
           526 => x"84",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"84",
           531 => x"82",
           532 => x"82",
           533 => x"82",
           534 => x"84",
           535 => x"82",
           536 => x"82",
           537 => x"82",
           538 => x"84",
           539 => x"82",
           540 => x"81",
           541 => x"82",
           542 => x"84",
           543 => x"82",
           544 => x"82",
           545 => x"82",
           546 => x"84",
           547 => x"82",
           548 => x"82",
           549 => x"82",
           550 => x"84",
           551 => x"82",
           552 => x"82",
           553 => x"82",
           554 => x"84",
           555 => x"82",
           556 => x"81",
           557 => x"82",
           558 => x"84",
           559 => x"82",
           560 => x"81",
           561 => x"82",
           562 => x"84",
           563 => x"82",
           564 => x"81",
           565 => x"82",
           566 => x"84",
           567 => x"82",
           568 => x"80",
           569 => x"82",
           570 => x"84",
           571 => x"82",
           572 => x"80",
           573 => x"82",
           574 => x"84",
           575 => x"82",
           576 => x"80",
           577 => x"82",
           578 => x"84",
           579 => x"82",
           580 => x"80",
           581 => x"82",
           582 => x"84",
           583 => x"82",
           584 => x"81",
           585 => x"82",
           586 => x"84",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"84",
           591 => x"82",
           592 => x"81",
           593 => x"82",
           594 => x"84",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"84",
           599 => x"3c",
           600 => x"10",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"51",
           609 => x"73",
           610 => x"73",
           611 => x"81",
           612 => x"10",
           613 => x"07",
           614 => x"0c",
           615 => x"72",
           616 => x"81",
           617 => x"09",
           618 => x"71",
           619 => x"0a",
           620 => x"72",
           621 => x"51",
           622 => x"82",
           623 => x"82",
           624 => x"8e",
           625 => x"70",
           626 => x"0c",
           627 => x"93",
           628 => x"81",
           629 => x"c8",
           630 => x"d5",
           631 => x"82",
           632 => x"fb",
           633 => x"d5",
           634 => x"05",
           635 => x"f0",
           636 => x"0c",
           637 => x"08",
           638 => x"54",
           639 => x"08",
           640 => x"53",
           641 => x"08",
           642 => x"9a",
           643 => x"e4",
           644 => x"d5",
           645 => x"05",
           646 => x"f0",
           647 => x"08",
           648 => x"e4",
           649 => x"87",
           650 => x"d5",
           651 => x"82",
           652 => x"02",
           653 => x"0c",
           654 => x"82",
           655 => x"90",
           656 => x"11",
           657 => x"32",
           658 => x"51",
           659 => x"71",
           660 => x"0b",
           661 => x"08",
           662 => x"25",
           663 => x"39",
           664 => x"d5",
           665 => x"05",
           666 => x"39",
           667 => x"08",
           668 => x"ff",
           669 => x"f0",
           670 => x"0c",
           671 => x"d5",
           672 => x"05",
           673 => x"f0",
           674 => x"08",
           675 => x"08",
           676 => x"82",
           677 => x"f8",
           678 => x"2e",
           679 => x"80",
           680 => x"f0",
           681 => x"08",
           682 => x"38",
           683 => x"08",
           684 => x"51",
           685 => x"82",
           686 => x"70",
           687 => x"08",
           688 => x"52",
           689 => x"08",
           690 => x"ff",
           691 => x"06",
           692 => x"0b",
           693 => x"08",
           694 => x"80",
           695 => x"d5",
           696 => x"05",
           697 => x"f0",
           698 => x"08",
           699 => x"73",
           700 => x"f0",
           701 => x"08",
           702 => x"d5",
           703 => x"05",
           704 => x"f0",
           705 => x"08",
           706 => x"d5",
           707 => x"05",
           708 => x"39",
           709 => x"08",
           710 => x"52",
           711 => x"82",
           712 => x"88",
           713 => x"82",
           714 => x"f4",
           715 => x"82",
           716 => x"f4",
           717 => x"d5",
           718 => x"3d",
           719 => x"f0",
           720 => x"d5",
           721 => x"82",
           722 => x"f4",
           723 => x"0b",
           724 => x"08",
           725 => x"82",
           726 => x"88",
           727 => x"d5",
           728 => x"05",
           729 => x"0b",
           730 => x"08",
           731 => x"82",
           732 => x"90",
           733 => x"d5",
           734 => x"05",
           735 => x"f0",
           736 => x"08",
           737 => x"f0",
           738 => x"08",
           739 => x"f0",
           740 => x"70",
           741 => x"81",
           742 => x"d5",
           743 => x"82",
           744 => x"dc",
           745 => x"d5",
           746 => x"05",
           747 => x"f0",
           748 => x"08",
           749 => x"80",
           750 => x"d5",
           751 => x"05",
           752 => x"d5",
           753 => x"8e",
           754 => x"d5",
           755 => x"82",
           756 => x"02",
           757 => x"0c",
           758 => x"82",
           759 => x"90",
           760 => x"d5",
           761 => x"05",
           762 => x"f0",
           763 => x"08",
           764 => x"f0",
           765 => x"08",
           766 => x"f0",
           767 => x"08",
           768 => x"3f",
           769 => x"08",
           770 => x"f0",
           771 => x"0c",
           772 => x"08",
           773 => x"70",
           774 => x"0c",
           775 => x"3d",
           776 => x"f0",
           777 => x"d5",
           778 => x"82",
           779 => x"ed",
           780 => x"0b",
           781 => x"08",
           782 => x"82",
           783 => x"88",
           784 => x"80",
           785 => x"0c",
           786 => x"08",
           787 => x"85",
           788 => x"81",
           789 => x"32",
           790 => x"51",
           791 => x"53",
           792 => x"8d",
           793 => x"82",
           794 => x"e0",
           795 => x"ac",
           796 => x"f0",
           797 => x"08",
           798 => x"53",
           799 => x"f0",
           800 => x"34",
           801 => x"06",
           802 => x"2e",
           803 => x"82",
           804 => x"8c",
           805 => x"05",
           806 => x"08",
           807 => x"82",
           808 => x"e4",
           809 => x"81",
           810 => x"72",
           811 => x"8b",
           812 => x"f0",
           813 => x"33",
           814 => x"27",
           815 => x"82",
           816 => x"f8",
           817 => x"72",
           818 => x"ee",
           819 => x"f0",
           820 => x"33",
           821 => x"2e",
           822 => x"80",
           823 => x"d5",
           824 => x"05",
           825 => x"2b",
           826 => x"51",
           827 => x"b2",
           828 => x"f0",
           829 => x"22",
           830 => x"70",
           831 => x"81",
           832 => x"51",
           833 => x"2e",
           834 => x"d5",
           835 => x"05",
           836 => x"80",
           837 => x"72",
           838 => x"08",
           839 => x"fe",
           840 => x"d5",
           841 => x"05",
           842 => x"2b",
           843 => x"70",
           844 => x"72",
           845 => x"51",
           846 => x"51",
           847 => x"82",
           848 => x"e8",
           849 => x"d5",
           850 => x"05",
           851 => x"d5",
           852 => x"05",
           853 => x"d0",
           854 => x"53",
           855 => x"f0",
           856 => x"34",
           857 => x"08",
           858 => x"70",
           859 => x"98",
           860 => x"53",
           861 => x"8b",
           862 => x"0b",
           863 => x"08",
           864 => x"82",
           865 => x"e4",
           866 => x"83",
           867 => x"06",
           868 => x"72",
           869 => x"82",
           870 => x"e8",
           871 => x"88",
           872 => x"2b",
           873 => x"70",
           874 => x"51",
           875 => x"72",
           876 => x"08",
           877 => x"fd",
           878 => x"d5",
           879 => x"05",
           880 => x"2a",
           881 => x"51",
           882 => x"80",
           883 => x"82",
           884 => x"e8",
           885 => x"98",
           886 => x"2c",
           887 => x"72",
           888 => x"0b",
           889 => x"08",
           890 => x"82",
           891 => x"f8",
           892 => x"11",
           893 => x"08",
           894 => x"53",
           895 => x"08",
           896 => x"80",
           897 => x"94",
           898 => x"f0",
           899 => x"08",
           900 => x"82",
           901 => x"70",
           902 => x"51",
           903 => x"82",
           904 => x"e4",
           905 => x"90",
           906 => x"72",
           907 => x"08",
           908 => x"82",
           909 => x"e4",
           910 => x"a0",
           911 => x"72",
           912 => x"08",
           913 => x"fc",
           914 => x"d5",
           915 => x"05",
           916 => x"80",
           917 => x"72",
           918 => x"08",
           919 => x"fc",
           920 => x"d5",
           921 => x"05",
           922 => x"c0",
           923 => x"72",
           924 => x"08",
           925 => x"fb",
           926 => x"d5",
           927 => x"05",
           928 => x"07",
           929 => x"82",
           930 => x"e4",
           931 => x"0b",
           932 => x"08",
           933 => x"fb",
           934 => x"d5",
           935 => x"05",
           936 => x"07",
           937 => x"82",
           938 => x"e4",
           939 => x"c1",
           940 => x"82",
           941 => x"fc",
           942 => x"d5",
           943 => x"05",
           944 => x"51",
           945 => x"d5",
           946 => x"05",
           947 => x"0b",
           948 => x"08",
           949 => x"8d",
           950 => x"d5",
           951 => x"05",
           952 => x"f0",
           953 => x"08",
           954 => x"d5",
           955 => x"05",
           956 => x"51",
           957 => x"d5",
           958 => x"05",
           959 => x"f0",
           960 => x"22",
           961 => x"53",
           962 => x"f0",
           963 => x"23",
           964 => x"82",
           965 => x"90",
           966 => x"d5",
           967 => x"05",
           968 => x"82",
           969 => x"90",
           970 => x"08",
           971 => x"08",
           972 => x"82",
           973 => x"e4",
           974 => x"83",
           975 => x"06",
           976 => x"53",
           977 => x"ab",
           978 => x"f0",
           979 => x"33",
           980 => x"53",
           981 => x"53",
           982 => x"08",
           983 => x"52",
           984 => x"3f",
           985 => x"08",
           986 => x"d5",
           987 => x"05",
           988 => x"82",
           989 => x"fc",
           990 => x"9d",
           991 => x"d5",
           992 => x"72",
           993 => x"08",
           994 => x"82",
           995 => x"ec",
           996 => x"82",
           997 => x"f4",
           998 => x"71",
           999 => x"72",
          1000 => x"08",
          1001 => x"8b",
          1002 => x"d5",
          1003 => x"05",
          1004 => x"f0",
          1005 => x"08",
          1006 => x"d5",
          1007 => x"05",
          1008 => x"82",
          1009 => x"fc",
          1010 => x"d5",
          1011 => x"05",
          1012 => x"2a",
          1013 => x"51",
          1014 => x"72",
          1015 => x"38",
          1016 => x"08",
          1017 => x"70",
          1018 => x"72",
          1019 => x"82",
          1020 => x"fc",
          1021 => x"53",
          1022 => x"82",
          1023 => x"53",
          1024 => x"f0",
          1025 => x"23",
          1026 => x"d5",
          1027 => x"05",
          1028 => x"f3",
          1029 => x"e4",
          1030 => x"82",
          1031 => x"f4",
          1032 => x"d5",
          1033 => x"05",
          1034 => x"d5",
          1035 => x"05",
          1036 => x"31",
          1037 => x"82",
          1038 => x"ec",
          1039 => x"c1",
          1040 => x"f0",
          1041 => x"22",
          1042 => x"70",
          1043 => x"51",
          1044 => x"2e",
          1045 => x"d5",
          1046 => x"05",
          1047 => x"f0",
          1048 => x"08",
          1049 => x"d5",
          1050 => x"05",
          1051 => x"82",
          1052 => x"dc",
          1053 => x"a2",
          1054 => x"f0",
          1055 => x"08",
          1056 => x"08",
          1057 => x"84",
          1058 => x"f0",
          1059 => x"0c",
          1060 => x"d5",
          1061 => x"05",
          1062 => x"d5",
          1063 => x"05",
          1064 => x"f0",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"80",
          1068 => x"82",
          1069 => x"e4",
          1070 => x"82",
          1071 => x"72",
          1072 => x"08",
          1073 => x"82",
          1074 => x"fc",
          1075 => x"82",
          1076 => x"fc",
          1077 => x"d5",
          1078 => x"05",
          1079 => x"bf",
          1080 => x"72",
          1081 => x"08",
          1082 => x"81",
          1083 => x"0b",
          1084 => x"08",
          1085 => x"a9",
          1086 => x"f0",
          1087 => x"22",
          1088 => x"07",
          1089 => x"82",
          1090 => x"e4",
          1091 => x"f8",
          1092 => x"f0",
          1093 => x"34",
          1094 => x"d5",
          1095 => x"05",
          1096 => x"f0",
          1097 => x"22",
          1098 => x"70",
          1099 => x"51",
          1100 => x"2e",
          1101 => x"d5",
          1102 => x"05",
          1103 => x"f0",
          1104 => x"08",
          1105 => x"d5",
          1106 => x"05",
          1107 => x"82",
          1108 => x"d8",
          1109 => x"a2",
          1110 => x"f0",
          1111 => x"08",
          1112 => x"08",
          1113 => x"84",
          1114 => x"f0",
          1115 => x"0c",
          1116 => x"d5",
          1117 => x"05",
          1118 => x"d5",
          1119 => x"05",
          1120 => x"f0",
          1121 => x"0c",
          1122 => x"08",
          1123 => x"70",
          1124 => x"53",
          1125 => x"f0",
          1126 => x"23",
          1127 => x"0b",
          1128 => x"08",
          1129 => x"82",
          1130 => x"f0",
          1131 => x"d5",
          1132 => x"05",
          1133 => x"f0",
          1134 => x"08",
          1135 => x"54",
          1136 => x"a5",
          1137 => x"d5",
          1138 => x"72",
          1139 => x"d5",
          1140 => x"05",
          1141 => x"f0",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"70",
          1145 => x"89",
          1146 => x"38",
          1147 => x"08",
          1148 => x"53",
          1149 => x"82",
          1150 => x"f8",
          1151 => x"15",
          1152 => x"51",
          1153 => x"d5",
          1154 => x"05",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"72",
          1158 => x"51",
          1159 => x"d5",
          1160 => x"05",
          1161 => x"f0",
          1162 => x"08",
          1163 => x"f0",
          1164 => x"33",
          1165 => x"d5",
          1166 => x"05",
          1167 => x"82",
          1168 => x"f0",
          1169 => x"d5",
          1170 => x"05",
          1171 => x"82",
          1172 => x"fc",
          1173 => x"53",
          1174 => x"82",
          1175 => x"70",
          1176 => x"08",
          1177 => x"53",
          1178 => x"08",
          1179 => x"80",
          1180 => x"fe",
          1181 => x"d5",
          1182 => x"05",
          1183 => x"f4",
          1184 => x"54",
          1185 => x"31",
          1186 => x"82",
          1187 => x"fc",
          1188 => x"d5",
          1189 => x"05",
          1190 => x"06",
          1191 => x"80",
          1192 => x"82",
          1193 => x"ec",
          1194 => x"11",
          1195 => x"82",
          1196 => x"ec",
          1197 => x"d5",
          1198 => x"05",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"80",
          1202 => x"38",
          1203 => x"08",
          1204 => x"70",
          1205 => x"d5",
          1206 => x"05",
          1207 => x"f0",
          1208 => x"08",
          1209 => x"d5",
          1210 => x"05",
          1211 => x"f0",
          1212 => x"22",
          1213 => x"90",
          1214 => x"06",
          1215 => x"d5",
          1216 => x"05",
          1217 => x"53",
          1218 => x"f0",
          1219 => x"23",
          1220 => x"d5",
          1221 => x"05",
          1222 => x"53",
          1223 => x"f0",
          1224 => x"23",
          1225 => x"08",
          1226 => x"82",
          1227 => x"ec",
          1228 => x"d5",
          1229 => x"05",
          1230 => x"2a",
          1231 => x"51",
          1232 => x"80",
          1233 => x"38",
          1234 => x"08",
          1235 => x"70",
          1236 => x"98",
          1237 => x"f0",
          1238 => x"33",
          1239 => x"53",
          1240 => x"97",
          1241 => x"f0",
          1242 => x"22",
          1243 => x"51",
          1244 => x"d5",
          1245 => x"05",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"82",
          1249 => x"fc",
          1250 => x"71",
          1251 => x"72",
          1252 => x"08",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"83",
          1256 => x"06",
          1257 => x"72",
          1258 => x"38",
          1259 => x"08",
          1260 => x"70",
          1261 => x"90",
          1262 => x"2c",
          1263 => x"51",
          1264 => x"53",
          1265 => x"d5",
          1266 => x"05",
          1267 => x"31",
          1268 => x"82",
          1269 => x"ec",
          1270 => x"39",
          1271 => x"08",
          1272 => x"70",
          1273 => x"90",
          1274 => x"2c",
          1275 => x"51",
          1276 => x"53",
          1277 => x"d5",
          1278 => x"05",
          1279 => x"31",
          1280 => x"82",
          1281 => x"ec",
          1282 => x"d5",
          1283 => x"05",
          1284 => x"80",
          1285 => x"72",
          1286 => x"d5",
          1287 => x"05",
          1288 => x"54",
          1289 => x"d5",
          1290 => x"05",
          1291 => x"2b",
          1292 => x"51",
          1293 => x"25",
          1294 => x"d5",
          1295 => x"05",
          1296 => x"51",
          1297 => x"d2",
          1298 => x"f0",
          1299 => x"22",
          1300 => x"70",
          1301 => x"51",
          1302 => x"2e",
          1303 => x"d5",
          1304 => x"05",
          1305 => x"51",
          1306 => x"80",
          1307 => x"d5",
          1308 => x"05",
          1309 => x"2a",
          1310 => x"51",
          1311 => x"80",
          1312 => x"82",
          1313 => x"88",
          1314 => x"ab",
          1315 => x"3f",
          1316 => x"d5",
          1317 => x"05",
          1318 => x"2a",
          1319 => x"51",
          1320 => x"80",
          1321 => x"82",
          1322 => x"88",
          1323 => x"a0",
          1324 => x"3f",
          1325 => x"08",
          1326 => x"70",
          1327 => x"81",
          1328 => x"53",
          1329 => x"b1",
          1330 => x"f0",
          1331 => x"08",
          1332 => x"89",
          1333 => x"d5",
          1334 => x"05",
          1335 => x"90",
          1336 => x"06",
          1337 => x"d5",
          1338 => x"05",
          1339 => x"d5",
          1340 => x"05",
          1341 => x"bc",
          1342 => x"f0",
          1343 => x"22",
          1344 => x"70",
          1345 => x"51",
          1346 => x"2e",
          1347 => x"d5",
          1348 => x"05",
          1349 => x"54",
          1350 => x"d5",
          1351 => x"05",
          1352 => x"2b",
          1353 => x"51",
          1354 => x"25",
          1355 => x"d5",
          1356 => x"05",
          1357 => x"51",
          1358 => x"d2",
          1359 => x"f0",
          1360 => x"22",
          1361 => x"70",
          1362 => x"51",
          1363 => x"2e",
          1364 => x"d5",
          1365 => x"05",
          1366 => x"54",
          1367 => x"d5",
          1368 => x"05",
          1369 => x"2b",
          1370 => x"51",
          1371 => x"25",
          1372 => x"d5",
          1373 => x"05",
          1374 => x"51",
          1375 => x"d2",
          1376 => x"f0",
          1377 => x"22",
          1378 => x"70",
          1379 => x"51",
          1380 => x"38",
          1381 => x"08",
          1382 => x"ff",
          1383 => x"72",
          1384 => x"08",
          1385 => x"73",
          1386 => x"90",
          1387 => x"80",
          1388 => x"38",
          1389 => x"08",
          1390 => x"52",
          1391 => x"f4",
          1392 => x"82",
          1393 => x"f8",
          1394 => x"72",
          1395 => x"09",
          1396 => x"38",
          1397 => x"08",
          1398 => x"52",
          1399 => x"08",
          1400 => x"51",
          1401 => x"81",
          1402 => x"d5",
          1403 => x"05",
          1404 => x"80",
          1405 => x"81",
          1406 => x"38",
          1407 => x"08",
          1408 => x"ff",
          1409 => x"72",
          1410 => x"08",
          1411 => x"72",
          1412 => x"06",
          1413 => x"ff",
          1414 => x"bb",
          1415 => x"f0",
          1416 => x"08",
          1417 => x"f0",
          1418 => x"08",
          1419 => x"82",
          1420 => x"fc",
          1421 => x"05",
          1422 => x"08",
          1423 => x"53",
          1424 => x"ff",
          1425 => x"d5",
          1426 => x"05",
          1427 => x"80",
          1428 => x"81",
          1429 => x"38",
          1430 => x"08",
          1431 => x"ff",
          1432 => x"72",
          1433 => x"08",
          1434 => x"72",
          1435 => x"06",
          1436 => x"ff",
          1437 => x"df",
          1438 => x"f0",
          1439 => x"08",
          1440 => x"f0",
          1441 => x"08",
          1442 => x"53",
          1443 => x"82",
          1444 => x"fc",
          1445 => x"05",
          1446 => x"08",
          1447 => x"ff",
          1448 => x"d5",
          1449 => x"05",
          1450 => x"f4",
          1451 => x"82",
          1452 => x"88",
          1453 => x"82",
          1454 => x"f0",
          1455 => x"05",
          1456 => x"08",
          1457 => x"82",
          1458 => x"f0",
          1459 => x"33",
          1460 => x"e0",
          1461 => x"82",
          1462 => x"e4",
          1463 => x"87",
          1464 => x"06",
          1465 => x"72",
          1466 => x"c3",
          1467 => x"f0",
          1468 => x"22",
          1469 => x"54",
          1470 => x"f0",
          1471 => x"23",
          1472 => x"70",
          1473 => x"53",
          1474 => x"a3",
          1475 => x"f0",
          1476 => x"08",
          1477 => x"85",
          1478 => x"39",
          1479 => x"08",
          1480 => x"52",
          1481 => x"08",
          1482 => x"51",
          1483 => x"80",
          1484 => x"f0",
          1485 => x"23",
          1486 => x"82",
          1487 => x"f8",
          1488 => x"72",
          1489 => x"81",
          1490 => x"81",
          1491 => x"f0",
          1492 => x"23",
          1493 => x"d5",
          1494 => x"05",
          1495 => x"82",
          1496 => x"e8",
          1497 => x"0b",
          1498 => x"08",
          1499 => x"ea",
          1500 => x"d5",
          1501 => x"05",
          1502 => x"d5",
          1503 => x"05",
          1504 => x"b0",
          1505 => x"39",
          1506 => x"08",
          1507 => x"8c",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"53",
          1511 => x"08",
          1512 => x"82",
          1513 => x"95",
          1514 => x"d5",
          1515 => x"82",
          1516 => x"02",
          1517 => x"0c",
          1518 => x"82",
          1519 => x"53",
          1520 => x"08",
          1521 => x"52",
          1522 => x"08",
          1523 => x"51",
          1524 => x"82",
          1525 => x"70",
          1526 => x"0c",
          1527 => x"0d",
          1528 => x"0c",
          1529 => x"f0",
          1530 => x"d5",
          1531 => x"3d",
          1532 => x"82",
          1533 => x"f8",
          1534 => x"f1",
          1535 => x"11",
          1536 => x"2a",
          1537 => x"70",
          1538 => x"51",
          1539 => x"72",
          1540 => x"38",
          1541 => x"d5",
          1542 => x"05",
          1543 => x"39",
          1544 => x"08",
          1545 => x"53",
          1546 => x"d5",
          1547 => x"05",
          1548 => x"82",
          1549 => x"88",
          1550 => x"72",
          1551 => x"08",
          1552 => x"72",
          1553 => x"53",
          1554 => x"b0",
          1555 => x"c8",
          1556 => x"c8",
          1557 => x"d5",
          1558 => x"05",
          1559 => x"11",
          1560 => x"72",
          1561 => x"e4",
          1562 => x"80",
          1563 => x"38",
          1564 => x"d5",
          1565 => x"05",
          1566 => x"39",
          1567 => x"08",
          1568 => x"08",
          1569 => x"51",
          1570 => x"53",
          1571 => x"d5",
          1572 => x"72",
          1573 => x"38",
          1574 => x"d5",
          1575 => x"05",
          1576 => x"f0",
          1577 => x"08",
          1578 => x"f0",
          1579 => x"0c",
          1580 => x"f0",
          1581 => x"08",
          1582 => x"0c",
          1583 => x"82",
          1584 => x"04",
          1585 => x"08",
          1586 => x"f0",
          1587 => x"0d",
          1588 => x"d5",
          1589 => x"05",
          1590 => x"f0",
          1591 => x"08",
          1592 => x"70",
          1593 => x"81",
          1594 => x"06",
          1595 => x"51",
          1596 => x"2e",
          1597 => x"0b",
          1598 => x"08",
          1599 => x"80",
          1600 => x"d5",
          1601 => x"05",
          1602 => x"33",
          1603 => x"08",
          1604 => x"81",
          1605 => x"f0",
          1606 => x"0c",
          1607 => x"d5",
          1608 => x"05",
          1609 => x"ff",
          1610 => x"80",
          1611 => x"82",
          1612 => x"8c",
          1613 => x"d5",
          1614 => x"05",
          1615 => x"d5",
          1616 => x"05",
          1617 => x"11",
          1618 => x"72",
          1619 => x"e4",
          1620 => x"80",
          1621 => x"38",
          1622 => x"d5",
          1623 => x"05",
          1624 => x"39",
          1625 => x"08",
          1626 => x"70",
          1627 => x"08",
          1628 => x"53",
          1629 => x"08",
          1630 => x"82",
          1631 => x"87",
          1632 => x"d5",
          1633 => x"82",
          1634 => x"02",
          1635 => x"0c",
          1636 => x"82",
          1637 => x"52",
          1638 => x"08",
          1639 => x"51",
          1640 => x"d5",
          1641 => x"82",
          1642 => x"53",
          1643 => x"82",
          1644 => x"04",
          1645 => x"08",
          1646 => x"f0",
          1647 => x"0d",
          1648 => x"08",
          1649 => x"85",
          1650 => x"81",
          1651 => x"32",
          1652 => x"51",
          1653 => x"53",
          1654 => x"8d",
          1655 => x"82",
          1656 => x"fc",
          1657 => x"cb",
          1658 => x"f0",
          1659 => x"08",
          1660 => x"70",
          1661 => x"81",
          1662 => x"51",
          1663 => x"2e",
          1664 => x"82",
          1665 => x"8c",
          1666 => x"d5",
          1667 => x"05",
          1668 => x"8c",
          1669 => x"14",
          1670 => x"38",
          1671 => x"08",
          1672 => x"70",
          1673 => x"d5",
          1674 => x"05",
          1675 => x"54",
          1676 => x"34",
          1677 => x"05",
          1678 => x"d5",
          1679 => x"05",
          1680 => x"08",
          1681 => x"12",
          1682 => x"f0",
          1683 => x"08",
          1684 => x"f0",
          1685 => x"0c",
          1686 => x"d7",
          1687 => x"f0",
          1688 => x"08",
          1689 => x"08",
          1690 => x"53",
          1691 => x"08",
          1692 => x"70",
          1693 => x"53",
          1694 => x"51",
          1695 => x"2d",
          1696 => x"08",
          1697 => x"38",
          1698 => x"08",
          1699 => x"8c",
          1700 => x"05",
          1701 => x"82",
          1702 => x"88",
          1703 => x"82",
          1704 => x"fc",
          1705 => x"53",
          1706 => x"0b",
          1707 => x"08",
          1708 => x"82",
          1709 => x"fc",
          1710 => x"d5",
          1711 => x"3d",
          1712 => x"f0",
          1713 => x"d5",
          1714 => x"82",
          1715 => x"f9",
          1716 => x"d5",
          1717 => x"05",
          1718 => x"33",
          1719 => x"70",
          1720 => x"51",
          1721 => x"80",
          1722 => x"ff",
          1723 => x"f0",
          1724 => x"0c",
          1725 => x"82",
          1726 => x"88",
          1727 => x"11",
          1728 => x"2a",
          1729 => x"51",
          1730 => x"71",
          1731 => x"c5",
          1732 => x"f0",
          1733 => x"08",
          1734 => x"08",
          1735 => x"53",
          1736 => x"33",
          1737 => x"06",
          1738 => x"85",
          1739 => x"d5",
          1740 => x"05",
          1741 => x"08",
          1742 => x"12",
          1743 => x"f0",
          1744 => x"08",
          1745 => x"70",
          1746 => x"08",
          1747 => x"51",
          1748 => x"b6",
          1749 => x"f0",
          1750 => x"08",
          1751 => x"70",
          1752 => x"81",
          1753 => x"51",
          1754 => x"2e",
          1755 => x"82",
          1756 => x"88",
          1757 => x"08",
          1758 => x"d5",
          1759 => x"05",
          1760 => x"82",
          1761 => x"fc",
          1762 => x"38",
          1763 => x"08",
          1764 => x"82",
          1765 => x"88",
          1766 => x"53",
          1767 => x"70",
          1768 => x"52",
          1769 => x"34",
          1770 => x"d5",
          1771 => x"05",
          1772 => x"39",
          1773 => x"08",
          1774 => x"70",
          1775 => x"71",
          1776 => x"a1",
          1777 => x"f0",
          1778 => x"08",
          1779 => x"08",
          1780 => x"52",
          1781 => x"51",
          1782 => x"82",
          1783 => x"70",
          1784 => x"08",
          1785 => x"52",
          1786 => x"08",
          1787 => x"80",
          1788 => x"38",
          1789 => x"08",
          1790 => x"82",
          1791 => x"f4",
          1792 => x"d5",
          1793 => x"05",
          1794 => x"33",
          1795 => x"08",
          1796 => x"52",
          1797 => x"08",
          1798 => x"ff",
          1799 => x"06",
          1800 => x"d5",
          1801 => x"05",
          1802 => x"52",
          1803 => x"f0",
          1804 => x"34",
          1805 => x"d5",
          1806 => x"05",
          1807 => x"52",
          1808 => x"f0",
          1809 => x"34",
          1810 => x"08",
          1811 => x"52",
          1812 => x"08",
          1813 => x"85",
          1814 => x"0b",
          1815 => x"08",
          1816 => x"a6",
          1817 => x"f0",
          1818 => x"08",
          1819 => x"81",
          1820 => x"0c",
          1821 => x"08",
          1822 => x"70",
          1823 => x"70",
          1824 => x"08",
          1825 => x"51",
          1826 => x"d5",
          1827 => x"05",
          1828 => x"e4",
          1829 => x"0d",
          1830 => x"0c",
          1831 => x"f0",
          1832 => x"d5",
          1833 => x"3d",
          1834 => x"f0",
          1835 => x"08",
          1836 => x"08",
          1837 => x"82",
          1838 => x"8c",
          1839 => x"d5",
          1840 => x"05",
          1841 => x"f0",
          1842 => x"08",
          1843 => x"a2",
          1844 => x"f0",
          1845 => x"08",
          1846 => x"08",
          1847 => x"26",
          1848 => x"82",
          1849 => x"f8",
          1850 => x"d5",
          1851 => x"05",
          1852 => x"82",
          1853 => x"fc",
          1854 => x"27",
          1855 => x"82",
          1856 => x"fc",
          1857 => x"d5",
          1858 => x"05",
          1859 => x"d5",
          1860 => x"05",
          1861 => x"f0",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"08",
          1866 => x"82",
          1867 => x"90",
          1868 => x"05",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"05",
          1873 => x"08",
          1874 => x"82",
          1875 => x"90",
          1876 => x"2e",
          1877 => x"82",
          1878 => x"fc",
          1879 => x"05",
          1880 => x"08",
          1881 => x"82",
          1882 => x"f8",
          1883 => x"05",
          1884 => x"08",
          1885 => x"82",
          1886 => x"fc",
          1887 => x"d5",
          1888 => x"05",
          1889 => x"71",
          1890 => x"ff",
          1891 => x"d5",
          1892 => x"05",
          1893 => x"82",
          1894 => x"90",
          1895 => x"d5",
          1896 => x"05",
          1897 => x"82",
          1898 => x"90",
          1899 => x"d5",
          1900 => x"05",
          1901 => x"ba",
          1902 => x"f0",
          1903 => x"08",
          1904 => x"82",
          1905 => x"f8",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"fc",
          1910 => x"52",
          1911 => x"82",
          1912 => x"fc",
          1913 => x"05",
          1914 => x"08",
          1915 => x"ff",
          1916 => x"d5",
          1917 => x"05",
          1918 => x"d5",
          1919 => x"85",
          1920 => x"d5",
          1921 => x"82",
          1922 => x"02",
          1923 => x"0c",
          1924 => x"82",
          1925 => x"88",
          1926 => x"d5",
          1927 => x"05",
          1928 => x"f0",
          1929 => x"08",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"05",
          1933 => x"08",
          1934 => x"70",
          1935 => x"51",
          1936 => x"2e",
          1937 => x"39",
          1938 => x"08",
          1939 => x"ff",
          1940 => x"f0",
          1941 => x"0c",
          1942 => x"08",
          1943 => x"82",
          1944 => x"88",
          1945 => x"70",
          1946 => x"0c",
          1947 => x"0d",
          1948 => x"0c",
          1949 => x"f0",
          1950 => x"d5",
          1951 => x"3d",
          1952 => x"f0",
          1953 => x"08",
          1954 => x"08",
          1955 => x"82",
          1956 => x"8c",
          1957 => x"71",
          1958 => x"f0",
          1959 => x"08",
          1960 => x"d5",
          1961 => x"05",
          1962 => x"f0",
          1963 => x"08",
          1964 => x"72",
          1965 => x"f0",
          1966 => x"08",
          1967 => x"d5",
          1968 => x"05",
          1969 => x"ff",
          1970 => x"80",
          1971 => x"ff",
          1972 => x"d5",
          1973 => x"05",
          1974 => x"d5",
          1975 => x"84",
          1976 => x"d5",
          1977 => x"82",
          1978 => x"02",
          1979 => x"0c",
          1980 => x"82",
          1981 => x"88",
          1982 => x"d5",
          1983 => x"05",
          1984 => x"f0",
          1985 => x"08",
          1986 => x"08",
          1987 => x"82",
          1988 => x"90",
          1989 => x"2e",
          1990 => x"82",
          1991 => x"90",
          1992 => x"05",
          1993 => x"08",
          1994 => x"82",
          1995 => x"90",
          1996 => x"05",
          1997 => x"08",
          1998 => x"82",
          1999 => x"90",
          2000 => x"2e",
          2001 => x"d5",
          2002 => x"05",
          2003 => x"33",
          2004 => x"08",
          2005 => x"81",
          2006 => x"f0",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"52",
          2010 => x"34",
          2011 => x"08",
          2012 => x"81",
          2013 => x"f0",
          2014 => x"0c",
          2015 => x"82",
          2016 => x"88",
          2017 => x"82",
          2018 => x"51",
          2019 => x"82",
          2020 => x"04",
          2021 => x"08",
          2022 => x"f0",
          2023 => x"0d",
          2024 => x"08",
          2025 => x"80",
          2026 => x"38",
          2027 => x"08",
          2028 => x"52",
          2029 => x"d5",
          2030 => x"05",
          2031 => x"82",
          2032 => x"8c",
          2033 => x"d5",
          2034 => x"05",
          2035 => x"72",
          2036 => x"53",
          2037 => x"71",
          2038 => x"38",
          2039 => x"82",
          2040 => x"88",
          2041 => x"71",
          2042 => x"f0",
          2043 => x"08",
          2044 => x"d5",
          2045 => x"05",
          2046 => x"ff",
          2047 => x"70",
          2048 => x"0b",
          2049 => x"08",
          2050 => x"81",
          2051 => x"d5",
          2052 => x"05",
          2053 => x"82",
          2054 => x"90",
          2055 => x"d5",
          2056 => x"05",
          2057 => x"84",
          2058 => x"39",
          2059 => x"08",
          2060 => x"80",
          2061 => x"38",
          2062 => x"08",
          2063 => x"70",
          2064 => x"70",
          2065 => x"0b",
          2066 => x"08",
          2067 => x"80",
          2068 => x"d5",
          2069 => x"05",
          2070 => x"82",
          2071 => x"8c",
          2072 => x"d5",
          2073 => x"05",
          2074 => x"52",
          2075 => x"38",
          2076 => x"d5",
          2077 => x"05",
          2078 => x"82",
          2079 => x"88",
          2080 => x"33",
          2081 => x"08",
          2082 => x"70",
          2083 => x"31",
          2084 => x"f0",
          2085 => x"0c",
          2086 => x"52",
          2087 => x"80",
          2088 => x"f0",
          2089 => x"0c",
          2090 => x"08",
          2091 => x"82",
          2092 => x"85",
          2093 => x"d5",
          2094 => x"82",
          2095 => x"02",
          2096 => x"0c",
          2097 => x"82",
          2098 => x"8c",
          2099 => x"82",
          2100 => x"88",
          2101 => x"81",
          2102 => x"d5",
          2103 => x"82",
          2104 => x"f8",
          2105 => x"d5",
          2106 => x"05",
          2107 => x"70",
          2108 => x"80",
          2109 => x"82",
          2110 => x"70",
          2111 => x"08",
          2112 => x"54",
          2113 => x"08",
          2114 => x"8c",
          2115 => x"82",
          2116 => x"f4",
          2117 => x"39",
          2118 => x"08",
          2119 => x"82",
          2120 => x"f8",
          2121 => x"54",
          2122 => x"82",
          2123 => x"f8",
          2124 => x"82",
          2125 => x"88",
          2126 => x"82",
          2127 => x"fc",
          2128 => x"fb",
          2129 => x"d5",
          2130 => x"82",
          2131 => x"f4",
          2132 => x"82",
          2133 => x"f4",
          2134 => x"d5",
          2135 => x"3d",
          2136 => x"f0",
          2137 => x"d5",
          2138 => x"82",
          2139 => x"fd",
          2140 => x"d5",
          2141 => x"05",
          2142 => x"f0",
          2143 => x"0c",
          2144 => x"08",
          2145 => x"8d",
          2146 => x"82",
          2147 => x"fc",
          2148 => x"ec",
          2149 => x"f0",
          2150 => x"08",
          2151 => x"82",
          2152 => x"f8",
          2153 => x"05",
          2154 => x"08",
          2155 => x"70",
          2156 => x"51",
          2157 => x"2e",
          2158 => x"d5",
          2159 => x"05",
          2160 => x"82",
          2161 => x"8c",
          2162 => x"d5",
          2163 => x"05",
          2164 => x"84",
          2165 => x"39",
          2166 => x"08",
          2167 => x"ff",
          2168 => x"f0",
          2169 => x"0c",
          2170 => x"08",
          2171 => x"82",
          2172 => x"88",
          2173 => x"70",
          2174 => x"08",
          2175 => x"51",
          2176 => x"08",
          2177 => x"82",
          2178 => x"85",
          2179 => x"d5",
          2180 => x"82",
          2181 => x"02",
          2182 => x"0c",
          2183 => x"82",
          2184 => x"88",
          2185 => x"d5",
          2186 => x"05",
          2187 => x"f0",
          2188 => x"08",
          2189 => x"d4",
          2190 => x"f0",
          2191 => x"08",
          2192 => x"d5",
          2193 => x"05",
          2194 => x"f0",
          2195 => x"08",
          2196 => x"d5",
          2197 => x"05",
          2198 => x"f0",
          2199 => x"08",
          2200 => x"38",
          2201 => x"08",
          2202 => x"51",
          2203 => x"f0",
          2204 => x"08",
          2205 => x"71",
          2206 => x"f0",
          2207 => x"08",
          2208 => x"d5",
          2209 => x"05",
          2210 => x"39",
          2211 => x"08",
          2212 => x"70",
          2213 => x"0c",
          2214 => x"0d",
          2215 => x"0c",
          2216 => x"f0",
          2217 => x"d5",
          2218 => x"3d",
          2219 => x"82",
          2220 => x"fc",
          2221 => x"d5",
          2222 => x"05",
          2223 => x"b9",
          2224 => x"f0",
          2225 => x"08",
          2226 => x"f0",
          2227 => x"0c",
          2228 => x"d5",
          2229 => x"05",
          2230 => x"f0",
          2231 => x"08",
          2232 => x"0b",
          2233 => x"08",
          2234 => x"82",
          2235 => x"f4",
          2236 => x"d5",
          2237 => x"05",
          2238 => x"f0",
          2239 => x"08",
          2240 => x"38",
          2241 => x"08",
          2242 => x"30",
          2243 => x"08",
          2244 => x"80",
          2245 => x"f0",
          2246 => x"0c",
          2247 => x"08",
          2248 => x"8a",
          2249 => x"82",
          2250 => x"f0",
          2251 => x"d5",
          2252 => x"05",
          2253 => x"f0",
          2254 => x"0c",
          2255 => x"d5",
          2256 => x"05",
          2257 => x"d5",
          2258 => x"05",
          2259 => x"c5",
          2260 => x"e4",
          2261 => x"d5",
          2262 => x"05",
          2263 => x"d5",
          2264 => x"05",
          2265 => x"90",
          2266 => x"f0",
          2267 => x"08",
          2268 => x"f0",
          2269 => x"0c",
          2270 => x"08",
          2271 => x"70",
          2272 => x"0c",
          2273 => x"0d",
          2274 => x"0c",
          2275 => x"f0",
          2276 => x"d5",
          2277 => x"3d",
          2278 => x"82",
          2279 => x"fc",
          2280 => x"d5",
          2281 => x"05",
          2282 => x"99",
          2283 => x"f0",
          2284 => x"08",
          2285 => x"f0",
          2286 => x"0c",
          2287 => x"d5",
          2288 => x"05",
          2289 => x"f0",
          2290 => x"08",
          2291 => x"38",
          2292 => x"08",
          2293 => x"30",
          2294 => x"08",
          2295 => x"81",
          2296 => x"f0",
          2297 => x"08",
          2298 => x"f0",
          2299 => x"08",
          2300 => x"3f",
          2301 => x"08",
          2302 => x"f0",
          2303 => x"0c",
          2304 => x"f0",
          2305 => x"08",
          2306 => x"38",
          2307 => x"08",
          2308 => x"30",
          2309 => x"08",
          2310 => x"82",
          2311 => x"f8",
          2312 => x"82",
          2313 => x"54",
          2314 => x"82",
          2315 => x"04",
          2316 => x"08",
          2317 => x"f0",
          2318 => x"0d",
          2319 => x"d5",
          2320 => x"05",
          2321 => x"d5",
          2322 => x"05",
          2323 => x"c5",
          2324 => x"e4",
          2325 => x"d5",
          2326 => x"85",
          2327 => x"d5",
          2328 => x"82",
          2329 => x"02",
          2330 => x"0c",
          2331 => x"81",
          2332 => x"f0",
          2333 => x"08",
          2334 => x"f0",
          2335 => x"08",
          2336 => x"82",
          2337 => x"70",
          2338 => x"0c",
          2339 => x"0d",
          2340 => x"0c",
          2341 => x"f0",
          2342 => x"d5",
          2343 => x"3d",
          2344 => x"82",
          2345 => x"fc",
          2346 => x"0b",
          2347 => x"08",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"d5",
          2351 => x"05",
          2352 => x"38",
          2353 => x"08",
          2354 => x"80",
          2355 => x"80",
          2356 => x"f0",
          2357 => x"08",
          2358 => x"82",
          2359 => x"8c",
          2360 => x"82",
          2361 => x"8c",
          2362 => x"d5",
          2363 => x"05",
          2364 => x"d5",
          2365 => x"05",
          2366 => x"39",
          2367 => x"08",
          2368 => x"80",
          2369 => x"38",
          2370 => x"08",
          2371 => x"82",
          2372 => x"88",
          2373 => x"ad",
          2374 => x"f0",
          2375 => x"08",
          2376 => x"08",
          2377 => x"31",
          2378 => x"08",
          2379 => x"82",
          2380 => x"f8",
          2381 => x"d5",
          2382 => x"05",
          2383 => x"d5",
          2384 => x"05",
          2385 => x"f0",
          2386 => x"08",
          2387 => x"d5",
          2388 => x"05",
          2389 => x"f0",
          2390 => x"08",
          2391 => x"d5",
          2392 => x"05",
          2393 => x"39",
          2394 => x"08",
          2395 => x"80",
          2396 => x"82",
          2397 => x"88",
          2398 => x"82",
          2399 => x"f4",
          2400 => x"91",
          2401 => x"f0",
          2402 => x"08",
          2403 => x"f0",
          2404 => x"0c",
          2405 => x"f0",
          2406 => x"08",
          2407 => x"0c",
          2408 => x"82",
          2409 => x"04",
          2410 => x"08",
          2411 => x"f0",
          2412 => x"0d",
          2413 => x"d5",
          2414 => x"05",
          2415 => x"f0",
          2416 => x"08",
          2417 => x"0c",
          2418 => x"08",
          2419 => x"70",
          2420 => x"72",
          2421 => x"82",
          2422 => x"f8",
          2423 => x"81",
          2424 => x"72",
          2425 => x"81",
          2426 => x"82",
          2427 => x"88",
          2428 => x"08",
          2429 => x"0c",
          2430 => x"82",
          2431 => x"f8",
          2432 => x"72",
          2433 => x"81",
          2434 => x"81",
          2435 => x"f0",
          2436 => x"34",
          2437 => x"08",
          2438 => x"70",
          2439 => x"71",
          2440 => x"51",
          2441 => x"82",
          2442 => x"f8",
          2443 => x"d5",
          2444 => x"05",
          2445 => x"b0",
          2446 => x"06",
          2447 => x"82",
          2448 => x"88",
          2449 => x"08",
          2450 => x"0c",
          2451 => x"53",
          2452 => x"d5",
          2453 => x"05",
          2454 => x"f0",
          2455 => x"33",
          2456 => x"08",
          2457 => x"82",
          2458 => x"e8",
          2459 => x"e2",
          2460 => x"82",
          2461 => x"e8",
          2462 => x"f8",
          2463 => x"80",
          2464 => x"0b",
          2465 => x"08",
          2466 => x"82",
          2467 => x"88",
          2468 => x"08",
          2469 => x"0c",
          2470 => x"53",
          2471 => x"d5",
          2472 => x"05",
          2473 => x"39",
          2474 => x"d5",
          2475 => x"05",
          2476 => x"f0",
          2477 => x"08",
          2478 => x"05",
          2479 => x"08",
          2480 => x"33",
          2481 => x"08",
          2482 => x"80",
          2483 => x"d5",
          2484 => x"05",
          2485 => x"a0",
          2486 => x"81",
          2487 => x"f0",
          2488 => x"0c",
          2489 => x"82",
          2490 => x"f8",
          2491 => x"af",
          2492 => x"38",
          2493 => x"08",
          2494 => x"53",
          2495 => x"83",
          2496 => x"80",
          2497 => x"f0",
          2498 => x"0c",
          2499 => x"88",
          2500 => x"f0",
          2501 => x"34",
          2502 => x"d5",
          2503 => x"05",
          2504 => x"73",
          2505 => x"82",
          2506 => x"f8",
          2507 => x"72",
          2508 => x"38",
          2509 => x"0b",
          2510 => x"08",
          2511 => x"82",
          2512 => x"0b",
          2513 => x"08",
          2514 => x"80",
          2515 => x"f0",
          2516 => x"0c",
          2517 => x"08",
          2518 => x"53",
          2519 => x"81",
          2520 => x"d5",
          2521 => x"05",
          2522 => x"e0",
          2523 => x"38",
          2524 => x"08",
          2525 => x"e0",
          2526 => x"72",
          2527 => x"08",
          2528 => x"82",
          2529 => x"f8",
          2530 => x"11",
          2531 => x"82",
          2532 => x"f8",
          2533 => x"d5",
          2534 => x"05",
          2535 => x"73",
          2536 => x"82",
          2537 => x"f8",
          2538 => x"11",
          2539 => x"82",
          2540 => x"f8",
          2541 => x"d5",
          2542 => x"05",
          2543 => x"89",
          2544 => x"80",
          2545 => x"f0",
          2546 => x"0c",
          2547 => x"82",
          2548 => x"f8",
          2549 => x"d5",
          2550 => x"05",
          2551 => x"72",
          2552 => x"38",
          2553 => x"d5",
          2554 => x"05",
          2555 => x"39",
          2556 => x"08",
          2557 => x"70",
          2558 => x"08",
          2559 => x"29",
          2560 => x"08",
          2561 => x"70",
          2562 => x"f0",
          2563 => x"0c",
          2564 => x"08",
          2565 => x"70",
          2566 => x"71",
          2567 => x"51",
          2568 => x"53",
          2569 => x"d5",
          2570 => x"05",
          2571 => x"39",
          2572 => x"08",
          2573 => x"53",
          2574 => x"90",
          2575 => x"f0",
          2576 => x"08",
          2577 => x"f0",
          2578 => x"0c",
          2579 => x"08",
          2580 => x"82",
          2581 => x"fc",
          2582 => x"0c",
          2583 => x"82",
          2584 => x"ec",
          2585 => x"d5",
          2586 => x"05",
          2587 => x"e4",
          2588 => x"0d",
          2589 => x"0c",
          2590 => x"f0",
          2591 => x"d5",
          2592 => x"3d",
          2593 => x"82",
          2594 => x"f0",
          2595 => x"d5",
          2596 => x"05",
          2597 => x"73",
          2598 => x"f0",
          2599 => x"08",
          2600 => x"53",
          2601 => x"72",
          2602 => x"08",
          2603 => x"72",
          2604 => x"53",
          2605 => x"09",
          2606 => x"38",
          2607 => x"08",
          2608 => x"70",
          2609 => x"71",
          2610 => x"39",
          2611 => x"08",
          2612 => x"53",
          2613 => x"09",
          2614 => x"38",
          2615 => x"d5",
          2616 => x"05",
          2617 => x"f0",
          2618 => x"08",
          2619 => x"05",
          2620 => x"08",
          2621 => x"33",
          2622 => x"08",
          2623 => x"82",
          2624 => x"f8",
          2625 => x"72",
          2626 => x"81",
          2627 => x"38",
          2628 => x"08",
          2629 => x"70",
          2630 => x"71",
          2631 => x"51",
          2632 => x"82",
          2633 => x"f8",
          2634 => x"d5",
          2635 => x"05",
          2636 => x"f0",
          2637 => x"0c",
          2638 => x"08",
          2639 => x"80",
          2640 => x"38",
          2641 => x"08",
          2642 => x"80",
          2643 => x"38",
          2644 => x"90",
          2645 => x"f0",
          2646 => x"34",
          2647 => x"08",
          2648 => x"70",
          2649 => x"71",
          2650 => x"51",
          2651 => x"82",
          2652 => x"f8",
          2653 => x"a4",
          2654 => x"82",
          2655 => x"f4",
          2656 => x"d5",
          2657 => x"05",
          2658 => x"81",
          2659 => x"70",
          2660 => x"72",
          2661 => x"f0",
          2662 => x"34",
          2663 => x"82",
          2664 => x"f8",
          2665 => x"72",
          2666 => x"38",
          2667 => x"d5",
          2668 => x"05",
          2669 => x"39",
          2670 => x"08",
          2671 => x"53",
          2672 => x"90",
          2673 => x"f0",
          2674 => x"33",
          2675 => x"26",
          2676 => x"39",
          2677 => x"d5",
          2678 => x"05",
          2679 => x"39",
          2680 => x"d5",
          2681 => x"05",
          2682 => x"82",
          2683 => x"f8",
          2684 => x"af",
          2685 => x"38",
          2686 => x"08",
          2687 => x"53",
          2688 => x"83",
          2689 => x"80",
          2690 => x"f0",
          2691 => x"0c",
          2692 => x"8a",
          2693 => x"f0",
          2694 => x"34",
          2695 => x"d5",
          2696 => x"05",
          2697 => x"f0",
          2698 => x"33",
          2699 => x"27",
          2700 => x"82",
          2701 => x"f8",
          2702 => x"80",
          2703 => x"94",
          2704 => x"f0",
          2705 => x"33",
          2706 => x"53",
          2707 => x"f0",
          2708 => x"34",
          2709 => x"08",
          2710 => x"d0",
          2711 => x"72",
          2712 => x"08",
          2713 => x"82",
          2714 => x"f8",
          2715 => x"90",
          2716 => x"38",
          2717 => x"08",
          2718 => x"f9",
          2719 => x"72",
          2720 => x"08",
          2721 => x"82",
          2722 => x"f8",
          2723 => x"72",
          2724 => x"38",
          2725 => x"d5",
          2726 => x"05",
          2727 => x"39",
          2728 => x"08",
          2729 => x"82",
          2730 => x"f4",
          2731 => x"54",
          2732 => x"8d",
          2733 => x"82",
          2734 => x"ec",
          2735 => x"f7",
          2736 => x"f0",
          2737 => x"33",
          2738 => x"f0",
          2739 => x"08",
          2740 => x"f0",
          2741 => x"33",
          2742 => x"d5",
          2743 => x"05",
          2744 => x"f0",
          2745 => x"08",
          2746 => x"05",
          2747 => x"08",
          2748 => x"55",
          2749 => x"82",
          2750 => x"f8",
          2751 => x"a5",
          2752 => x"f0",
          2753 => x"33",
          2754 => x"2e",
          2755 => x"d5",
          2756 => x"05",
          2757 => x"d5",
          2758 => x"05",
          2759 => x"f0",
          2760 => x"08",
          2761 => x"08",
          2762 => x"71",
          2763 => x"0b",
          2764 => x"08",
          2765 => x"82",
          2766 => x"ec",
          2767 => x"d5",
          2768 => x"3d",
          2769 => x"f0",
          2770 => x"3d",
          2771 => x"08",
          2772 => x"59",
          2773 => x"80",
          2774 => x"39",
          2775 => x"0c",
          2776 => x"54",
          2777 => x"74",
          2778 => x"a0",
          2779 => x"06",
          2780 => x"15",
          2781 => x"80",
          2782 => x"29",
          2783 => x"05",
          2784 => x"56",
          2785 => x"82",
          2786 => x"82",
          2787 => x"54",
          2788 => x"08",
          2789 => x"fc",
          2790 => x"e4",
          2791 => x"84",
          2792 => x"73",
          2793 => x"b4",
          2794 => x"70",
          2795 => x"58",
          2796 => x"27",
          2797 => x"54",
          2798 => x"e4",
          2799 => x"0d",
          2800 => x"0d",
          2801 => x"93",
          2802 => x"38",
          2803 => x"82",
          2804 => x"52",
          2805 => x"82",
          2806 => x"81",
          2807 => x"b3",
          2808 => x"f9",
          2809 => x"b8",
          2810 => x"39",
          2811 => x"51",
          2812 => x"82",
          2813 => x"80",
          2814 => x"b3",
          2815 => x"dd",
          2816 => x"fc",
          2817 => x"39",
          2818 => x"51",
          2819 => x"82",
          2820 => x"80",
          2821 => x"b4",
          2822 => x"c1",
          2823 => x"d4",
          2824 => x"82",
          2825 => x"b5",
          2826 => x"84",
          2827 => x"82",
          2828 => x"a9",
          2829 => x"bc",
          2830 => x"82",
          2831 => x"9d",
          2832 => x"ec",
          2833 => x"82",
          2834 => x"91",
          2835 => x"9c",
          2836 => x"82",
          2837 => x"85",
          2838 => x"c0",
          2839 => x"3f",
          2840 => x"04",
          2841 => x"77",
          2842 => x"74",
          2843 => x"8a",
          2844 => x"75",
          2845 => x"51",
          2846 => x"e8",
          2847 => x"ef",
          2848 => x"d5",
          2849 => x"75",
          2850 => x"3f",
          2851 => x"08",
          2852 => x"75",
          2853 => x"d0",
          2854 => x"be",
          2855 => x"0d",
          2856 => x"0d",
          2857 => x"05",
          2858 => x"33",
          2859 => x"68",
          2860 => x"7a",
          2861 => x"51",
          2862 => x"78",
          2863 => x"ff",
          2864 => x"81",
          2865 => x"07",
          2866 => x"06",
          2867 => x"56",
          2868 => x"38",
          2869 => x"52",
          2870 => x"52",
          2871 => x"f9",
          2872 => x"e4",
          2873 => x"d5",
          2874 => x"38",
          2875 => x"08",
          2876 => x"88",
          2877 => x"e4",
          2878 => x"3d",
          2879 => x"84",
          2880 => x"52",
          2881 => x"96",
          2882 => x"d5",
          2883 => x"82",
          2884 => x"90",
          2885 => x"74",
          2886 => x"38",
          2887 => x"19",
          2888 => x"39",
          2889 => x"05",
          2890 => x"ad",
          2891 => x"70",
          2892 => x"25",
          2893 => x"9f",
          2894 => x"51",
          2895 => x"74",
          2896 => x"38",
          2897 => x"53",
          2898 => x"88",
          2899 => x"51",
          2900 => x"76",
          2901 => x"d5",
          2902 => x"3d",
          2903 => x"3d",
          2904 => x"84",
          2905 => x"33",
          2906 => x"58",
          2907 => x"52",
          2908 => x"ad",
          2909 => x"e4",
          2910 => x"76",
          2911 => x"38",
          2912 => x"9c",
          2913 => x"82",
          2914 => x"61",
          2915 => x"82",
          2916 => x"7f",
          2917 => x"78",
          2918 => x"e4",
          2919 => x"39",
          2920 => x"82",
          2921 => x"8a",
          2922 => x"f3",
          2923 => x"61",
          2924 => x"05",
          2925 => x"33",
          2926 => x"68",
          2927 => x"5c",
          2928 => x"7a",
          2929 => x"fc",
          2930 => x"8e",
          2931 => x"84",
          2932 => x"86",
          2933 => x"74",
          2934 => x"80",
          2935 => x"2e",
          2936 => x"a0",
          2937 => x"80",
          2938 => x"18",
          2939 => x"27",
          2940 => x"22",
          2941 => x"88",
          2942 => x"de",
          2943 => x"82",
          2944 => x"ff",
          2945 => x"82",
          2946 => x"c3",
          2947 => x"53",
          2948 => x"8e",
          2949 => x"52",
          2950 => x"51",
          2951 => x"3f",
          2952 => x"b7",
          2953 => x"b7",
          2954 => x"15",
          2955 => x"74",
          2956 => x"7a",
          2957 => x"72",
          2958 => x"b7",
          2959 => x"b7",
          2960 => x"39",
          2961 => x"51",
          2962 => x"3f",
          2963 => x"82",
          2964 => x"52",
          2965 => x"dc",
          2966 => x"39",
          2967 => x"51",
          2968 => x"3f",
          2969 => x"79",
          2970 => x"38",
          2971 => x"33",
          2972 => x"56",
          2973 => x"83",
          2974 => x"80",
          2975 => x"27",
          2976 => x"53",
          2977 => x"70",
          2978 => x"51",
          2979 => x"2e",
          2980 => x"80",
          2981 => x"38",
          2982 => x"08",
          2983 => x"88",
          2984 => x"c8",
          2985 => x"51",
          2986 => x"81",
          2987 => x"b6",
          2988 => x"ac",
          2989 => x"3f",
          2990 => x"1c",
          2991 => x"8a",
          2992 => x"e4",
          2993 => x"70",
          2994 => x"57",
          2995 => x"09",
          2996 => x"38",
          2997 => x"82",
          2998 => x"98",
          2999 => x"2c",
          3000 => x"70",
          3001 => x"32",
          3002 => x"72",
          3003 => x"07",
          3004 => x"58",
          3005 => x"57",
          3006 => x"d8",
          3007 => x"2e",
          3008 => x"85",
          3009 => x"8c",
          3010 => x"53",
          3011 => x"fd",
          3012 => x"53",
          3013 => x"e4",
          3014 => x"0d",
          3015 => x"0d",
          3016 => x"33",
          3017 => x"53",
          3018 => x"52",
          3019 => x"aa",
          3020 => x"b4",
          3021 => x"e3",
          3022 => x"c0",
          3023 => x"cc",
          3024 => x"b5",
          3025 => x"b7",
          3026 => x"b5",
          3027 => x"80",
          3028 => x"a1",
          3029 => x"3d",
          3030 => x"3d",
          3031 => x"96",
          3032 => x"a5",
          3033 => x"51",
          3034 => x"82",
          3035 => x"99",
          3036 => x"51",
          3037 => x"72",
          3038 => x"81",
          3039 => x"71",
          3040 => x"38",
          3041 => x"af",
          3042 => x"88",
          3043 => x"3f",
          3044 => x"a3",
          3045 => x"2a",
          3046 => x"51",
          3047 => x"2e",
          3048 => x"51",
          3049 => x"82",
          3050 => x"99",
          3051 => x"51",
          3052 => x"72",
          3053 => x"81",
          3054 => x"71",
          3055 => x"38",
          3056 => x"f3",
          3057 => x"a8",
          3058 => x"3f",
          3059 => x"e7",
          3060 => x"2a",
          3061 => x"51",
          3062 => x"2e",
          3063 => x"51",
          3064 => x"82",
          3065 => x"98",
          3066 => x"51",
          3067 => x"72",
          3068 => x"81",
          3069 => x"71",
          3070 => x"38",
          3071 => x"b7",
          3072 => x"d0",
          3073 => x"3f",
          3074 => x"ab",
          3075 => x"2a",
          3076 => x"51",
          3077 => x"2e",
          3078 => x"51",
          3079 => x"82",
          3080 => x"98",
          3081 => x"51",
          3082 => x"72",
          3083 => x"81",
          3084 => x"71",
          3085 => x"38",
          3086 => x"fb",
          3087 => x"f8",
          3088 => x"3f",
          3089 => x"ef",
          3090 => x"2a",
          3091 => x"51",
          3092 => x"2e",
          3093 => x"51",
          3094 => x"82",
          3095 => x"97",
          3096 => x"51",
          3097 => x"a4",
          3098 => x"3d",
          3099 => x"3d",
          3100 => x"84",
          3101 => x"33",
          3102 => x"56",
          3103 => x"51",
          3104 => x"0b",
          3105 => x"d8",
          3106 => x"a9",
          3107 => x"82",
          3108 => x"82",
          3109 => x"81",
          3110 => x"82",
          3111 => x"30",
          3112 => x"e4",
          3113 => x"25",
          3114 => x"51",
          3115 => x"0b",
          3116 => x"d8",
          3117 => x"82",
          3118 => x"54",
          3119 => x"09",
          3120 => x"38",
          3121 => x"53",
          3122 => x"51",
          3123 => x"3f",
          3124 => x"08",
          3125 => x"38",
          3126 => x"08",
          3127 => x"3f",
          3128 => x"ec",
          3129 => x"96",
          3130 => x"0b",
          3131 => x"d0",
          3132 => x"0b",
          3133 => x"33",
          3134 => x"2e",
          3135 => x"8c",
          3136 => x"d8",
          3137 => x"75",
          3138 => x"3f",
          3139 => x"d5",
          3140 => x"3d",
          3141 => x"3d",
          3142 => x"41",
          3143 => x"82",
          3144 => x"5f",
          3145 => x"51",
          3146 => x"3f",
          3147 => x"08",
          3148 => x"59",
          3149 => x"09",
          3150 => x"38",
          3151 => x"83",
          3152 => x"e4",
          3153 => x"db",
          3154 => x"53",
          3155 => x"d7",
          3156 => x"88",
          3157 => x"d5",
          3158 => x"2e",
          3159 => x"b9",
          3160 => x"df",
          3161 => x"41",
          3162 => x"a0",
          3163 => x"ea",
          3164 => x"70",
          3165 => x"f8",
          3166 => x"fd",
          3167 => x"3d",
          3168 => x"51",
          3169 => x"82",
          3170 => x"90",
          3171 => x"2c",
          3172 => x"80",
          3173 => x"a3",
          3174 => x"c2",
          3175 => x"78",
          3176 => x"d2",
          3177 => x"24",
          3178 => x"80",
          3179 => x"38",
          3180 => x"80",
          3181 => x"d6",
          3182 => x"c0",
          3183 => x"38",
          3184 => x"24",
          3185 => x"78",
          3186 => x"8c",
          3187 => x"39",
          3188 => x"2e",
          3189 => x"78",
          3190 => x"92",
          3191 => x"c3",
          3192 => x"38",
          3193 => x"2e",
          3194 => x"8a",
          3195 => x"81",
          3196 => x"88",
          3197 => x"83",
          3198 => x"78",
          3199 => x"89",
          3200 => x"8a",
          3201 => x"85",
          3202 => x"38",
          3203 => x"b5",
          3204 => x"11",
          3205 => x"05",
          3206 => x"3f",
          3207 => x"08",
          3208 => x"c5",
          3209 => x"fe",
          3210 => x"ff",
          3211 => x"ec",
          3212 => x"d5",
          3213 => x"2e",
          3214 => x"b5",
          3215 => x"11",
          3216 => x"05",
          3217 => x"3f",
          3218 => x"08",
          3219 => x"d5",
          3220 => x"82",
          3221 => x"ff",
          3222 => x"64",
          3223 => x"79",
          3224 => x"ec",
          3225 => x"78",
          3226 => x"05",
          3227 => x"7a",
          3228 => x"81",
          3229 => x"3d",
          3230 => x"53",
          3231 => x"51",
          3232 => x"82",
          3233 => x"80",
          3234 => x"38",
          3235 => x"fc",
          3236 => x"84",
          3237 => x"e1",
          3238 => x"e4",
          3239 => x"fd",
          3240 => x"3d",
          3241 => x"53",
          3242 => x"51",
          3243 => x"82",
          3244 => x"80",
          3245 => x"38",
          3246 => x"51",
          3247 => x"3f",
          3248 => x"64",
          3249 => x"38",
          3250 => x"70",
          3251 => x"33",
          3252 => x"81",
          3253 => x"39",
          3254 => x"80",
          3255 => x"84",
          3256 => x"95",
          3257 => x"e4",
          3258 => x"fc",
          3259 => x"3d",
          3260 => x"53",
          3261 => x"51",
          3262 => x"82",
          3263 => x"80",
          3264 => x"38",
          3265 => x"f8",
          3266 => x"84",
          3267 => x"e9",
          3268 => x"e4",
          3269 => x"fc",
          3270 => x"ba",
          3271 => x"ad",
          3272 => x"5a",
          3273 => x"a8",
          3274 => x"33",
          3275 => x"5a",
          3276 => x"2e",
          3277 => x"55",
          3278 => x"33",
          3279 => x"82",
          3280 => x"ff",
          3281 => x"81",
          3282 => x"05",
          3283 => x"39",
          3284 => x"b3",
          3285 => x"39",
          3286 => x"80",
          3287 => x"84",
          3288 => x"95",
          3289 => x"e4",
          3290 => x"38",
          3291 => x"33",
          3292 => x"2e",
          3293 => x"d4",
          3294 => x"80",
          3295 => x"d4",
          3296 => x"78",
          3297 => x"38",
          3298 => x"08",
          3299 => x"82",
          3300 => x"59",
          3301 => x"88",
          3302 => x"90",
          3303 => x"39",
          3304 => x"33",
          3305 => x"2e",
          3306 => x"d4",
          3307 => x"9a",
          3308 => x"c6",
          3309 => x"80",
          3310 => x"82",
          3311 => x"45",
          3312 => x"d4",
          3313 => x"80",
          3314 => x"3d",
          3315 => x"53",
          3316 => x"51",
          3317 => x"82",
          3318 => x"80",
          3319 => x"d4",
          3320 => x"78",
          3321 => x"38",
          3322 => x"08",
          3323 => x"39",
          3324 => x"33",
          3325 => x"2e",
          3326 => x"d4",
          3327 => x"bb",
          3328 => x"ca",
          3329 => x"80",
          3330 => x"82",
          3331 => x"44",
          3332 => x"d4",
          3333 => x"78",
          3334 => x"38",
          3335 => x"08",
          3336 => x"82",
          3337 => x"59",
          3338 => x"88",
          3339 => x"a4",
          3340 => x"39",
          3341 => x"08",
          3342 => x"b5",
          3343 => x"11",
          3344 => x"05",
          3345 => x"3f",
          3346 => x"08",
          3347 => x"38",
          3348 => x"5c",
          3349 => x"83",
          3350 => x"7a",
          3351 => x"30",
          3352 => x"9f",
          3353 => x"06",
          3354 => x"5a",
          3355 => x"88",
          3356 => x"2e",
          3357 => x"43",
          3358 => x"51",
          3359 => x"a0",
          3360 => x"62",
          3361 => x"64",
          3362 => x"3f",
          3363 => x"51",
          3364 => x"b5",
          3365 => x"11",
          3366 => x"05",
          3367 => x"3f",
          3368 => x"08",
          3369 => x"c1",
          3370 => x"fe",
          3371 => x"ff",
          3372 => x"e7",
          3373 => x"d5",
          3374 => x"2e",
          3375 => x"59",
          3376 => x"05",
          3377 => x"64",
          3378 => x"b5",
          3379 => x"11",
          3380 => x"05",
          3381 => x"3f",
          3382 => x"08",
          3383 => x"89",
          3384 => x"33",
          3385 => x"bb",
          3386 => x"a9",
          3387 => x"f1",
          3388 => x"80",
          3389 => x"51",
          3390 => x"3f",
          3391 => x"33",
          3392 => x"2e",
          3393 => x"9f",
          3394 => x"38",
          3395 => x"fc",
          3396 => x"84",
          3397 => x"e1",
          3398 => x"e4",
          3399 => x"91",
          3400 => x"02",
          3401 => x"33",
          3402 => x"81",
          3403 => x"b1",
          3404 => x"90",
          3405 => x"3f",
          3406 => x"b5",
          3407 => x"11",
          3408 => x"05",
          3409 => x"3f",
          3410 => x"08",
          3411 => x"99",
          3412 => x"fe",
          3413 => x"ff",
          3414 => x"e0",
          3415 => x"d5",
          3416 => x"2e",
          3417 => x"59",
          3418 => x"05",
          3419 => x"82",
          3420 => x"78",
          3421 => x"fe",
          3422 => x"ff",
          3423 => x"e0",
          3424 => x"d5",
          3425 => x"38",
          3426 => x"61",
          3427 => x"52",
          3428 => x"51",
          3429 => x"3f",
          3430 => x"08",
          3431 => x"52",
          3432 => x"a9",
          3433 => x"46",
          3434 => x"78",
          3435 => x"b9",
          3436 => x"26",
          3437 => x"82",
          3438 => x"39",
          3439 => x"f0",
          3440 => x"84",
          3441 => x"e0",
          3442 => x"e4",
          3443 => x"93",
          3444 => x"02",
          3445 => x"22",
          3446 => x"05",
          3447 => x"42",
          3448 => x"82",
          3449 => x"c3",
          3450 => x"9f",
          3451 => x"fe",
          3452 => x"ff",
          3453 => x"df",
          3454 => x"d5",
          3455 => x"2e",
          3456 => x"b5",
          3457 => x"11",
          3458 => x"05",
          3459 => x"3f",
          3460 => x"08",
          3461 => x"38",
          3462 => x"0c",
          3463 => x"05",
          3464 => x"fe",
          3465 => x"ff",
          3466 => x"de",
          3467 => x"d5",
          3468 => x"38",
          3469 => x"61",
          3470 => x"52",
          3471 => x"51",
          3472 => x"3f",
          3473 => x"08",
          3474 => x"52",
          3475 => x"a7",
          3476 => x"46",
          3477 => x"78",
          3478 => x"8d",
          3479 => x"27",
          3480 => x"3d",
          3481 => x"53",
          3482 => x"51",
          3483 => x"82",
          3484 => x"80",
          3485 => x"61",
          3486 => x"59",
          3487 => x"42",
          3488 => x"82",
          3489 => x"c2",
          3490 => x"ab",
          3491 => x"ff",
          3492 => x"ff",
          3493 => x"e3",
          3494 => x"d5",
          3495 => x"2e",
          3496 => x"64",
          3497 => x"b0",
          3498 => x"ae",
          3499 => x"78",
          3500 => x"ff",
          3501 => x"ff",
          3502 => x"e3",
          3503 => x"d5",
          3504 => x"2e",
          3505 => x"64",
          3506 => x"cc",
          3507 => x"8a",
          3508 => x"78",
          3509 => x"e4",
          3510 => x"f5",
          3511 => x"d5",
          3512 => x"82",
          3513 => x"ff",
          3514 => x"f4",
          3515 => x"bc",
          3516 => x"f1",
          3517 => x"c3",
          3518 => x"39",
          3519 => x"51",
          3520 => x"80",
          3521 => x"39",
          3522 => x"f4",
          3523 => x"3d",
          3524 => x"80",
          3525 => x"38",
          3526 => x"79",
          3527 => x"3f",
          3528 => x"08",
          3529 => x"e4",
          3530 => x"82",
          3531 => x"d5",
          3532 => x"b5",
          3533 => x"05",
          3534 => x"3f",
          3535 => x"08",
          3536 => x"5a",
          3537 => x"2e",
          3538 => x"82",
          3539 => x"51",
          3540 => x"82",
          3541 => x"8f",
          3542 => x"38",
          3543 => x"82",
          3544 => x"7a",
          3545 => x"38",
          3546 => x"8c",
          3547 => x"39",
          3548 => x"ad",
          3549 => x"39",
          3550 => x"56",
          3551 => x"bc",
          3552 => x"53",
          3553 => x"52",
          3554 => x"b0",
          3555 => x"a7",
          3556 => x"39",
          3557 => x"3d",
          3558 => x"51",
          3559 => x"ab",
          3560 => x"82",
          3561 => x"80",
          3562 => x"cc",
          3563 => x"ff",
          3564 => x"ff",
          3565 => x"93",
          3566 => x"80",
          3567 => x"d8",
          3568 => x"ff",
          3569 => x"ff",
          3570 => x"82",
          3571 => x"82",
          3572 => x"7c",
          3573 => x"80",
          3574 => x"80",
          3575 => x"80",
          3576 => x"ff",
          3577 => x"ea",
          3578 => x"d5",
          3579 => x"d5",
          3580 => x"70",
          3581 => x"07",
          3582 => x"5b",
          3583 => x"5a",
          3584 => x"83",
          3585 => x"78",
          3586 => x"78",
          3587 => x"38",
          3588 => x"81",
          3589 => x"59",
          3590 => x"38",
          3591 => x"7e",
          3592 => x"59",
          3593 => x"7e",
          3594 => x"81",
          3595 => x"82",
          3596 => x"ff",
          3597 => x"7c",
          3598 => x"3f",
          3599 => x"82",
          3600 => x"ff",
          3601 => x"f2",
          3602 => x"3d",
          3603 => x"82",
          3604 => x"87",
          3605 => x"70",
          3606 => x"87",
          3607 => x"72",
          3608 => x"3f",
          3609 => x"08",
          3610 => x"08",
          3611 => x"84",
          3612 => x"51",
          3613 => x"72",
          3614 => x"08",
          3615 => x"87",
          3616 => x"70",
          3617 => x"87",
          3618 => x"72",
          3619 => x"3f",
          3620 => x"08",
          3621 => x"08",
          3622 => x"84",
          3623 => x"51",
          3624 => x"72",
          3625 => x"08",
          3626 => x"8c",
          3627 => x"87",
          3628 => x"0c",
          3629 => x"0b",
          3630 => x"94",
          3631 => x"cd",
          3632 => x"b9",
          3633 => x"84",
          3634 => x"34",
          3635 => x"f1",
          3636 => x"3d",
          3637 => x"0c",
          3638 => x"82",
          3639 => x"54",
          3640 => x"92",
          3641 => x"bd",
          3642 => x"bd",
          3643 => x"bd",
          3644 => x"bd",
          3645 => x"de",
          3646 => x"e3",
          3647 => x"ec",
          3648 => x"92",
          3649 => x"fe",
          3650 => x"52",
          3651 => x"88",
          3652 => x"d8",
          3653 => x"e4",
          3654 => x"06",
          3655 => x"14",
          3656 => x"80",
          3657 => x"71",
          3658 => x"0c",
          3659 => x"04",
          3660 => x"76",
          3661 => x"55",
          3662 => x"54",
          3663 => x"81",
          3664 => x"33",
          3665 => x"2e",
          3666 => x"86",
          3667 => x"53",
          3668 => x"33",
          3669 => x"2e",
          3670 => x"86",
          3671 => x"53",
          3672 => x"52",
          3673 => x"09",
          3674 => x"38",
          3675 => x"12",
          3676 => x"33",
          3677 => x"a2",
          3678 => x"81",
          3679 => x"2e",
          3680 => x"ea",
          3681 => x"81",
          3682 => x"72",
          3683 => x"70",
          3684 => x"38",
          3685 => x"80",
          3686 => x"73",
          3687 => x"72",
          3688 => x"70",
          3689 => x"81",
          3690 => x"81",
          3691 => x"32",
          3692 => x"80",
          3693 => x"51",
          3694 => x"80",
          3695 => x"80",
          3696 => x"05",
          3697 => x"75",
          3698 => x"70",
          3699 => x"0c",
          3700 => x"04",
          3701 => x"76",
          3702 => x"80",
          3703 => x"86",
          3704 => x"52",
          3705 => x"c0",
          3706 => x"e4",
          3707 => x"80",
          3708 => x"74",
          3709 => x"d5",
          3710 => x"3d",
          3711 => x"3d",
          3712 => x"11",
          3713 => x"52",
          3714 => x"70",
          3715 => x"98",
          3716 => x"33",
          3717 => x"82",
          3718 => x"26",
          3719 => x"84",
          3720 => x"83",
          3721 => x"26",
          3722 => x"85",
          3723 => x"84",
          3724 => x"26",
          3725 => x"86",
          3726 => x"85",
          3727 => x"26",
          3728 => x"88",
          3729 => x"86",
          3730 => x"e7",
          3731 => x"38",
          3732 => x"54",
          3733 => x"87",
          3734 => x"cc",
          3735 => x"87",
          3736 => x"0c",
          3737 => x"c0",
          3738 => x"82",
          3739 => x"c0",
          3740 => x"83",
          3741 => x"c0",
          3742 => x"84",
          3743 => x"c0",
          3744 => x"85",
          3745 => x"c0",
          3746 => x"86",
          3747 => x"c0",
          3748 => x"74",
          3749 => x"a4",
          3750 => x"c0",
          3751 => x"80",
          3752 => x"98",
          3753 => x"52",
          3754 => x"e4",
          3755 => x"0d",
          3756 => x"0d",
          3757 => x"c0",
          3758 => x"81",
          3759 => x"c0",
          3760 => x"5e",
          3761 => x"87",
          3762 => x"08",
          3763 => x"1c",
          3764 => x"98",
          3765 => x"79",
          3766 => x"87",
          3767 => x"08",
          3768 => x"1c",
          3769 => x"98",
          3770 => x"79",
          3771 => x"87",
          3772 => x"08",
          3773 => x"1c",
          3774 => x"98",
          3775 => x"7b",
          3776 => x"87",
          3777 => x"08",
          3778 => x"1c",
          3779 => x"0c",
          3780 => x"ff",
          3781 => x"83",
          3782 => x"58",
          3783 => x"57",
          3784 => x"56",
          3785 => x"55",
          3786 => x"54",
          3787 => x"53",
          3788 => x"ff",
          3789 => x"bd",
          3790 => x"9d",
          3791 => x"3d",
          3792 => x"3d",
          3793 => x"05",
          3794 => x"fc",
          3795 => x"ff",
          3796 => x"55",
          3797 => x"84",
          3798 => x"2e",
          3799 => x"c0",
          3800 => x"70",
          3801 => x"2a",
          3802 => x"53",
          3803 => x"80",
          3804 => x"71",
          3805 => x"81",
          3806 => x"70",
          3807 => x"81",
          3808 => x"06",
          3809 => x"80",
          3810 => x"71",
          3811 => x"81",
          3812 => x"70",
          3813 => x"73",
          3814 => x"51",
          3815 => x"80",
          3816 => x"2e",
          3817 => x"c0",
          3818 => x"74",
          3819 => x"82",
          3820 => x"87",
          3821 => x"ff",
          3822 => x"8f",
          3823 => x"30",
          3824 => x"51",
          3825 => x"82",
          3826 => x"83",
          3827 => x"f9",
          3828 => x"a7",
          3829 => x"77",
          3830 => x"81",
          3831 => x"7a",
          3832 => x"eb",
          3833 => x"fc",
          3834 => x"ff",
          3835 => x"87",
          3836 => x"53",
          3837 => x"86",
          3838 => x"94",
          3839 => x"08",
          3840 => x"70",
          3841 => x"56",
          3842 => x"2e",
          3843 => x"91",
          3844 => x"06",
          3845 => x"d7",
          3846 => x"32",
          3847 => x"51",
          3848 => x"2e",
          3849 => x"93",
          3850 => x"06",
          3851 => x"ff",
          3852 => x"81",
          3853 => x"87",
          3854 => x"54",
          3855 => x"86",
          3856 => x"94",
          3857 => x"74",
          3858 => x"82",
          3859 => x"89",
          3860 => x"f9",
          3861 => x"54",
          3862 => x"70",
          3863 => x"53",
          3864 => x"77",
          3865 => x"38",
          3866 => x"06",
          3867 => x"d3",
          3868 => x"81",
          3869 => x"57",
          3870 => x"c0",
          3871 => x"75",
          3872 => x"38",
          3873 => x"94",
          3874 => x"70",
          3875 => x"81",
          3876 => x"52",
          3877 => x"8c",
          3878 => x"2a",
          3879 => x"51",
          3880 => x"38",
          3881 => x"70",
          3882 => x"51",
          3883 => x"8d",
          3884 => x"2a",
          3885 => x"51",
          3886 => x"be",
          3887 => x"ff",
          3888 => x"c0",
          3889 => x"70",
          3890 => x"38",
          3891 => x"90",
          3892 => x"0c",
          3893 => x"33",
          3894 => x"06",
          3895 => x"70",
          3896 => x"76",
          3897 => x"0c",
          3898 => x"04",
          3899 => x"82",
          3900 => x"70",
          3901 => x"54",
          3902 => x"94",
          3903 => x"80",
          3904 => x"87",
          3905 => x"51",
          3906 => x"82",
          3907 => x"06",
          3908 => x"70",
          3909 => x"38",
          3910 => x"06",
          3911 => x"94",
          3912 => x"80",
          3913 => x"87",
          3914 => x"52",
          3915 => x"81",
          3916 => x"d5",
          3917 => x"84",
          3918 => x"ff",
          3919 => x"d5",
          3920 => x"ff",
          3921 => x"e4",
          3922 => x"3d",
          3923 => x"fc",
          3924 => x"ff",
          3925 => x"87",
          3926 => x"52",
          3927 => x"86",
          3928 => x"94",
          3929 => x"08",
          3930 => x"70",
          3931 => x"51",
          3932 => x"70",
          3933 => x"38",
          3934 => x"06",
          3935 => x"94",
          3936 => x"80",
          3937 => x"87",
          3938 => x"52",
          3939 => x"98",
          3940 => x"2c",
          3941 => x"71",
          3942 => x"0c",
          3943 => x"04",
          3944 => x"87",
          3945 => x"08",
          3946 => x"8a",
          3947 => x"70",
          3948 => x"b4",
          3949 => x"9e",
          3950 => x"d4",
          3951 => x"c0",
          3952 => x"82",
          3953 => x"87",
          3954 => x"08",
          3955 => x"0c",
          3956 => x"98",
          3957 => x"8c",
          3958 => x"9e",
          3959 => x"d4",
          3960 => x"c0",
          3961 => x"82",
          3962 => x"87",
          3963 => x"08",
          3964 => x"0c",
          3965 => x"b0",
          3966 => x"9c",
          3967 => x"9e",
          3968 => x"d4",
          3969 => x"c0",
          3970 => x"82",
          3971 => x"87",
          3972 => x"08",
          3973 => x"0c",
          3974 => x"c0",
          3975 => x"ac",
          3976 => x"9e",
          3977 => x"d4",
          3978 => x"c0",
          3979 => x"51",
          3980 => x"b4",
          3981 => x"9e",
          3982 => x"d4",
          3983 => x"c0",
          3984 => x"82",
          3985 => x"87",
          3986 => x"08",
          3987 => x"0c",
          3988 => x"d4",
          3989 => x"0b",
          3990 => x"90",
          3991 => x"80",
          3992 => x"52",
          3993 => x"2e",
          3994 => x"52",
          3995 => x"c5",
          3996 => x"87",
          3997 => x"08",
          3998 => x"0a",
          3999 => x"52",
          4000 => x"83",
          4001 => x"71",
          4002 => x"34",
          4003 => x"c0",
          4004 => x"70",
          4005 => x"06",
          4006 => x"70",
          4007 => x"38",
          4008 => x"82",
          4009 => x"80",
          4010 => x"9e",
          4011 => x"88",
          4012 => x"51",
          4013 => x"80",
          4014 => x"81",
          4015 => x"d4",
          4016 => x"0b",
          4017 => x"90",
          4018 => x"80",
          4019 => x"52",
          4020 => x"2e",
          4021 => x"52",
          4022 => x"c9",
          4023 => x"87",
          4024 => x"08",
          4025 => x"80",
          4026 => x"52",
          4027 => x"83",
          4028 => x"71",
          4029 => x"34",
          4030 => x"c0",
          4031 => x"70",
          4032 => x"06",
          4033 => x"70",
          4034 => x"38",
          4035 => x"82",
          4036 => x"80",
          4037 => x"9e",
          4038 => x"82",
          4039 => x"51",
          4040 => x"80",
          4041 => x"81",
          4042 => x"d4",
          4043 => x"0b",
          4044 => x"90",
          4045 => x"80",
          4046 => x"52",
          4047 => x"2e",
          4048 => x"52",
          4049 => x"cd",
          4050 => x"87",
          4051 => x"08",
          4052 => x"80",
          4053 => x"52",
          4054 => x"83",
          4055 => x"71",
          4056 => x"34",
          4057 => x"c0",
          4058 => x"70",
          4059 => x"51",
          4060 => x"80",
          4061 => x"81",
          4062 => x"d4",
          4063 => x"c0",
          4064 => x"70",
          4065 => x"70",
          4066 => x"51",
          4067 => x"d4",
          4068 => x"0b",
          4069 => x"90",
          4070 => x"80",
          4071 => x"52",
          4072 => x"83",
          4073 => x"71",
          4074 => x"34",
          4075 => x"90",
          4076 => x"f0",
          4077 => x"2a",
          4078 => x"70",
          4079 => x"34",
          4080 => x"c0",
          4081 => x"70",
          4082 => x"52",
          4083 => x"2e",
          4084 => x"52",
          4085 => x"d3",
          4086 => x"9e",
          4087 => x"87",
          4088 => x"70",
          4089 => x"34",
          4090 => x"04",
          4091 => x"82",
          4092 => x"ff",
          4093 => x"82",
          4094 => x"54",
          4095 => x"89",
          4096 => x"ec",
          4097 => x"d2",
          4098 => x"80",
          4099 => x"d5",
          4100 => x"c6",
          4101 => x"80",
          4102 => x"82",
          4103 => x"82",
          4104 => x"11",
          4105 => x"be",
          4106 => x"93",
          4107 => x"d4",
          4108 => x"73",
          4109 => x"38",
          4110 => x"08",
          4111 => x"08",
          4112 => x"82",
          4113 => x"ff",
          4114 => x"82",
          4115 => x"54",
          4116 => x"94",
          4117 => x"80",
          4118 => x"84",
          4119 => x"52",
          4120 => x"51",
          4121 => x"3f",
          4122 => x"33",
          4123 => x"2e",
          4124 => x"d4",
          4125 => x"d4",
          4126 => x"54",
          4127 => x"ec",
          4128 => x"d6",
          4129 => x"ca",
          4130 => x"80",
          4131 => x"82",
          4132 => x"82",
          4133 => x"11",
          4134 => x"bf",
          4135 => x"92",
          4136 => x"d4",
          4137 => x"73",
          4138 => x"38",
          4139 => x"33",
          4140 => x"a4",
          4141 => x"a2",
          4142 => x"d3",
          4143 => x"80",
          4144 => x"82",
          4145 => x"52",
          4146 => x"51",
          4147 => x"3f",
          4148 => x"33",
          4149 => x"2e",
          4150 => x"d4",
          4151 => x"82",
          4152 => x"ff",
          4153 => x"82",
          4154 => x"54",
          4155 => x"89",
          4156 => x"84",
          4157 => x"ed",
          4158 => x"c7",
          4159 => x"80",
          4160 => x"82",
          4161 => x"ff",
          4162 => x"82",
          4163 => x"54",
          4164 => x"89",
          4165 => x"a4",
          4166 => x"c9",
          4167 => x"cd",
          4168 => x"80",
          4169 => x"82",
          4170 => x"ff",
          4171 => x"82",
          4172 => x"54",
          4173 => x"89",
          4174 => x"b8",
          4175 => x"a5",
          4176 => x"c0",
          4177 => x"9d",
          4178 => x"a8",
          4179 => x"c0",
          4180 => x"91",
          4181 => x"d4",
          4182 => x"82",
          4183 => x"ff",
          4184 => x"82",
          4185 => x"52",
          4186 => x"51",
          4187 => x"3f",
          4188 => x"51",
          4189 => x"3f",
          4190 => x"22",
          4191 => x"cc",
          4192 => x"d6",
          4193 => x"b8",
          4194 => x"84",
          4195 => x"51",
          4196 => x"82",
          4197 => x"bd",
          4198 => x"76",
          4199 => x"54",
          4200 => x"08",
          4201 => x"f4",
          4202 => x"ae",
          4203 => x"cb",
          4204 => x"80",
          4205 => x"82",
          4206 => x"56",
          4207 => x"52",
          4208 => x"ec",
          4209 => x"e4",
          4210 => x"c0",
          4211 => x"31",
          4212 => x"d5",
          4213 => x"82",
          4214 => x"ff",
          4215 => x"82",
          4216 => x"54",
          4217 => x"a9",
          4218 => x"c0",
          4219 => x"84",
          4220 => x"51",
          4221 => x"82",
          4222 => x"bd",
          4223 => x"76",
          4224 => x"54",
          4225 => x"08",
          4226 => x"cc",
          4227 => x"ca",
          4228 => x"ff",
          4229 => x"87",
          4230 => x"fe",
          4231 => x"92",
          4232 => x"05",
          4233 => x"26",
          4234 => x"84",
          4235 => x"fc",
          4236 => x"08",
          4237 => x"f8",
          4238 => x"82",
          4239 => x"97",
          4240 => x"88",
          4241 => x"82",
          4242 => x"8b",
          4243 => x"94",
          4244 => x"82",
          4245 => x"ff",
          4246 => x"84",
          4247 => x"71",
          4248 => x"04",
          4249 => x"c0",
          4250 => x"04",
          4251 => x"08",
          4252 => x"84",
          4253 => x"3d",
          4254 => x"2b",
          4255 => x"79",
          4256 => x"98",
          4257 => x"13",
          4258 => x"51",
          4259 => x"51",
          4260 => x"82",
          4261 => x"33",
          4262 => x"74",
          4263 => x"82",
          4264 => x"08",
          4265 => x"05",
          4266 => x"71",
          4267 => x"52",
          4268 => x"09",
          4269 => x"38",
          4270 => x"82",
          4271 => x"85",
          4272 => x"fb",
          4273 => x"02",
          4274 => x"05",
          4275 => x"55",
          4276 => x"80",
          4277 => x"82",
          4278 => x"52",
          4279 => x"ad",
          4280 => x"f1",
          4281 => x"a0",
          4282 => x"c8",
          4283 => x"c8",
          4284 => x"51",
          4285 => x"3f",
          4286 => x"05",
          4287 => x"34",
          4288 => x"06",
          4289 => x"77",
          4290 => x"ce",
          4291 => x"34",
          4292 => x"04",
          4293 => x"7c",
          4294 => x"b7",
          4295 => x"88",
          4296 => x"33",
          4297 => x"33",
          4298 => x"82",
          4299 => x"70",
          4300 => x"59",
          4301 => x"74",
          4302 => x"38",
          4303 => x"fb",
          4304 => x"b4",
          4305 => x"29",
          4306 => x"05",
          4307 => x"54",
          4308 => x"9d",
          4309 => x"d5",
          4310 => x"0c",
          4311 => x"33",
          4312 => x"82",
          4313 => x"70",
          4314 => x"5a",
          4315 => x"a7",
          4316 => x"78",
          4317 => x"ff",
          4318 => x"82",
          4319 => x"81",
          4320 => x"82",
          4321 => x"74",
          4322 => x"55",
          4323 => x"87",
          4324 => x"82",
          4325 => x"77",
          4326 => x"38",
          4327 => x"08",
          4328 => x"2e",
          4329 => x"d5",
          4330 => x"74",
          4331 => x"3d",
          4332 => x"76",
          4333 => x"75",
          4334 => x"82",
          4335 => x"b0",
          4336 => x"51",
          4337 => x"3f",
          4338 => x"08",
          4339 => x"e6",
          4340 => x"0d",
          4341 => x"0d",
          4342 => x"53",
          4343 => x"08",
          4344 => x"2e",
          4345 => x"51",
          4346 => x"80",
          4347 => x"14",
          4348 => x"54",
          4349 => x"e6",
          4350 => x"82",
          4351 => x"82",
          4352 => x"52",
          4353 => x"95",
          4354 => x"80",
          4355 => x"82",
          4356 => x"51",
          4357 => x"80",
          4358 => x"b0",
          4359 => x"0d",
          4360 => x"0d",
          4361 => x"52",
          4362 => x"08",
          4363 => x"e7",
          4364 => x"e4",
          4365 => x"38",
          4366 => x"08",
          4367 => x"52",
          4368 => x"52",
          4369 => x"bf",
          4370 => x"e4",
          4371 => x"ba",
          4372 => x"ff",
          4373 => x"82",
          4374 => x"55",
          4375 => x"d5",
          4376 => x"9d",
          4377 => x"e4",
          4378 => x"70",
          4379 => x"80",
          4380 => x"53",
          4381 => x"17",
          4382 => x"52",
          4383 => x"da",
          4384 => x"2e",
          4385 => x"ff",
          4386 => x"3d",
          4387 => x"3d",
          4388 => x"08",
          4389 => x"5a",
          4390 => x"58",
          4391 => x"82",
          4392 => x"51",
          4393 => x"3f",
          4394 => x"08",
          4395 => x"ff",
          4396 => x"b0",
          4397 => x"80",
          4398 => x"3d",
          4399 => x"81",
          4400 => x"82",
          4401 => x"80",
          4402 => x"75",
          4403 => x"b7",
          4404 => x"e4",
          4405 => x"58",
          4406 => x"82",
          4407 => x"25",
          4408 => x"d5",
          4409 => x"05",
          4410 => x"55",
          4411 => x"74",
          4412 => x"70",
          4413 => x"2a",
          4414 => x"78",
          4415 => x"38",
          4416 => x"38",
          4417 => x"08",
          4418 => x"53",
          4419 => x"87",
          4420 => x"e4",
          4421 => x"89",
          4422 => x"a4",
          4423 => x"ba",
          4424 => x"2e",
          4425 => x"9b",
          4426 => x"79",
          4427 => x"c5",
          4428 => x"ff",
          4429 => x"ab",
          4430 => x"82",
          4431 => x"74",
          4432 => x"77",
          4433 => x"0c",
          4434 => x"04",
          4435 => x"7c",
          4436 => x"71",
          4437 => x"59",
          4438 => x"a0",
          4439 => x"06",
          4440 => x"33",
          4441 => x"77",
          4442 => x"38",
          4443 => x"5b",
          4444 => x"56",
          4445 => x"a0",
          4446 => x"06",
          4447 => x"75",
          4448 => x"80",
          4449 => x"29",
          4450 => x"05",
          4451 => x"55",
          4452 => x"3f",
          4453 => x"08",
          4454 => x"74",
          4455 => x"b3",
          4456 => x"d5",
          4457 => x"c5",
          4458 => x"33",
          4459 => x"2e",
          4460 => x"82",
          4461 => x"b5",
          4462 => x"3f",
          4463 => x"1a",
          4464 => x"fc",
          4465 => x"05",
          4466 => x"3f",
          4467 => x"08",
          4468 => x"38",
          4469 => x"78",
          4470 => x"fd",
          4471 => x"d5",
          4472 => x"ff",
          4473 => x"85",
          4474 => x"91",
          4475 => x"70",
          4476 => x"51",
          4477 => x"27",
          4478 => x"80",
          4479 => x"d5",
          4480 => x"3d",
          4481 => x"3d",
          4482 => x"08",
          4483 => x"b4",
          4484 => x"5f",
          4485 => x"af",
          4486 => x"d5",
          4487 => x"d5",
          4488 => x"5b",
          4489 => x"38",
          4490 => x"ac",
          4491 => x"73",
          4492 => x"55",
          4493 => x"81",
          4494 => x"70",
          4495 => x"56",
          4496 => x"81",
          4497 => x"51",
          4498 => x"82",
          4499 => x"82",
          4500 => x"82",
          4501 => x"80",
          4502 => x"38",
          4503 => x"52",
          4504 => x"08",
          4505 => x"f1",
          4506 => x"e4",
          4507 => x"8c",
          4508 => x"d0",
          4509 => x"ed",
          4510 => x"39",
          4511 => x"08",
          4512 => x"b0",
          4513 => x"f8",
          4514 => x"70",
          4515 => x"9a",
          4516 => x"d5",
          4517 => x"82",
          4518 => x"74",
          4519 => x"06",
          4520 => x"82",
          4521 => x"51",
          4522 => x"3f",
          4523 => x"08",
          4524 => x"82",
          4525 => x"25",
          4526 => x"d5",
          4527 => x"05",
          4528 => x"55",
          4529 => x"80",
          4530 => x"ff",
          4531 => x"51",
          4532 => x"81",
          4533 => x"ff",
          4534 => x"93",
          4535 => x"38",
          4536 => x"ff",
          4537 => x"06",
          4538 => x"86",
          4539 => x"d5",
          4540 => x"8c",
          4541 => x"b0",
          4542 => x"84",
          4543 => x"3f",
          4544 => x"ec",
          4545 => x"d5",
          4546 => x"2b",
          4547 => x"51",
          4548 => x"2e",
          4549 => x"81",
          4550 => x"ed",
          4551 => x"98",
          4552 => x"2c",
          4553 => x"33",
          4554 => x"70",
          4555 => x"98",
          4556 => x"84",
          4557 => x"a4",
          4558 => x"15",
          4559 => x"51",
          4560 => x"59",
          4561 => x"58",
          4562 => x"78",
          4563 => x"38",
          4564 => x"b4",
          4565 => x"80",
          4566 => x"ff",
          4567 => x"98",
          4568 => x"80",
          4569 => x"ce",
          4570 => x"74",
          4571 => x"f6",
          4572 => x"d5",
          4573 => x"ff",
          4574 => x"80",
          4575 => x"74",
          4576 => x"34",
          4577 => x"39",
          4578 => x"0a",
          4579 => x"0a",
          4580 => x"2c",
          4581 => x"06",
          4582 => x"73",
          4583 => x"38",
          4584 => x"52",
          4585 => x"ce",
          4586 => x"e4",
          4587 => x"06",
          4588 => x"38",
          4589 => x"56",
          4590 => x"80",
          4591 => x"1c",
          4592 => x"ed",
          4593 => x"98",
          4594 => x"2c",
          4595 => x"33",
          4596 => x"70",
          4597 => x"10",
          4598 => x"2b",
          4599 => x"11",
          4600 => x"51",
          4601 => x"51",
          4602 => x"2e",
          4603 => x"fe",
          4604 => x"c3",
          4605 => x"7d",
          4606 => x"82",
          4607 => x"80",
          4608 => x"9c",
          4609 => x"75",
          4610 => x"34",
          4611 => x"9c",
          4612 => x"3d",
          4613 => x"0c",
          4614 => x"95",
          4615 => x"38",
          4616 => x"82",
          4617 => x"54",
          4618 => x"82",
          4619 => x"54",
          4620 => x"fd",
          4621 => x"ed",
          4622 => x"73",
          4623 => x"38",
          4624 => x"70",
          4625 => x"55",
          4626 => x"9e",
          4627 => x"54",
          4628 => x"15",
          4629 => x"80",
          4630 => x"ff",
          4631 => x"98",
          4632 => x"a8",
          4633 => x"55",
          4634 => x"ed",
          4635 => x"11",
          4636 => x"82",
          4637 => x"73",
          4638 => x"3d",
          4639 => x"82",
          4640 => x"54",
          4641 => x"89",
          4642 => x"54",
          4643 => x"a4",
          4644 => x"a8",
          4645 => x"80",
          4646 => x"ff",
          4647 => x"98",
          4648 => x"a4",
          4649 => x"56",
          4650 => x"25",
          4651 => x"f1",
          4652 => x"74",
          4653 => x"52",
          4654 => x"f8",
          4655 => x"80",
          4656 => x"80",
          4657 => x"98",
          4658 => x"a4",
          4659 => x"55",
          4660 => x"da",
          4661 => x"a8",
          4662 => x"2b",
          4663 => x"82",
          4664 => x"5a",
          4665 => x"74",
          4666 => x"94",
          4667 => x"c8",
          4668 => x"51",
          4669 => x"3f",
          4670 => x"0a",
          4671 => x"0a",
          4672 => x"2c",
          4673 => x"33",
          4674 => x"73",
          4675 => x"38",
          4676 => x"83",
          4677 => x"0b",
          4678 => x"82",
          4679 => x"80",
          4680 => x"f0",
          4681 => x"3f",
          4682 => x"82",
          4683 => x"70",
          4684 => x"55",
          4685 => x"2e",
          4686 => x"82",
          4687 => x"ff",
          4688 => x"82",
          4689 => x"ff",
          4690 => x"82",
          4691 => x"82",
          4692 => x"52",
          4693 => x"a0",
          4694 => x"ed",
          4695 => x"98",
          4696 => x"2c",
          4697 => x"33",
          4698 => x"57",
          4699 => x"ad",
          4700 => x"54",
          4701 => x"74",
          4702 => x"c8",
          4703 => x"33",
          4704 => x"b0",
          4705 => x"80",
          4706 => x"80",
          4707 => x"98",
          4708 => x"a4",
          4709 => x"55",
          4710 => x"d5",
          4711 => x"c8",
          4712 => x"51",
          4713 => x"3f",
          4714 => x"33",
          4715 => x"70",
          4716 => x"ed",
          4717 => x"51",
          4718 => x"74",
          4719 => x"38",
          4720 => x"08",
          4721 => x"ff",
          4722 => x"74",
          4723 => x"29",
          4724 => x"05",
          4725 => x"82",
          4726 => x"58",
          4727 => x"75",
          4728 => x"fa",
          4729 => x"ed",
          4730 => x"05",
          4731 => x"34",
          4732 => x"08",
          4733 => x"ff",
          4734 => x"82",
          4735 => x"79",
          4736 => x"3f",
          4737 => x"08",
          4738 => x"54",
          4739 => x"82",
          4740 => x"54",
          4741 => x"8f",
          4742 => x"73",
          4743 => x"f1",
          4744 => x"39",
          4745 => x"80",
          4746 => x"a8",
          4747 => x"82",
          4748 => x"79",
          4749 => x"0c",
          4750 => x"04",
          4751 => x"33",
          4752 => x"2e",
          4753 => x"82",
          4754 => x"52",
          4755 => x"9e",
          4756 => x"ed",
          4757 => x"05",
          4758 => x"ed",
          4759 => x"81",
          4760 => x"dd",
          4761 => x"a8",
          4762 => x"a4",
          4763 => x"73",
          4764 => x"8c",
          4765 => x"54",
          4766 => x"a4",
          4767 => x"2b",
          4768 => x"75",
          4769 => x"56",
          4770 => x"74",
          4771 => x"74",
          4772 => x"14",
          4773 => x"82",
          4774 => x"52",
          4775 => x"ff",
          4776 => x"74",
          4777 => x"29",
          4778 => x"05",
          4779 => x"82",
          4780 => x"58",
          4781 => x"75",
          4782 => x"82",
          4783 => x"52",
          4784 => x"9d",
          4785 => x"ed",
          4786 => x"98",
          4787 => x"2c",
          4788 => x"33",
          4789 => x"57",
          4790 => x"f8",
          4791 => x"f1",
          4792 => x"88",
          4793 => x"cc",
          4794 => x"80",
          4795 => x"80",
          4796 => x"98",
          4797 => x"a4",
          4798 => x"55",
          4799 => x"de",
          4800 => x"39",
          4801 => x"33",
          4802 => x"06",
          4803 => x"33",
          4804 => x"74",
          4805 => x"e8",
          4806 => x"c8",
          4807 => x"14",
          4808 => x"ed",
          4809 => x"1a",
          4810 => x"54",
          4811 => x"3f",
          4812 => x"33",
          4813 => x"06",
          4814 => x"33",
          4815 => x"75",
          4816 => x"38",
          4817 => x"82",
          4818 => x"80",
          4819 => x"f0",
          4820 => x"3f",
          4821 => x"ed",
          4822 => x"0b",
          4823 => x"34",
          4824 => x"7a",
          4825 => x"d5",
          4826 => x"74",
          4827 => x"38",
          4828 => x"a5",
          4829 => x"d5",
          4830 => x"ed",
          4831 => x"d5",
          4832 => x"ff",
          4833 => x"53",
          4834 => x"51",
          4835 => x"3f",
          4836 => x"c0",
          4837 => x"29",
          4838 => x"05",
          4839 => x"56",
          4840 => x"2e",
          4841 => x"51",
          4842 => x"3f",
          4843 => x"08",
          4844 => x"34",
          4845 => x"08",
          4846 => x"81",
          4847 => x"52",
          4848 => x"a6",
          4849 => x"1b",
          4850 => x"39",
          4851 => x"74",
          4852 => x"ac",
          4853 => x"ff",
          4854 => x"99",
          4855 => x"2e",
          4856 => x"ae",
          4857 => x"dc",
          4858 => x"80",
          4859 => x"74",
          4860 => x"93",
          4861 => x"e4",
          4862 => x"a4",
          4863 => x"e4",
          4864 => x"06",
          4865 => x"74",
          4866 => x"ff",
          4867 => x"80",
          4868 => x"84",
          4869 => x"e0",
          4870 => x"56",
          4871 => x"2e",
          4872 => x"51",
          4873 => x"3f",
          4874 => x"08",
          4875 => x"34",
          4876 => x"08",
          4877 => x"81",
          4878 => x"52",
          4879 => x"a5",
          4880 => x"1b",
          4881 => x"ff",
          4882 => x"39",
          4883 => x"a4",
          4884 => x"34",
          4885 => x"53",
          4886 => x"33",
          4887 => x"ec",
          4888 => x"9c",
          4889 => x"a8",
          4890 => x"ff",
          4891 => x"a4",
          4892 => x"54",
          4893 => x"f5",
          4894 => x"f1",
          4895 => x"81",
          4896 => x"82",
          4897 => x"74",
          4898 => x"52",
          4899 => x"a4",
          4900 => x"39",
          4901 => x"33",
          4902 => x"2e",
          4903 => x"82",
          4904 => x"52",
          4905 => x"9a",
          4906 => x"ed",
          4907 => x"05",
          4908 => x"ed",
          4909 => x"c8",
          4910 => x"0d",
          4911 => x"0b",
          4912 => x"0c",
          4913 => x"82",
          4914 => x"82",
          4915 => x"80",
          4916 => x"f4",
          4917 => x"bb",
          4918 => x"d4",
          4919 => x"58",
          4920 => x"81",
          4921 => x"15",
          4922 => x"d4",
          4923 => x"84",
          4924 => x"85",
          4925 => x"d5",
          4926 => x"77",
          4927 => x"76",
          4928 => x"82",
          4929 => x"82",
          4930 => x"ff",
          4931 => x"80",
          4932 => x"ff",
          4933 => x"88",
          4934 => x"55",
          4935 => x"17",
          4936 => x"17",
          4937 => x"d0",
          4938 => x"29",
          4939 => x"08",
          4940 => x"51",
          4941 => x"82",
          4942 => x"83",
          4943 => x"3d",
          4944 => x"3d",
          4945 => x"81",
          4946 => x"27",
          4947 => x"12",
          4948 => x"11",
          4949 => x"ff",
          4950 => x"51",
          4951 => x"e4",
          4952 => x"0d",
          4953 => x"0d",
          4954 => x"22",
          4955 => x"aa",
          4956 => x"05",
          4957 => x"08",
          4958 => x"71",
          4959 => x"2b",
          4960 => x"33",
          4961 => x"71",
          4962 => x"02",
          4963 => x"05",
          4964 => x"ff",
          4965 => x"70",
          4966 => x"51",
          4967 => x"5b",
          4968 => x"54",
          4969 => x"34",
          4970 => x"34",
          4971 => x"08",
          4972 => x"2a",
          4973 => x"82",
          4974 => x"83",
          4975 => x"d5",
          4976 => x"17",
          4977 => x"12",
          4978 => x"2b",
          4979 => x"2b",
          4980 => x"06",
          4981 => x"52",
          4982 => x"83",
          4983 => x"70",
          4984 => x"54",
          4985 => x"12",
          4986 => x"ff",
          4987 => x"83",
          4988 => x"d5",
          4989 => x"56",
          4990 => x"72",
          4991 => x"89",
          4992 => x"fb",
          4993 => x"d5",
          4994 => x"84",
          4995 => x"22",
          4996 => x"72",
          4997 => x"33",
          4998 => x"71",
          4999 => x"83",
          5000 => x"5b",
          5001 => x"52",
          5002 => x"12",
          5003 => x"33",
          5004 => x"07",
          5005 => x"54",
          5006 => x"70",
          5007 => x"73",
          5008 => x"82",
          5009 => x"70",
          5010 => x"33",
          5011 => x"71",
          5012 => x"83",
          5013 => x"59",
          5014 => x"05",
          5015 => x"87",
          5016 => x"88",
          5017 => x"88",
          5018 => x"56",
          5019 => x"13",
          5020 => x"13",
          5021 => x"d4",
          5022 => x"33",
          5023 => x"71",
          5024 => x"70",
          5025 => x"06",
          5026 => x"53",
          5027 => x"53",
          5028 => x"70",
          5029 => x"87",
          5030 => x"fa",
          5031 => x"a2",
          5032 => x"d5",
          5033 => x"83",
          5034 => x"70",
          5035 => x"33",
          5036 => x"07",
          5037 => x"15",
          5038 => x"12",
          5039 => x"2b",
          5040 => x"07",
          5041 => x"55",
          5042 => x"57",
          5043 => x"80",
          5044 => x"38",
          5045 => x"ab",
          5046 => x"d4",
          5047 => x"70",
          5048 => x"33",
          5049 => x"71",
          5050 => x"74",
          5051 => x"81",
          5052 => x"88",
          5053 => x"83",
          5054 => x"f8",
          5055 => x"54",
          5056 => x"58",
          5057 => x"74",
          5058 => x"52",
          5059 => x"34",
          5060 => x"34",
          5061 => x"08",
          5062 => x"33",
          5063 => x"71",
          5064 => x"83",
          5065 => x"59",
          5066 => x"05",
          5067 => x"12",
          5068 => x"2b",
          5069 => x"ff",
          5070 => x"88",
          5071 => x"52",
          5072 => x"74",
          5073 => x"15",
          5074 => x"0d",
          5075 => x"0d",
          5076 => x"08",
          5077 => x"9e",
          5078 => x"83",
          5079 => x"82",
          5080 => x"12",
          5081 => x"2b",
          5082 => x"07",
          5083 => x"52",
          5084 => x"05",
          5085 => x"13",
          5086 => x"2b",
          5087 => x"05",
          5088 => x"71",
          5089 => x"2a",
          5090 => x"53",
          5091 => x"34",
          5092 => x"34",
          5093 => x"08",
          5094 => x"33",
          5095 => x"71",
          5096 => x"83",
          5097 => x"59",
          5098 => x"05",
          5099 => x"83",
          5100 => x"88",
          5101 => x"88",
          5102 => x"56",
          5103 => x"13",
          5104 => x"13",
          5105 => x"d4",
          5106 => x"11",
          5107 => x"33",
          5108 => x"07",
          5109 => x"0c",
          5110 => x"3d",
          5111 => x"3d",
          5112 => x"d5",
          5113 => x"83",
          5114 => x"ff",
          5115 => x"53",
          5116 => x"a7",
          5117 => x"d4",
          5118 => x"2b",
          5119 => x"11",
          5120 => x"33",
          5121 => x"71",
          5122 => x"75",
          5123 => x"81",
          5124 => x"98",
          5125 => x"2b",
          5126 => x"40",
          5127 => x"58",
          5128 => x"72",
          5129 => x"38",
          5130 => x"52",
          5131 => x"9d",
          5132 => x"39",
          5133 => x"85",
          5134 => x"8b",
          5135 => x"2b",
          5136 => x"79",
          5137 => x"51",
          5138 => x"76",
          5139 => x"75",
          5140 => x"56",
          5141 => x"34",
          5142 => x"08",
          5143 => x"12",
          5144 => x"33",
          5145 => x"07",
          5146 => x"54",
          5147 => x"53",
          5148 => x"34",
          5149 => x"34",
          5150 => x"08",
          5151 => x"0b",
          5152 => x"80",
          5153 => x"34",
          5154 => x"08",
          5155 => x"14",
          5156 => x"14",
          5157 => x"d4",
          5158 => x"33",
          5159 => x"71",
          5160 => x"70",
          5161 => x"07",
          5162 => x"53",
          5163 => x"54",
          5164 => x"72",
          5165 => x"8b",
          5166 => x"ff",
          5167 => x"52",
          5168 => x"08",
          5169 => x"f1",
          5170 => x"2e",
          5171 => x"51",
          5172 => x"83",
          5173 => x"f5",
          5174 => x"7e",
          5175 => x"e2",
          5176 => x"e4",
          5177 => x"ff",
          5178 => x"d4",
          5179 => x"33",
          5180 => x"71",
          5181 => x"70",
          5182 => x"58",
          5183 => x"ff",
          5184 => x"2e",
          5185 => x"75",
          5186 => x"70",
          5187 => x"33",
          5188 => x"07",
          5189 => x"ff",
          5190 => x"70",
          5191 => x"06",
          5192 => x"52",
          5193 => x"59",
          5194 => x"27",
          5195 => x"80",
          5196 => x"75",
          5197 => x"84",
          5198 => x"16",
          5199 => x"2b",
          5200 => x"75",
          5201 => x"81",
          5202 => x"85",
          5203 => x"59",
          5204 => x"83",
          5205 => x"d4",
          5206 => x"33",
          5207 => x"71",
          5208 => x"70",
          5209 => x"06",
          5210 => x"56",
          5211 => x"75",
          5212 => x"81",
          5213 => x"79",
          5214 => x"cc",
          5215 => x"74",
          5216 => x"c4",
          5217 => x"2e",
          5218 => x"89",
          5219 => x"f8",
          5220 => x"ac",
          5221 => x"80",
          5222 => x"75",
          5223 => x"3f",
          5224 => x"08",
          5225 => x"11",
          5226 => x"33",
          5227 => x"71",
          5228 => x"53",
          5229 => x"74",
          5230 => x"70",
          5231 => x"06",
          5232 => x"5c",
          5233 => x"78",
          5234 => x"76",
          5235 => x"57",
          5236 => x"34",
          5237 => x"08",
          5238 => x"71",
          5239 => x"86",
          5240 => x"12",
          5241 => x"2b",
          5242 => x"2a",
          5243 => x"53",
          5244 => x"73",
          5245 => x"75",
          5246 => x"82",
          5247 => x"70",
          5248 => x"33",
          5249 => x"71",
          5250 => x"83",
          5251 => x"5d",
          5252 => x"05",
          5253 => x"15",
          5254 => x"15",
          5255 => x"d4",
          5256 => x"71",
          5257 => x"33",
          5258 => x"71",
          5259 => x"70",
          5260 => x"5a",
          5261 => x"54",
          5262 => x"34",
          5263 => x"34",
          5264 => x"08",
          5265 => x"54",
          5266 => x"e4",
          5267 => x"0d",
          5268 => x"0d",
          5269 => x"d5",
          5270 => x"38",
          5271 => x"71",
          5272 => x"2e",
          5273 => x"51",
          5274 => x"82",
          5275 => x"53",
          5276 => x"e4",
          5277 => x"0d",
          5278 => x"0d",
          5279 => x"5c",
          5280 => x"40",
          5281 => x"08",
          5282 => x"81",
          5283 => x"f4",
          5284 => x"8e",
          5285 => x"ff",
          5286 => x"d5",
          5287 => x"83",
          5288 => x"8b",
          5289 => x"fc",
          5290 => x"54",
          5291 => x"7e",
          5292 => x"3f",
          5293 => x"08",
          5294 => x"06",
          5295 => x"08",
          5296 => x"83",
          5297 => x"ff",
          5298 => x"83",
          5299 => x"70",
          5300 => x"33",
          5301 => x"07",
          5302 => x"70",
          5303 => x"06",
          5304 => x"fc",
          5305 => x"29",
          5306 => x"81",
          5307 => x"88",
          5308 => x"90",
          5309 => x"4e",
          5310 => x"52",
          5311 => x"41",
          5312 => x"5b",
          5313 => x"8f",
          5314 => x"ff",
          5315 => x"31",
          5316 => x"ff",
          5317 => x"82",
          5318 => x"17",
          5319 => x"2b",
          5320 => x"29",
          5321 => x"81",
          5322 => x"98",
          5323 => x"2b",
          5324 => x"45",
          5325 => x"73",
          5326 => x"38",
          5327 => x"70",
          5328 => x"06",
          5329 => x"7b",
          5330 => x"38",
          5331 => x"73",
          5332 => x"81",
          5333 => x"78",
          5334 => x"3f",
          5335 => x"ff",
          5336 => x"e5",
          5337 => x"38",
          5338 => x"89",
          5339 => x"f6",
          5340 => x"a5",
          5341 => x"55",
          5342 => x"80",
          5343 => x"1d",
          5344 => x"83",
          5345 => x"88",
          5346 => x"57",
          5347 => x"3f",
          5348 => x"51",
          5349 => x"82",
          5350 => x"83",
          5351 => x"7e",
          5352 => x"70",
          5353 => x"d5",
          5354 => x"84",
          5355 => x"59",
          5356 => x"3f",
          5357 => x"08",
          5358 => x"75",
          5359 => x"06",
          5360 => x"85",
          5361 => x"54",
          5362 => x"80",
          5363 => x"51",
          5364 => x"82",
          5365 => x"1d",
          5366 => x"83",
          5367 => x"88",
          5368 => x"43",
          5369 => x"3f",
          5370 => x"51",
          5371 => x"82",
          5372 => x"83",
          5373 => x"7e",
          5374 => x"70",
          5375 => x"d5",
          5376 => x"84",
          5377 => x"59",
          5378 => x"3f",
          5379 => x"08",
          5380 => x"60",
          5381 => x"55",
          5382 => x"ff",
          5383 => x"a9",
          5384 => x"52",
          5385 => x"3f",
          5386 => x"08",
          5387 => x"e4",
          5388 => x"93",
          5389 => x"73",
          5390 => x"e4",
          5391 => x"95",
          5392 => x"51",
          5393 => x"7a",
          5394 => x"27",
          5395 => x"53",
          5396 => x"51",
          5397 => x"7a",
          5398 => x"82",
          5399 => x"05",
          5400 => x"f6",
          5401 => x"54",
          5402 => x"e4",
          5403 => x"0d",
          5404 => x"0d",
          5405 => x"70",
          5406 => x"d5",
          5407 => x"e4",
          5408 => x"d5",
          5409 => x"2e",
          5410 => x"53",
          5411 => x"d5",
          5412 => x"ff",
          5413 => x"74",
          5414 => x"0c",
          5415 => x"04",
          5416 => x"02",
          5417 => x"51",
          5418 => x"72",
          5419 => x"82",
          5420 => x"33",
          5421 => x"d5",
          5422 => x"3d",
          5423 => x"3d",
          5424 => x"05",
          5425 => x"05",
          5426 => x"56",
          5427 => x"72",
          5428 => x"e0",
          5429 => x"2b",
          5430 => x"8c",
          5431 => x"88",
          5432 => x"2e",
          5433 => x"88",
          5434 => x"0c",
          5435 => x"8c",
          5436 => x"71",
          5437 => x"87",
          5438 => x"0c",
          5439 => x"08",
          5440 => x"51",
          5441 => x"2e",
          5442 => x"c0",
          5443 => x"51",
          5444 => x"71",
          5445 => x"80",
          5446 => x"92",
          5447 => x"98",
          5448 => x"70",
          5449 => x"38",
          5450 => x"e0",
          5451 => x"d5",
          5452 => x"51",
          5453 => x"e4",
          5454 => x"0d",
          5455 => x"0d",
          5456 => x"02",
          5457 => x"05",
          5458 => x"58",
          5459 => x"52",
          5460 => x"3f",
          5461 => x"08",
          5462 => x"54",
          5463 => x"be",
          5464 => x"75",
          5465 => x"c0",
          5466 => x"87",
          5467 => x"12",
          5468 => x"84",
          5469 => x"40",
          5470 => x"85",
          5471 => x"98",
          5472 => x"7d",
          5473 => x"0c",
          5474 => x"85",
          5475 => x"06",
          5476 => x"71",
          5477 => x"38",
          5478 => x"71",
          5479 => x"05",
          5480 => x"19",
          5481 => x"a2",
          5482 => x"71",
          5483 => x"38",
          5484 => x"83",
          5485 => x"38",
          5486 => x"8a",
          5487 => x"98",
          5488 => x"71",
          5489 => x"c0",
          5490 => x"52",
          5491 => x"87",
          5492 => x"80",
          5493 => x"81",
          5494 => x"c0",
          5495 => x"53",
          5496 => x"82",
          5497 => x"71",
          5498 => x"1a",
          5499 => x"84",
          5500 => x"19",
          5501 => x"06",
          5502 => x"79",
          5503 => x"38",
          5504 => x"80",
          5505 => x"87",
          5506 => x"26",
          5507 => x"73",
          5508 => x"06",
          5509 => x"2e",
          5510 => x"52",
          5511 => x"82",
          5512 => x"8f",
          5513 => x"f3",
          5514 => x"62",
          5515 => x"05",
          5516 => x"57",
          5517 => x"83",
          5518 => x"52",
          5519 => x"3f",
          5520 => x"08",
          5521 => x"54",
          5522 => x"2e",
          5523 => x"81",
          5524 => x"74",
          5525 => x"c0",
          5526 => x"87",
          5527 => x"12",
          5528 => x"84",
          5529 => x"5f",
          5530 => x"0b",
          5531 => x"8c",
          5532 => x"0c",
          5533 => x"80",
          5534 => x"70",
          5535 => x"81",
          5536 => x"54",
          5537 => x"8c",
          5538 => x"81",
          5539 => x"7c",
          5540 => x"58",
          5541 => x"70",
          5542 => x"52",
          5543 => x"8a",
          5544 => x"98",
          5545 => x"71",
          5546 => x"c0",
          5547 => x"52",
          5548 => x"87",
          5549 => x"80",
          5550 => x"81",
          5551 => x"c0",
          5552 => x"53",
          5553 => x"82",
          5554 => x"71",
          5555 => x"19",
          5556 => x"81",
          5557 => x"ff",
          5558 => x"19",
          5559 => x"78",
          5560 => x"38",
          5561 => x"80",
          5562 => x"87",
          5563 => x"26",
          5564 => x"73",
          5565 => x"06",
          5566 => x"2e",
          5567 => x"52",
          5568 => x"82",
          5569 => x"8f",
          5570 => x"fa",
          5571 => x"02",
          5572 => x"05",
          5573 => x"05",
          5574 => x"71",
          5575 => x"57",
          5576 => x"82",
          5577 => x"81",
          5578 => x"54",
          5579 => x"38",
          5580 => x"c0",
          5581 => x"81",
          5582 => x"2e",
          5583 => x"71",
          5584 => x"38",
          5585 => x"87",
          5586 => x"11",
          5587 => x"80",
          5588 => x"80",
          5589 => x"83",
          5590 => x"38",
          5591 => x"72",
          5592 => x"2a",
          5593 => x"51",
          5594 => x"80",
          5595 => x"87",
          5596 => x"08",
          5597 => x"38",
          5598 => x"8c",
          5599 => x"96",
          5600 => x"0c",
          5601 => x"8c",
          5602 => x"08",
          5603 => x"51",
          5604 => x"38",
          5605 => x"56",
          5606 => x"80",
          5607 => x"85",
          5608 => x"77",
          5609 => x"83",
          5610 => x"75",
          5611 => x"d5",
          5612 => x"3d",
          5613 => x"3d",
          5614 => x"11",
          5615 => x"71",
          5616 => x"82",
          5617 => x"53",
          5618 => x"0d",
          5619 => x"0d",
          5620 => x"33",
          5621 => x"71",
          5622 => x"88",
          5623 => x"14",
          5624 => x"07",
          5625 => x"33",
          5626 => x"d5",
          5627 => x"53",
          5628 => x"52",
          5629 => x"04",
          5630 => x"73",
          5631 => x"92",
          5632 => x"52",
          5633 => x"81",
          5634 => x"70",
          5635 => x"70",
          5636 => x"3d",
          5637 => x"3d",
          5638 => x"52",
          5639 => x"70",
          5640 => x"34",
          5641 => x"51",
          5642 => x"81",
          5643 => x"70",
          5644 => x"70",
          5645 => x"05",
          5646 => x"88",
          5647 => x"72",
          5648 => x"0d",
          5649 => x"0d",
          5650 => x"54",
          5651 => x"80",
          5652 => x"71",
          5653 => x"53",
          5654 => x"81",
          5655 => x"ff",
          5656 => x"39",
          5657 => x"04",
          5658 => x"75",
          5659 => x"52",
          5660 => x"70",
          5661 => x"34",
          5662 => x"70",
          5663 => x"3d",
          5664 => x"3d",
          5665 => x"79",
          5666 => x"74",
          5667 => x"56",
          5668 => x"81",
          5669 => x"71",
          5670 => x"16",
          5671 => x"52",
          5672 => x"86",
          5673 => x"2e",
          5674 => x"82",
          5675 => x"86",
          5676 => x"fe",
          5677 => x"76",
          5678 => x"39",
          5679 => x"8a",
          5680 => x"51",
          5681 => x"71",
          5682 => x"33",
          5683 => x"0c",
          5684 => x"04",
          5685 => x"d5",
          5686 => x"fb",
          5687 => x"70",
          5688 => x"81",
          5689 => x"70",
          5690 => x"56",
          5691 => x"55",
          5692 => x"08",
          5693 => x"80",
          5694 => x"83",
          5695 => x"51",
          5696 => x"3f",
          5697 => x"08",
          5698 => x"06",
          5699 => x"2e",
          5700 => x"76",
          5701 => x"74",
          5702 => x"0c",
          5703 => x"04",
          5704 => x"7b",
          5705 => x"83",
          5706 => x"5a",
          5707 => x"80",
          5708 => x"54",
          5709 => x"53",
          5710 => x"53",
          5711 => x"52",
          5712 => x"3f",
          5713 => x"08",
          5714 => x"81",
          5715 => x"82",
          5716 => x"83",
          5717 => x"16",
          5718 => x"18",
          5719 => x"18",
          5720 => x"58",
          5721 => x"9f",
          5722 => x"33",
          5723 => x"2e",
          5724 => x"93",
          5725 => x"76",
          5726 => x"52",
          5727 => x"51",
          5728 => x"83",
          5729 => x"79",
          5730 => x"0c",
          5731 => x"04",
          5732 => x"78",
          5733 => x"80",
          5734 => x"17",
          5735 => x"38",
          5736 => x"fc",
          5737 => x"e4",
          5738 => x"d5",
          5739 => x"38",
          5740 => x"53",
          5741 => x"81",
          5742 => x"f7",
          5743 => x"d5",
          5744 => x"2e",
          5745 => x"55",
          5746 => x"b4",
          5747 => x"82",
          5748 => x"88",
          5749 => x"f8",
          5750 => x"70",
          5751 => x"c0",
          5752 => x"e4",
          5753 => x"d5",
          5754 => x"91",
          5755 => x"55",
          5756 => x"09",
          5757 => x"f0",
          5758 => x"33",
          5759 => x"2e",
          5760 => x"80",
          5761 => x"80",
          5762 => x"e4",
          5763 => x"17",
          5764 => x"fc",
          5765 => x"d4",
          5766 => x"b6",
          5767 => x"d8",
          5768 => x"85",
          5769 => x"75",
          5770 => x"3f",
          5771 => x"e4",
          5772 => x"9c",
          5773 => x"de",
          5774 => x"08",
          5775 => x"17",
          5776 => x"3f",
          5777 => x"52",
          5778 => x"51",
          5779 => x"a4",
          5780 => x"05",
          5781 => x"0c",
          5782 => x"75",
          5783 => x"33",
          5784 => x"3f",
          5785 => x"34",
          5786 => x"52",
          5787 => x"51",
          5788 => x"82",
          5789 => x"80",
          5790 => x"81",
          5791 => x"d5",
          5792 => x"3d",
          5793 => x"3d",
          5794 => x"1a",
          5795 => x"fe",
          5796 => x"54",
          5797 => x"73",
          5798 => x"8a",
          5799 => x"71",
          5800 => x"08",
          5801 => x"75",
          5802 => x"0c",
          5803 => x"04",
          5804 => x"7a",
          5805 => x"56",
          5806 => x"77",
          5807 => x"38",
          5808 => x"08",
          5809 => x"38",
          5810 => x"54",
          5811 => x"2e",
          5812 => x"72",
          5813 => x"38",
          5814 => x"8d",
          5815 => x"39",
          5816 => x"81",
          5817 => x"b6",
          5818 => x"2a",
          5819 => x"2a",
          5820 => x"05",
          5821 => x"55",
          5822 => x"82",
          5823 => x"81",
          5824 => x"83",
          5825 => x"b8",
          5826 => x"17",
          5827 => x"a8",
          5828 => x"55",
          5829 => x"57",
          5830 => x"3f",
          5831 => x"08",
          5832 => x"74",
          5833 => x"14",
          5834 => x"70",
          5835 => x"07",
          5836 => x"71",
          5837 => x"52",
          5838 => x"72",
          5839 => x"75",
          5840 => x"58",
          5841 => x"76",
          5842 => x"15",
          5843 => x"73",
          5844 => x"3f",
          5845 => x"08",
          5846 => x"76",
          5847 => x"06",
          5848 => x"05",
          5849 => x"3f",
          5850 => x"08",
          5851 => x"06",
          5852 => x"76",
          5853 => x"15",
          5854 => x"73",
          5855 => x"3f",
          5856 => x"08",
          5857 => x"82",
          5858 => x"06",
          5859 => x"05",
          5860 => x"3f",
          5861 => x"08",
          5862 => x"58",
          5863 => x"58",
          5864 => x"e4",
          5865 => x"0d",
          5866 => x"0d",
          5867 => x"5a",
          5868 => x"59",
          5869 => x"82",
          5870 => x"9c",
          5871 => x"82",
          5872 => x"33",
          5873 => x"2e",
          5874 => x"72",
          5875 => x"38",
          5876 => x"8d",
          5877 => x"39",
          5878 => x"81",
          5879 => x"f7",
          5880 => x"2a",
          5881 => x"2a",
          5882 => x"05",
          5883 => x"55",
          5884 => x"82",
          5885 => x"59",
          5886 => x"08",
          5887 => x"74",
          5888 => x"16",
          5889 => x"16",
          5890 => x"59",
          5891 => x"53",
          5892 => x"8f",
          5893 => x"2b",
          5894 => x"74",
          5895 => x"71",
          5896 => x"72",
          5897 => x"0b",
          5898 => x"74",
          5899 => x"17",
          5900 => x"75",
          5901 => x"3f",
          5902 => x"08",
          5903 => x"e4",
          5904 => x"38",
          5905 => x"06",
          5906 => x"78",
          5907 => x"54",
          5908 => x"77",
          5909 => x"33",
          5910 => x"71",
          5911 => x"51",
          5912 => x"34",
          5913 => x"76",
          5914 => x"17",
          5915 => x"75",
          5916 => x"3f",
          5917 => x"08",
          5918 => x"e4",
          5919 => x"38",
          5920 => x"ff",
          5921 => x"10",
          5922 => x"76",
          5923 => x"51",
          5924 => x"be",
          5925 => x"2a",
          5926 => x"05",
          5927 => x"f9",
          5928 => x"d5",
          5929 => x"82",
          5930 => x"ab",
          5931 => x"0a",
          5932 => x"2b",
          5933 => x"70",
          5934 => x"70",
          5935 => x"54",
          5936 => x"82",
          5937 => x"8f",
          5938 => x"07",
          5939 => x"f6",
          5940 => x"0b",
          5941 => x"78",
          5942 => x"0c",
          5943 => x"04",
          5944 => x"7a",
          5945 => x"08",
          5946 => x"59",
          5947 => x"a4",
          5948 => x"17",
          5949 => x"38",
          5950 => x"aa",
          5951 => x"73",
          5952 => x"fd",
          5953 => x"d5",
          5954 => x"82",
          5955 => x"80",
          5956 => x"39",
          5957 => x"eb",
          5958 => x"80",
          5959 => x"d5",
          5960 => x"80",
          5961 => x"52",
          5962 => x"84",
          5963 => x"e4",
          5964 => x"d5",
          5965 => x"2e",
          5966 => x"82",
          5967 => x"81",
          5968 => x"82",
          5969 => x"ff",
          5970 => x"80",
          5971 => x"75",
          5972 => x"3f",
          5973 => x"08",
          5974 => x"16",
          5975 => x"94",
          5976 => x"55",
          5977 => x"27",
          5978 => x"15",
          5979 => x"84",
          5980 => x"07",
          5981 => x"17",
          5982 => x"76",
          5983 => x"a6",
          5984 => x"73",
          5985 => x"0c",
          5986 => x"04",
          5987 => x"7c",
          5988 => x"59",
          5989 => x"95",
          5990 => x"08",
          5991 => x"2e",
          5992 => x"17",
          5993 => x"b2",
          5994 => x"ae",
          5995 => x"7a",
          5996 => x"3f",
          5997 => x"82",
          5998 => x"27",
          5999 => x"82",
          6000 => x"55",
          6001 => x"08",
          6002 => x"d2",
          6003 => x"08",
          6004 => x"08",
          6005 => x"38",
          6006 => x"17",
          6007 => x"54",
          6008 => x"82",
          6009 => x"7a",
          6010 => x"06",
          6011 => x"81",
          6012 => x"17",
          6013 => x"83",
          6014 => x"75",
          6015 => x"f9",
          6016 => x"59",
          6017 => x"08",
          6018 => x"81",
          6019 => x"82",
          6020 => x"59",
          6021 => x"08",
          6022 => x"70",
          6023 => x"25",
          6024 => x"82",
          6025 => x"54",
          6026 => x"55",
          6027 => x"38",
          6028 => x"08",
          6029 => x"38",
          6030 => x"54",
          6031 => x"90",
          6032 => x"18",
          6033 => x"38",
          6034 => x"39",
          6035 => x"38",
          6036 => x"16",
          6037 => x"08",
          6038 => x"38",
          6039 => x"78",
          6040 => x"38",
          6041 => x"51",
          6042 => x"82",
          6043 => x"80",
          6044 => x"80",
          6045 => x"e4",
          6046 => x"09",
          6047 => x"38",
          6048 => x"08",
          6049 => x"e4",
          6050 => x"30",
          6051 => x"80",
          6052 => x"07",
          6053 => x"55",
          6054 => x"38",
          6055 => x"09",
          6056 => x"ae",
          6057 => x"80",
          6058 => x"53",
          6059 => x"51",
          6060 => x"82",
          6061 => x"82",
          6062 => x"30",
          6063 => x"e4",
          6064 => x"25",
          6065 => x"79",
          6066 => x"38",
          6067 => x"8f",
          6068 => x"79",
          6069 => x"f9",
          6070 => x"d5",
          6071 => x"74",
          6072 => x"90",
          6073 => x"17",
          6074 => x"94",
          6075 => x"54",
          6076 => x"86",
          6077 => x"94",
          6078 => x"17",
          6079 => x"54",
          6080 => x"34",
          6081 => x"56",
          6082 => x"90",
          6083 => x"80",
          6084 => x"82",
          6085 => x"55",
          6086 => x"56",
          6087 => x"82",
          6088 => x"8c",
          6089 => x"f8",
          6090 => x"70",
          6091 => x"f0",
          6092 => x"e4",
          6093 => x"56",
          6094 => x"08",
          6095 => x"7b",
          6096 => x"f6",
          6097 => x"d5",
          6098 => x"d5",
          6099 => x"17",
          6100 => x"80",
          6101 => x"b8",
          6102 => x"57",
          6103 => x"77",
          6104 => x"81",
          6105 => x"15",
          6106 => x"78",
          6107 => x"81",
          6108 => x"53",
          6109 => x"15",
          6110 => x"ab",
          6111 => x"e4",
          6112 => x"df",
          6113 => x"22",
          6114 => x"30",
          6115 => x"70",
          6116 => x"51",
          6117 => x"82",
          6118 => x"8a",
          6119 => x"f8",
          6120 => x"7c",
          6121 => x"56",
          6122 => x"80",
          6123 => x"f1",
          6124 => x"06",
          6125 => x"e9",
          6126 => x"18",
          6127 => x"08",
          6128 => x"38",
          6129 => x"82",
          6130 => x"38",
          6131 => x"54",
          6132 => x"74",
          6133 => x"82",
          6134 => x"22",
          6135 => x"79",
          6136 => x"38",
          6137 => x"98",
          6138 => x"cd",
          6139 => x"22",
          6140 => x"54",
          6141 => x"26",
          6142 => x"52",
          6143 => x"b0",
          6144 => x"e4",
          6145 => x"d5",
          6146 => x"2e",
          6147 => x"0b",
          6148 => x"08",
          6149 => x"9c",
          6150 => x"d5",
          6151 => x"85",
          6152 => x"bd",
          6153 => x"31",
          6154 => x"73",
          6155 => x"f4",
          6156 => x"d5",
          6157 => x"18",
          6158 => x"18",
          6159 => x"08",
          6160 => x"72",
          6161 => x"38",
          6162 => x"58",
          6163 => x"89",
          6164 => x"18",
          6165 => x"ff",
          6166 => x"05",
          6167 => x"80",
          6168 => x"d5",
          6169 => x"3d",
          6170 => x"3d",
          6171 => x"08",
          6172 => x"a0",
          6173 => x"54",
          6174 => x"77",
          6175 => x"80",
          6176 => x"0c",
          6177 => x"53",
          6178 => x"80",
          6179 => x"38",
          6180 => x"06",
          6181 => x"b5",
          6182 => x"98",
          6183 => x"14",
          6184 => x"92",
          6185 => x"2a",
          6186 => x"56",
          6187 => x"26",
          6188 => x"80",
          6189 => x"16",
          6190 => x"77",
          6191 => x"53",
          6192 => x"38",
          6193 => x"51",
          6194 => x"82",
          6195 => x"53",
          6196 => x"0b",
          6197 => x"08",
          6198 => x"38",
          6199 => x"d5",
          6200 => x"2e",
          6201 => x"9c",
          6202 => x"d5",
          6203 => x"80",
          6204 => x"8a",
          6205 => x"15",
          6206 => x"80",
          6207 => x"14",
          6208 => x"51",
          6209 => x"82",
          6210 => x"53",
          6211 => x"d5",
          6212 => x"2e",
          6213 => x"82",
          6214 => x"e4",
          6215 => x"ba",
          6216 => x"82",
          6217 => x"ff",
          6218 => x"82",
          6219 => x"52",
          6220 => x"f3",
          6221 => x"e4",
          6222 => x"72",
          6223 => x"72",
          6224 => x"f2",
          6225 => x"d5",
          6226 => x"15",
          6227 => x"15",
          6228 => x"b8",
          6229 => x"0c",
          6230 => x"82",
          6231 => x"8a",
          6232 => x"f7",
          6233 => x"7d",
          6234 => x"5b",
          6235 => x"76",
          6236 => x"3f",
          6237 => x"08",
          6238 => x"e4",
          6239 => x"38",
          6240 => x"08",
          6241 => x"08",
          6242 => x"f0",
          6243 => x"d5",
          6244 => x"82",
          6245 => x"80",
          6246 => x"d5",
          6247 => x"18",
          6248 => x"51",
          6249 => x"81",
          6250 => x"81",
          6251 => x"81",
          6252 => x"e4",
          6253 => x"83",
          6254 => x"77",
          6255 => x"72",
          6256 => x"38",
          6257 => x"75",
          6258 => x"81",
          6259 => x"a5",
          6260 => x"e4",
          6261 => x"52",
          6262 => x"8e",
          6263 => x"e4",
          6264 => x"d5",
          6265 => x"2e",
          6266 => x"73",
          6267 => x"81",
          6268 => x"87",
          6269 => x"d5",
          6270 => x"3d",
          6271 => x"3d",
          6272 => x"11",
          6273 => x"ae",
          6274 => x"e4",
          6275 => x"ff",
          6276 => x"33",
          6277 => x"71",
          6278 => x"81",
          6279 => x"94",
          6280 => x"92",
          6281 => x"e4",
          6282 => x"73",
          6283 => x"82",
          6284 => x"85",
          6285 => x"fc",
          6286 => x"79",
          6287 => x"ff",
          6288 => x"12",
          6289 => x"eb",
          6290 => x"70",
          6291 => x"72",
          6292 => x"81",
          6293 => x"73",
          6294 => x"94",
          6295 => x"98",
          6296 => x"0d",
          6297 => x"0d",
          6298 => x"51",
          6299 => x"81",
          6300 => x"80",
          6301 => x"70",
          6302 => x"33",
          6303 => x"81",
          6304 => x"16",
          6305 => x"51",
          6306 => x"70",
          6307 => x"0c",
          6308 => x"04",
          6309 => x"60",
          6310 => x"84",
          6311 => x"5b",
          6312 => x"5d",
          6313 => x"08",
          6314 => x"80",
          6315 => x"08",
          6316 => x"ed",
          6317 => x"d5",
          6318 => x"82",
          6319 => x"82",
          6320 => x"19",
          6321 => x"55",
          6322 => x"38",
          6323 => x"dc",
          6324 => x"33",
          6325 => x"81",
          6326 => x"53",
          6327 => x"34",
          6328 => x"08",
          6329 => x"e5",
          6330 => x"06",
          6331 => x"56",
          6332 => x"08",
          6333 => x"2e",
          6334 => x"83",
          6335 => x"75",
          6336 => x"72",
          6337 => x"d5",
          6338 => x"df",
          6339 => x"72",
          6340 => x"81",
          6341 => x"81",
          6342 => x"2e",
          6343 => x"ff",
          6344 => x"39",
          6345 => x"09",
          6346 => x"ca",
          6347 => x"2a",
          6348 => x"51",
          6349 => x"2e",
          6350 => x"15",
          6351 => x"bf",
          6352 => x"1c",
          6353 => x"0c",
          6354 => x"73",
          6355 => x"81",
          6356 => x"38",
          6357 => x"53",
          6358 => x"09",
          6359 => x"8f",
          6360 => x"08",
          6361 => x"5a",
          6362 => x"82",
          6363 => x"83",
          6364 => x"53",
          6365 => x"38",
          6366 => x"81",
          6367 => x"29",
          6368 => x"54",
          6369 => x"58",
          6370 => x"17",
          6371 => x"51",
          6372 => x"82",
          6373 => x"83",
          6374 => x"56",
          6375 => x"96",
          6376 => x"fe",
          6377 => x"38",
          6378 => x"76",
          6379 => x"73",
          6380 => x"54",
          6381 => x"83",
          6382 => x"09",
          6383 => x"38",
          6384 => x"8c",
          6385 => x"38",
          6386 => x"86",
          6387 => x"06",
          6388 => x"72",
          6389 => x"38",
          6390 => x"26",
          6391 => x"10",
          6392 => x"73",
          6393 => x"70",
          6394 => x"51",
          6395 => x"81",
          6396 => x"5c",
          6397 => x"93",
          6398 => x"fc",
          6399 => x"d5",
          6400 => x"ff",
          6401 => x"7d",
          6402 => x"ff",
          6403 => x"0c",
          6404 => x"52",
          6405 => x"d2",
          6406 => x"e4",
          6407 => x"d5",
          6408 => x"38",
          6409 => x"fd",
          6410 => x"39",
          6411 => x"1a",
          6412 => x"d5",
          6413 => x"3d",
          6414 => x"3d",
          6415 => x"08",
          6416 => x"52",
          6417 => x"d7",
          6418 => x"e4",
          6419 => x"d5",
          6420 => x"a4",
          6421 => x"70",
          6422 => x"0b",
          6423 => x"98",
          6424 => x"7e",
          6425 => x"3f",
          6426 => x"08",
          6427 => x"e4",
          6428 => x"38",
          6429 => x"70",
          6430 => x"75",
          6431 => x"58",
          6432 => x"8b",
          6433 => x"06",
          6434 => x"06",
          6435 => x"86",
          6436 => x"81",
          6437 => x"c3",
          6438 => x"2a",
          6439 => x"51",
          6440 => x"2e",
          6441 => x"82",
          6442 => x"8f",
          6443 => x"06",
          6444 => x"ab",
          6445 => x"86",
          6446 => x"06",
          6447 => x"73",
          6448 => x"75",
          6449 => x"81",
          6450 => x"73",
          6451 => x"38",
          6452 => x"76",
          6453 => x"70",
          6454 => x"ac",
          6455 => x"5d",
          6456 => x"2e",
          6457 => x"81",
          6458 => x"17",
          6459 => x"76",
          6460 => x"06",
          6461 => x"8c",
          6462 => x"18",
          6463 => x"b6",
          6464 => x"e4",
          6465 => x"ff",
          6466 => x"81",
          6467 => x"33",
          6468 => x"8d",
          6469 => x"59",
          6470 => x"5c",
          6471 => x"e4",
          6472 => x"05",
          6473 => x"3f",
          6474 => x"08",
          6475 => x"06",
          6476 => x"2e",
          6477 => x"81",
          6478 => x"e6",
          6479 => x"80",
          6480 => x"82",
          6481 => x"78",
          6482 => x"22",
          6483 => x"19",
          6484 => x"e1",
          6485 => x"82",
          6486 => x"2e",
          6487 => x"80",
          6488 => x"5a",
          6489 => x"83",
          6490 => x"09",
          6491 => x"38",
          6492 => x"8c",
          6493 => x"a5",
          6494 => x"70",
          6495 => x"81",
          6496 => x"57",
          6497 => x"90",
          6498 => x"2e",
          6499 => x"10",
          6500 => x"51",
          6501 => x"38",
          6502 => x"81",
          6503 => x"54",
          6504 => x"ff",
          6505 => x"bb",
          6506 => x"38",
          6507 => x"b5",
          6508 => x"e4",
          6509 => x"06",
          6510 => x"2e",
          6511 => x"19",
          6512 => x"54",
          6513 => x"8b",
          6514 => x"52",
          6515 => x"51",
          6516 => x"82",
          6517 => x"80",
          6518 => x"81",
          6519 => x"0b",
          6520 => x"80",
          6521 => x"f5",
          6522 => x"d5",
          6523 => x"82",
          6524 => x"80",
          6525 => x"38",
          6526 => x"e4",
          6527 => x"0d",
          6528 => x"0d",
          6529 => x"ab",
          6530 => x"a0",
          6531 => x"5a",
          6532 => x"85",
          6533 => x"8c",
          6534 => x"22",
          6535 => x"73",
          6536 => x"38",
          6537 => x"10",
          6538 => x"51",
          6539 => x"39",
          6540 => x"1a",
          6541 => x"3d",
          6542 => x"59",
          6543 => x"02",
          6544 => x"33",
          6545 => x"73",
          6546 => x"a8",
          6547 => x"0b",
          6548 => x"81",
          6549 => x"08",
          6550 => x"8b",
          6551 => x"78",
          6552 => x"3f",
          6553 => x"80",
          6554 => x"56",
          6555 => x"83",
          6556 => x"55",
          6557 => x"2e",
          6558 => x"83",
          6559 => x"82",
          6560 => x"8f",
          6561 => x"06",
          6562 => x"75",
          6563 => x"90",
          6564 => x"06",
          6565 => x"56",
          6566 => x"87",
          6567 => x"a0",
          6568 => x"ff",
          6569 => x"80",
          6570 => x"c0",
          6571 => x"87",
          6572 => x"bf",
          6573 => x"74",
          6574 => x"06",
          6575 => x"27",
          6576 => x"14",
          6577 => x"34",
          6578 => x"18",
          6579 => x"57",
          6580 => x"e3",
          6581 => x"ec",
          6582 => x"80",
          6583 => x"80",
          6584 => x"38",
          6585 => x"73",
          6586 => x"38",
          6587 => x"33",
          6588 => x"e0",
          6589 => x"e4",
          6590 => x"8c",
          6591 => x"54",
          6592 => x"94",
          6593 => x"55",
          6594 => x"74",
          6595 => x"38",
          6596 => x"33",
          6597 => x"39",
          6598 => x"05",
          6599 => x"78",
          6600 => x"56",
          6601 => x"76",
          6602 => x"38",
          6603 => x"15",
          6604 => x"55",
          6605 => x"34",
          6606 => x"e3",
          6607 => x"f9",
          6608 => x"d5",
          6609 => x"38",
          6610 => x"80",
          6611 => x"fe",
          6612 => x"55",
          6613 => x"2e",
          6614 => x"82",
          6615 => x"55",
          6616 => x"08",
          6617 => x"81",
          6618 => x"38",
          6619 => x"05",
          6620 => x"34",
          6621 => x"05",
          6622 => x"2a",
          6623 => x"51",
          6624 => x"59",
          6625 => x"90",
          6626 => x"8c",
          6627 => x"f9",
          6628 => x"d5",
          6629 => x"59",
          6630 => x"51",
          6631 => x"82",
          6632 => x"57",
          6633 => x"08",
          6634 => x"ff",
          6635 => x"80",
          6636 => x"38",
          6637 => x"90",
          6638 => x"31",
          6639 => x"51",
          6640 => x"82",
          6641 => x"57",
          6642 => x"08",
          6643 => x"a0",
          6644 => x"91",
          6645 => x"e4",
          6646 => x"06",
          6647 => x"08",
          6648 => x"e3",
          6649 => x"d5",
          6650 => x"82",
          6651 => x"81",
          6652 => x"1c",
          6653 => x"08",
          6654 => x"06",
          6655 => x"7c",
          6656 => x"8f",
          6657 => x"34",
          6658 => x"08",
          6659 => x"82",
          6660 => x"52",
          6661 => x"df",
          6662 => x"8d",
          6663 => x"77",
          6664 => x"83",
          6665 => x"8b",
          6666 => x"1b",
          6667 => x"17",
          6668 => x"73",
          6669 => x"e4",
          6670 => x"05",
          6671 => x"3f",
          6672 => x"83",
          6673 => x"81",
          6674 => x"77",
          6675 => x"73",
          6676 => x"2e",
          6677 => x"10",
          6678 => x"51",
          6679 => x"38",
          6680 => x"07",
          6681 => x"34",
          6682 => x"1d",
          6683 => x"79",
          6684 => x"3f",
          6685 => x"08",
          6686 => x"e4",
          6687 => x"38",
          6688 => x"78",
          6689 => x"98",
          6690 => x"7b",
          6691 => x"3f",
          6692 => x"08",
          6693 => x"e4",
          6694 => x"a0",
          6695 => x"e4",
          6696 => x"1a",
          6697 => x"c0",
          6698 => x"a0",
          6699 => x"1a",
          6700 => x"91",
          6701 => x"08",
          6702 => x"98",
          6703 => x"73",
          6704 => x"81",
          6705 => x"34",
          6706 => x"82",
          6707 => x"94",
          6708 => x"fa",
          6709 => x"70",
          6710 => x"08",
          6711 => x"56",
          6712 => x"72",
          6713 => x"38",
          6714 => x"51",
          6715 => x"82",
          6716 => x"54",
          6717 => x"08",
          6718 => x"98",
          6719 => x"75",
          6720 => x"3f",
          6721 => x"08",
          6722 => x"e4",
          6723 => x"9c",
          6724 => x"e5",
          6725 => x"0b",
          6726 => x"90",
          6727 => x"27",
          6728 => x"d5",
          6729 => x"74",
          6730 => x"3f",
          6731 => x"08",
          6732 => x"e4",
          6733 => x"c3",
          6734 => x"2e",
          6735 => x"83",
          6736 => x"73",
          6737 => x"0c",
          6738 => x"04",
          6739 => x"7e",
          6740 => x"5f",
          6741 => x"0b",
          6742 => x"98",
          6743 => x"2e",
          6744 => x"ac",
          6745 => x"2e",
          6746 => x"80",
          6747 => x"8c",
          6748 => x"22",
          6749 => x"5c",
          6750 => x"2e",
          6751 => x"78",
          6752 => x"22",
          6753 => x"56",
          6754 => x"38",
          6755 => x"15",
          6756 => x"ff",
          6757 => x"72",
          6758 => x"86",
          6759 => x"80",
          6760 => x"18",
          6761 => x"ff",
          6762 => x"5b",
          6763 => x"52",
          6764 => x"75",
          6765 => x"d7",
          6766 => x"d5",
          6767 => x"ff",
          6768 => x"81",
          6769 => x"95",
          6770 => x"27",
          6771 => x"88",
          6772 => x"7a",
          6773 => x"15",
          6774 => x"9f",
          6775 => x"76",
          6776 => x"07",
          6777 => x"80",
          6778 => x"54",
          6779 => x"2e",
          6780 => x"57",
          6781 => x"7a",
          6782 => x"74",
          6783 => x"5b",
          6784 => x"79",
          6785 => x"22",
          6786 => x"72",
          6787 => x"7a",
          6788 => x"25",
          6789 => x"06",
          6790 => x"77",
          6791 => x"53",
          6792 => x"14",
          6793 => x"89",
          6794 => x"57",
          6795 => x"19",
          6796 => x"1b",
          6797 => x"74",
          6798 => x"38",
          6799 => x"09",
          6800 => x"38",
          6801 => x"78",
          6802 => x"30",
          6803 => x"80",
          6804 => x"54",
          6805 => x"90",
          6806 => x"2e",
          6807 => x"76",
          6808 => x"58",
          6809 => x"57",
          6810 => x"81",
          6811 => x"81",
          6812 => x"79",
          6813 => x"38",
          6814 => x"05",
          6815 => x"81",
          6816 => x"18",
          6817 => x"81",
          6818 => x"8b",
          6819 => x"96",
          6820 => x"57",
          6821 => x"72",
          6822 => x"33",
          6823 => x"72",
          6824 => x"d3",
          6825 => x"89",
          6826 => x"73",
          6827 => x"11",
          6828 => x"99",
          6829 => x"9c",
          6830 => x"11",
          6831 => x"88",
          6832 => x"38",
          6833 => x"53",
          6834 => x"83",
          6835 => x"81",
          6836 => x"80",
          6837 => x"a0",
          6838 => x"ff",
          6839 => x"53",
          6840 => x"81",
          6841 => x"81",
          6842 => x"81",
          6843 => x"56",
          6844 => x"72",
          6845 => x"77",
          6846 => x"53",
          6847 => x"14",
          6848 => x"08",
          6849 => x"51",
          6850 => x"38",
          6851 => x"34",
          6852 => x"53",
          6853 => x"88",
          6854 => x"1c",
          6855 => x"52",
          6856 => x"3f",
          6857 => x"08",
          6858 => x"13",
          6859 => x"3f",
          6860 => x"08",
          6861 => x"98",
          6862 => x"fa",
          6863 => x"e4",
          6864 => x"23",
          6865 => x"04",
          6866 => x"62",
          6867 => x"5e",
          6868 => x"33",
          6869 => x"73",
          6870 => x"38",
          6871 => x"80",
          6872 => x"38",
          6873 => x"8d",
          6874 => x"05",
          6875 => x"0c",
          6876 => x"15",
          6877 => x"70",
          6878 => x"56",
          6879 => x"09",
          6880 => x"38",
          6881 => x"80",
          6882 => x"30",
          6883 => x"78",
          6884 => x"54",
          6885 => x"73",
          6886 => x"63",
          6887 => x"54",
          6888 => x"96",
          6889 => x"0b",
          6890 => x"80",
          6891 => x"e7",
          6892 => x"d5",
          6893 => x"87",
          6894 => x"41",
          6895 => x"11",
          6896 => x"80",
          6897 => x"fc",
          6898 => x"8f",
          6899 => x"e4",
          6900 => x"82",
          6901 => x"ff",
          6902 => x"d5",
          6903 => x"92",
          6904 => x"1a",
          6905 => x"08",
          6906 => x"55",
          6907 => x"81",
          6908 => x"d5",
          6909 => x"ff",
          6910 => x"af",
          6911 => x"9f",
          6912 => x"80",
          6913 => x"51",
          6914 => x"b4",
          6915 => x"dc",
          6916 => x"75",
          6917 => x"91",
          6918 => x"82",
          6919 => x"d9",
          6920 => x"d5",
          6921 => x"de",
          6922 => x"fe",
          6923 => x"38",
          6924 => x"54",
          6925 => x"81",
          6926 => x"89",
          6927 => x"41",
          6928 => x"33",
          6929 => x"73",
          6930 => x"81",
          6931 => x"81",
          6932 => x"dc",
          6933 => x"70",
          6934 => x"07",
          6935 => x"73",
          6936 => x"44",
          6937 => x"82",
          6938 => x"81",
          6939 => x"06",
          6940 => x"22",
          6941 => x"2e",
          6942 => x"d2",
          6943 => x"2e",
          6944 => x"80",
          6945 => x"1a",
          6946 => x"ae",
          6947 => x"06",
          6948 => x"79",
          6949 => x"ae",
          6950 => x"06",
          6951 => x"10",
          6952 => x"74",
          6953 => x"a0",
          6954 => x"ae",
          6955 => x"26",
          6956 => x"54",
          6957 => x"81",
          6958 => x"81",
          6959 => x"78",
          6960 => x"76",
          6961 => x"73",
          6962 => x"84",
          6963 => x"80",
          6964 => x"78",
          6965 => x"05",
          6966 => x"fe",
          6967 => x"a0",
          6968 => x"70",
          6969 => x"51",
          6970 => x"54",
          6971 => x"84",
          6972 => x"38",
          6973 => x"78",
          6974 => x"19",
          6975 => x"56",
          6976 => x"78",
          6977 => x"56",
          6978 => x"76",
          6979 => x"83",
          6980 => x"7a",
          6981 => x"ff",
          6982 => x"56",
          6983 => x"2e",
          6984 => x"93",
          6985 => x"70",
          6986 => x"22",
          6987 => x"73",
          6988 => x"38",
          6989 => x"74",
          6990 => x"06",
          6991 => x"2e",
          6992 => x"85",
          6993 => x"07",
          6994 => x"2e",
          6995 => x"16",
          6996 => x"22",
          6997 => x"ae",
          6998 => x"78",
          6999 => x"05",
          7000 => x"59",
          7001 => x"8f",
          7002 => x"70",
          7003 => x"73",
          7004 => x"81",
          7005 => x"8b",
          7006 => x"a0",
          7007 => x"e8",
          7008 => x"59",
          7009 => x"7c",
          7010 => x"22",
          7011 => x"57",
          7012 => x"2e",
          7013 => x"75",
          7014 => x"38",
          7015 => x"70",
          7016 => x"25",
          7017 => x"7c",
          7018 => x"38",
          7019 => x"89",
          7020 => x"07",
          7021 => x"80",
          7022 => x"7e",
          7023 => x"38",
          7024 => x"79",
          7025 => x"70",
          7026 => x"25",
          7027 => x"51",
          7028 => x"73",
          7029 => x"38",
          7030 => x"fe",
          7031 => x"79",
          7032 => x"76",
          7033 => x"7c",
          7034 => x"be",
          7035 => x"88",
          7036 => x"82",
          7037 => x"06",
          7038 => x"8b",
          7039 => x"76",
          7040 => x"76",
          7041 => x"83",
          7042 => x"51",
          7043 => x"3f",
          7044 => x"08",
          7045 => x"06",
          7046 => x"70",
          7047 => x"55",
          7048 => x"2e",
          7049 => x"80",
          7050 => x"c7",
          7051 => x"57",
          7052 => x"76",
          7053 => x"ff",
          7054 => x"78",
          7055 => x"76",
          7056 => x"59",
          7057 => x"39",
          7058 => x"05",
          7059 => x"55",
          7060 => x"34",
          7061 => x"80",
          7062 => x"80",
          7063 => x"75",
          7064 => x"8c",
          7065 => x"3f",
          7066 => x"08",
          7067 => x"38",
          7068 => x"83",
          7069 => x"a4",
          7070 => x"16",
          7071 => x"26",
          7072 => x"82",
          7073 => x"9f",
          7074 => x"99",
          7075 => x"7b",
          7076 => x"17",
          7077 => x"ff",
          7078 => x"5c",
          7079 => x"05",
          7080 => x"34",
          7081 => x"fd",
          7082 => x"1e",
          7083 => x"81",
          7084 => x"81",
          7085 => x"85",
          7086 => x"34",
          7087 => x"09",
          7088 => x"38",
          7089 => x"81",
          7090 => x"7b",
          7091 => x"73",
          7092 => x"38",
          7093 => x"54",
          7094 => x"09",
          7095 => x"38",
          7096 => x"57",
          7097 => x"70",
          7098 => x"54",
          7099 => x"7b",
          7100 => x"73",
          7101 => x"38",
          7102 => x"57",
          7103 => x"70",
          7104 => x"54",
          7105 => x"85",
          7106 => x"07",
          7107 => x"1f",
          7108 => x"ea",
          7109 => x"d5",
          7110 => x"1f",
          7111 => x"82",
          7112 => x"80",
          7113 => x"82",
          7114 => x"84",
          7115 => x"06",
          7116 => x"74",
          7117 => x"81",
          7118 => x"2a",
          7119 => x"73",
          7120 => x"38",
          7121 => x"54",
          7122 => x"f8",
          7123 => x"80",
          7124 => x"34",
          7125 => x"c2",
          7126 => x"06",
          7127 => x"38",
          7128 => x"39",
          7129 => x"70",
          7130 => x"54",
          7131 => x"86",
          7132 => x"84",
          7133 => x"06",
          7134 => x"73",
          7135 => x"38",
          7136 => x"83",
          7137 => x"05",
          7138 => x"7f",
          7139 => x"3f",
          7140 => x"08",
          7141 => x"f8",
          7142 => x"82",
          7143 => x"92",
          7144 => x"f6",
          7145 => x"5b",
          7146 => x"70",
          7147 => x"59",
          7148 => x"73",
          7149 => x"c6",
          7150 => x"81",
          7151 => x"70",
          7152 => x"52",
          7153 => x"8d",
          7154 => x"38",
          7155 => x"09",
          7156 => x"a5",
          7157 => x"d0",
          7158 => x"ff",
          7159 => x"53",
          7160 => x"91",
          7161 => x"73",
          7162 => x"d0",
          7163 => x"71",
          7164 => x"f7",
          7165 => x"82",
          7166 => x"55",
          7167 => x"55",
          7168 => x"81",
          7169 => x"74",
          7170 => x"56",
          7171 => x"12",
          7172 => x"70",
          7173 => x"38",
          7174 => x"81",
          7175 => x"51",
          7176 => x"51",
          7177 => x"89",
          7178 => x"70",
          7179 => x"53",
          7180 => x"70",
          7181 => x"51",
          7182 => x"09",
          7183 => x"38",
          7184 => x"38",
          7185 => x"77",
          7186 => x"70",
          7187 => x"2a",
          7188 => x"07",
          7189 => x"51",
          7190 => x"8f",
          7191 => x"84",
          7192 => x"83",
          7193 => x"94",
          7194 => x"74",
          7195 => x"38",
          7196 => x"0c",
          7197 => x"86",
          7198 => x"c0",
          7199 => x"82",
          7200 => x"8c",
          7201 => x"fa",
          7202 => x"56",
          7203 => x"17",
          7204 => x"b4",
          7205 => x"52",
          7206 => x"f4",
          7207 => x"82",
          7208 => x"81",
          7209 => x"b6",
          7210 => x"8a",
          7211 => x"e4",
          7212 => x"ff",
          7213 => x"55",
          7214 => x"d5",
          7215 => x"06",
          7216 => x"80",
          7217 => x"33",
          7218 => x"81",
          7219 => x"81",
          7220 => x"81",
          7221 => x"eb",
          7222 => x"70",
          7223 => x"07",
          7224 => x"73",
          7225 => x"81",
          7226 => x"81",
          7227 => x"83",
          7228 => x"94",
          7229 => x"16",
          7230 => x"3f",
          7231 => x"08",
          7232 => x"e4",
          7233 => x"9d",
          7234 => x"82",
          7235 => x"81",
          7236 => x"ce",
          7237 => x"d5",
          7238 => x"82",
          7239 => x"80",
          7240 => x"82",
          7241 => x"d5",
          7242 => x"3d",
          7243 => x"3d",
          7244 => x"84",
          7245 => x"05",
          7246 => x"80",
          7247 => x"51",
          7248 => x"82",
          7249 => x"58",
          7250 => x"0b",
          7251 => x"08",
          7252 => x"38",
          7253 => x"08",
          7254 => x"ed",
          7255 => x"08",
          7256 => x"56",
          7257 => x"87",
          7258 => x"75",
          7259 => x"fe",
          7260 => x"54",
          7261 => x"2e",
          7262 => x"14",
          7263 => x"a0",
          7264 => x"e4",
          7265 => x"06",
          7266 => x"54",
          7267 => x"38",
          7268 => x"87",
          7269 => x"82",
          7270 => x"06",
          7271 => x"56",
          7272 => x"38",
          7273 => x"80",
          7274 => x"18",
          7275 => x"d8",
          7276 => x"15",
          7277 => x"81",
          7278 => x"c6",
          7279 => x"d5",
          7280 => x"ff",
          7281 => x"06",
          7282 => x"56",
          7283 => x"38",
          7284 => x"8f",
          7285 => x"2a",
          7286 => x"51",
          7287 => x"72",
          7288 => x"80",
          7289 => x"52",
          7290 => x"3f",
          7291 => x"08",
          7292 => x"57",
          7293 => x"93",
          7294 => x"26",
          7295 => x"82",
          7296 => x"33",
          7297 => x"2e",
          7298 => x"8c",
          7299 => x"59",
          7300 => x"fa",
          7301 => x"58",
          7302 => x"2e",
          7303 => x"fe",
          7304 => x"a9",
          7305 => x"e4",
          7306 => x"79",
          7307 => x"5b",
          7308 => x"90",
          7309 => x"75",
          7310 => x"38",
          7311 => x"d5",
          7312 => x"70",
          7313 => x"2a",
          7314 => x"95",
          7315 => x"29",
          7316 => x"5a",
          7317 => x"57",
          7318 => x"5b",
          7319 => x"80",
          7320 => x"7a",
          7321 => x"fc",
          7322 => x"d5",
          7323 => x"ff",
          7324 => x"0b",
          7325 => x"1a",
          7326 => x"72",
          7327 => x"81",
          7328 => x"81",
          7329 => x"27",
          7330 => x"80",
          7331 => x"81",
          7332 => x"56",
          7333 => x"27",
          7334 => x"56",
          7335 => x"84",
          7336 => x"56",
          7337 => x"84",
          7338 => x"c3",
          7339 => x"86",
          7340 => x"e4",
          7341 => x"ff",
          7342 => x"84",
          7343 => x"81",
          7344 => x"38",
          7345 => x"51",
          7346 => x"82",
          7347 => x"83",
          7348 => x"58",
          7349 => x"80",
          7350 => x"c9",
          7351 => x"d5",
          7352 => x"77",
          7353 => x"80",
          7354 => x"82",
          7355 => x"c8",
          7356 => x"11",
          7357 => x"06",
          7358 => x"8d",
          7359 => x"26",
          7360 => x"74",
          7361 => x"78",
          7362 => x"c5",
          7363 => x"59",
          7364 => x"15",
          7365 => x"2e",
          7366 => x"13",
          7367 => x"72",
          7368 => x"38",
          7369 => x"f2",
          7370 => x"14",
          7371 => x"3f",
          7372 => x"08",
          7373 => x"e4",
          7374 => x"23",
          7375 => x"57",
          7376 => x"83",
          7377 => x"cb",
          7378 => x"ea",
          7379 => x"e4",
          7380 => x"ff",
          7381 => x"8d",
          7382 => x"14",
          7383 => x"3f",
          7384 => x"08",
          7385 => x"14",
          7386 => x"3f",
          7387 => x"08",
          7388 => x"06",
          7389 => x"72",
          7390 => x"9e",
          7391 => x"22",
          7392 => x"84",
          7393 => x"5a",
          7394 => x"83",
          7395 => x"14",
          7396 => x"79",
          7397 => x"e1",
          7398 => x"d5",
          7399 => x"82",
          7400 => x"80",
          7401 => x"38",
          7402 => x"08",
          7403 => x"ff",
          7404 => x"38",
          7405 => x"83",
          7406 => x"83",
          7407 => x"74",
          7408 => x"85",
          7409 => x"89",
          7410 => x"76",
          7411 => x"ca",
          7412 => x"70",
          7413 => x"7b",
          7414 => x"73",
          7415 => x"17",
          7416 => x"b0",
          7417 => x"55",
          7418 => x"09",
          7419 => x"38",
          7420 => x"51",
          7421 => x"82",
          7422 => x"83",
          7423 => x"53",
          7424 => x"82",
          7425 => x"82",
          7426 => x"e4",
          7427 => x"bd",
          7428 => x"e4",
          7429 => x"0c",
          7430 => x"53",
          7431 => x"56",
          7432 => x"81",
          7433 => x"13",
          7434 => x"74",
          7435 => x"82",
          7436 => x"74",
          7437 => x"81",
          7438 => x"06",
          7439 => x"83",
          7440 => x"2a",
          7441 => x"72",
          7442 => x"26",
          7443 => x"ff",
          7444 => x"0c",
          7445 => x"15",
          7446 => x"0b",
          7447 => x"76",
          7448 => x"81",
          7449 => x"38",
          7450 => x"51",
          7451 => x"82",
          7452 => x"83",
          7453 => x"53",
          7454 => x"09",
          7455 => x"f9",
          7456 => x"52",
          7457 => x"88",
          7458 => x"e4",
          7459 => x"38",
          7460 => x"08",
          7461 => x"84",
          7462 => x"c6",
          7463 => x"d5",
          7464 => x"ff",
          7465 => x"72",
          7466 => x"2e",
          7467 => x"80",
          7468 => x"14",
          7469 => x"3f",
          7470 => x"08",
          7471 => x"a4",
          7472 => x"81",
          7473 => x"84",
          7474 => x"c6",
          7475 => x"d5",
          7476 => x"8a",
          7477 => x"2e",
          7478 => x"9d",
          7479 => x"14",
          7480 => x"3f",
          7481 => x"08",
          7482 => x"84",
          7483 => x"c5",
          7484 => x"d5",
          7485 => x"15",
          7486 => x"34",
          7487 => x"22",
          7488 => x"72",
          7489 => x"23",
          7490 => x"23",
          7491 => x"0b",
          7492 => x"80",
          7493 => x"0c",
          7494 => x"82",
          7495 => x"90",
          7496 => x"fb",
          7497 => x"54",
          7498 => x"80",
          7499 => x"73",
          7500 => x"80",
          7501 => x"72",
          7502 => x"80",
          7503 => x"86",
          7504 => x"15",
          7505 => x"71",
          7506 => x"81",
          7507 => x"81",
          7508 => x"ff",
          7509 => x"82",
          7510 => x"81",
          7511 => x"88",
          7512 => x"08",
          7513 => x"39",
          7514 => x"73",
          7515 => x"74",
          7516 => x"0c",
          7517 => x"04",
          7518 => x"02",
          7519 => x"7a",
          7520 => x"fc",
          7521 => x"f4",
          7522 => x"54",
          7523 => x"d5",
          7524 => x"bc",
          7525 => x"e4",
          7526 => x"82",
          7527 => x"70",
          7528 => x"73",
          7529 => x"38",
          7530 => x"78",
          7531 => x"2e",
          7532 => x"74",
          7533 => x"0c",
          7534 => x"80",
          7535 => x"80",
          7536 => x"70",
          7537 => x"51",
          7538 => x"82",
          7539 => x"54",
          7540 => x"e4",
          7541 => x"0d",
          7542 => x"0d",
          7543 => x"05",
          7544 => x"33",
          7545 => x"54",
          7546 => x"84",
          7547 => x"bf",
          7548 => x"99",
          7549 => x"53",
          7550 => x"05",
          7551 => x"ae",
          7552 => x"e4",
          7553 => x"d5",
          7554 => x"a4",
          7555 => x"69",
          7556 => x"70",
          7557 => x"b0",
          7558 => x"e4",
          7559 => x"d5",
          7560 => x"38",
          7561 => x"05",
          7562 => x"2b",
          7563 => x"80",
          7564 => x"86",
          7565 => x"06",
          7566 => x"2e",
          7567 => x"74",
          7568 => x"38",
          7569 => x"09",
          7570 => x"38",
          7571 => x"b1",
          7572 => x"e4",
          7573 => x"39",
          7574 => x"33",
          7575 => x"73",
          7576 => x"77",
          7577 => x"81",
          7578 => x"73",
          7579 => x"38",
          7580 => x"bc",
          7581 => x"07",
          7582 => x"b4",
          7583 => x"2a",
          7584 => x"51",
          7585 => x"2e",
          7586 => x"62",
          7587 => x"d6",
          7588 => x"d5",
          7589 => x"82",
          7590 => x"52",
          7591 => x"51",
          7592 => x"62",
          7593 => x"8b",
          7594 => x"53",
          7595 => x"51",
          7596 => x"80",
          7597 => x"05",
          7598 => x"3f",
          7599 => x"0b",
          7600 => x"75",
          7601 => x"f1",
          7602 => x"11",
          7603 => x"80",
          7604 => x"98",
          7605 => x"51",
          7606 => x"82",
          7607 => x"55",
          7608 => x"08",
          7609 => x"b7",
          7610 => x"c4",
          7611 => x"05",
          7612 => x"2a",
          7613 => x"51",
          7614 => x"80",
          7615 => x"84",
          7616 => x"39",
          7617 => x"70",
          7618 => x"54",
          7619 => x"a9",
          7620 => x"06",
          7621 => x"2e",
          7622 => x"55",
          7623 => x"73",
          7624 => x"c4",
          7625 => x"d5",
          7626 => x"ff",
          7627 => x"0c",
          7628 => x"d5",
          7629 => x"f8",
          7630 => x"2a",
          7631 => x"51",
          7632 => x"2e",
          7633 => x"80",
          7634 => x"7a",
          7635 => x"a0",
          7636 => x"a4",
          7637 => x"53",
          7638 => x"d5",
          7639 => x"d5",
          7640 => x"d5",
          7641 => x"1b",
          7642 => x"05",
          7643 => x"dd",
          7644 => x"e4",
          7645 => x"e4",
          7646 => x"0c",
          7647 => x"56",
          7648 => x"84",
          7649 => x"90",
          7650 => x"0b",
          7651 => x"80",
          7652 => x"0c",
          7653 => x"1a",
          7654 => x"2a",
          7655 => x"51",
          7656 => x"2e",
          7657 => x"82",
          7658 => x"80",
          7659 => x"38",
          7660 => x"08",
          7661 => x"8a",
          7662 => x"89",
          7663 => x"59",
          7664 => x"76",
          7665 => x"c5",
          7666 => x"d5",
          7667 => x"82",
          7668 => x"81",
          7669 => x"82",
          7670 => x"e4",
          7671 => x"09",
          7672 => x"38",
          7673 => x"78",
          7674 => x"30",
          7675 => x"80",
          7676 => x"77",
          7677 => x"38",
          7678 => x"06",
          7679 => x"c3",
          7680 => x"1a",
          7681 => x"38",
          7682 => x"06",
          7683 => x"2e",
          7684 => x"52",
          7685 => x"ee",
          7686 => x"e4",
          7687 => x"82",
          7688 => x"75",
          7689 => x"d5",
          7690 => x"9c",
          7691 => x"39",
          7692 => x"74",
          7693 => x"d5",
          7694 => x"3d",
          7695 => x"3d",
          7696 => x"65",
          7697 => x"5d",
          7698 => x"0c",
          7699 => x"05",
          7700 => x"f9",
          7701 => x"d5",
          7702 => x"82",
          7703 => x"8a",
          7704 => x"33",
          7705 => x"2e",
          7706 => x"56",
          7707 => x"90",
          7708 => x"06",
          7709 => x"74",
          7710 => x"b9",
          7711 => x"82",
          7712 => x"34",
          7713 => x"ad",
          7714 => x"91",
          7715 => x"56",
          7716 => x"8c",
          7717 => x"1a",
          7718 => x"74",
          7719 => x"38",
          7720 => x"80",
          7721 => x"38",
          7722 => x"70",
          7723 => x"56",
          7724 => x"b4",
          7725 => x"11",
          7726 => x"77",
          7727 => x"5b",
          7728 => x"38",
          7729 => x"88",
          7730 => x"8f",
          7731 => x"08",
          7732 => x"c3",
          7733 => x"d5",
          7734 => x"81",
          7735 => x"9f",
          7736 => x"2e",
          7737 => x"74",
          7738 => x"98",
          7739 => x"7e",
          7740 => x"3f",
          7741 => x"08",
          7742 => x"83",
          7743 => x"e4",
          7744 => x"89",
          7745 => x"77",
          7746 => x"d8",
          7747 => x"7f",
          7748 => x"58",
          7749 => x"75",
          7750 => x"75",
          7751 => x"77",
          7752 => x"7c",
          7753 => x"33",
          7754 => x"91",
          7755 => x"e4",
          7756 => x"38",
          7757 => x"33",
          7758 => x"80",
          7759 => x"b4",
          7760 => x"31",
          7761 => x"27",
          7762 => x"80",
          7763 => x"52",
          7764 => x"77",
          7765 => x"7d",
          7766 => x"bd",
          7767 => x"89",
          7768 => x"39",
          7769 => x"0c",
          7770 => x"83",
          7771 => x"80",
          7772 => x"55",
          7773 => x"83",
          7774 => x"9c",
          7775 => x"7e",
          7776 => x"3f",
          7777 => x"08",
          7778 => x"75",
          7779 => x"08",
          7780 => x"1f",
          7781 => x"7c",
          7782 => x"a9",
          7783 => x"31",
          7784 => x"7f",
          7785 => x"94",
          7786 => x"94",
          7787 => x"5c",
          7788 => x"80",
          7789 => x"d5",
          7790 => x"3d",
          7791 => x"3d",
          7792 => x"65",
          7793 => x"5d",
          7794 => x"0c",
          7795 => x"05",
          7796 => x"f6",
          7797 => x"d5",
          7798 => x"82",
          7799 => x"8a",
          7800 => x"33",
          7801 => x"2e",
          7802 => x"56",
          7803 => x"90",
          7804 => x"81",
          7805 => x"06",
          7806 => x"87",
          7807 => x"2e",
          7808 => x"95",
          7809 => x"91",
          7810 => x"56",
          7811 => x"81",
          7812 => x"34",
          7813 => x"95",
          7814 => x"08",
          7815 => x"56",
          7816 => x"84",
          7817 => x"5c",
          7818 => x"82",
          7819 => x"18",
          7820 => x"ff",
          7821 => x"74",
          7822 => x"7e",
          7823 => x"ff",
          7824 => x"2a",
          7825 => x"7a",
          7826 => x"8c",
          7827 => x"08",
          7828 => x"38",
          7829 => x"39",
          7830 => x"52",
          7831 => x"ac",
          7832 => x"e4",
          7833 => x"d5",
          7834 => x"2e",
          7835 => x"74",
          7836 => x"91",
          7837 => x"2e",
          7838 => x"74",
          7839 => x"88",
          7840 => x"38",
          7841 => x"0c",
          7842 => x"15",
          7843 => x"08",
          7844 => x"06",
          7845 => x"51",
          7846 => x"3f",
          7847 => x"08",
          7848 => x"98",
          7849 => x"7e",
          7850 => x"da",
          7851 => x"e4",
          7852 => x"fe",
          7853 => x"d5",
          7854 => x"7c",
          7855 => x"57",
          7856 => x"80",
          7857 => x"1b",
          7858 => x"22",
          7859 => x"75",
          7860 => x"38",
          7861 => x"59",
          7862 => x"53",
          7863 => x"1a",
          7864 => x"b6",
          7865 => x"d5",
          7866 => x"a3",
          7867 => x"11",
          7868 => x"56",
          7869 => x"27",
          7870 => x"80",
          7871 => x"08",
          7872 => x"2b",
          7873 => x"b8",
          7874 => x"ba",
          7875 => x"55",
          7876 => x"16",
          7877 => x"2b",
          7878 => x"39",
          7879 => x"94",
          7880 => x"94",
          7881 => x"ff",
          7882 => x"82",
          7883 => x"fd",
          7884 => x"77",
          7885 => x"55",
          7886 => x"0c",
          7887 => x"83",
          7888 => x"80",
          7889 => x"55",
          7890 => x"83",
          7891 => x"9c",
          7892 => x"7e",
          7893 => x"b8",
          7894 => x"e4",
          7895 => x"38",
          7896 => x"52",
          7897 => x"83",
          7898 => x"b8",
          7899 => x"b9",
          7900 => x"55",
          7901 => x"16",
          7902 => x"31",
          7903 => x"7f",
          7904 => x"94",
          7905 => x"70",
          7906 => x"8c",
          7907 => x"58",
          7908 => x"76",
          7909 => x"75",
          7910 => x"19",
          7911 => x"39",
          7912 => x"80",
          7913 => x"74",
          7914 => x"80",
          7915 => x"d5",
          7916 => x"3d",
          7917 => x"3d",
          7918 => x"3d",
          7919 => x"70",
          7920 => x"df",
          7921 => x"e4",
          7922 => x"d5",
          7923 => x"80",
          7924 => x"33",
          7925 => x"70",
          7926 => x"55",
          7927 => x"2e",
          7928 => x"a0",
          7929 => x"78",
          7930 => x"a4",
          7931 => x"e4",
          7932 => x"d5",
          7933 => x"d8",
          7934 => x"08",
          7935 => x"a0",
          7936 => x"73",
          7937 => x"88",
          7938 => x"74",
          7939 => x"51",
          7940 => x"8c",
          7941 => x"9c",
          7942 => x"b7",
          7943 => x"88",
          7944 => x"96",
          7945 => x"b7",
          7946 => x"52",
          7947 => x"ff",
          7948 => x"78",
          7949 => x"83",
          7950 => x"51",
          7951 => x"3f",
          7952 => x"08",
          7953 => x"81",
          7954 => x"57",
          7955 => x"34",
          7956 => x"e4",
          7957 => x"0d",
          7958 => x"0d",
          7959 => x"54",
          7960 => x"82",
          7961 => x"53",
          7962 => x"08",
          7963 => x"3d",
          7964 => x"73",
          7965 => x"3f",
          7966 => x"08",
          7967 => x"e4",
          7968 => x"82",
          7969 => x"74",
          7970 => x"d5",
          7971 => x"3d",
          7972 => x"3d",
          7973 => x"51",
          7974 => x"8b",
          7975 => x"82",
          7976 => x"24",
          7977 => x"d5",
          7978 => x"ed",
          7979 => x"52",
          7980 => x"e4",
          7981 => x"0d",
          7982 => x"0d",
          7983 => x"3d",
          7984 => x"95",
          7985 => x"e6",
          7986 => x"e4",
          7987 => x"d5",
          7988 => x"e0",
          7989 => x"64",
          7990 => x"d0",
          7991 => x"e8",
          7992 => x"e4",
          7993 => x"d5",
          7994 => x"38",
          7995 => x"05",
          7996 => x"2b",
          7997 => x"80",
          7998 => x"76",
          7999 => x"0c",
          8000 => x"02",
          8001 => x"70",
          8002 => x"81",
          8003 => x"56",
          8004 => x"9e",
          8005 => x"53",
          8006 => x"c9",
          8007 => x"d5",
          8008 => x"15",
          8009 => x"82",
          8010 => x"84",
          8011 => x"06",
          8012 => x"55",
          8013 => x"e4",
          8014 => x"0d",
          8015 => x"3d",
          8016 => x"3d",
          8017 => x"3d",
          8018 => x"80",
          8019 => x"53",
          8020 => x"fd",
          8021 => x"80",
          8022 => x"e7",
          8023 => x"d5",
          8024 => x"82",
          8025 => x"83",
          8026 => x"80",
          8027 => x"7a",
          8028 => x"08",
          8029 => x"0c",
          8030 => x"d5",
          8031 => x"73",
          8032 => x"83",
          8033 => x"80",
          8034 => x"52",
          8035 => x"3f",
          8036 => x"08",
          8037 => x"e4",
          8038 => x"38",
          8039 => x"08",
          8040 => x"ff",
          8041 => x"82",
          8042 => x"57",
          8043 => x"08",
          8044 => x"80",
          8045 => x"52",
          8046 => x"c2",
          8047 => x"e4",
          8048 => x"3d",
          8049 => x"74",
          8050 => x"3f",
          8051 => x"08",
          8052 => x"e4",
          8053 => x"38",
          8054 => x"51",
          8055 => x"82",
          8056 => x"57",
          8057 => x"08",
          8058 => x"da",
          8059 => x"7b",
          8060 => x"3f",
          8061 => x"e4",
          8062 => x"38",
          8063 => x"51",
          8064 => x"82",
          8065 => x"57",
          8066 => x"08",
          8067 => x"38",
          8068 => x"09",
          8069 => x"38",
          8070 => x"ee",
          8071 => x"ea",
          8072 => x"3d",
          8073 => x"52",
          8074 => x"a0",
          8075 => x"3d",
          8076 => x"11",
          8077 => x"5a",
          8078 => x"2e",
          8079 => x"80",
          8080 => x"81",
          8081 => x"70",
          8082 => x"56",
          8083 => x"81",
          8084 => x"78",
          8085 => x"38",
          8086 => x"9c",
          8087 => x"82",
          8088 => x"18",
          8089 => x"08",
          8090 => x"ff",
          8091 => x"55",
          8092 => x"74",
          8093 => x"38",
          8094 => x"e1",
          8095 => x"55",
          8096 => x"34",
          8097 => x"77",
          8098 => x"81",
          8099 => x"ff",
          8100 => x"3d",
          8101 => x"58",
          8102 => x"80",
          8103 => x"c0",
          8104 => x"29",
          8105 => x"05",
          8106 => x"33",
          8107 => x"56",
          8108 => x"2e",
          8109 => x"16",
          8110 => x"33",
          8111 => x"73",
          8112 => x"16",
          8113 => x"26",
          8114 => x"55",
          8115 => x"91",
          8116 => x"54",
          8117 => x"70",
          8118 => x"34",
          8119 => x"ec",
          8120 => x"70",
          8121 => x"34",
          8122 => x"09",
          8123 => x"38",
          8124 => x"39",
          8125 => x"08",
          8126 => x"59",
          8127 => x"7a",
          8128 => x"5c",
          8129 => x"26",
          8130 => x"7a",
          8131 => x"d5",
          8132 => x"df",
          8133 => x"f7",
          8134 => x"7d",
          8135 => x"05",
          8136 => x"57",
          8137 => x"3f",
          8138 => x"08",
          8139 => x"e4",
          8140 => x"38",
          8141 => x"53",
          8142 => x"38",
          8143 => x"54",
          8144 => x"92",
          8145 => x"33",
          8146 => x"70",
          8147 => x"54",
          8148 => x"38",
          8149 => x"15",
          8150 => x"70",
          8151 => x"58",
          8152 => x"82",
          8153 => x"8a",
          8154 => x"89",
          8155 => x"53",
          8156 => x"b7",
          8157 => x"ff",
          8158 => x"c9",
          8159 => x"d5",
          8160 => x"15",
          8161 => x"53",
          8162 => x"c9",
          8163 => x"d5",
          8164 => x"26",
          8165 => x"30",
          8166 => x"70",
          8167 => x"77",
          8168 => x"18",
          8169 => x"51",
          8170 => x"88",
          8171 => x"73",
          8172 => x"52",
          8173 => x"bb",
          8174 => x"d5",
          8175 => x"82",
          8176 => x"81",
          8177 => x"38",
          8178 => x"08",
          8179 => x"9e",
          8180 => x"e4",
          8181 => x"0c",
          8182 => x"0c",
          8183 => x"81",
          8184 => x"76",
          8185 => x"38",
          8186 => x"94",
          8187 => x"94",
          8188 => x"16",
          8189 => x"2a",
          8190 => x"51",
          8191 => x"72",
          8192 => x"38",
          8193 => x"51",
          8194 => x"3f",
          8195 => x"08",
          8196 => x"e4",
          8197 => x"82",
          8198 => x"56",
          8199 => x"52",
          8200 => x"b5",
          8201 => x"d5",
          8202 => x"73",
          8203 => x"38",
          8204 => x"b0",
          8205 => x"73",
          8206 => x"27",
          8207 => x"98",
          8208 => x"9e",
          8209 => x"08",
          8210 => x"0c",
          8211 => x"06",
          8212 => x"2e",
          8213 => x"52",
          8214 => x"b4",
          8215 => x"d5",
          8216 => x"38",
          8217 => x"16",
          8218 => x"80",
          8219 => x"0b",
          8220 => x"81",
          8221 => x"75",
          8222 => x"d5",
          8223 => x"58",
          8224 => x"54",
          8225 => x"74",
          8226 => x"73",
          8227 => x"90",
          8228 => x"c0",
          8229 => x"90",
          8230 => x"83",
          8231 => x"72",
          8232 => x"38",
          8233 => x"08",
          8234 => x"77",
          8235 => x"80",
          8236 => x"d5",
          8237 => x"3d",
          8238 => x"3d",
          8239 => x"89",
          8240 => x"2e",
          8241 => x"80",
          8242 => x"fc",
          8243 => x"3d",
          8244 => x"e0",
          8245 => x"d5",
          8246 => x"82",
          8247 => x"80",
          8248 => x"76",
          8249 => x"75",
          8250 => x"3f",
          8251 => x"08",
          8252 => x"e4",
          8253 => x"38",
          8254 => x"70",
          8255 => x"57",
          8256 => x"a2",
          8257 => x"33",
          8258 => x"70",
          8259 => x"55",
          8260 => x"2e",
          8261 => x"16",
          8262 => x"51",
          8263 => x"82",
          8264 => x"88",
          8265 => x"54",
          8266 => x"84",
          8267 => x"52",
          8268 => x"bc",
          8269 => x"d5",
          8270 => x"74",
          8271 => x"81",
          8272 => x"85",
          8273 => x"74",
          8274 => x"38",
          8275 => x"74",
          8276 => x"d5",
          8277 => x"3d",
          8278 => x"3d",
          8279 => x"3d",
          8280 => x"70",
          8281 => x"bb",
          8282 => x"e4",
          8283 => x"82",
          8284 => x"73",
          8285 => x"0d",
          8286 => x"0d",
          8287 => x"3d",
          8288 => x"71",
          8289 => x"e7",
          8290 => x"d5",
          8291 => x"82",
          8292 => x"80",
          8293 => x"94",
          8294 => x"e4",
          8295 => x"51",
          8296 => x"3f",
          8297 => x"08",
          8298 => x"39",
          8299 => x"08",
          8300 => x"c1",
          8301 => x"d5",
          8302 => x"82",
          8303 => x"84",
          8304 => x"06",
          8305 => x"53",
          8306 => x"d5",
          8307 => x"38",
          8308 => x"51",
          8309 => x"72",
          8310 => x"ff",
          8311 => x"82",
          8312 => x"84",
          8313 => x"70",
          8314 => x"2c",
          8315 => x"e4",
          8316 => x"51",
          8317 => x"82",
          8318 => x"87",
          8319 => x"ed",
          8320 => x"57",
          8321 => x"3d",
          8322 => x"3d",
          8323 => x"9e",
          8324 => x"e4",
          8325 => x"d5",
          8326 => x"38",
          8327 => x"51",
          8328 => x"82",
          8329 => x"55",
          8330 => x"08",
          8331 => x"80",
          8332 => x"70",
          8333 => x"58",
          8334 => x"85",
          8335 => x"8d",
          8336 => x"2e",
          8337 => x"52",
          8338 => x"80",
          8339 => x"d5",
          8340 => x"3d",
          8341 => x"3d",
          8342 => x"55",
          8343 => x"92",
          8344 => x"52",
          8345 => x"dd",
          8346 => x"d5",
          8347 => x"82",
          8348 => x"82",
          8349 => x"74",
          8350 => x"9c",
          8351 => x"11",
          8352 => x"59",
          8353 => x"75",
          8354 => x"38",
          8355 => x"81",
          8356 => x"5b",
          8357 => x"82",
          8358 => x"39",
          8359 => x"08",
          8360 => x"59",
          8361 => x"09",
          8362 => x"c0",
          8363 => x"5f",
          8364 => x"92",
          8365 => x"51",
          8366 => x"3f",
          8367 => x"08",
          8368 => x"38",
          8369 => x"08",
          8370 => x"38",
          8371 => x"08",
          8372 => x"d5",
          8373 => x"80",
          8374 => x"81",
          8375 => x"59",
          8376 => x"14",
          8377 => x"c9",
          8378 => x"39",
          8379 => x"82",
          8380 => x"57",
          8381 => x"38",
          8382 => x"18",
          8383 => x"ff",
          8384 => x"82",
          8385 => x"5b",
          8386 => x"08",
          8387 => x"7c",
          8388 => x"12",
          8389 => x"52",
          8390 => x"82",
          8391 => x"06",
          8392 => x"14",
          8393 => x"8e",
          8394 => x"e4",
          8395 => x"ff",
          8396 => x"70",
          8397 => x"82",
          8398 => x"51",
          8399 => x"b8",
          8400 => x"a9",
          8401 => x"d5",
          8402 => x"0a",
          8403 => x"70",
          8404 => x"84",
          8405 => x"51",
          8406 => x"ff",
          8407 => x"56",
          8408 => x"38",
          8409 => x"7c",
          8410 => x"0c",
          8411 => x"81",
          8412 => x"74",
          8413 => x"7a",
          8414 => x"0c",
          8415 => x"04",
          8416 => x"79",
          8417 => x"05",
          8418 => x"57",
          8419 => x"82",
          8420 => x"56",
          8421 => x"08",
          8422 => x"91",
          8423 => x"75",
          8424 => x"90",
          8425 => x"81",
          8426 => x"06",
          8427 => x"87",
          8428 => x"2e",
          8429 => x"94",
          8430 => x"73",
          8431 => x"27",
          8432 => x"73",
          8433 => x"d5",
          8434 => x"88",
          8435 => x"76",
          8436 => x"8c",
          8437 => x"e4",
          8438 => x"19",
          8439 => x"ca",
          8440 => x"08",
          8441 => x"ff",
          8442 => x"82",
          8443 => x"ff",
          8444 => x"06",
          8445 => x"56",
          8446 => x"08",
          8447 => x"81",
          8448 => x"82",
          8449 => x"75",
          8450 => x"54",
          8451 => x"08",
          8452 => x"27",
          8453 => x"17",
          8454 => x"d5",
          8455 => x"76",
          8456 => x"bc",
          8457 => x"e4",
          8458 => x"17",
          8459 => x"0c",
          8460 => x"80",
          8461 => x"73",
          8462 => x"75",
          8463 => x"38",
          8464 => x"34",
          8465 => x"82",
          8466 => x"89",
          8467 => x"e0",
          8468 => x"53",
          8469 => x"9c",
          8470 => x"3d",
          8471 => x"3f",
          8472 => x"08",
          8473 => x"e4",
          8474 => x"38",
          8475 => x"3d",
          8476 => x"3d",
          8477 => x"cd",
          8478 => x"d5",
          8479 => x"82",
          8480 => x"81",
          8481 => x"80",
          8482 => x"70",
          8483 => x"81",
          8484 => x"56",
          8485 => x"81",
          8486 => x"98",
          8487 => x"74",
          8488 => x"38",
          8489 => x"05",
          8490 => x"06",
          8491 => x"55",
          8492 => x"38",
          8493 => x"51",
          8494 => x"3f",
          8495 => x"08",
          8496 => x"70",
          8497 => x"55",
          8498 => x"2e",
          8499 => x"78",
          8500 => x"e4",
          8501 => x"08",
          8502 => x"38",
          8503 => x"d5",
          8504 => x"76",
          8505 => x"70",
          8506 => x"b5",
          8507 => x"d5",
          8508 => x"82",
          8509 => x"80",
          8510 => x"d5",
          8511 => x"73",
          8512 => x"90",
          8513 => x"e4",
          8514 => x"d5",
          8515 => x"38",
          8516 => x"d0",
          8517 => x"e4",
          8518 => x"88",
          8519 => x"e4",
          8520 => x"38",
          8521 => x"ab",
          8522 => x"e4",
          8523 => x"e4",
          8524 => x"82",
          8525 => x"07",
          8526 => x"55",
          8527 => x"2e",
          8528 => x"80",
          8529 => x"80",
          8530 => x"77",
          8531 => x"90",
          8532 => x"e4",
          8533 => x"8c",
          8534 => x"ff",
          8535 => x"82",
          8536 => x"55",
          8537 => x"e4",
          8538 => x"0d",
          8539 => x"0d",
          8540 => x"3d",
          8541 => x"52",
          8542 => x"d7",
          8543 => x"d5",
          8544 => x"82",
          8545 => x"82",
          8546 => x"5e",
          8547 => x"3d",
          8548 => x"cb",
          8549 => x"d5",
          8550 => x"82",
          8551 => x"86",
          8552 => x"82",
          8553 => x"d5",
          8554 => x"2e",
          8555 => x"82",
          8556 => x"80",
          8557 => x"70",
          8558 => x"06",
          8559 => x"54",
          8560 => x"38",
          8561 => x"52",
          8562 => x"52",
          8563 => x"bc",
          8564 => x"e4",
          8565 => x"56",
          8566 => x"08",
          8567 => x"54",
          8568 => x"08",
          8569 => x"81",
          8570 => x"82",
          8571 => x"e4",
          8572 => x"09",
          8573 => x"38",
          8574 => x"ba",
          8575 => x"b6",
          8576 => x"e4",
          8577 => x"51",
          8578 => x"3f",
          8579 => x"08",
          8580 => x"e4",
          8581 => x"38",
          8582 => x"52",
          8583 => x"ff",
          8584 => x"78",
          8585 => x"b8",
          8586 => x"54",
          8587 => x"c3",
          8588 => x"88",
          8589 => x"80",
          8590 => x"ff",
          8591 => x"75",
          8592 => x"11",
          8593 => x"b7",
          8594 => x"53",
          8595 => x"53",
          8596 => x"51",
          8597 => x"3f",
          8598 => x"0b",
          8599 => x"34",
          8600 => x"80",
          8601 => x"51",
          8602 => x"3f",
          8603 => x"0b",
          8604 => x"77",
          8605 => x"89",
          8606 => x"e4",
          8607 => x"d5",
          8608 => x"38",
          8609 => x"0a",
          8610 => x"05",
          8611 => x"86",
          8612 => x"64",
          8613 => x"ff",
          8614 => x"64",
          8615 => x"8b",
          8616 => x"54",
          8617 => x"15",
          8618 => x"ff",
          8619 => x"82",
          8620 => x"54",
          8621 => x"53",
          8622 => x"51",
          8623 => x"3f",
          8624 => x"e4",
          8625 => x"0d",
          8626 => x"0d",
          8627 => x"05",
          8628 => x"3f",
          8629 => x"3d",
          8630 => x"52",
          8631 => x"d4",
          8632 => x"d5",
          8633 => x"82",
          8634 => x"82",
          8635 => x"4e",
          8636 => x"52",
          8637 => x"52",
          8638 => x"3f",
          8639 => x"08",
          8640 => x"e4",
          8641 => x"38",
          8642 => x"05",
          8643 => x"06",
          8644 => x"73",
          8645 => x"a0",
          8646 => x"08",
          8647 => x"ff",
          8648 => x"ff",
          8649 => x"b0",
          8650 => x"92",
          8651 => x"54",
          8652 => x"3f",
          8653 => x"52",
          8654 => x"8c",
          8655 => x"e4",
          8656 => x"d5",
          8657 => x"38",
          8658 => x"08",
          8659 => x"06",
          8660 => x"a3",
          8661 => x"92",
          8662 => x"81",
          8663 => x"d5",
          8664 => x"2e",
          8665 => x"81",
          8666 => x"51",
          8667 => x"3f",
          8668 => x"08",
          8669 => x"e4",
          8670 => x"38",
          8671 => x"53",
          8672 => x"8d",
          8673 => x"16",
          8674 => x"b9",
          8675 => x"05",
          8676 => x"34",
          8677 => x"70",
          8678 => x"81",
          8679 => x"55",
          8680 => x"74",
          8681 => x"73",
          8682 => x"78",
          8683 => x"83",
          8684 => x"16",
          8685 => x"2a",
          8686 => x"51",
          8687 => x"80",
          8688 => x"38",
          8689 => x"80",
          8690 => x"52",
          8691 => x"b4",
          8692 => x"d5",
          8693 => x"78",
          8694 => x"aa",
          8695 => x"82",
          8696 => x"80",
          8697 => x"38",
          8698 => x"08",
          8699 => x"ff",
          8700 => x"82",
          8701 => x"79",
          8702 => x"58",
          8703 => x"d5",
          8704 => x"c1",
          8705 => x"33",
          8706 => x"2e",
          8707 => x"9a",
          8708 => x"75",
          8709 => x"ff",
          8710 => x"78",
          8711 => x"83",
          8712 => x"39",
          8713 => x"08",
          8714 => x"51",
          8715 => x"82",
          8716 => x"55",
          8717 => x"08",
          8718 => x"51",
          8719 => x"3f",
          8720 => x"08",
          8721 => x"d5",
          8722 => x"3d",
          8723 => x"3d",
          8724 => x"df",
          8725 => x"84",
          8726 => x"05",
          8727 => x"82",
          8728 => x"cc",
          8729 => x"3d",
          8730 => x"3f",
          8731 => x"08",
          8732 => x"e4",
          8733 => x"38",
          8734 => x"52",
          8735 => x"05",
          8736 => x"3f",
          8737 => x"08",
          8738 => x"e4",
          8739 => x"02",
          8740 => x"33",
          8741 => x"54",
          8742 => x"aa",
          8743 => x"06",
          8744 => x"8b",
          8745 => x"06",
          8746 => x"07",
          8747 => x"56",
          8748 => x"34",
          8749 => x"0b",
          8750 => x"78",
          8751 => x"97",
          8752 => x"e4",
          8753 => x"82",
          8754 => x"96",
          8755 => x"ee",
          8756 => x"56",
          8757 => x"3d",
          8758 => x"95",
          8759 => x"ce",
          8760 => x"e4",
          8761 => x"d5",
          8762 => x"cb",
          8763 => x"64",
          8764 => x"d0",
          8765 => x"d0",
          8766 => x"e4",
          8767 => x"d5",
          8768 => x"38",
          8769 => x"05",
          8770 => x"06",
          8771 => x"73",
          8772 => x"16",
          8773 => x"22",
          8774 => x"07",
          8775 => x"1f",
          8776 => x"f2",
          8777 => x"81",
          8778 => x"34",
          8779 => x"a1",
          8780 => x"d5",
          8781 => x"74",
          8782 => x"0c",
          8783 => x"04",
          8784 => x"6a",
          8785 => x"80",
          8786 => x"cc",
          8787 => x"3d",
          8788 => x"3f",
          8789 => x"08",
          8790 => x"08",
          8791 => x"d5",
          8792 => x"80",
          8793 => x"57",
          8794 => x"81",
          8795 => x"70",
          8796 => x"55",
          8797 => x"80",
          8798 => x"5d",
          8799 => x"52",
          8800 => x"52",
          8801 => x"97",
          8802 => x"e4",
          8803 => x"d5",
          8804 => x"d2",
          8805 => x"73",
          8806 => x"f8",
          8807 => x"e4",
          8808 => x"d5",
          8809 => x"38",
          8810 => x"08",
          8811 => x"08",
          8812 => x"56",
          8813 => x"19",
          8814 => x"59",
          8815 => x"74",
          8816 => x"56",
          8817 => x"ec",
          8818 => x"75",
          8819 => x"74",
          8820 => x"2e",
          8821 => x"16",
          8822 => x"33",
          8823 => x"73",
          8824 => x"38",
          8825 => x"84",
          8826 => x"06",
          8827 => x"7a",
          8828 => x"76",
          8829 => x"07",
          8830 => x"54",
          8831 => x"80",
          8832 => x"80",
          8833 => x"7b",
          8834 => x"53",
          8835 => x"80",
          8836 => x"e4",
          8837 => x"d5",
          8838 => x"38",
          8839 => x"55",
          8840 => x"56",
          8841 => x"8b",
          8842 => x"56",
          8843 => x"83",
          8844 => x"75",
          8845 => x"51",
          8846 => x"3f",
          8847 => x"08",
          8848 => x"82",
          8849 => x"99",
          8850 => x"e6",
          8851 => x"53",
          8852 => x"b4",
          8853 => x"3d",
          8854 => x"3f",
          8855 => x"08",
          8856 => x"08",
          8857 => x"d5",
          8858 => x"dd",
          8859 => x"a0",
          8860 => x"70",
          8861 => x"9b",
          8862 => x"6d",
          8863 => x"55",
          8864 => x"27",
          8865 => x"77",
          8866 => x"51",
          8867 => x"3f",
          8868 => x"08",
          8869 => x"26",
          8870 => x"82",
          8871 => x"51",
          8872 => x"83",
          8873 => x"d5",
          8874 => x"95",
          8875 => x"d5",
          8876 => x"ff",
          8877 => x"74",
          8878 => x"38",
          8879 => x"c8",
          8880 => x"9b",
          8881 => x"d5",
          8882 => x"38",
          8883 => x"27",
          8884 => x"89",
          8885 => x"8b",
          8886 => x"27",
          8887 => x"55",
          8888 => x"81",
          8889 => x"8f",
          8890 => x"2a",
          8891 => x"70",
          8892 => x"34",
          8893 => x"74",
          8894 => x"05",
          8895 => x"16",
          8896 => x"51",
          8897 => x"9f",
          8898 => x"38",
          8899 => x"54",
          8900 => x"81",
          8901 => x"b1",
          8902 => x"2e",
          8903 => x"a3",
          8904 => x"15",
          8905 => x"54",
          8906 => x"09",
          8907 => x"38",
          8908 => x"75",
          8909 => x"40",
          8910 => x"52",
          8911 => x"52",
          8912 => x"db",
          8913 => x"e4",
          8914 => x"d5",
          8915 => x"f7",
          8916 => x"74",
          8917 => x"bc",
          8918 => x"e4",
          8919 => x"d5",
          8920 => x"38",
          8921 => x"38",
          8922 => x"74",
          8923 => x"39",
          8924 => x"08",
          8925 => x"81",
          8926 => x"38",
          8927 => x"74",
          8928 => x"38",
          8929 => x"51",
          8930 => x"3f",
          8931 => x"08",
          8932 => x"e4",
          8933 => x"a0",
          8934 => x"e4",
          8935 => x"51",
          8936 => x"3f",
          8937 => x"0b",
          8938 => x"8b",
          8939 => x"66",
          8940 => x"91",
          8941 => x"81",
          8942 => x"34",
          8943 => x"9c",
          8944 => x"d5",
          8945 => x"73",
          8946 => x"d5",
          8947 => x"3d",
          8948 => x"3d",
          8949 => x"02",
          8950 => x"cb",
          8951 => x"3d",
          8952 => x"72",
          8953 => x"5a",
          8954 => x"82",
          8955 => x"58",
          8956 => x"08",
          8957 => x"91",
          8958 => x"77",
          8959 => x"7c",
          8960 => x"38",
          8961 => x"59",
          8962 => x"90",
          8963 => x"81",
          8964 => x"06",
          8965 => x"73",
          8966 => x"54",
          8967 => x"82",
          8968 => x"39",
          8969 => x"8b",
          8970 => x"11",
          8971 => x"2b",
          8972 => x"54",
          8973 => x"fe",
          8974 => x"ff",
          8975 => x"70",
          8976 => x"07",
          8977 => x"d5",
          8978 => x"90",
          8979 => x"40",
          8980 => x"55",
          8981 => x"88",
          8982 => x"08",
          8983 => x"38",
          8984 => x"77",
          8985 => x"56",
          8986 => x"51",
          8987 => x"3f",
          8988 => x"55",
          8989 => x"08",
          8990 => x"38",
          8991 => x"d5",
          8992 => x"2e",
          8993 => x"82",
          8994 => x"ff",
          8995 => x"38",
          8996 => x"08",
          8997 => x"16",
          8998 => x"2e",
          8999 => x"87",
          9000 => x"74",
          9001 => x"74",
          9002 => x"81",
          9003 => x"38",
          9004 => x"ff",
          9005 => x"2e",
          9006 => x"7b",
          9007 => x"80",
          9008 => x"81",
          9009 => x"81",
          9010 => x"06",
          9011 => x"56",
          9012 => x"52",
          9013 => x"9d",
          9014 => x"d5",
          9015 => x"82",
          9016 => x"80",
          9017 => x"81",
          9018 => x"56",
          9019 => x"d3",
          9020 => x"ff",
          9021 => x"7c",
          9022 => x"55",
          9023 => x"b3",
          9024 => x"1b",
          9025 => x"1b",
          9026 => x"33",
          9027 => x"54",
          9028 => x"34",
          9029 => x"fe",
          9030 => x"08",
          9031 => x"74",
          9032 => x"75",
          9033 => x"16",
          9034 => x"33",
          9035 => x"73",
          9036 => x"77",
          9037 => x"d5",
          9038 => x"3d",
          9039 => x"3d",
          9040 => x"02",
          9041 => x"ef",
          9042 => x"3d",
          9043 => x"59",
          9044 => x"8b",
          9045 => x"82",
          9046 => x"24",
          9047 => x"82",
          9048 => x"84",
          9049 => x"ac",
          9050 => x"51",
          9051 => x"2e",
          9052 => x"75",
          9053 => x"e4",
          9054 => x"e4",
          9055 => x"d5",
          9056 => x"82",
          9057 => x"33",
          9058 => x"81",
          9059 => x"ff",
          9060 => x"82",
          9061 => x"81",
          9062 => x"81",
          9063 => x"83",
          9064 => x"da",
          9065 => x"2a",
          9066 => x"51",
          9067 => x"74",
          9068 => x"9a",
          9069 => x"53",
          9070 => x"51",
          9071 => x"3f",
          9072 => x"08",
          9073 => x"55",
          9074 => x"92",
          9075 => x"80",
          9076 => x"38",
          9077 => x"06",
          9078 => x"2e",
          9079 => x"49",
          9080 => x"87",
          9081 => x"79",
          9082 => x"78",
          9083 => x"26",
          9084 => x"19",
          9085 => x"74",
          9086 => x"38",
          9087 => x"fe",
          9088 => x"2a",
          9089 => x"70",
          9090 => x"59",
          9091 => x"7a",
          9092 => x"56",
          9093 => x"80",
          9094 => x"51",
          9095 => x"74",
          9096 => x"64",
          9097 => x"e0",
          9098 => x"74",
          9099 => x"7f",
          9100 => x"89",
          9101 => x"82",
          9102 => x"8b",
          9103 => x"fe",
          9104 => x"92",
          9105 => x"d5",
          9106 => x"ff",
          9107 => x"8e",
          9108 => x"d4",
          9109 => x"81",
          9110 => x"38",
          9111 => x"1b",
          9112 => x"33",
          9113 => x"80",
          9114 => x"38",
          9115 => x"51",
          9116 => x"3f",
          9117 => x"08",
          9118 => x"52",
          9119 => x"cd",
          9120 => x"e4",
          9121 => x"39",
          9122 => x"05",
          9123 => x"7f",
          9124 => x"f7",
          9125 => x"82",
          9126 => x"8a",
          9127 => x"83",
          9128 => x"06",
          9129 => x"08",
          9130 => x"74",
          9131 => x"5f",
          9132 => x"56",
          9133 => x"8a",
          9134 => x"7f",
          9135 => x"56",
          9136 => x"27",
          9137 => x"93",
          9138 => x"80",
          9139 => x"38",
          9140 => x"70",
          9141 => x"44",
          9142 => x"95",
          9143 => x"06",
          9144 => x"2e",
          9145 => x"62",
          9146 => x"74",
          9147 => x"83",
          9148 => x"06",
          9149 => x"82",
          9150 => x"2e",
          9151 => x"78",
          9152 => x"2e",
          9153 => x"80",
          9154 => x"ae",
          9155 => x"2a",
          9156 => x"82",
          9157 => x"56",
          9158 => x"2e",
          9159 => x"77",
          9160 => x"82",
          9161 => x"79",
          9162 => x"70",
          9163 => x"5a",
          9164 => x"86",
          9165 => x"27",
          9166 => x"52",
          9167 => x"a9",
          9168 => x"d5",
          9169 => x"29",
          9170 => x"70",
          9171 => x"55",
          9172 => x"0b",
          9173 => x"08",
          9174 => x"05",
          9175 => x"ff",
          9176 => x"27",
          9177 => x"89",
          9178 => x"ae",
          9179 => x"2a",
          9180 => x"82",
          9181 => x"56",
          9182 => x"2e",
          9183 => x"77",
          9184 => x"82",
          9185 => x"79",
          9186 => x"70",
          9187 => x"5a",
          9188 => x"86",
          9189 => x"27",
          9190 => x"52",
          9191 => x"a9",
          9192 => x"d5",
          9193 => x"84",
          9194 => x"d5",
          9195 => x"f5",
          9196 => x"81",
          9197 => x"e4",
          9198 => x"d5",
          9199 => x"71",
          9200 => x"83",
          9201 => x"5e",
          9202 => x"89",
          9203 => x"5c",
          9204 => x"1f",
          9205 => x"05",
          9206 => x"ff",
          9207 => x"70",
          9208 => x"31",
          9209 => x"57",
          9210 => x"83",
          9211 => x"06",
          9212 => x"1c",
          9213 => x"5c",
          9214 => x"1d",
          9215 => x"29",
          9216 => x"31",
          9217 => x"55",
          9218 => x"87",
          9219 => x"7c",
          9220 => x"7a",
          9221 => x"31",
          9222 => x"a8",
          9223 => x"d5",
          9224 => x"7d",
          9225 => x"81",
          9226 => x"82",
          9227 => x"83",
          9228 => x"80",
          9229 => x"87",
          9230 => x"81",
          9231 => x"fd",
          9232 => x"ad",
          9233 => x"2e",
          9234 => x"80",
          9235 => x"ff",
          9236 => x"d5",
          9237 => x"a0",
          9238 => x"38",
          9239 => x"74",
          9240 => x"86",
          9241 => x"fd",
          9242 => x"81",
          9243 => x"80",
          9244 => x"83",
          9245 => x"39",
          9246 => x"08",
          9247 => x"92",
          9248 => x"ed",
          9249 => x"59",
          9250 => x"27",
          9251 => x"86",
          9252 => x"55",
          9253 => x"09",
          9254 => x"38",
          9255 => x"f5",
          9256 => x"38",
          9257 => x"55",
          9258 => x"86",
          9259 => x"80",
          9260 => x"7a",
          9261 => x"b0",
          9262 => x"82",
          9263 => x"7a",
          9264 => x"81",
          9265 => x"52",
          9266 => x"ff",
          9267 => x"79",
          9268 => x"7b",
          9269 => x"06",
          9270 => x"51",
          9271 => x"3f",
          9272 => x"1c",
          9273 => x"32",
          9274 => x"96",
          9275 => x"06",
          9276 => x"91",
          9277 => x"8d",
          9278 => x"55",
          9279 => x"ff",
          9280 => x"74",
          9281 => x"06",
          9282 => x"51",
          9283 => x"3f",
          9284 => x"52",
          9285 => x"ff",
          9286 => x"f8",
          9287 => x"34",
          9288 => x"1b",
          9289 => x"d0",
          9290 => x"52",
          9291 => x"ff",
          9292 => x"7e",
          9293 => x"51",
          9294 => x"3f",
          9295 => x"09",
          9296 => x"cb",
          9297 => x"b2",
          9298 => x"c3",
          9299 => x"8d",
          9300 => x"52",
          9301 => x"ff",
          9302 => x"82",
          9303 => x"51",
          9304 => x"3f",
          9305 => x"1b",
          9306 => x"8c",
          9307 => x"b2",
          9308 => x"8d",
          9309 => x"80",
          9310 => x"1c",
          9311 => x"80",
          9312 => x"93",
          9313 => x"ac",
          9314 => x"1b",
          9315 => x"82",
          9316 => x"52",
          9317 => x"ff",
          9318 => x"7c",
          9319 => x"06",
          9320 => x"51",
          9321 => x"3f",
          9322 => x"a4",
          9323 => x"0b",
          9324 => x"93",
          9325 => x"c0",
          9326 => x"51",
          9327 => x"3f",
          9328 => x"52",
          9329 => x"70",
          9330 => x"8c",
          9331 => x"54",
          9332 => x"52",
          9333 => x"88",
          9334 => x"56",
          9335 => x"08",
          9336 => x"7d",
          9337 => x"81",
          9338 => x"38",
          9339 => x"1f",
          9340 => x"7f",
          9341 => x"af",
          9342 => x"53",
          9343 => x"51",
          9344 => x"3f",
          9345 => x"a4",
          9346 => x"51",
          9347 => x"3f",
          9348 => x"e4",
          9349 => x"e4",
          9350 => x"8b",
          9351 => x"18",
          9352 => x"1b",
          9353 => x"ee",
          9354 => x"83",
          9355 => x"ff",
          9356 => x"82",
          9357 => x"78",
          9358 => x"bc",
          9359 => x"87",
          9360 => x"52",
          9361 => x"87",
          9362 => x"54",
          9363 => x"7a",
          9364 => x"ff",
          9365 => x"66",
          9366 => x"7a",
          9367 => x"88",
          9368 => x"80",
          9369 => x"2e",
          9370 => x"9a",
          9371 => x"7a",
          9372 => x"a2",
          9373 => x"84",
          9374 => x"8b",
          9375 => x"0a",
          9376 => x"51",
          9377 => x"ff",
          9378 => x"7d",
          9379 => x"38",
          9380 => x"52",
          9381 => x"8a",
          9382 => x"55",
          9383 => x"62",
          9384 => x"74",
          9385 => x"75",
          9386 => x"7f",
          9387 => x"f7",
          9388 => x"e4",
          9389 => x"38",
          9390 => x"82",
          9391 => x"52",
          9392 => x"8b",
          9393 => x"16",
          9394 => x"56",
          9395 => x"38",
          9396 => x"77",
          9397 => x"8d",
          9398 => x"7d",
          9399 => x"38",
          9400 => x"57",
          9401 => x"83",
          9402 => x"76",
          9403 => x"7a",
          9404 => x"ff",
          9405 => x"82",
          9406 => x"81",
          9407 => x"16",
          9408 => x"56",
          9409 => x"38",
          9410 => x"83",
          9411 => x"86",
          9412 => x"ff",
          9413 => x"38",
          9414 => x"82",
          9415 => x"81",
          9416 => x"2e",
          9417 => x"54",
          9418 => x"52",
          9419 => x"84",
          9420 => x"56",
          9421 => x"08",
          9422 => x"64",
          9423 => x"55",
          9424 => x"16",
          9425 => x"82",
          9426 => x"53",
          9427 => x"51",
          9428 => x"3f",
          9429 => x"62",
          9430 => x"06",
          9431 => x"fd",
          9432 => x"53",
          9433 => x"51",
          9434 => x"3f",
          9435 => x"52",
          9436 => x"89",
          9437 => x"be",
          9438 => x"75",
          9439 => x"81",
          9440 => x"0b",
          9441 => x"77",
          9442 => x"76",
          9443 => x"67",
          9444 => x"fd",
          9445 => x"51",
          9446 => x"3f",
          9447 => x"16",
          9448 => x"e4",
          9449 => x"bf",
          9450 => x"86",
          9451 => x"d5",
          9452 => x"16",
          9453 => x"83",
          9454 => x"ff",
          9455 => x"67",
          9456 => x"1b",
          9457 => x"ce",
          9458 => x"77",
          9459 => x"7f",
          9460 => x"d3",
          9461 => x"82",
          9462 => x"a2",
          9463 => x"80",
          9464 => x"ff",
          9465 => x"81",
          9466 => x"e4",
          9467 => x"89",
          9468 => x"8a",
          9469 => x"86",
          9470 => x"e4",
          9471 => x"82",
          9472 => x"9a",
          9473 => x"f5",
          9474 => x"60",
          9475 => x"79",
          9476 => x"5a",
          9477 => x"78",
          9478 => x"8d",
          9479 => x"55",
          9480 => x"fc",
          9481 => x"51",
          9482 => x"7a",
          9483 => x"81",
          9484 => x"8c",
          9485 => x"74",
          9486 => x"38",
          9487 => x"81",
          9488 => x"81",
          9489 => x"8a",
          9490 => x"06",
          9491 => x"76",
          9492 => x"76",
          9493 => x"55",
          9494 => x"e4",
          9495 => x"0d",
          9496 => x"0d",
          9497 => x"05",
          9498 => x"59",
          9499 => x"2e",
          9500 => x"87",
          9501 => x"76",
          9502 => x"84",
          9503 => x"80",
          9504 => x"38",
          9505 => x"77",
          9506 => x"56",
          9507 => x"34",
          9508 => x"bb",
          9509 => x"38",
          9510 => x"05",
          9511 => x"8c",
          9512 => x"08",
          9513 => x"3f",
          9514 => x"70",
          9515 => x"07",
          9516 => x"30",
          9517 => x"56",
          9518 => x"0c",
          9519 => x"18",
          9520 => x"0d",
          9521 => x"0d",
          9522 => x"08",
          9523 => x"75",
          9524 => x"89",
          9525 => x"54",
          9526 => x"16",
          9527 => x"51",
          9528 => x"82",
          9529 => x"91",
          9530 => x"08",
          9531 => x"81",
          9532 => x"88",
          9533 => x"83",
          9534 => x"74",
          9535 => x"0c",
          9536 => x"04",
          9537 => x"75",
          9538 => x"53",
          9539 => x"51",
          9540 => x"3f",
          9541 => x"85",
          9542 => x"ea",
          9543 => x"80",
          9544 => x"6a",
          9545 => x"70",
          9546 => x"d8",
          9547 => x"72",
          9548 => x"3f",
          9549 => x"8d",
          9550 => x"0d",
          9551 => x"0d",
          9552 => x"05",
          9553 => x"55",
          9554 => x"72",
          9555 => x"8a",
          9556 => x"ff",
          9557 => x"80",
          9558 => x"ff",
          9559 => x"51",
          9560 => x"2e",
          9561 => x"b4",
          9562 => x"2e",
          9563 => x"c9",
          9564 => x"72",
          9565 => x"38",
          9566 => x"83",
          9567 => x"53",
          9568 => x"ff",
          9569 => x"71",
          9570 => x"a8",
          9571 => x"51",
          9572 => x"81",
          9573 => x"81",
          9574 => x"51",
          9575 => x"e4",
          9576 => x"0d",
          9577 => x"0d",
          9578 => x"22",
          9579 => x"96",
          9580 => x"51",
          9581 => x"80",
          9582 => x"38",
          9583 => x"39",
          9584 => x"2e",
          9585 => x"91",
          9586 => x"ff",
          9587 => x"70",
          9588 => x"a8",
          9589 => x"54",
          9590 => x"d5",
          9591 => x"3d",
          9592 => x"3d",
          9593 => x"70",
          9594 => x"26",
          9595 => x"70",
          9596 => x"06",
          9597 => x"57",
          9598 => x"72",
          9599 => x"82",
          9600 => x"75",
          9601 => x"57",
          9602 => x"70",
          9603 => x"75",
          9604 => x"52",
          9605 => x"fb",
          9606 => x"82",
          9607 => x"70",
          9608 => x"81",
          9609 => x"18",
          9610 => x"53",
          9611 => x"80",
          9612 => x"88",
          9613 => x"38",
          9614 => x"82",
          9615 => x"51",
          9616 => x"71",
          9617 => x"76",
          9618 => x"54",
          9619 => x"c3",
          9620 => x"31",
          9621 => x"71",
          9622 => x"a4",
          9623 => x"51",
          9624 => x"12",
          9625 => x"d0",
          9626 => x"39",
          9627 => x"90",
          9628 => x"51",
          9629 => x"b0",
          9630 => x"39",
          9631 => x"51",
          9632 => x"ff",
          9633 => x"39",
          9634 => x"38",
          9635 => x"56",
          9636 => x"71",
          9637 => x"d5",
          9638 => x"3d",
          9639 => x"ff",
          9640 => x"00",
          9641 => x"ff",
          9642 => x"ff",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"69",
          9789 => x"00",
          9790 => x"69",
          9791 => x"6c",
          9792 => x"69",
          9793 => x"00",
          9794 => x"6c",
          9795 => x"00",
          9796 => x"65",
          9797 => x"00",
          9798 => x"63",
          9799 => x"72",
          9800 => x"63",
          9801 => x"00",
          9802 => x"64",
          9803 => x"00",
          9804 => x"64",
          9805 => x"00",
          9806 => x"65",
          9807 => x"65",
          9808 => x"65",
          9809 => x"69",
          9810 => x"69",
          9811 => x"66",
          9812 => x"66",
          9813 => x"61",
          9814 => x"00",
          9815 => x"6d",
          9816 => x"65",
          9817 => x"72",
          9818 => x"65",
          9819 => x"00",
          9820 => x"6e",
          9821 => x"00",
          9822 => x"65",
          9823 => x"00",
          9824 => x"62",
          9825 => x"63",
          9826 => x"62",
          9827 => x"63",
          9828 => x"69",
          9829 => x"00",
          9830 => x"64",
          9831 => x"69",
          9832 => x"45",
          9833 => x"72",
          9834 => x"6e",
          9835 => x"6e",
          9836 => x"65",
          9837 => x"72",
          9838 => x"69",
          9839 => x"6e",
          9840 => x"72",
          9841 => x"79",
          9842 => x"6f",
          9843 => x"6c",
          9844 => x"6f",
          9845 => x"2e",
          9846 => x"6f",
          9847 => x"74",
          9848 => x"6f",
          9849 => x"2e",
          9850 => x"6e",
          9851 => x"69",
          9852 => x"69",
          9853 => x"61",
          9854 => x"00",
          9855 => x"63",
          9856 => x"73",
          9857 => x"6e",
          9858 => x"2e",
          9859 => x"69",
          9860 => x"61",
          9861 => x"61",
          9862 => x"65",
          9863 => x"74",
          9864 => x"00",
          9865 => x"69",
          9866 => x"68",
          9867 => x"6c",
          9868 => x"6e",
          9869 => x"69",
          9870 => x"00",
          9871 => x"44",
          9872 => x"20",
          9873 => x"74",
          9874 => x"72",
          9875 => x"63",
          9876 => x"2e",
          9877 => x"72",
          9878 => x"20",
          9879 => x"62",
          9880 => x"69",
          9881 => x"6e",
          9882 => x"69",
          9883 => x"00",
          9884 => x"69",
          9885 => x"6e",
          9886 => x"65",
          9887 => x"6c",
          9888 => x"00",
          9889 => x"6f",
          9890 => x"6d",
          9891 => x"69",
          9892 => x"20",
          9893 => x"65",
          9894 => x"74",
          9895 => x"66",
          9896 => x"64",
          9897 => x"20",
          9898 => x"6b",
          9899 => x"6f",
          9900 => x"74",
          9901 => x"6f",
          9902 => x"64",
          9903 => x"69",
          9904 => x"75",
          9905 => x"6f",
          9906 => x"61",
          9907 => x"6e",
          9908 => x"6e",
          9909 => x"6c",
          9910 => x"00",
          9911 => x"69",
          9912 => x"69",
          9913 => x"6f",
          9914 => x"64",
          9915 => x"6e",
          9916 => x"66",
          9917 => x"65",
          9918 => x"6d",
          9919 => x"72",
          9920 => x"00",
          9921 => x"6f",
          9922 => x"61",
          9923 => x"6f",
          9924 => x"20",
          9925 => x"65",
          9926 => x"00",
          9927 => x"61",
          9928 => x"65",
          9929 => x"73",
          9930 => x"63",
          9931 => x"65",
          9932 => x"00",
          9933 => x"75",
          9934 => x"73",
          9935 => x"00",
          9936 => x"6e",
          9937 => x"77",
          9938 => x"72",
          9939 => x"2e",
          9940 => x"25",
          9941 => x"62",
          9942 => x"73",
          9943 => x"20",
          9944 => x"25",
          9945 => x"62",
          9946 => x"73",
          9947 => x"63",
          9948 => x"00",
          9949 => x"65",
          9950 => x"00",
          9951 => x"30",
          9952 => x"00",
          9953 => x"20",
          9954 => x"30",
          9955 => x"00",
          9956 => x"20",
          9957 => x"20",
          9958 => x"00",
          9959 => x"30",
          9960 => x"00",
          9961 => x"20",
          9962 => x"7c",
          9963 => x"00",
          9964 => x"4f",
          9965 => x"2a",
          9966 => x"73",
          9967 => x"00",
          9968 => x"31",
          9969 => x"2f",
          9970 => x"30",
          9971 => x"31",
          9972 => x"00",
          9973 => x"5a",
          9974 => x"20",
          9975 => x"20",
          9976 => x"78",
          9977 => x"73",
          9978 => x"20",
          9979 => x"0a",
          9980 => x"50",
          9981 => x"6e",
          9982 => x"72",
          9983 => x"20",
          9984 => x"64",
          9985 => x"00",
          9986 => x"69",
          9987 => x"20",
          9988 => x"65",
          9989 => x"70",
          9990 => x"53",
          9991 => x"6e",
          9992 => x"72",
          9993 => x"00",
          9994 => x"4f",
          9995 => x"20",
          9996 => x"69",
          9997 => x"72",
          9998 => x"74",
          9999 => x"4f",
         10000 => x"20",
         10001 => x"69",
         10002 => x"72",
         10003 => x"74",
         10004 => x"41",
         10005 => x"20",
         10006 => x"69",
         10007 => x"72",
         10008 => x"74",
         10009 => x"41",
         10010 => x"20",
         10011 => x"69",
         10012 => x"72",
         10013 => x"74",
         10014 => x"41",
         10015 => x"20",
         10016 => x"69",
         10017 => x"72",
         10018 => x"74",
         10019 => x"41",
         10020 => x"20",
         10021 => x"69",
         10022 => x"72",
         10023 => x"74",
         10024 => x"65",
         10025 => x"6e",
         10026 => x"70",
         10027 => x"6d",
         10028 => x"2e",
         10029 => x"6e",
         10030 => x"69",
         10031 => x"74",
         10032 => x"72",
         10033 => x"00",
         10034 => x"75",
         10035 => x"78",
         10036 => x"62",
         10037 => x"00",
         10038 => x"4f",
         10039 => x"70",
         10040 => x"73",
         10041 => x"3a",
         10042 => x"61",
         10043 => x"64",
         10044 => x"20",
         10045 => x"74",
         10046 => x"69",
         10047 => x"73",
         10048 => x"61",
         10049 => x"30",
         10050 => x"6c",
         10051 => x"65",
         10052 => x"69",
         10053 => x"61",
         10054 => x"6c",
         10055 => x"00",
         10056 => x"20",
         10057 => x"6c",
         10058 => x"69",
         10059 => x"2e",
         10060 => x"00",
         10061 => x"6f",
         10062 => x"6e",
         10063 => x"2e",
         10064 => x"6f",
         10065 => x"72",
         10066 => x"2e",
         10067 => x"00",
         10068 => x"30",
         10069 => x"28",
         10070 => x"78",
         10071 => x"25",
         10072 => x"78",
         10073 => x"38",
         10074 => x"00",
         10075 => x"75",
         10076 => x"4d",
         10077 => x"72",
         10078 => x"43",
         10079 => x"6c",
         10080 => x"2e",
         10081 => x"30",
         10082 => x"20",
         10083 => x"58",
         10084 => x"3f",
         10085 => x"30",
         10086 => x"20",
         10087 => x"58",
         10088 => x"30",
         10089 => x"20",
         10090 => x"6c",
         10091 => x"00",
         10092 => x"78",
         10093 => x"74",
         10094 => x"20",
         10095 => x"65",
         10096 => x"25",
         10097 => x"78",
         10098 => x"2e",
         10099 => x"61",
         10100 => x"6e",
         10101 => x"6f",
         10102 => x"40",
         10103 => x"38",
         10104 => x"2e",
         10105 => x"00",
         10106 => x"61",
         10107 => x"72",
         10108 => x"72",
         10109 => x"20",
         10110 => x"65",
         10111 => x"64",
         10112 => x"00",
         10113 => x"65",
         10114 => x"72",
         10115 => x"67",
         10116 => x"70",
         10117 => x"61",
         10118 => x"6e",
         10119 => x"00",
         10120 => x"6f",
         10121 => x"72",
         10122 => x"6f",
         10123 => x"67",
         10124 => x"00",
         10125 => x"50",
         10126 => x"69",
         10127 => x"64",
         10128 => x"73",
         10129 => x"2e",
         10130 => x"00",
         10131 => x"64",
         10132 => x"73",
         10133 => x"00",
         10134 => x"64",
         10135 => x"73",
         10136 => x"61",
         10137 => x"6f",
         10138 => x"6e",
         10139 => x"00",
         10140 => x"65",
         10141 => x"79",
         10142 => x"68",
         10143 => x"74",
         10144 => x"20",
         10145 => x"6e",
         10146 => x"70",
         10147 => x"65",
         10148 => x"63",
         10149 => x"61",
         10150 => x"00",
         10151 => x"75",
         10152 => x"6e",
         10153 => x"2e",
         10154 => x"6e",
         10155 => x"69",
         10156 => x"69",
         10157 => x"72",
         10158 => x"74",
         10159 => x"2e",
         10160 => x"64",
         10161 => x"2f",
         10162 => x"25",
         10163 => x"64",
         10164 => x"2e",
         10165 => x"64",
         10166 => x"6f",
         10167 => x"6f",
         10168 => x"67",
         10169 => x"74",
         10170 => x"00",
         10171 => x"28",
         10172 => x"6d",
         10173 => x"43",
         10174 => x"6e",
         10175 => x"29",
         10176 => x"0a",
         10177 => x"69",
         10178 => x"20",
         10179 => x"6c",
         10180 => x"6e",
         10181 => x"3a",
         10182 => x"20",
         10183 => x"42",
         10184 => x"52",
         10185 => x"20",
         10186 => x"38",
         10187 => x"30",
         10188 => x"2e",
         10189 => x"20",
         10190 => x"44",
         10191 => x"20",
         10192 => x"20",
         10193 => x"38",
         10194 => x"30",
         10195 => x"2e",
         10196 => x"20",
         10197 => x"4e",
         10198 => x"42",
         10199 => x"20",
         10200 => x"38",
         10201 => x"30",
         10202 => x"2e",
         10203 => x"20",
         10204 => x"52",
         10205 => x"20",
         10206 => x"20",
         10207 => x"38",
         10208 => x"30",
         10209 => x"2e",
         10210 => x"20",
         10211 => x"41",
         10212 => x"20",
         10213 => x"20",
         10214 => x"38",
         10215 => x"30",
         10216 => x"2e",
         10217 => x"20",
         10218 => x"44",
         10219 => x"52",
         10220 => x"20",
         10221 => x"76",
         10222 => x"73",
         10223 => x"30",
         10224 => x"2e",
         10225 => x"20",
         10226 => x"49",
         10227 => x"31",
         10228 => x"20",
         10229 => x"6d",
         10230 => x"20",
         10231 => x"30",
         10232 => x"2e",
         10233 => x"20",
         10234 => x"4e",
         10235 => x"43",
         10236 => x"20",
         10237 => x"61",
         10238 => x"6c",
         10239 => x"30",
         10240 => x"2e",
         10241 => x"20",
         10242 => x"49",
         10243 => x"4f",
         10244 => x"42",
         10245 => x"00",
         10246 => x"20",
         10247 => x"42",
         10248 => x"43",
         10249 => x"20",
         10250 => x"4f",
         10251 => x"00",
         10252 => x"20",
         10253 => x"53",
         10254 => x"20",
         10255 => x"50",
         10256 => x"64",
         10257 => x"73",
         10258 => x"3a",
         10259 => x"20",
         10260 => x"50",
         10261 => x"65",
         10262 => x"20",
         10263 => x"74",
         10264 => x"41",
         10265 => x"65",
         10266 => x"3d",
         10267 => x"38",
         10268 => x"00",
         10269 => x"20",
         10270 => x"50",
         10271 => x"65",
         10272 => x"79",
         10273 => x"61",
         10274 => x"41",
         10275 => x"65",
         10276 => x"3d",
         10277 => x"38",
         10278 => x"00",
         10279 => x"20",
         10280 => x"74",
         10281 => x"20",
         10282 => x"72",
         10283 => x"64",
         10284 => x"73",
         10285 => x"20",
         10286 => x"3d",
         10287 => x"38",
         10288 => x"00",
         10289 => x"69",
         10290 => x"00",
         10291 => x"20",
         10292 => x"50",
         10293 => x"64",
         10294 => x"20",
         10295 => x"20",
         10296 => x"20",
         10297 => x"20",
         10298 => x"3d",
         10299 => x"34",
         10300 => x"00",
         10301 => x"20",
         10302 => x"79",
         10303 => x"6d",
         10304 => x"6f",
         10305 => x"46",
         10306 => x"20",
         10307 => x"20",
         10308 => x"3d",
         10309 => x"2e",
         10310 => x"64",
         10311 => x"0a",
         10312 => x"20",
         10313 => x"44",
         10314 => x"20",
         10315 => x"63",
         10316 => x"72",
         10317 => x"20",
         10318 => x"20",
         10319 => x"3d",
         10320 => x"2e",
         10321 => x"64",
         10322 => x"0a",
         10323 => x"20",
         10324 => x"69",
         10325 => x"6f",
         10326 => x"53",
         10327 => x"4d",
         10328 => x"6f",
         10329 => x"46",
         10330 => x"3d",
         10331 => x"2e",
         10332 => x"64",
         10333 => x"0a",
         10334 => x"6d",
         10335 => x"00",
         10336 => x"65",
         10337 => x"6d",
         10338 => x"6c",
         10339 => x"00",
         10340 => x"56",
         10341 => x"56",
         10342 => x"00",
         10343 => x"6e",
         10344 => x"77",
         10345 => x"00",
         10346 => x"00",
         10347 => x"00",
         10348 => x"00",
         10349 => x"00",
         10350 => x"00",
         10351 => x"00",
         10352 => x"00",
         10353 => x"00",
         10354 => x"00",
         10355 => x"00",
         10356 => x"00",
         10357 => x"00",
         10358 => x"00",
         10359 => x"00",
         10360 => x"00",
         10361 => x"00",
         10362 => x"00",
         10363 => x"00",
         10364 => x"00",
         10365 => x"00",
         10366 => x"00",
         10367 => x"00",
         10368 => x"00",
         10369 => x"00",
         10370 => x"00",
         10371 => x"00",
         10372 => x"00",
         10373 => x"00",
         10374 => x"00",
         10375 => x"00",
         10376 => x"00",
         10377 => x"00",
         10378 => x"00",
         10379 => x"00",
         10380 => x"00",
         10381 => x"00",
         10382 => x"00",
         10383 => x"00",
         10384 => x"00",
         10385 => x"00",
         10386 => x"00",
         10387 => x"00",
         10388 => x"00",
         10389 => x"00",
         10390 => x"00",
         10391 => x"00",
         10392 => x"00",
         10393 => x"00",
         10394 => x"00",
         10395 => x"00",
         10396 => x"00",
         10397 => x"00",
         10398 => x"00",
         10399 => x"00",
         10400 => x"00",
         10401 => x"00",
         10402 => x"00",
         10403 => x"00",
         10404 => x"00",
         10405 => x"00",
         10406 => x"00",
         10407 => x"00",
         10408 => x"00",
         10409 => x"00",
         10410 => x"00",
         10411 => x"5b",
         10412 => x"5b",
         10413 => x"5b",
         10414 => x"5b",
         10415 => x"5b",
         10416 => x"5b",
         10417 => x"5b",
         10418 => x"30",
         10419 => x"5b",
         10420 => x"5b",
         10421 => x"5b",
         10422 => x"00",
         10423 => x"00",
         10424 => x"00",
         10425 => x"00",
         10426 => x"00",
         10427 => x"00",
         10428 => x"00",
         10429 => x"00",
         10430 => x"00",
         10431 => x"00",
         10432 => x"00",
         10433 => x"69",
         10434 => x"72",
         10435 => x"69",
         10436 => x"00",
         10437 => x"00",
         10438 => x"30",
         10439 => x"20",
         10440 => x"0a",
         10441 => x"61",
         10442 => x"64",
         10443 => x"20",
         10444 => x"65",
         10445 => x"68",
         10446 => x"69",
         10447 => x"72",
         10448 => x"69",
         10449 => x"74",
         10450 => x"4f",
         10451 => x"00",
         10452 => x"61",
         10453 => x"74",
         10454 => x"65",
         10455 => x"72",
         10456 => x"65",
         10457 => x"73",
         10458 => x"79",
         10459 => x"6c",
         10460 => x"64",
         10461 => x"62",
         10462 => x"67",
         10463 => x"44",
         10464 => x"2a",
         10465 => x"3f",
         10466 => x"00",
         10467 => x"2c",
         10468 => x"5d",
         10469 => x"41",
         10470 => x"41",
         10471 => x"00",
         10472 => x"fe",
         10473 => x"44",
         10474 => x"2e",
         10475 => x"4f",
         10476 => x"4d",
         10477 => x"20",
         10478 => x"54",
         10479 => x"20",
         10480 => x"4f",
         10481 => x"4d",
         10482 => x"20",
         10483 => x"54",
         10484 => x"20",
         10485 => x"00",
         10486 => x"00",
         10487 => x"00",
         10488 => x"00",
         10489 => x"03",
         10490 => x"0e",
         10491 => x"16",
         10492 => x"00",
         10493 => x"9a",
         10494 => x"41",
         10495 => x"45",
         10496 => x"49",
         10497 => x"92",
         10498 => x"4f",
         10499 => x"99",
         10500 => x"9d",
         10501 => x"49",
         10502 => x"a5",
         10503 => x"a9",
         10504 => x"ad",
         10505 => x"b1",
         10506 => x"b5",
         10507 => x"b9",
         10508 => x"bd",
         10509 => x"c1",
         10510 => x"c5",
         10511 => x"c9",
         10512 => x"cd",
         10513 => x"d1",
         10514 => x"d5",
         10515 => x"d9",
         10516 => x"dd",
         10517 => x"e1",
         10518 => x"e5",
         10519 => x"e9",
         10520 => x"ed",
         10521 => x"f1",
         10522 => x"f5",
         10523 => x"f9",
         10524 => x"fd",
         10525 => x"2e",
         10526 => x"5b",
         10527 => x"22",
         10528 => x"3e",
         10529 => x"00",
         10530 => x"01",
         10531 => x"10",
         10532 => x"00",
         10533 => x"00",
         10534 => x"01",
         10535 => x"04",
         10536 => x"10",
         10537 => x"00",
         10538 => x"c7",
         10539 => x"e9",
         10540 => x"e4",
         10541 => x"e5",
         10542 => x"ea",
         10543 => x"e8",
         10544 => x"ee",
         10545 => x"c4",
         10546 => x"c9",
         10547 => x"c6",
         10548 => x"f6",
         10549 => x"fb",
         10550 => x"ff",
         10551 => x"dc",
         10552 => x"a3",
         10553 => x"a7",
         10554 => x"e1",
         10555 => x"f3",
         10556 => x"f1",
         10557 => x"aa",
         10558 => x"bf",
         10559 => x"ac",
         10560 => x"bc",
         10561 => x"ab",
         10562 => x"91",
         10563 => x"93",
         10564 => x"24",
         10565 => x"62",
         10566 => x"55",
         10567 => x"51",
         10568 => x"5d",
         10569 => x"5b",
         10570 => x"14",
         10571 => x"2c",
         10572 => x"00",
         10573 => x"5e",
         10574 => x"5a",
         10575 => x"69",
         10576 => x"60",
         10577 => x"6c",
         10578 => x"68",
         10579 => x"65",
         10580 => x"58",
         10581 => x"53",
         10582 => x"6a",
         10583 => x"0c",
         10584 => x"84",
         10585 => x"90",
         10586 => x"b1",
         10587 => x"93",
         10588 => x"a3",
         10589 => x"b5",
         10590 => x"a6",
         10591 => x"a9",
         10592 => x"1e",
         10593 => x"b5",
         10594 => x"61",
         10595 => x"65",
         10596 => x"20",
         10597 => x"f7",
         10598 => x"b0",
         10599 => x"b7",
         10600 => x"7f",
         10601 => x"a0",
         10602 => x"61",
         10603 => x"e0",
         10604 => x"f8",
         10605 => x"ff",
         10606 => x"78",
         10607 => x"30",
         10608 => x"06",
         10609 => x"10",
         10610 => x"2e",
         10611 => x"06",
         10612 => x"4d",
         10613 => x"81",
         10614 => x"82",
         10615 => x"84",
         10616 => x"87",
         10617 => x"89",
         10618 => x"8b",
         10619 => x"8d",
         10620 => x"8f",
         10621 => x"91",
         10622 => x"93",
         10623 => x"f6",
         10624 => x"97",
         10625 => x"98",
         10626 => x"9b",
         10627 => x"9d",
         10628 => x"9f",
         10629 => x"a0",
         10630 => x"a2",
         10631 => x"a4",
         10632 => x"a7",
         10633 => x"a9",
         10634 => x"ab",
         10635 => x"ac",
         10636 => x"af",
         10637 => x"b1",
         10638 => x"b3",
         10639 => x"b5",
         10640 => x"b7",
         10641 => x"b8",
         10642 => x"bb",
         10643 => x"bc",
         10644 => x"f7",
         10645 => x"c1",
         10646 => x"c3",
         10647 => x"c5",
         10648 => x"c7",
         10649 => x"c7",
         10650 => x"cb",
         10651 => x"cd",
         10652 => x"dd",
         10653 => x"8e",
         10654 => x"12",
         10655 => x"03",
         10656 => x"f4",
         10657 => x"f8",
         10658 => x"22",
         10659 => x"3a",
         10660 => x"65",
         10661 => x"3b",
         10662 => x"66",
         10663 => x"40",
         10664 => x"41",
         10665 => x"0a",
         10666 => x"40",
         10667 => x"86",
         10668 => x"89",
         10669 => x"58",
         10670 => x"5a",
         10671 => x"5c",
         10672 => x"5e",
         10673 => x"93",
         10674 => x"62",
         10675 => x"64",
         10676 => x"66",
         10677 => x"97",
         10678 => x"6a",
         10679 => x"6c",
         10680 => x"6e",
         10681 => x"70",
         10682 => x"9d",
         10683 => x"74",
         10684 => x"76",
         10685 => x"78",
         10686 => x"7a",
         10687 => x"7c",
         10688 => x"7e",
         10689 => x"a6",
         10690 => x"82",
         10691 => x"84",
         10692 => x"86",
         10693 => x"ae",
         10694 => x"b1",
         10695 => x"45",
         10696 => x"8e",
         10697 => x"90",
         10698 => x"b7",
         10699 => x"03",
         10700 => x"fe",
         10701 => x"ac",
         10702 => x"86",
         10703 => x"89",
         10704 => x"b1",
         10705 => x"c2",
         10706 => x"a3",
         10707 => x"c4",
         10708 => x"cc",
         10709 => x"8c",
         10710 => x"8f",
         10711 => x"18",
         10712 => x"0a",
         10713 => x"f3",
         10714 => x"f5",
         10715 => x"f7",
         10716 => x"f9",
         10717 => x"fa",
         10718 => x"20",
         10719 => x"10",
         10720 => x"22",
         10721 => x"36",
         10722 => x"0e",
         10723 => x"01",
         10724 => x"d0",
         10725 => x"61",
         10726 => x"00",
         10727 => x"7d",
         10728 => x"63",
         10729 => x"96",
         10730 => x"5a",
         10731 => x"08",
         10732 => x"06",
         10733 => x"08",
         10734 => x"08",
         10735 => x"06",
         10736 => x"07",
         10737 => x"52",
         10738 => x"54",
         10739 => x"56",
         10740 => x"60",
         10741 => x"70",
         10742 => x"ba",
         10743 => x"c8",
         10744 => x"ca",
         10745 => x"da",
         10746 => x"f8",
         10747 => x"ea",
         10748 => x"fa",
         10749 => x"80",
         10750 => x"90",
         10751 => x"a0",
         10752 => x"b0",
         10753 => x"b8",
         10754 => x"b2",
         10755 => x"cc",
         10756 => x"c3",
         10757 => x"02",
         10758 => x"02",
         10759 => x"01",
         10760 => x"f3",
         10761 => x"fc",
         10762 => x"01",
         10763 => x"70",
         10764 => x"84",
         10765 => x"83",
         10766 => x"1a",
         10767 => x"2f",
         10768 => x"02",
         10769 => x"06",
         10770 => x"02",
         10771 => x"64",
         10772 => x"26",
         10773 => x"1a",
         10774 => x"00",
         10775 => x"00",
         10776 => x"02",
         10777 => x"00",
         10778 => x"00",
         10779 => x"00",
         10780 => x"04",
         10781 => x"00",
         10782 => x"00",
         10783 => x"00",
         10784 => x"14",
         10785 => x"00",
         10786 => x"00",
         10787 => x"00",
         10788 => x"2b",
         10789 => x"00",
         10790 => x"00",
         10791 => x"00",
         10792 => x"30",
         10793 => x"00",
         10794 => x"00",
         10795 => x"00",
         10796 => x"3c",
         10797 => x"00",
         10798 => x"00",
         10799 => x"00",
         10800 => x"3d",
         10801 => x"00",
         10802 => x"00",
         10803 => x"00",
         10804 => x"3f",
         10805 => x"00",
         10806 => x"00",
         10807 => x"00",
         10808 => x"40",
         10809 => x"00",
         10810 => x"00",
         10811 => x"00",
         10812 => x"41",
         10813 => x"00",
         10814 => x"00",
         10815 => x"00",
         10816 => x"42",
         10817 => x"00",
         10818 => x"00",
         10819 => x"00",
         10820 => x"43",
         10821 => x"00",
         10822 => x"00",
         10823 => x"00",
         10824 => x"50",
         10825 => x"00",
         10826 => x"00",
         10827 => x"00",
         10828 => x"51",
         10829 => x"00",
         10830 => x"00",
         10831 => x"00",
         10832 => x"54",
         10833 => x"00",
         10834 => x"00",
         10835 => x"00",
         10836 => x"55",
         10837 => x"00",
         10838 => x"00",
         10839 => x"00",
         10840 => x"79",
         10841 => x"00",
         10842 => x"00",
         10843 => x"00",
         10844 => x"78",
         10845 => x"00",
         10846 => x"00",
         10847 => x"00",
         10848 => x"82",
         10849 => x"00",
         10850 => x"00",
         10851 => x"00",
         10852 => x"83",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"85",
         10857 => x"00",
         10858 => x"00",
         10859 => x"00",
         10860 => x"87",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"8c",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"8d",
         10869 => x"00",
         10870 => x"00",
         10871 => x"00",
         10872 => x"8e",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"8f",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"01",
         10885 => x"00",
         10886 => x"01",
         10887 => x"81",
         10888 => x"00",
         10889 => x"7f",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"f5",
         10895 => x"f5",
         10896 => x"f5",
         10897 => x"00",
         10898 => x"01",
         10899 => x"01",
         10900 => x"01",
         10901 => x"00",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"00",
         10927 => x"00",
         10928 => x"00",
         10929 => x"00",
         10930 => x"00",
         10931 => x"00",
         10932 => x"00",
         10933 => x"00",
         10934 => x"01",
         10935 => x"03",
         10936 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"9d",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"9c",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"9f",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"8b",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"95",
           269 => x"0b",
           270 => x"0b",
           271 => x"b3",
           272 => x"0b",
           273 => x"0b",
           274 => x"d1",
           275 => x"0b",
           276 => x"0b",
           277 => x"f0",
           278 => x"0b",
           279 => x"0b",
           280 => x"8f",
           281 => x"0b",
           282 => x"0b",
           283 => x"ad",
           284 => x"0b",
           285 => x"0b",
           286 => x"cd",
           287 => x"0b",
           288 => x"0b",
           289 => x"ed",
           290 => x"0b",
           291 => x"0b",
           292 => x"8d",
           293 => x"0b",
           294 => x"0b",
           295 => x"ad",
           296 => x"0b",
           297 => x"0b",
           298 => x"cd",
           299 => x"0b",
           300 => x"0b",
           301 => x"ed",
           302 => x"0b",
           303 => x"0b",
           304 => x"8d",
           305 => x"0b",
           306 => x"0b",
           307 => x"ad",
           308 => x"0b",
           309 => x"0b",
           310 => x"cd",
           311 => x"0b",
           312 => x"0b",
           313 => x"ed",
           314 => x"0b",
           315 => x"0b",
           316 => x"8d",
           317 => x"0b",
           318 => x"0b",
           319 => x"ad",
           320 => x"0b",
           321 => x"0b",
           322 => x"cd",
           323 => x"0b",
           324 => x"0b",
           325 => x"ed",
           326 => x"0b",
           327 => x"0b",
           328 => x"8d",
           329 => x"0b",
           330 => x"0b",
           331 => x"ad",
           332 => x"0b",
           333 => x"0b",
           334 => x"cd",
           335 => x"0b",
           336 => x"0b",
           337 => x"ed",
           338 => x"0b",
           339 => x"0b",
           340 => x"8d",
           341 => x"0b",
           342 => x"0b",
           343 => x"ad",
           344 => x"0b",
           345 => x"0b",
           346 => x"cd",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"84",
           393 => x"82",
           394 => x"af",
           395 => x"d5",
           396 => x"80",
           397 => x"d5",
           398 => x"ad",
           399 => x"f0",
           400 => x"90",
           401 => x"f0",
           402 => x"2d",
           403 => x"08",
           404 => x"04",
           405 => x"0c",
           406 => x"82",
           407 => x"84",
           408 => x"82",
           409 => x"80",
           410 => x"82",
           411 => x"84",
           412 => x"82",
           413 => x"80",
           414 => x"82",
           415 => x"84",
           416 => x"82",
           417 => x"93",
           418 => x"d5",
           419 => x"80",
           420 => x"d5",
           421 => x"c0",
           422 => x"f0",
           423 => x"90",
           424 => x"f0",
           425 => x"2d",
           426 => x"08",
           427 => x"04",
           428 => x"0c",
           429 => x"2d",
           430 => x"08",
           431 => x"04",
           432 => x"0c",
           433 => x"2d",
           434 => x"08",
           435 => x"04",
           436 => x"0c",
           437 => x"2d",
           438 => x"08",
           439 => x"04",
           440 => x"0c",
           441 => x"2d",
           442 => x"08",
           443 => x"04",
           444 => x"0c",
           445 => x"2d",
           446 => x"08",
           447 => x"04",
           448 => x"0c",
           449 => x"2d",
           450 => x"08",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"04",
           468 => x"0c",
           469 => x"2d",
           470 => x"08",
           471 => x"04",
           472 => x"0c",
           473 => x"2d",
           474 => x"08",
           475 => x"04",
           476 => x"0c",
           477 => x"2d",
           478 => x"08",
           479 => x"04",
           480 => x"0c",
           481 => x"2d",
           482 => x"08",
           483 => x"04",
           484 => x"0c",
           485 => x"2d",
           486 => x"08",
           487 => x"04",
           488 => x"0c",
           489 => x"2d",
           490 => x"08",
           491 => x"04",
           492 => x"0c",
           493 => x"2d",
           494 => x"08",
           495 => x"04",
           496 => x"0c",
           497 => x"2d",
           498 => x"08",
           499 => x"04",
           500 => x"0c",
           501 => x"2d",
           502 => x"08",
           503 => x"04",
           504 => x"0c",
           505 => x"2d",
           506 => x"08",
           507 => x"04",
           508 => x"0c",
           509 => x"2d",
           510 => x"08",
           511 => x"04",
           512 => x"0c",
           513 => x"2d",
           514 => x"08",
           515 => x"04",
           516 => x"0c",
           517 => x"2d",
           518 => x"08",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"04",
           536 => x"0c",
           537 => x"2d",
           538 => x"08",
           539 => x"04",
           540 => x"0c",
           541 => x"2d",
           542 => x"08",
           543 => x"04",
           544 => x"0c",
           545 => x"2d",
           546 => x"08",
           547 => x"04",
           548 => x"0c",
           549 => x"2d",
           550 => x"08",
           551 => x"04",
           552 => x"0c",
           553 => x"2d",
           554 => x"08",
           555 => x"04",
           556 => x"0c",
           557 => x"2d",
           558 => x"08",
           559 => x"04",
           560 => x"0c",
           561 => x"2d",
           562 => x"08",
           563 => x"04",
           564 => x"0c",
           565 => x"2d",
           566 => x"08",
           567 => x"04",
           568 => x"0c",
           569 => x"2d",
           570 => x"08",
           571 => x"04",
           572 => x"0c",
           573 => x"2d",
           574 => x"08",
           575 => x"04",
           576 => x"0c",
           577 => x"2d",
           578 => x"08",
           579 => x"04",
           580 => x"0c",
           581 => x"2d",
           582 => x"08",
           583 => x"04",
           584 => x"0c",
           585 => x"2d",
           586 => x"08",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"04",
           600 => x"00",
           601 => x"10",
           602 => x"10",
           603 => x"10",
           604 => x"10",
           605 => x"10",
           606 => x"10",
           607 => x"10",
           608 => x"53",
           609 => x"00",
           610 => x"06",
           611 => x"09",
           612 => x"05",
           613 => x"2b",
           614 => x"06",
           615 => x"04",
           616 => x"72",
           617 => x"05",
           618 => x"05",
           619 => x"72",
           620 => x"53",
           621 => x"51",
           622 => x"04",
           623 => x"70",
           624 => x"27",
           625 => x"71",
           626 => x"53",
           627 => x"0b",
           628 => x"8c",
           629 => x"f0",
           630 => x"82",
           631 => x"02",
           632 => x"0c",
           633 => x"82",
           634 => x"8c",
           635 => x"d5",
           636 => x"05",
           637 => x"f0",
           638 => x"08",
           639 => x"f0",
           640 => x"08",
           641 => x"c8",
           642 => x"84",
           643 => x"d5",
           644 => x"82",
           645 => x"f8",
           646 => x"d5",
           647 => x"05",
           648 => x"d5",
           649 => x"54",
           650 => x"82",
           651 => x"04",
           652 => x"08",
           653 => x"f0",
           654 => x"0d",
           655 => x"08",
           656 => x"85",
           657 => x"81",
           658 => x"06",
           659 => x"52",
           660 => x"80",
           661 => x"f0",
           662 => x"08",
           663 => x"8d",
           664 => x"82",
           665 => x"f4",
           666 => x"c4",
           667 => x"f0",
           668 => x"08",
           669 => x"d5",
           670 => x"05",
           671 => x"82",
           672 => x"f8",
           673 => x"d5",
           674 => x"05",
           675 => x"f0",
           676 => x"0c",
           677 => x"08",
           678 => x"8a",
           679 => x"38",
           680 => x"d5",
           681 => x"05",
           682 => x"e9",
           683 => x"f0",
           684 => x"08",
           685 => x"3f",
           686 => x"08",
           687 => x"f0",
           688 => x"0c",
           689 => x"f0",
           690 => x"08",
           691 => x"81",
           692 => x"80",
           693 => x"f0",
           694 => x"0c",
           695 => x"82",
           696 => x"fc",
           697 => x"d5",
           698 => x"05",
           699 => x"71",
           700 => x"d5",
           701 => x"05",
           702 => x"82",
           703 => x"8c",
           704 => x"d5",
           705 => x"05",
           706 => x"82",
           707 => x"fc",
           708 => x"80",
           709 => x"f0",
           710 => x"08",
           711 => x"34",
           712 => x"08",
           713 => x"70",
           714 => x"08",
           715 => x"52",
           716 => x"08",
           717 => x"82",
           718 => x"87",
           719 => x"d5",
           720 => x"82",
           721 => x"02",
           722 => x"0c",
           723 => x"86",
           724 => x"f0",
           725 => x"34",
           726 => x"08",
           727 => x"82",
           728 => x"e0",
           729 => x"0a",
           730 => x"f0",
           731 => x"0c",
           732 => x"08",
           733 => x"82",
           734 => x"fc",
           735 => x"d5",
           736 => x"05",
           737 => x"d5",
           738 => x"05",
           739 => x"d5",
           740 => x"05",
           741 => x"54",
           742 => x"82",
           743 => x"70",
           744 => x"08",
           745 => x"82",
           746 => x"ec",
           747 => x"d5",
           748 => x"05",
           749 => x"54",
           750 => x"82",
           751 => x"dc",
           752 => x"82",
           753 => x"54",
           754 => x"82",
           755 => x"04",
           756 => x"08",
           757 => x"f0",
           758 => x"0d",
           759 => x"08",
           760 => x"82",
           761 => x"fc",
           762 => x"d5",
           763 => x"05",
           764 => x"d5",
           765 => x"05",
           766 => x"d5",
           767 => x"05",
           768 => x"a3",
           769 => x"e4",
           770 => x"d5",
           771 => x"05",
           772 => x"f0",
           773 => x"08",
           774 => x"e4",
           775 => x"87",
           776 => x"d5",
           777 => x"82",
           778 => x"02",
           779 => x"0c",
           780 => x"80",
           781 => x"f0",
           782 => x"23",
           783 => x"08",
           784 => x"53",
           785 => x"14",
           786 => x"f0",
           787 => x"08",
           788 => x"70",
           789 => x"81",
           790 => x"06",
           791 => x"51",
           792 => x"2e",
           793 => x"0b",
           794 => x"08",
           795 => x"96",
           796 => x"d5",
           797 => x"05",
           798 => x"33",
           799 => x"d5",
           800 => x"05",
           801 => x"ff",
           802 => x"80",
           803 => x"38",
           804 => x"08",
           805 => x"81",
           806 => x"f0",
           807 => x"0c",
           808 => x"08",
           809 => x"70",
           810 => x"53",
           811 => x"95",
           812 => x"d5",
           813 => x"05",
           814 => x"73",
           815 => x"38",
           816 => x"08",
           817 => x"53",
           818 => x"81",
           819 => x"d5",
           820 => x"05",
           821 => x"b0",
           822 => x"06",
           823 => x"82",
           824 => x"e8",
           825 => x"98",
           826 => x"2c",
           827 => x"72",
           828 => x"d5",
           829 => x"05",
           830 => x"2a",
           831 => x"70",
           832 => x"51",
           833 => x"80",
           834 => x"82",
           835 => x"e4",
           836 => x"82",
           837 => x"53",
           838 => x"f0",
           839 => x"23",
           840 => x"82",
           841 => x"e8",
           842 => x"98",
           843 => x"2c",
           844 => x"2b",
           845 => x"11",
           846 => x"53",
           847 => x"72",
           848 => x"08",
           849 => x"82",
           850 => x"e8",
           851 => x"82",
           852 => x"f8",
           853 => x"15",
           854 => x"51",
           855 => x"d5",
           856 => x"05",
           857 => x"f0",
           858 => x"33",
           859 => x"70",
           860 => x"51",
           861 => x"25",
           862 => x"ff",
           863 => x"f0",
           864 => x"34",
           865 => x"08",
           866 => x"70",
           867 => x"81",
           868 => x"53",
           869 => x"38",
           870 => x"08",
           871 => x"70",
           872 => x"90",
           873 => x"2c",
           874 => x"51",
           875 => x"53",
           876 => x"f0",
           877 => x"23",
           878 => x"82",
           879 => x"e4",
           880 => x"83",
           881 => x"06",
           882 => x"72",
           883 => x"38",
           884 => x"08",
           885 => x"70",
           886 => x"98",
           887 => x"53",
           888 => x"81",
           889 => x"f0",
           890 => x"34",
           891 => x"08",
           892 => x"e0",
           893 => x"f0",
           894 => x"0c",
           895 => x"f0",
           896 => x"08",
           897 => x"92",
           898 => x"d5",
           899 => x"05",
           900 => x"2b",
           901 => x"11",
           902 => x"51",
           903 => x"04",
           904 => x"08",
           905 => x"70",
           906 => x"53",
           907 => x"f0",
           908 => x"23",
           909 => x"08",
           910 => x"70",
           911 => x"53",
           912 => x"f0",
           913 => x"23",
           914 => x"82",
           915 => x"e4",
           916 => x"81",
           917 => x"53",
           918 => x"f0",
           919 => x"23",
           920 => x"82",
           921 => x"e4",
           922 => x"80",
           923 => x"53",
           924 => x"f0",
           925 => x"23",
           926 => x"82",
           927 => x"e4",
           928 => x"88",
           929 => x"72",
           930 => x"08",
           931 => x"80",
           932 => x"f0",
           933 => x"34",
           934 => x"82",
           935 => x"e4",
           936 => x"84",
           937 => x"72",
           938 => x"08",
           939 => x"fb",
           940 => x"0b",
           941 => x"08",
           942 => x"82",
           943 => x"ec",
           944 => x"11",
           945 => x"82",
           946 => x"ec",
           947 => x"e3",
           948 => x"f0",
           949 => x"34",
           950 => x"82",
           951 => x"90",
           952 => x"d5",
           953 => x"05",
           954 => x"82",
           955 => x"90",
           956 => x"08",
           957 => x"82",
           958 => x"fc",
           959 => x"d5",
           960 => x"05",
           961 => x"51",
           962 => x"d5",
           963 => x"05",
           964 => x"39",
           965 => x"08",
           966 => x"82",
           967 => x"90",
           968 => x"05",
           969 => x"08",
           970 => x"70",
           971 => x"f0",
           972 => x"0c",
           973 => x"08",
           974 => x"70",
           975 => x"81",
           976 => x"51",
           977 => x"2e",
           978 => x"d5",
           979 => x"05",
           980 => x"2b",
           981 => x"2c",
           982 => x"f0",
           983 => x"08",
           984 => x"83",
           985 => x"e4",
           986 => x"82",
           987 => x"f4",
           988 => x"39",
           989 => x"08",
           990 => x"51",
           991 => x"82",
           992 => x"53",
           993 => x"f0",
           994 => x"23",
           995 => x"08",
           996 => x"53",
           997 => x"08",
           998 => x"73",
           999 => x"54",
          1000 => x"f0",
          1001 => x"23",
          1002 => x"82",
          1003 => x"90",
          1004 => x"d5",
          1005 => x"05",
          1006 => x"82",
          1007 => x"90",
          1008 => x"08",
          1009 => x"08",
          1010 => x"82",
          1011 => x"e4",
          1012 => x"83",
          1013 => x"06",
          1014 => x"53",
          1015 => x"ab",
          1016 => x"f0",
          1017 => x"33",
          1018 => x"53",
          1019 => x"53",
          1020 => x"08",
          1021 => x"52",
          1022 => x"3f",
          1023 => x"08",
          1024 => x"d5",
          1025 => x"05",
          1026 => x"82",
          1027 => x"fc",
          1028 => x"9b",
          1029 => x"d5",
          1030 => x"72",
          1031 => x"08",
          1032 => x"82",
          1033 => x"ec",
          1034 => x"82",
          1035 => x"f4",
          1036 => x"71",
          1037 => x"72",
          1038 => x"08",
          1039 => x"8a",
          1040 => x"d5",
          1041 => x"05",
          1042 => x"2a",
          1043 => x"51",
          1044 => x"80",
          1045 => x"82",
          1046 => x"90",
          1047 => x"d5",
          1048 => x"05",
          1049 => x"82",
          1050 => x"90",
          1051 => x"08",
          1052 => x"08",
          1053 => x"53",
          1054 => x"d5",
          1055 => x"05",
          1056 => x"f0",
          1057 => x"08",
          1058 => x"d5",
          1059 => x"05",
          1060 => x"82",
          1061 => x"dc",
          1062 => x"82",
          1063 => x"dc",
          1064 => x"d5",
          1065 => x"05",
          1066 => x"f0",
          1067 => x"08",
          1068 => x"38",
          1069 => x"08",
          1070 => x"70",
          1071 => x"53",
          1072 => x"f0",
          1073 => x"23",
          1074 => x"08",
          1075 => x"30",
          1076 => x"08",
          1077 => x"82",
          1078 => x"e4",
          1079 => x"ff",
          1080 => x"53",
          1081 => x"f0",
          1082 => x"23",
          1083 => x"88",
          1084 => x"f0",
          1085 => x"23",
          1086 => x"d5",
          1087 => x"05",
          1088 => x"c0",
          1089 => x"72",
          1090 => x"08",
          1091 => x"80",
          1092 => x"d5",
          1093 => x"05",
          1094 => x"82",
          1095 => x"f4",
          1096 => x"d5",
          1097 => x"05",
          1098 => x"2a",
          1099 => x"51",
          1100 => x"80",
          1101 => x"82",
          1102 => x"90",
          1103 => x"d5",
          1104 => x"05",
          1105 => x"82",
          1106 => x"90",
          1107 => x"08",
          1108 => x"08",
          1109 => x"53",
          1110 => x"d5",
          1111 => x"05",
          1112 => x"f0",
          1113 => x"08",
          1114 => x"d5",
          1115 => x"05",
          1116 => x"82",
          1117 => x"d8",
          1118 => x"82",
          1119 => x"d8",
          1120 => x"d5",
          1121 => x"05",
          1122 => x"f0",
          1123 => x"22",
          1124 => x"51",
          1125 => x"d5",
          1126 => x"05",
          1127 => x"f4",
          1128 => x"f0",
          1129 => x"0c",
          1130 => x"08",
          1131 => x"82",
          1132 => x"f4",
          1133 => x"d5",
          1134 => x"05",
          1135 => x"70",
          1136 => x"55",
          1137 => x"82",
          1138 => x"53",
          1139 => x"82",
          1140 => x"f0",
          1141 => x"d5",
          1142 => x"05",
          1143 => x"f0",
          1144 => x"08",
          1145 => x"53",
          1146 => x"a4",
          1147 => x"f0",
          1148 => x"08",
          1149 => x"54",
          1150 => x"08",
          1151 => x"70",
          1152 => x"51",
          1153 => x"82",
          1154 => x"d0",
          1155 => x"39",
          1156 => x"08",
          1157 => x"53",
          1158 => x"11",
          1159 => x"82",
          1160 => x"d0",
          1161 => x"d5",
          1162 => x"05",
          1163 => x"d5",
          1164 => x"05",
          1165 => x"82",
          1166 => x"f0",
          1167 => x"05",
          1168 => x"08",
          1169 => x"82",
          1170 => x"f4",
          1171 => x"53",
          1172 => x"08",
          1173 => x"52",
          1174 => x"3f",
          1175 => x"08",
          1176 => x"f0",
          1177 => x"0c",
          1178 => x"f0",
          1179 => x"08",
          1180 => x"38",
          1181 => x"82",
          1182 => x"f0",
          1183 => x"d5",
          1184 => x"72",
          1185 => x"75",
          1186 => x"72",
          1187 => x"08",
          1188 => x"82",
          1189 => x"e4",
          1190 => x"b2",
          1191 => x"72",
          1192 => x"38",
          1193 => x"08",
          1194 => x"ff",
          1195 => x"72",
          1196 => x"08",
          1197 => x"82",
          1198 => x"e4",
          1199 => x"86",
          1200 => x"06",
          1201 => x"72",
          1202 => x"e7",
          1203 => x"f0",
          1204 => x"22",
          1205 => x"82",
          1206 => x"cc",
          1207 => x"d5",
          1208 => x"05",
          1209 => x"82",
          1210 => x"cc",
          1211 => x"d5",
          1212 => x"05",
          1213 => x"72",
          1214 => x"81",
          1215 => x"82",
          1216 => x"cc",
          1217 => x"05",
          1218 => x"d5",
          1219 => x"05",
          1220 => x"82",
          1221 => x"cc",
          1222 => x"05",
          1223 => x"d5",
          1224 => x"05",
          1225 => x"f0",
          1226 => x"22",
          1227 => x"08",
          1228 => x"82",
          1229 => x"e4",
          1230 => x"83",
          1231 => x"06",
          1232 => x"72",
          1233 => x"d0",
          1234 => x"f0",
          1235 => x"33",
          1236 => x"70",
          1237 => x"d5",
          1238 => x"05",
          1239 => x"51",
          1240 => x"24",
          1241 => x"d5",
          1242 => x"05",
          1243 => x"06",
          1244 => x"82",
          1245 => x"e4",
          1246 => x"39",
          1247 => x"08",
          1248 => x"53",
          1249 => x"08",
          1250 => x"73",
          1251 => x"54",
          1252 => x"f0",
          1253 => x"34",
          1254 => x"08",
          1255 => x"70",
          1256 => x"81",
          1257 => x"53",
          1258 => x"b1",
          1259 => x"f0",
          1260 => x"33",
          1261 => x"70",
          1262 => x"90",
          1263 => x"2c",
          1264 => x"51",
          1265 => x"82",
          1266 => x"ec",
          1267 => x"75",
          1268 => x"72",
          1269 => x"08",
          1270 => x"af",
          1271 => x"f0",
          1272 => x"33",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"82",
          1278 => x"ec",
          1279 => x"75",
          1280 => x"72",
          1281 => x"08",
          1282 => x"82",
          1283 => x"e4",
          1284 => x"83",
          1285 => x"53",
          1286 => x"82",
          1287 => x"ec",
          1288 => x"11",
          1289 => x"82",
          1290 => x"ec",
          1291 => x"90",
          1292 => x"2c",
          1293 => x"73",
          1294 => x"82",
          1295 => x"88",
          1296 => x"a0",
          1297 => x"3f",
          1298 => x"d5",
          1299 => x"05",
          1300 => x"2a",
          1301 => x"51",
          1302 => x"80",
          1303 => x"82",
          1304 => x"88",
          1305 => x"ad",
          1306 => x"3f",
          1307 => x"82",
          1308 => x"e4",
          1309 => x"84",
          1310 => x"06",
          1311 => x"72",
          1312 => x"38",
          1313 => x"08",
          1314 => x"52",
          1315 => x"a5",
          1316 => x"82",
          1317 => x"e4",
          1318 => x"85",
          1319 => x"06",
          1320 => x"72",
          1321 => x"38",
          1322 => x"08",
          1323 => x"52",
          1324 => x"81",
          1325 => x"f0",
          1326 => x"22",
          1327 => x"70",
          1328 => x"51",
          1329 => x"2e",
          1330 => x"d5",
          1331 => x"05",
          1332 => x"51",
          1333 => x"82",
          1334 => x"f4",
          1335 => x"72",
          1336 => x"81",
          1337 => x"82",
          1338 => x"88",
          1339 => x"82",
          1340 => x"f8",
          1341 => x"89",
          1342 => x"d5",
          1343 => x"05",
          1344 => x"2a",
          1345 => x"51",
          1346 => x"80",
          1347 => x"82",
          1348 => x"ec",
          1349 => x"11",
          1350 => x"82",
          1351 => x"ec",
          1352 => x"90",
          1353 => x"2c",
          1354 => x"73",
          1355 => x"82",
          1356 => x"88",
          1357 => x"b0",
          1358 => x"3f",
          1359 => x"d5",
          1360 => x"05",
          1361 => x"2a",
          1362 => x"51",
          1363 => x"80",
          1364 => x"82",
          1365 => x"e8",
          1366 => x"11",
          1367 => x"82",
          1368 => x"e8",
          1369 => x"98",
          1370 => x"2c",
          1371 => x"73",
          1372 => x"82",
          1373 => x"88",
          1374 => x"b0",
          1375 => x"3f",
          1376 => x"d5",
          1377 => x"05",
          1378 => x"2a",
          1379 => x"51",
          1380 => x"b0",
          1381 => x"f0",
          1382 => x"22",
          1383 => x"54",
          1384 => x"f0",
          1385 => x"23",
          1386 => x"70",
          1387 => x"53",
          1388 => x"90",
          1389 => x"f0",
          1390 => x"08",
          1391 => x"87",
          1392 => x"39",
          1393 => x"08",
          1394 => x"53",
          1395 => x"2e",
          1396 => x"97",
          1397 => x"f0",
          1398 => x"08",
          1399 => x"f0",
          1400 => x"33",
          1401 => x"3f",
          1402 => x"82",
          1403 => x"f8",
          1404 => x"72",
          1405 => x"09",
          1406 => x"cb",
          1407 => x"f0",
          1408 => x"22",
          1409 => x"53",
          1410 => x"f0",
          1411 => x"23",
          1412 => x"ff",
          1413 => x"83",
          1414 => x"81",
          1415 => x"d5",
          1416 => x"05",
          1417 => x"d5",
          1418 => x"05",
          1419 => x"52",
          1420 => x"08",
          1421 => x"81",
          1422 => x"f0",
          1423 => x"0c",
          1424 => x"3f",
          1425 => x"82",
          1426 => x"f8",
          1427 => x"72",
          1428 => x"09",
          1429 => x"cb",
          1430 => x"f0",
          1431 => x"22",
          1432 => x"53",
          1433 => x"f0",
          1434 => x"23",
          1435 => x"ff",
          1436 => x"83",
          1437 => x"80",
          1438 => x"d5",
          1439 => x"05",
          1440 => x"d5",
          1441 => x"05",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"81",
          1446 => x"f0",
          1447 => x"0c",
          1448 => x"82",
          1449 => x"f0",
          1450 => x"d5",
          1451 => x"38",
          1452 => x"08",
          1453 => x"52",
          1454 => x"08",
          1455 => x"ff",
          1456 => x"f0",
          1457 => x"0c",
          1458 => x"08",
          1459 => x"70",
          1460 => x"85",
          1461 => x"39",
          1462 => x"08",
          1463 => x"70",
          1464 => x"81",
          1465 => x"53",
          1466 => x"80",
          1467 => x"d5",
          1468 => x"05",
          1469 => x"54",
          1470 => x"d5",
          1471 => x"05",
          1472 => x"2b",
          1473 => x"51",
          1474 => x"25",
          1475 => x"d5",
          1476 => x"05",
          1477 => x"51",
          1478 => x"d2",
          1479 => x"f0",
          1480 => x"08",
          1481 => x"f0",
          1482 => x"33",
          1483 => x"3f",
          1484 => x"d5",
          1485 => x"05",
          1486 => x"39",
          1487 => x"08",
          1488 => x"53",
          1489 => x"09",
          1490 => x"38",
          1491 => x"d5",
          1492 => x"05",
          1493 => x"82",
          1494 => x"ec",
          1495 => x"0b",
          1496 => x"08",
          1497 => x"8a",
          1498 => x"f0",
          1499 => x"23",
          1500 => x"82",
          1501 => x"88",
          1502 => x"82",
          1503 => x"f8",
          1504 => x"84",
          1505 => x"ea",
          1506 => x"f0",
          1507 => x"08",
          1508 => x"70",
          1509 => x"08",
          1510 => x"51",
          1511 => x"f0",
          1512 => x"08",
          1513 => x"0c",
          1514 => x"82",
          1515 => x"04",
          1516 => x"08",
          1517 => x"f0",
          1518 => x"0d",
          1519 => x"08",
          1520 => x"f0",
          1521 => x"08",
          1522 => x"f0",
          1523 => x"08",
          1524 => x"3f",
          1525 => x"08",
          1526 => x"e4",
          1527 => x"3d",
          1528 => x"f0",
          1529 => x"d5",
          1530 => x"82",
          1531 => x"fb",
          1532 => x"0b",
          1533 => x"08",
          1534 => x"82",
          1535 => x"85",
          1536 => x"81",
          1537 => x"32",
          1538 => x"51",
          1539 => x"53",
          1540 => x"8d",
          1541 => x"82",
          1542 => x"f4",
          1543 => x"92",
          1544 => x"f0",
          1545 => x"08",
          1546 => x"82",
          1547 => x"88",
          1548 => x"05",
          1549 => x"08",
          1550 => x"53",
          1551 => x"f0",
          1552 => x"34",
          1553 => x"06",
          1554 => x"2e",
          1555 => x"f1",
          1556 => x"f1",
          1557 => x"82",
          1558 => x"fc",
          1559 => x"90",
          1560 => x"53",
          1561 => x"d5",
          1562 => x"72",
          1563 => x"b1",
          1564 => x"82",
          1565 => x"f8",
          1566 => x"a5",
          1567 => x"c8",
          1568 => x"c8",
          1569 => x"8a",
          1570 => x"08",
          1571 => x"82",
          1572 => x"53",
          1573 => x"8a",
          1574 => x"82",
          1575 => x"f8",
          1576 => x"d5",
          1577 => x"05",
          1578 => x"d5",
          1579 => x"05",
          1580 => x"d5",
          1581 => x"05",
          1582 => x"e4",
          1583 => x"0d",
          1584 => x"0c",
          1585 => x"f0",
          1586 => x"d5",
          1587 => x"3d",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"d5",
          1591 => x"05",
          1592 => x"33",
          1593 => x"70",
          1594 => x"81",
          1595 => x"51",
          1596 => x"80",
          1597 => x"ff",
          1598 => x"f0",
          1599 => x"0c",
          1600 => x"82",
          1601 => x"88",
          1602 => x"72",
          1603 => x"f0",
          1604 => x"08",
          1605 => x"d5",
          1606 => x"05",
          1607 => x"82",
          1608 => x"fc",
          1609 => x"81",
          1610 => x"72",
          1611 => x"38",
          1612 => x"08",
          1613 => x"82",
          1614 => x"8c",
          1615 => x"82",
          1616 => x"fc",
          1617 => x"90",
          1618 => x"53",
          1619 => x"d5",
          1620 => x"72",
          1621 => x"ab",
          1622 => x"82",
          1623 => x"f8",
          1624 => x"9f",
          1625 => x"f0",
          1626 => x"08",
          1627 => x"f0",
          1628 => x"0c",
          1629 => x"f0",
          1630 => x"08",
          1631 => x"0c",
          1632 => x"82",
          1633 => x"04",
          1634 => x"08",
          1635 => x"f0",
          1636 => x"0d",
          1637 => x"08",
          1638 => x"f0",
          1639 => x"08",
          1640 => x"82",
          1641 => x"70",
          1642 => x"0c",
          1643 => x"0d",
          1644 => x"0c",
          1645 => x"f0",
          1646 => x"d5",
          1647 => x"3d",
          1648 => x"f0",
          1649 => x"08",
          1650 => x"70",
          1651 => x"81",
          1652 => x"06",
          1653 => x"51",
          1654 => x"2e",
          1655 => x"0b",
          1656 => x"08",
          1657 => x"81",
          1658 => x"d5",
          1659 => x"05",
          1660 => x"33",
          1661 => x"70",
          1662 => x"51",
          1663 => x"80",
          1664 => x"38",
          1665 => x"08",
          1666 => x"82",
          1667 => x"8c",
          1668 => x"54",
          1669 => x"88",
          1670 => x"9f",
          1671 => x"f0",
          1672 => x"08",
          1673 => x"82",
          1674 => x"88",
          1675 => x"57",
          1676 => x"75",
          1677 => x"81",
          1678 => x"82",
          1679 => x"8c",
          1680 => x"11",
          1681 => x"8c",
          1682 => x"d5",
          1683 => x"05",
          1684 => x"d5",
          1685 => x"05",
          1686 => x"80",
          1687 => x"d5",
          1688 => x"05",
          1689 => x"f0",
          1690 => x"08",
          1691 => x"f0",
          1692 => x"08",
          1693 => x"06",
          1694 => x"08",
          1695 => x"72",
          1696 => x"e4",
          1697 => x"a3",
          1698 => x"f0",
          1699 => x"08",
          1700 => x"81",
          1701 => x"0c",
          1702 => x"08",
          1703 => x"70",
          1704 => x"08",
          1705 => x"51",
          1706 => x"ff",
          1707 => x"f0",
          1708 => x"0c",
          1709 => x"08",
          1710 => x"82",
          1711 => x"87",
          1712 => x"d5",
          1713 => x"82",
          1714 => x"02",
          1715 => x"0c",
          1716 => x"82",
          1717 => x"88",
          1718 => x"11",
          1719 => x"32",
          1720 => x"51",
          1721 => x"71",
          1722 => x"38",
          1723 => x"d5",
          1724 => x"05",
          1725 => x"39",
          1726 => x"08",
          1727 => x"85",
          1728 => x"86",
          1729 => x"06",
          1730 => x"52",
          1731 => x"80",
          1732 => x"d5",
          1733 => x"05",
          1734 => x"f0",
          1735 => x"08",
          1736 => x"12",
          1737 => x"bf",
          1738 => x"71",
          1739 => x"82",
          1740 => x"88",
          1741 => x"11",
          1742 => x"8c",
          1743 => x"d5",
          1744 => x"05",
          1745 => x"33",
          1746 => x"f0",
          1747 => x"0c",
          1748 => x"82",
          1749 => x"d5",
          1750 => x"05",
          1751 => x"33",
          1752 => x"70",
          1753 => x"51",
          1754 => x"80",
          1755 => x"38",
          1756 => x"08",
          1757 => x"70",
          1758 => x"82",
          1759 => x"fc",
          1760 => x"52",
          1761 => x"08",
          1762 => x"a9",
          1763 => x"f0",
          1764 => x"08",
          1765 => x"08",
          1766 => x"53",
          1767 => x"33",
          1768 => x"51",
          1769 => x"14",
          1770 => x"82",
          1771 => x"f8",
          1772 => x"d7",
          1773 => x"f0",
          1774 => x"08",
          1775 => x"05",
          1776 => x"81",
          1777 => x"d5",
          1778 => x"05",
          1779 => x"f0",
          1780 => x"08",
          1781 => x"08",
          1782 => x"2d",
          1783 => x"08",
          1784 => x"f0",
          1785 => x"0c",
          1786 => x"f0",
          1787 => x"08",
          1788 => x"f2",
          1789 => x"f0",
          1790 => x"08",
          1791 => x"08",
          1792 => x"82",
          1793 => x"88",
          1794 => x"11",
          1795 => x"f0",
          1796 => x"0c",
          1797 => x"f0",
          1798 => x"08",
          1799 => x"81",
          1800 => x"82",
          1801 => x"f0",
          1802 => x"07",
          1803 => x"d5",
          1804 => x"05",
          1805 => x"82",
          1806 => x"f0",
          1807 => x"07",
          1808 => x"d5",
          1809 => x"05",
          1810 => x"f0",
          1811 => x"08",
          1812 => x"f0",
          1813 => x"33",
          1814 => x"ff",
          1815 => x"f0",
          1816 => x"0c",
          1817 => x"d5",
          1818 => x"05",
          1819 => x"08",
          1820 => x"12",
          1821 => x"f0",
          1822 => x"08",
          1823 => x"06",
          1824 => x"f0",
          1825 => x"0c",
          1826 => x"82",
          1827 => x"f8",
          1828 => x"d5",
          1829 => x"3d",
          1830 => x"f0",
          1831 => x"d5",
          1832 => x"82",
          1833 => x"fd",
          1834 => x"d5",
          1835 => x"05",
          1836 => x"f0",
          1837 => x"0c",
          1838 => x"08",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"d5",
          1842 => x"05",
          1843 => x"82",
          1844 => x"d5",
          1845 => x"05",
          1846 => x"f0",
          1847 => x"08",
          1848 => x"38",
          1849 => x"08",
          1850 => x"82",
          1851 => x"90",
          1852 => x"51",
          1853 => x"08",
          1854 => x"71",
          1855 => x"38",
          1856 => x"08",
          1857 => x"82",
          1858 => x"90",
          1859 => x"82",
          1860 => x"fc",
          1861 => x"d5",
          1862 => x"05",
          1863 => x"f0",
          1864 => x"08",
          1865 => x"f0",
          1866 => x"0c",
          1867 => x"08",
          1868 => x"81",
          1869 => x"f0",
          1870 => x"0c",
          1871 => x"08",
          1872 => x"ff",
          1873 => x"f0",
          1874 => x"0c",
          1875 => x"08",
          1876 => x"80",
          1877 => x"38",
          1878 => x"08",
          1879 => x"ff",
          1880 => x"f0",
          1881 => x"0c",
          1882 => x"08",
          1883 => x"ff",
          1884 => x"f0",
          1885 => x"0c",
          1886 => x"08",
          1887 => x"82",
          1888 => x"f8",
          1889 => x"51",
          1890 => x"34",
          1891 => x"82",
          1892 => x"90",
          1893 => x"05",
          1894 => x"08",
          1895 => x"82",
          1896 => x"90",
          1897 => x"05",
          1898 => x"08",
          1899 => x"82",
          1900 => x"90",
          1901 => x"2e",
          1902 => x"d5",
          1903 => x"05",
          1904 => x"33",
          1905 => x"08",
          1906 => x"81",
          1907 => x"f0",
          1908 => x"0c",
          1909 => x"08",
          1910 => x"52",
          1911 => x"34",
          1912 => x"08",
          1913 => x"81",
          1914 => x"f0",
          1915 => x"0c",
          1916 => x"82",
          1917 => x"88",
          1918 => x"82",
          1919 => x"51",
          1920 => x"82",
          1921 => x"04",
          1922 => x"08",
          1923 => x"f0",
          1924 => x"0d",
          1925 => x"08",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"d5",
          1929 => x"05",
          1930 => x"33",
          1931 => x"08",
          1932 => x"81",
          1933 => x"f0",
          1934 => x"0c",
          1935 => x"06",
          1936 => x"80",
          1937 => x"da",
          1938 => x"f0",
          1939 => x"08",
          1940 => x"d5",
          1941 => x"05",
          1942 => x"f0",
          1943 => x"08",
          1944 => x"08",
          1945 => x"31",
          1946 => x"e4",
          1947 => x"3d",
          1948 => x"f0",
          1949 => x"d5",
          1950 => x"82",
          1951 => x"fe",
          1952 => x"d5",
          1953 => x"05",
          1954 => x"f0",
          1955 => x"0c",
          1956 => x"08",
          1957 => x"52",
          1958 => x"d5",
          1959 => x"05",
          1960 => x"82",
          1961 => x"8c",
          1962 => x"d5",
          1963 => x"05",
          1964 => x"70",
          1965 => x"d5",
          1966 => x"05",
          1967 => x"82",
          1968 => x"fc",
          1969 => x"81",
          1970 => x"70",
          1971 => x"38",
          1972 => x"82",
          1973 => x"88",
          1974 => x"82",
          1975 => x"51",
          1976 => x"82",
          1977 => x"04",
          1978 => x"08",
          1979 => x"f0",
          1980 => x"0d",
          1981 => x"08",
          1982 => x"82",
          1983 => x"fc",
          1984 => x"d5",
          1985 => x"05",
          1986 => x"f0",
          1987 => x"0c",
          1988 => x"08",
          1989 => x"80",
          1990 => x"38",
          1991 => x"08",
          1992 => x"81",
          1993 => x"f0",
          1994 => x"0c",
          1995 => x"08",
          1996 => x"ff",
          1997 => x"f0",
          1998 => x"0c",
          1999 => x"08",
          2000 => x"80",
          2001 => x"82",
          2002 => x"f8",
          2003 => x"70",
          2004 => x"f0",
          2005 => x"08",
          2006 => x"d5",
          2007 => x"05",
          2008 => x"f0",
          2009 => x"08",
          2010 => x"71",
          2011 => x"f0",
          2012 => x"08",
          2013 => x"d5",
          2014 => x"05",
          2015 => x"39",
          2016 => x"08",
          2017 => x"70",
          2018 => x"0c",
          2019 => x"0d",
          2020 => x"0c",
          2021 => x"f0",
          2022 => x"d5",
          2023 => x"3d",
          2024 => x"f0",
          2025 => x"08",
          2026 => x"f4",
          2027 => x"f0",
          2028 => x"08",
          2029 => x"82",
          2030 => x"8c",
          2031 => x"05",
          2032 => x"08",
          2033 => x"82",
          2034 => x"88",
          2035 => x"33",
          2036 => x"06",
          2037 => x"51",
          2038 => x"84",
          2039 => x"39",
          2040 => x"08",
          2041 => x"52",
          2042 => x"d5",
          2043 => x"05",
          2044 => x"82",
          2045 => x"88",
          2046 => x"81",
          2047 => x"51",
          2048 => x"80",
          2049 => x"f0",
          2050 => x"0c",
          2051 => x"82",
          2052 => x"90",
          2053 => x"05",
          2054 => x"08",
          2055 => x"82",
          2056 => x"90",
          2057 => x"2e",
          2058 => x"81",
          2059 => x"f0",
          2060 => x"08",
          2061 => x"e8",
          2062 => x"f0",
          2063 => x"08",
          2064 => x"53",
          2065 => x"ff",
          2066 => x"f0",
          2067 => x"0c",
          2068 => x"82",
          2069 => x"8c",
          2070 => x"05",
          2071 => x"08",
          2072 => x"82",
          2073 => x"8c",
          2074 => x"33",
          2075 => x"8c",
          2076 => x"82",
          2077 => x"fc",
          2078 => x"39",
          2079 => x"08",
          2080 => x"70",
          2081 => x"f0",
          2082 => x"08",
          2083 => x"71",
          2084 => x"d5",
          2085 => x"05",
          2086 => x"52",
          2087 => x"39",
          2088 => x"d5",
          2089 => x"05",
          2090 => x"f0",
          2091 => x"08",
          2092 => x"0c",
          2093 => x"82",
          2094 => x"04",
          2095 => x"08",
          2096 => x"f0",
          2097 => x"0d",
          2098 => x"08",
          2099 => x"52",
          2100 => x"08",
          2101 => x"51",
          2102 => x"82",
          2103 => x"70",
          2104 => x"08",
          2105 => x"82",
          2106 => x"f8",
          2107 => x"05",
          2108 => x"54",
          2109 => x"3f",
          2110 => x"08",
          2111 => x"f0",
          2112 => x"0c",
          2113 => x"f0",
          2114 => x"08",
          2115 => x"0b",
          2116 => x"08",
          2117 => x"bc",
          2118 => x"f0",
          2119 => x"08",
          2120 => x"08",
          2121 => x"05",
          2122 => x"34",
          2123 => x"08",
          2124 => x"53",
          2125 => x"08",
          2126 => x"52",
          2127 => x"08",
          2128 => x"51",
          2129 => x"82",
          2130 => x"70",
          2131 => x"08",
          2132 => x"54",
          2133 => x"08",
          2134 => x"82",
          2135 => x"88",
          2136 => x"d5",
          2137 => x"82",
          2138 => x"02",
          2139 => x"0c",
          2140 => x"82",
          2141 => x"88",
          2142 => x"d5",
          2143 => x"05",
          2144 => x"f0",
          2145 => x"08",
          2146 => x"0b",
          2147 => x"08",
          2148 => x"80",
          2149 => x"d5",
          2150 => x"05",
          2151 => x"33",
          2152 => x"08",
          2153 => x"81",
          2154 => x"f0",
          2155 => x"0c",
          2156 => x"06",
          2157 => x"80",
          2158 => x"82",
          2159 => x"8c",
          2160 => x"05",
          2161 => x"08",
          2162 => x"82",
          2163 => x"8c",
          2164 => x"2e",
          2165 => x"be",
          2166 => x"f0",
          2167 => x"08",
          2168 => x"d5",
          2169 => x"05",
          2170 => x"f0",
          2171 => x"08",
          2172 => x"08",
          2173 => x"31",
          2174 => x"f0",
          2175 => x"0c",
          2176 => x"f0",
          2177 => x"08",
          2178 => x"0c",
          2179 => x"82",
          2180 => x"04",
          2181 => x"08",
          2182 => x"f0",
          2183 => x"0d",
          2184 => x"08",
          2185 => x"82",
          2186 => x"fc",
          2187 => x"d5",
          2188 => x"05",
          2189 => x"80",
          2190 => x"d5",
          2191 => x"05",
          2192 => x"82",
          2193 => x"90",
          2194 => x"d5",
          2195 => x"05",
          2196 => x"82",
          2197 => x"90",
          2198 => x"d5",
          2199 => x"05",
          2200 => x"a9",
          2201 => x"f0",
          2202 => x"08",
          2203 => x"d5",
          2204 => x"05",
          2205 => x"71",
          2206 => x"d5",
          2207 => x"05",
          2208 => x"82",
          2209 => x"fc",
          2210 => x"be",
          2211 => x"f0",
          2212 => x"08",
          2213 => x"e4",
          2214 => x"3d",
          2215 => x"f0",
          2216 => x"d5",
          2217 => x"82",
          2218 => x"f9",
          2219 => x"0b",
          2220 => x"08",
          2221 => x"82",
          2222 => x"88",
          2223 => x"25",
          2224 => x"d5",
          2225 => x"05",
          2226 => x"d5",
          2227 => x"05",
          2228 => x"82",
          2229 => x"f4",
          2230 => x"d5",
          2231 => x"05",
          2232 => x"81",
          2233 => x"f0",
          2234 => x"0c",
          2235 => x"08",
          2236 => x"82",
          2237 => x"fc",
          2238 => x"d5",
          2239 => x"05",
          2240 => x"b9",
          2241 => x"f0",
          2242 => x"08",
          2243 => x"f0",
          2244 => x"0c",
          2245 => x"d5",
          2246 => x"05",
          2247 => x"f0",
          2248 => x"08",
          2249 => x"0b",
          2250 => x"08",
          2251 => x"82",
          2252 => x"f0",
          2253 => x"d5",
          2254 => x"05",
          2255 => x"82",
          2256 => x"8c",
          2257 => x"82",
          2258 => x"88",
          2259 => x"82",
          2260 => x"d5",
          2261 => x"82",
          2262 => x"f8",
          2263 => x"82",
          2264 => x"fc",
          2265 => x"2e",
          2266 => x"d5",
          2267 => x"05",
          2268 => x"d5",
          2269 => x"05",
          2270 => x"f0",
          2271 => x"08",
          2272 => x"e4",
          2273 => x"3d",
          2274 => x"f0",
          2275 => x"d5",
          2276 => x"82",
          2277 => x"fb",
          2278 => x"0b",
          2279 => x"08",
          2280 => x"82",
          2281 => x"88",
          2282 => x"25",
          2283 => x"d5",
          2284 => x"05",
          2285 => x"d5",
          2286 => x"05",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"d5",
          2290 => x"05",
          2291 => x"90",
          2292 => x"f0",
          2293 => x"08",
          2294 => x"f0",
          2295 => x"0c",
          2296 => x"d5",
          2297 => x"05",
          2298 => x"d5",
          2299 => x"05",
          2300 => x"a2",
          2301 => x"e4",
          2302 => x"d5",
          2303 => x"05",
          2304 => x"d5",
          2305 => x"05",
          2306 => x"90",
          2307 => x"f0",
          2308 => x"08",
          2309 => x"f0",
          2310 => x"0c",
          2311 => x"08",
          2312 => x"70",
          2313 => x"0c",
          2314 => x"0d",
          2315 => x"0c",
          2316 => x"f0",
          2317 => x"d5",
          2318 => x"3d",
          2319 => x"82",
          2320 => x"8c",
          2321 => x"82",
          2322 => x"88",
          2323 => x"80",
          2324 => x"d5",
          2325 => x"82",
          2326 => x"54",
          2327 => x"82",
          2328 => x"04",
          2329 => x"08",
          2330 => x"f0",
          2331 => x"0d",
          2332 => x"d5",
          2333 => x"05",
          2334 => x"d5",
          2335 => x"05",
          2336 => x"3f",
          2337 => x"08",
          2338 => x"e4",
          2339 => x"3d",
          2340 => x"f0",
          2341 => x"d5",
          2342 => x"82",
          2343 => x"fd",
          2344 => x"0b",
          2345 => x"08",
          2346 => x"80",
          2347 => x"f0",
          2348 => x"0c",
          2349 => x"08",
          2350 => x"82",
          2351 => x"88",
          2352 => x"b9",
          2353 => x"f0",
          2354 => x"08",
          2355 => x"38",
          2356 => x"d5",
          2357 => x"05",
          2358 => x"38",
          2359 => x"08",
          2360 => x"10",
          2361 => x"08",
          2362 => x"82",
          2363 => x"fc",
          2364 => x"82",
          2365 => x"fc",
          2366 => x"b8",
          2367 => x"f0",
          2368 => x"08",
          2369 => x"e1",
          2370 => x"f0",
          2371 => x"08",
          2372 => x"08",
          2373 => x"26",
          2374 => x"d5",
          2375 => x"05",
          2376 => x"f0",
          2377 => x"08",
          2378 => x"f0",
          2379 => x"0c",
          2380 => x"08",
          2381 => x"82",
          2382 => x"fc",
          2383 => x"82",
          2384 => x"f8",
          2385 => x"d5",
          2386 => x"05",
          2387 => x"82",
          2388 => x"fc",
          2389 => x"d5",
          2390 => x"05",
          2391 => x"82",
          2392 => x"8c",
          2393 => x"95",
          2394 => x"f0",
          2395 => x"08",
          2396 => x"38",
          2397 => x"08",
          2398 => x"70",
          2399 => x"08",
          2400 => x"51",
          2401 => x"d5",
          2402 => x"05",
          2403 => x"d5",
          2404 => x"05",
          2405 => x"d5",
          2406 => x"05",
          2407 => x"e4",
          2408 => x"0d",
          2409 => x"0c",
          2410 => x"f0",
          2411 => x"d5",
          2412 => x"3d",
          2413 => x"82",
          2414 => x"f0",
          2415 => x"d5",
          2416 => x"05",
          2417 => x"73",
          2418 => x"f0",
          2419 => x"08",
          2420 => x"53",
          2421 => x"72",
          2422 => x"08",
          2423 => x"72",
          2424 => x"53",
          2425 => x"09",
          2426 => x"38",
          2427 => x"08",
          2428 => x"70",
          2429 => x"71",
          2430 => x"39",
          2431 => x"08",
          2432 => x"53",
          2433 => x"09",
          2434 => x"38",
          2435 => x"d5",
          2436 => x"05",
          2437 => x"f0",
          2438 => x"08",
          2439 => x"05",
          2440 => x"08",
          2441 => x"33",
          2442 => x"08",
          2443 => x"82",
          2444 => x"f8",
          2445 => x"72",
          2446 => x"81",
          2447 => x"38",
          2448 => x"08",
          2449 => x"70",
          2450 => x"71",
          2451 => x"51",
          2452 => x"82",
          2453 => x"f8",
          2454 => x"d5",
          2455 => x"05",
          2456 => x"f0",
          2457 => x"0c",
          2458 => x"08",
          2459 => x"80",
          2460 => x"38",
          2461 => x"08",
          2462 => x"80",
          2463 => x"38",
          2464 => x"90",
          2465 => x"f0",
          2466 => x"34",
          2467 => x"08",
          2468 => x"70",
          2469 => x"71",
          2470 => x"51",
          2471 => x"82",
          2472 => x"f8",
          2473 => x"a4",
          2474 => x"82",
          2475 => x"f4",
          2476 => x"d5",
          2477 => x"05",
          2478 => x"81",
          2479 => x"70",
          2480 => x"72",
          2481 => x"f0",
          2482 => x"34",
          2483 => x"82",
          2484 => x"f8",
          2485 => x"72",
          2486 => x"38",
          2487 => x"d5",
          2488 => x"05",
          2489 => x"39",
          2490 => x"08",
          2491 => x"53",
          2492 => x"90",
          2493 => x"f0",
          2494 => x"33",
          2495 => x"26",
          2496 => x"39",
          2497 => x"d5",
          2498 => x"05",
          2499 => x"39",
          2500 => x"d5",
          2501 => x"05",
          2502 => x"82",
          2503 => x"f8",
          2504 => x"af",
          2505 => x"38",
          2506 => x"08",
          2507 => x"53",
          2508 => x"83",
          2509 => x"80",
          2510 => x"f0",
          2511 => x"0c",
          2512 => x"8a",
          2513 => x"f0",
          2514 => x"34",
          2515 => x"d5",
          2516 => x"05",
          2517 => x"f0",
          2518 => x"33",
          2519 => x"27",
          2520 => x"82",
          2521 => x"f8",
          2522 => x"80",
          2523 => x"94",
          2524 => x"f0",
          2525 => x"33",
          2526 => x"53",
          2527 => x"f0",
          2528 => x"34",
          2529 => x"08",
          2530 => x"d0",
          2531 => x"72",
          2532 => x"08",
          2533 => x"82",
          2534 => x"f8",
          2535 => x"90",
          2536 => x"38",
          2537 => x"08",
          2538 => x"f9",
          2539 => x"72",
          2540 => x"08",
          2541 => x"82",
          2542 => x"f8",
          2543 => x"72",
          2544 => x"38",
          2545 => x"d5",
          2546 => x"05",
          2547 => x"39",
          2548 => x"08",
          2549 => x"82",
          2550 => x"f4",
          2551 => x"54",
          2552 => x"8d",
          2553 => x"82",
          2554 => x"ec",
          2555 => x"f7",
          2556 => x"f0",
          2557 => x"33",
          2558 => x"f0",
          2559 => x"08",
          2560 => x"f0",
          2561 => x"33",
          2562 => x"d5",
          2563 => x"05",
          2564 => x"f0",
          2565 => x"08",
          2566 => x"05",
          2567 => x"08",
          2568 => x"55",
          2569 => x"82",
          2570 => x"f8",
          2571 => x"a5",
          2572 => x"f0",
          2573 => x"33",
          2574 => x"2e",
          2575 => x"d5",
          2576 => x"05",
          2577 => x"d5",
          2578 => x"05",
          2579 => x"f0",
          2580 => x"08",
          2581 => x"08",
          2582 => x"71",
          2583 => x"0b",
          2584 => x"08",
          2585 => x"82",
          2586 => x"ec",
          2587 => x"d5",
          2588 => x"3d",
          2589 => x"f0",
          2590 => x"d5",
          2591 => x"82",
          2592 => x"f7",
          2593 => x"0b",
          2594 => x"08",
          2595 => x"82",
          2596 => x"8c",
          2597 => x"80",
          2598 => x"d5",
          2599 => x"05",
          2600 => x"51",
          2601 => x"53",
          2602 => x"f0",
          2603 => x"34",
          2604 => x"06",
          2605 => x"2e",
          2606 => x"91",
          2607 => x"f0",
          2608 => x"08",
          2609 => x"05",
          2610 => x"ce",
          2611 => x"f0",
          2612 => x"33",
          2613 => x"2e",
          2614 => x"a4",
          2615 => x"82",
          2616 => x"f0",
          2617 => x"d5",
          2618 => x"05",
          2619 => x"81",
          2620 => x"70",
          2621 => x"72",
          2622 => x"f0",
          2623 => x"34",
          2624 => x"08",
          2625 => x"53",
          2626 => x"09",
          2627 => x"dc",
          2628 => x"f0",
          2629 => x"08",
          2630 => x"05",
          2631 => x"08",
          2632 => x"33",
          2633 => x"08",
          2634 => x"82",
          2635 => x"f8",
          2636 => x"d5",
          2637 => x"05",
          2638 => x"f0",
          2639 => x"08",
          2640 => x"b6",
          2641 => x"f0",
          2642 => x"08",
          2643 => x"84",
          2644 => x"39",
          2645 => x"d5",
          2646 => x"05",
          2647 => x"f0",
          2648 => x"08",
          2649 => x"05",
          2650 => x"08",
          2651 => x"33",
          2652 => x"08",
          2653 => x"81",
          2654 => x"0b",
          2655 => x"08",
          2656 => x"82",
          2657 => x"88",
          2658 => x"08",
          2659 => x"0c",
          2660 => x"53",
          2661 => x"d5",
          2662 => x"05",
          2663 => x"39",
          2664 => x"08",
          2665 => x"53",
          2666 => x"8d",
          2667 => x"82",
          2668 => x"ec",
          2669 => x"80",
          2670 => x"f0",
          2671 => x"33",
          2672 => x"27",
          2673 => x"d5",
          2674 => x"05",
          2675 => x"b9",
          2676 => x"8d",
          2677 => x"82",
          2678 => x"ec",
          2679 => x"d8",
          2680 => x"82",
          2681 => x"f4",
          2682 => x"39",
          2683 => x"08",
          2684 => x"53",
          2685 => x"90",
          2686 => x"f0",
          2687 => x"33",
          2688 => x"26",
          2689 => x"39",
          2690 => x"d5",
          2691 => x"05",
          2692 => x"39",
          2693 => x"d5",
          2694 => x"05",
          2695 => x"82",
          2696 => x"fc",
          2697 => x"d5",
          2698 => x"05",
          2699 => x"73",
          2700 => x"38",
          2701 => x"08",
          2702 => x"53",
          2703 => x"27",
          2704 => x"d5",
          2705 => x"05",
          2706 => x"51",
          2707 => x"d5",
          2708 => x"05",
          2709 => x"f0",
          2710 => x"33",
          2711 => x"53",
          2712 => x"f0",
          2713 => x"34",
          2714 => x"08",
          2715 => x"53",
          2716 => x"ad",
          2717 => x"f0",
          2718 => x"33",
          2719 => x"53",
          2720 => x"f0",
          2721 => x"34",
          2722 => x"08",
          2723 => x"53",
          2724 => x"8d",
          2725 => x"82",
          2726 => x"ec",
          2727 => x"98",
          2728 => x"f0",
          2729 => x"33",
          2730 => x"08",
          2731 => x"54",
          2732 => x"26",
          2733 => x"0b",
          2734 => x"08",
          2735 => x"80",
          2736 => x"d5",
          2737 => x"05",
          2738 => x"d5",
          2739 => x"05",
          2740 => x"d5",
          2741 => x"05",
          2742 => x"82",
          2743 => x"fc",
          2744 => x"d5",
          2745 => x"05",
          2746 => x"81",
          2747 => x"70",
          2748 => x"52",
          2749 => x"33",
          2750 => x"08",
          2751 => x"fe",
          2752 => x"d5",
          2753 => x"05",
          2754 => x"80",
          2755 => x"82",
          2756 => x"fc",
          2757 => x"82",
          2758 => x"fc",
          2759 => x"d5",
          2760 => x"05",
          2761 => x"f0",
          2762 => x"08",
          2763 => x"81",
          2764 => x"f0",
          2765 => x"0c",
          2766 => x"08",
          2767 => x"82",
          2768 => x"8b",
          2769 => x"d5",
          2770 => x"f8",
          2771 => x"70",
          2772 => x"56",
          2773 => x"2e",
          2774 => x"8c",
          2775 => x"79",
          2776 => x"33",
          2777 => x"39",
          2778 => x"73",
          2779 => x"81",
          2780 => x"81",
          2781 => x"39",
          2782 => x"90",
          2783 => x"dc",
          2784 => x"52",
          2785 => x"3f",
          2786 => x"08",
          2787 => x"08",
          2788 => x"76",
          2789 => x"e7",
          2790 => x"d5",
          2791 => x"38",
          2792 => x"54",
          2793 => x"ff",
          2794 => x"17",
          2795 => x"06",
          2796 => x"77",
          2797 => x"ff",
          2798 => x"d5",
          2799 => x"3d",
          2800 => x"3d",
          2801 => x"71",
          2802 => x"8e",
          2803 => x"29",
          2804 => x"05",
          2805 => x"04",
          2806 => x"51",
          2807 => x"82",
          2808 => x"80",
          2809 => x"b3",
          2810 => x"f2",
          2811 => x"c8",
          2812 => x"39",
          2813 => x"51",
          2814 => x"82",
          2815 => x"80",
          2816 => x"b3",
          2817 => x"d6",
          2818 => x"8c",
          2819 => x"39",
          2820 => x"51",
          2821 => x"82",
          2822 => x"80",
          2823 => x"b4",
          2824 => x"39",
          2825 => x"51",
          2826 => x"b5",
          2827 => x"39",
          2828 => x"51",
          2829 => x"b5",
          2830 => x"39",
          2831 => x"51",
          2832 => x"b5",
          2833 => x"39",
          2834 => x"51",
          2835 => x"b6",
          2836 => x"39",
          2837 => x"51",
          2838 => x"b6",
          2839 => x"86",
          2840 => x"0d",
          2841 => x"0d",
          2842 => x"56",
          2843 => x"26",
          2844 => x"52",
          2845 => x"29",
          2846 => x"87",
          2847 => x"51",
          2848 => x"82",
          2849 => x"52",
          2850 => x"a5",
          2851 => x"e4",
          2852 => x"53",
          2853 => x"b6",
          2854 => x"ba",
          2855 => x"3d",
          2856 => x"3d",
          2857 => x"84",
          2858 => x"05",
          2859 => x"80",
          2860 => x"70",
          2861 => x"25",
          2862 => x"59",
          2863 => x"87",
          2864 => x"38",
          2865 => x"76",
          2866 => x"ff",
          2867 => x"93",
          2868 => x"82",
          2869 => x"76",
          2870 => x"70",
          2871 => x"91",
          2872 => x"d5",
          2873 => x"82",
          2874 => x"b9",
          2875 => x"e4",
          2876 => x"98",
          2877 => x"d5",
          2878 => x"96",
          2879 => x"54",
          2880 => x"77",
          2881 => x"81",
          2882 => x"82",
          2883 => x"57",
          2884 => x"08",
          2885 => x"55",
          2886 => x"89",
          2887 => x"75",
          2888 => x"d7",
          2889 => x"d8",
          2890 => x"9e",
          2891 => x"30",
          2892 => x"80",
          2893 => x"70",
          2894 => x"06",
          2895 => x"56",
          2896 => x"90",
          2897 => x"f4",
          2898 => x"98",
          2899 => x"78",
          2900 => x"3f",
          2901 => x"82",
          2902 => x"96",
          2903 => x"f8",
          2904 => x"02",
          2905 => x"05",
          2906 => x"ff",
          2907 => x"7b",
          2908 => x"fe",
          2909 => x"d5",
          2910 => x"38",
          2911 => x"88",
          2912 => x"2e",
          2913 => x"39",
          2914 => x"56",
          2915 => x"54",
          2916 => x"53",
          2917 => x"51",
          2918 => x"d5",
          2919 => x"83",
          2920 => x"77",
          2921 => x"0c",
          2922 => x"04",
          2923 => x"7f",
          2924 => x"8c",
          2925 => x"05",
          2926 => x"15",
          2927 => x"5c",
          2928 => x"5e",
          2929 => x"b6",
          2930 => x"b8",
          2931 => x"b7",
          2932 => x"b8",
          2933 => x"55",
          2934 => x"81",
          2935 => x"90",
          2936 => x"7b",
          2937 => x"38",
          2938 => x"74",
          2939 => x"7a",
          2940 => x"72",
          2941 => x"b7",
          2942 => x"b7",
          2943 => x"39",
          2944 => x"51",
          2945 => x"3f",
          2946 => x"80",
          2947 => x"18",
          2948 => x"27",
          2949 => x"08",
          2950 => x"fc",
          2951 => x"bb",
          2952 => x"82",
          2953 => x"ff",
          2954 => x"84",
          2955 => x"39",
          2956 => x"72",
          2957 => x"38",
          2958 => x"82",
          2959 => x"ff",
          2960 => x"89",
          2961 => x"a4",
          2962 => x"8f",
          2963 => x"55",
          2964 => x"08",
          2965 => x"d6",
          2966 => x"fc",
          2967 => x"a8",
          2968 => x"f7",
          2969 => x"74",
          2970 => x"c6",
          2971 => x"70",
          2972 => x"80",
          2973 => x"27",
          2974 => x"56",
          2975 => x"74",
          2976 => x"81",
          2977 => x"06",
          2978 => x"06",
          2979 => x"80",
          2980 => x"73",
          2981 => x"8a",
          2982 => x"c8",
          2983 => x"51",
          2984 => x"f1",
          2985 => x"a0",
          2986 => x"3f",
          2987 => x"ff",
          2988 => x"b7",
          2989 => x"ae",
          2990 => x"79",
          2991 => x"9d",
          2992 => x"d5",
          2993 => x"2b",
          2994 => x"51",
          2995 => x"2e",
          2996 => x"aa",
          2997 => x"3f",
          2998 => x"08",
          2999 => x"98",
          3000 => x"32",
          3001 => x"9b",
          3002 => x"70",
          3003 => x"75",
          3004 => x"58",
          3005 => x"51",
          3006 => x"24",
          3007 => x"9b",
          3008 => x"06",
          3009 => x"53",
          3010 => x"1e",
          3011 => x"26",
          3012 => x"ff",
          3013 => x"d5",
          3014 => x"3d",
          3015 => x"3d",
          3016 => x"05",
          3017 => x"b0",
          3018 => x"b4",
          3019 => x"b5",
          3020 => x"d4",
          3021 => x"a5",
          3022 => x"b7",
          3023 => x"b7",
          3024 => x"d4",
          3025 => x"82",
          3026 => x"ff",
          3027 => x"74",
          3028 => x"38",
          3029 => x"86",
          3030 => x"fe",
          3031 => x"c0",
          3032 => x"53",
          3033 => x"81",
          3034 => x"3f",
          3035 => x"51",
          3036 => x"80",
          3037 => x"3f",
          3038 => x"70",
          3039 => x"52",
          3040 => x"92",
          3041 => x"98",
          3042 => x"b8",
          3043 => x"c4",
          3044 => x"98",
          3045 => x"82",
          3046 => x"06",
          3047 => x"80",
          3048 => x"81",
          3049 => x"3f",
          3050 => x"51",
          3051 => x"80",
          3052 => x"3f",
          3053 => x"70",
          3054 => x"52",
          3055 => x"92",
          3056 => x"97",
          3057 => x"b8",
          3058 => x"88",
          3059 => x"97",
          3060 => x"84",
          3061 => x"06",
          3062 => x"80",
          3063 => x"81",
          3064 => x"3f",
          3065 => x"51",
          3066 => x"80",
          3067 => x"3f",
          3068 => x"70",
          3069 => x"52",
          3070 => x"92",
          3071 => x"97",
          3072 => x"b8",
          3073 => x"cc",
          3074 => x"97",
          3075 => x"86",
          3076 => x"06",
          3077 => x"80",
          3078 => x"81",
          3079 => x"3f",
          3080 => x"51",
          3081 => x"80",
          3082 => x"3f",
          3083 => x"70",
          3084 => x"52",
          3085 => x"92",
          3086 => x"96",
          3087 => x"b8",
          3088 => x"90",
          3089 => x"96",
          3090 => x"88",
          3091 => x"06",
          3092 => x"80",
          3093 => x"81",
          3094 => x"3f",
          3095 => x"51",
          3096 => x"80",
          3097 => x"3f",
          3098 => x"84",
          3099 => x"fb",
          3100 => x"02",
          3101 => x"05",
          3102 => x"56",
          3103 => x"75",
          3104 => x"3f",
          3105 => x"d0",
          3106 => x"73",
          3107 => x"53",
          3108 => x"52",
          3109 => x"51",
          3110 => x"3f",
          3111 => x"08",
          3112 => x"d5",
          3113 => x"80",
          3114 => x"31",
          3115 => x"73",
          3116 => x"d0",
          3117 => x"0b",
          3118 => x"33",
          3119 => x"2e",
          3120 => x"af",
          3121 => x"f4",
          3122 => x"75",
          3123 => x"b8",
          3124 => x"e4",
          3125 => x"8b",
          3126 => x"e4",
          3127 => x"86",
          3128 => x"82",
          3129 => x"81",
          3130 => x"82",
          3131 => x"82",
          3132 => x"0b",
          3133 => x"d8",
          3134 => x"82",
          3135 => x"06",
          3136 => x"b9",
          3137 => x"52",
          3138 => x"fb",
          3139 => x"82",
          3140 => x"87",
          3141 => x"cd",
          3142 => x"70",
          3143 => x"7e",
          3144 => x"0c",
          3145 => x"7d",
          3146 => x"93",
          3147 => x"e4",
          3148 => x"06",
          3149 => x"2e",
          3150 => x"a3",
          3151 => x"59",
          3152 => x"b9",
          3153 => x"51",
          3154 => x"7d",
          3155 => x"82",
          3156 => x"81",
          3157 => x"82",
          3158 => x"7e",
          3159 => x"82",
          3160 => x"8d",
          3161 => x"70",
          3162 => x"ba",
          3163 => x"b0",
          3164 => x"3d",
          3165 => x"80",
          3166 => x"51",
          3167 => x"b5",
          3168 => x"05",
          3169 => x"3f",
          3170 => x"08",
          3171 => x"90",
          3172 => x"78",
          3173 => x"87",
          3174 => x"80",
          3175 => x"38",
          3176 => x"81",
          3177 => x"bd",
          3178 => x"78",
          3179 => x"ba",
          3180 => x"2e",
          3181 => x"8a",
          3182 => x"80",
          3183 => x"99",
          3184 => x"c0",
          3185 => x"38",
          3186 => x"82",
          3187 => x"bf",
          3188 => x"f9",
          3189 => x"38",
          3190 => x"24",
          3191 => x"80",
          3192 => x"8a",
          3193 => x"f8",
          3194 => x"38",
          3195 => x"78",
          3196 => x"8a",
          3197 => x"81",
          3198 => x"38",
          3199 => x"2e",
          3200 => x"8a",
          3201 => x"81",
          3202 => x"fd",
          3203 => x"39",
          3204 => x"80",
          3205 => x"84",
          3206 => x"de",
          3207 => x"e4",
          3208 => x"fe",
          3209 => x"3d",
          3210 => x"53",
          3211 => x"51",
          3212 => x"82",
          3213 => x"80",
          3214 => x"38",
          3215 => x"f8",
          3216 => x"84",
          3217 => x"b2",
          3218 => x"e4",
          3219 => x"82",
          3220 => x"43",
          3221 => x"51",
          3222 => x"3f",
          3223 => x"5a",
          3224 => x"81",
          3225 => x"59",
          3226 => x"84",
          3227 => x"7a",
          3228 => x"38",
          3229 => x"b5",
          3230 => x"11",
          3231 => x"05",
          3232 => x"3f",
          3233 => x"08",
          3234 => x"de",
          3235 => x"fe",
          3236 => x"ff",
          3237 => x"eb",
          3238 => x"d5",
          3239 => x"2e",
          3240 => x"b5",
          3241 => x"11",
          3242 => x"05",
          3243 => x"3f",
          3244 => x"08",
          3245 => x"b2",
          3246 => x"b4",
          3247 => x"9b",
          3248 => x"79",
          3249 => x"89",
          3250 => x"79",
          3251 => x"5b",
          3252 => x"62",
          3253 => x"eb",
          3254 => x"ff",
          3255 => x"ff",
          3256 => x"eb",
          3257 => x"d5",
          3258 => x"2e",
          3259 => x"b5",
          3260 => x"11",
          3261 => x"05",
          3262 => x"3f",
          3263 => x"08",
          3264 => x"e6",
          3265 => x"fe",
          3266 => x"ff",
          3267 => x"ea",
          3268 => x"d5",
          3269 => x"2e",
          3270 => x"82",
          3271 => x"ff",
          3272 => x"64",
          3273 => x"27",
          3274 => x"70",
          3275 => x"5e",
          3276 => x"7c",
          3277 => x"78",
          3278 => x"79",
          3279 => x"52",
          3280 => x"51",
          3281 => x"3f",
          3282 => x"81",
          3283 => x"d5",
          3284 => x"cc",
          3285 => x"92",
          3286 => x"ff",
          3287 => x"ff",
          3288 => x"ea",
          3289 => x"d5",
          3290 => x"df",
          3291 => x"c8",
          3292 => x"80",
          3293 => x"82",
          3294 => x"45",
          3295 => x"82",
          3296 => x"59",
          3297 => x"88",
          3298 => x"88",
          3299 => x"39",
          3300 => x"33",
          3301 => x"2e",
          3302 => x"d4",
          3303 => x"ab",
          3304 => x"cb",
          3305 => x"80",
          3306 => x"82",
          3307 => x"45",
          3308 => x"d4",
          3309 => x"78",
          3310 => x"38",
          3311 => x"08",
          3312 => x"82",
          3313 => x"fc",
          3314 => x"b5",
          3315 => x"11",
          3316 => x"05",
          3317 => x"3f",
          3318 => x"08",
          3319 => x"82",
          3320 => x"59",
          3321 => x"89",
          3322 => x"84",
          3323 => x"cc",
          3324 => x"c9",
          3325 => x"80",
          3326 => x"82",
          3327 => x"44",
          3328 => x"d4",
          3329 => x"78",
          3330 => x"38",
          3331 => x"08",
          3332 => x"82",
          3333 => x"59",
          3334 => x"88",
          3335 => x"9c",
          3336 => x"39",
          3337 => x"33",
          3338 => x"2e",
          3339 => x"d4",
          3340 => x"88",
          3341 => x"b0",
          3342 => x"44",
          3343 => x"f8",
          3344 => x"84",
          3345 => x"b2",
          3346 => x"e4",
          3347 => x"a7",
          3348 => x"5c",
          3349 => x"2e",
          3350 => x"5c",
          3351 => x"70",
          3352 => x"07",
          3353 => x"7f",
          3354 => x"5a",
          3355 => x"2e",
          3356 => x"a0",
          3357 => x"88",
          3358 => x"ec",
          3359 => x"3f",
          3360 => x"54",
          3361 => x"52",
          3362 => x"a0",
          3363 => x"f8",
          3364 => x"39",
          3365 => x"80",
          3366 => x"84",
          3367 => x"da",
          3368 => x"e4",
          3369 => x"f9",
          3370 => x"3d",
          3371 => x"53",
          3372 => x"51",
          3373 => x"82",
          3374 => x"80",
          3375 => x"64",
          3376 => x"cf",
          3377 => x"34",
          3378 => x"45",
          3379 => x"fc",
          3380 => x"84",
          3381 => x"a2",
          3382 => x"e4",
          3383 => x"f9",
          3384 => x"70",
          3385 => x"82",
          3386 => x"ff",
          3387 => x"82",
          3388 => x"53",
          3389 => x"79",
          3390 => x"b4",
          3391 => x"79",
          3392 => x"ae",
          3393 => x"38",
          3394 => x"9f",
          3395 => x"fe",
          3396 => x"ff",
          3397 => x"e6",
          3398 => x"d5",
          3399 => x"2e",
          3400 => x"59",
          3401 => x"05",
          3402 => x"64",
          3403 => x"ff",
          3404 => x"bb",
          3405 => x"ae",
          3406 => x"39",
          3407 => x"f4",
          3408 => x"84",
          3409 => x"e1",
          3410 => x"e4",
          3411 => x"f8",
          3412 => x"3d",
          3413 => x"53",
          3414 => x"51",
          3415 => x"82",
          3416 => x"80",
          3417 => x"61",
          3418 => x"c2",
          3419 => x"70",
          3420 => x"23",
          3421 => x"3d",
          3422 => x"53",
          3423 => x"51",
          3424 => x"82",
          3425 => x"df",
          3426 => x"39",
          3427 => x"54",
          3428 => x"94",
          3429 => x"c3",
          3430 => x"c4",
          3431 => x"f8",
          3432 => x"ff",
          3433 => x"79",
          3434 => x"59",
          3435 => x"f7",
          3436 => x"9f",
          3437 => x"61",
          3438 => x"d0",
          3439 => x"fe",
          3440 => x"ff",
          3441 => x"df",
          3442 => x"d5",
          3443 => x"2e",
          3444 => x"59",
          3445 => x"05",
          3446 => x"82",
          3447 => x"78",
          3448 => x"39",
          3449 => x"51",
          3450 => x"ff",
          3451 => x"3d",
          3452 => x"53",
          3453 => x"51",
          3454 => x"82",
          3455 => x"80",
          3456 => x"38",
          3457 => x"f0",
          3458 => x"84",
          3459 => x"99",
          3460 => x"e4",
          3461 => x"a0",
          3462 => x"71",
          3463 => x"84",
          3464 => x"3d",
          3465 => x"53",
          3466 => x"51",
          3467 => x"82",
          3468 => x"e5",
          3469 => x"39",
          3470 => x"54",
          3471 => x"a0",
          3472 => x"97",
          3473 => x"c4",
          3474 => x"f8",
          3475 => x"ff",
          3476 => x"79",
          3477 => x"59",
          3478 => x"f6",
          3479 => x"79",
          3480 => x"b5",
          3481 => x"11",
          3482 => x"05",
          3483 => x"3f",
          3484 => x"08",
          3485 => x"38",
          3486 => x"0c",
          3487 => x"05",
          3488 => x"39",
          3489 => x"51",
          3490 => x"ff",
          3491 => x"3d",
          3492 => x"53",
          3493 => x"51",
          3494 => x"82",
          3495 => x"80",
          3496 => x"38",
          3497 => x"bb",
          3498 => x"a6",
          3499 => x"59",
          3500 => x"3d",
          3501 => x"53",
          3502 => x"51",
          3503 => x"82",
          3504 => x"80",
          3505 => x"38",
          3506 => x"bb",
          3507 => x"a6",
          3508 => x"59",
          3509 => x"d5",
          3510 => x"2e",
          3511 => x"82",
          3512 => x"52",
          3513 => x"51",
          3514 => x"3f",
          3515 => x"82",
          3516 => x"c1",
          3517 => x"a5",
          3518 => x"ee",
          3519 => x"a0",
          3520 => x"3f",
          3521 => x"a8",
          3522 => x"3f",
          3523 => x"97",
          3524 => x"78",
          3525 => x"d2",
          3526 => x"52",
          3527 => x"9c",
          3528 => x"e4",
          3529 => x"d5",
          3530 => x"2e",
          3531 => x"82",
          3532 => x"46",
          3533 => x"84",
          3534 => x"f5",
          3535 => x"e4",
          3536 => x"06",
          3537 => x"80",
          3538 => x"38",
          3539 => x"08",
          3540 => x"3f",
          3541 => x"08",
          3542 => x"c1",
          3543 => x"7a",
          3544 => x"38",
          3545 => x"89",
          3546 => x"2e",
          3547 => x"ca",
          3548 => x"2e",
          3549 => x"c2",
          3550 => x"b4",
          3551 => x"82",
          3552 => x"80",
          3553 => x"bc",
          3554 => x"ff",
          3555 => x"ff",
          3556 => x"b8",
          3557 => x"b5",
          3558 => x"05",
          3559 => x"3f",
          3560 => x"55",
          3561 => x"54",
          3562 => x"bc",
          3563 => x"3d",
          3564 => x"51",
          3565 => x"3f",
          3566 => x"54",
          3567 => x"bc",
          3568 => x"3d",
          3569 => x"51",
          3570 => x"3f",
          3571 => x"58",
          3572 => x"57",
          3573 => x"55",
          3574 => x"80",
          3575 => x"80",
          3576 => x"3d",
          3577 => x"51",
          3578 => x"82",
          3579 => x"82",
          3580 => x"09",
          3581 => x"72",
          3582 => x"51",
          3583 => x"80",
          3584 => x"26",
          3585 => x"5a",
          3586 => x"59",
          3587 => x"8d",
          3588 => x"70",
          3589 => x"5c",
          3590 => x"c3",
          3591 => x"32",
          3592 => x"07",
          3593 => x"38",
          3594 => x"09",
          3595 => x"38",
          3596 => x"51",
          3597 => x"3f",
          3598 => x"80",
          3599 => x"39",
          3600 => x"51",
          3601 => x"3f",
          3602 => x"f5",
          3603 => x"0b",
          3604 => x"34",
          3605 => x"8c",
          3606 => x"55",
          3607 => x"52",
          3608 => x"cd",
          3609 => x"e4",
          3610 => x"75",
          3611 => x"87",
          3612 => x"73",
          3613 => x"3f",
          3614 => x"e4",
          3615 => x"0c",
          3616 => x"9c",
          3617 => x"55",
          3618 => x"52",
          3619 => x"a1",
          3620 => x"e4",
          3621 => x"75",
          3622 => x"87",
          3623 => x"73",
          3624 => x"3f",
          3625 => x"e4",
          3626 => x"0c",
          3627 => x"0b",
          3628 => x"84",
          3629 => x"83",
          3630 => x"94",
          3631 => x"f7",
          3632 => x"fa",
          3633 => x"02",
          3634 => x"05",
          3635 => x"82",
          3636 => x"87",
          3637 => x"13",
          3638 => x"0c",
          3639 => x"0c",
          3640 => x"3f",
          3641 => x"82",
          3642 => x"ff",
          3643 => x"82",
          3644 => x"ff",
          3645 => x"80",
          3646 => x"92",
          3647 => x"51",
          3648 => x"f0",
          3649 => x"04",
          3650 => x"80",
          3651 => x"71",
          3652 => x"87",
          3653 => x"d5",
          3654 => x"ff",
          3655 => x"ff",
          3656 => x"72",
          3657 => x"38",
          3658 => x"e4",
          3659 => x"0d",
          3660 => x"0d",
          3661 => x"54",
          3662 => x"52",
          3663 => x"2e",
          3664 => x"72",
          3665 => x"a0",
          3666 => x"06",
          3667 => x"13",
          3668 => x"72",
          3669 => x"a2",
          3670 => x"06",
          3671 => x"13",
          3672 => x"72",
          3673 => x"2e",
          3674 => x"9f",
          3675 => x"81",
          3676 => x"72",
          3677 => x"70",
          3678 => x"38",
          3679 => x"80",
          3680 => x"73",
          3681 => x"39",
          3682 => x"80",
          3683 => x"54",
          3684 => x"83",
          3685 => x"70",
          3686 => x"38",
          3687 => x"80",
          3688 => x"54",
          3689 => x"09",
          3690 => x"38",
          3691 => x"a2",
          3692 => x"70",
          3693 => x"07",
          3694 => x"70",
          3695 => x"38",
          3696 => x"81",
          3697 => x"71",
          3698 => x"51",
          3699 => x"e4",
          3700 => x"0d",
          3701 => x"0d",
          3702 => x"08",
          3703 => x"38",
          3704 => x"05",
          3705 => x"d7",
          3706 => x"d5",
          3707 => x"38",
          3708 => x"39",
          3709 => x"82",
          3710 => x"86",
          3711 => x"fc",
          3712 => x"82",
          3713 => x"05",
          3714 => x"52",
          3715 => x"81",
          3716 => x"13",
          3717 => x"51",
          3718 => x"9e",
          3719 => x"38",
          3720 => x"51",
          3721 => x"97",
          3722 => x"38",
          3723 => x"51",
          3724 => x"bb",
          3725 => x"38",
          3726 => x"51",
          3727 => x"bb",
          3728 => x"38",
          3729 => x"55",
          3730 => x"87",
          3731 => x"d9",
          3732 => x"22",
          3733 => x"73",
          3734 => x"80",
          3735 => x"0b",
          3736 => x"9c",
          3737 => x"87",
          3738 => x"0c",
          3739 => x"87",
          3740 => x"0c",
          3741 => x"87",
          3742 => x"0c",
          3743 => x"87",
          3744 => x"0c",
          3745 => x"87",
          3746 => x"0c",
          3747 => x"87",
          3748 => x"0c",
          3749 => x"98",
          3750 => x"87",
          3751 => x"0c",
          3752 => x"c0",
          3753 => x"80",
          3754 => x"d5",
          3755 => x"3d",
          3756 => x"3d",
          3757 => x"87",
          3758 => x"5d",
          3759 => x"87",
          3760 => x"08",
          3761 => x"23",
          3762 => x"b8",
          3763 => x"82",
          3764 => x"c0",
          3765 => x"5a",
          3766 => x"34",
          3767 => x"b0",
          3768 => x"84",
          3769 => x"c0",
          3770 => x"5a",
          3771 => x"34",
          3772 => x"a8",
          3773 => x"86",
          3774 => x"c0",
          3775 => x"5c",
          3776 => x"23",
          3777 => x"a0",
          3778 => x"8a",
          3779 => x"7d",
          3780 => x"ff",
          3781 => x"7b",
          3782 => x"06",
          3783 => x"33",
          3784 => x"33",
          3785 => x"33",
          3786 => x"33",
          3787 => x"33",
          3788 => x"ff",
          3789 => x"82",
          3790 => x"ff",
          3791 => x"8f",
          3792 => x"fb",
          3793 => x"9f",
          3794 => x"d3",
          3795 => x"81",
          3796 => x"55",
          3797 => x"94",
          3798 => x"80",
          3799 => x"87",
          3800 => x"51",
          3801 => x"96",
          3802 => x"06",
          3803 => x"70",
          3804 => x"38",
          3805 => x"70",
          3806 => x"51",
          3807 => x"72",
          3808 => x"81",
          3809 => x"70",
          3810 => x"38",
          3811 => x"70",
          3812 => x"51",
          3813 => x"38",
          3814 => x"06",
          3815 => x"94",
          3816 => x"80",
          3817 => x"87",
          3818 => x"52",
          3819 => x"74",
          3820 => x"0c",
          3821 => x"04",
          3822 => x"02",
          3823 => x"70",
          3824 => x"2a",
          3825 => x"70",
          3826 => x"34",
          3827 => x"04",
          3828 => x"02",
          3829 => x"58",
          3830 => x"09",
          3831 => x"38",
          3832 => x"51",
          3833 => x"d3",
          3834 => x"81",
          3835 => x"56",
          3836 => x"84",
          3837 => x"2e",
          3838 => x"c0",
          3839 => x"72",
          3840 => x"2a",
          3841 => x"55",
          3842 => x"80",
          3843 => x"73",
          3844 => x"81",
          3845 => x"72",
          3846 => x"81",
          3847 => x"06",
          3848 => x"80",
          3849 => x"73",
          3850 => x"81",
          3851 => x"72",
          3852 => x"75",
          3853 => x"53",
          3854 => x"80",
          3855 => x"2e",
          3856 => x"c0",
          3857 => x"77",
          3858 => x"0b",
          3859 => x"0c",
          3860 => x"04",
          3861 => x"79",
          3862 => x"33",
          3863 => x"06",
          3864 => x"70",
          3865 => x"fc",
          3866 => x"ff",
          3867 => x"82",
          3868 => x"70",
          3869 => x"59",
          3870 => x"87",
          3871 => x"51",
          3872 => x"86",
          3873 => x"94",
          3874 => x"08",
          3875 => x"70",
          3876 => x"54",
          3877 => x"2e",
          3878 => x"91",
          3879 => x"06",
          3880 => x"d7",
          3881 => x"32",
          3882 => x"51",
          3883 => x"2e",
          3884 => x"93",
          3885 => x"06",
          3886 => x"ff",
          3887 => x"81",
          3888 => x"87",
          3889 => x"52",
          3890 => x"86",
          3891 => x"94",
          3892 => x"72",
          3893 => x"74",
          3894 => x"ff",
          3895 => x"57",
          3896 => x"38",
          3897 => x"e4",
          3898 => x"0d",
          3899 => x"0d",
          3900 => x"33",
          3901 => x"06",
          3902 => x"c0",
          3903 => x"72",
          3904 => x"38",
          3905 => x"94",
          3906 => x"70",
          3907 => x"81",
          3908 => x"51",
          3909 => x"e2",
          3910 => x"ff",
          3911 => x"c0",
          3912 => x"70",
          3913 => x"38",
          3914 => x"90",
          3915 => x"70",
          3916 => x"82",
          3917 => x"51",
          3918 => x"04",
          3919 => x"82",
          3920 => x"81",
          3921 => x"d5",
          3922 => x"fe",
          3923 => x"d3",
          3924 => x"81",
          3925 => x"53",
          3926 => x"84",
          3927 => x"2e",
          3928 => x"c0",
          3929 => x"71",
          3930 => x"2a",
          3931 => x"51",
          3932 => x"52",
          3933 => x"a0",
          3934 => x"ff",
          3935 => x"c0",
          3936 => x"70",
          3937 => x"38",
          3938 => x"90",
          3939 => x"70",
          3940 => x"98",
          3941 => x"51",
          3942 => x"e4",
          3943 => x"0d",
          3944 => x"0d",
          3945 => x"80",
          3946 => x"2a",
          3947 => x"51",
          3948 => x"84",
          3949 => x"c0",
          3950 => x"82",
          3951 => x"87",
          3952 => x"08",
          3953 => x"0c",
          3954 => x"94",
          3955 => x"88",
          3956 => x"9e",
          3957 => x"d4",
          3958 => x"c0",
          3959 => x"82",
          3960 => x"87",
          3961 => x"08",
          3962 => x"0c",
          3963 => x"ac",
          3964 => x"98",
          3965 => x"9e",
          3966 => x"d4",
          3967 => x"c0",
          3968 => x"82",
          3969 => x"87",
          3970 => x"08",
          3971 => x"0c",
          3972 => x"bc",
          3973 => x"a8",
          3974 => x"9e",
          3975 => x"d4",
          3976 => x"c0",
          3977 => x"82",
          3978 => x"87",
          3979 => x"08",
          3980 => x"d4",
          3981 => x"c0",
          3982 => x"82",
          3983 => x"87",
          3984 => x"08",
          3985 => x"0c",
          3986 => x"8c",
          3987 => x"c0",
          3988 => x"82",
          3989 => x"80",
          3990 => x"9e",
          3991 => x"84",
          3992 => x"51",
          3993 => x"80",
          3994 => x"81",
          3995 => x"d4",
          3996 => x"0b",
          3997 => x"90",
          3998 => x"80",
          3999 => x"52",
          4000 => x"2e",
          4001 => x"52",
          4002 => x"c6",
          4003 => x"87",
          4004 => x"08",
          4005 => x"0a",
          4006 => x"52",
          4007 => x"83",
          4008 => x"71",
          4009 => x"34",
          4010 => x"c0",
          4011 => x"70",
          4012 => x"06",
          4013 => x"70",
          4014 => x"38",
          4015 => x"82",
          4016 => x"80",
          4017 => x"9e",
          4018 => x"a0",
          4019 => x"51",
          4020 => x"80",
          4021 => x"81",
          4022 => x"d4",
          4023 => x"0b",
          4024 => x"90",
          4025 => x"80",
          4026 => x"52",
          4027 => x"2e",
          4028 => x"52",
          4029 => x"ca",
          4030 => x"87",
          4031 => x"08",
          4032 => x"80",
          4033 => x"52",
          4034 => x"83",
          4035 => x"71",
          4036 => x"34",
          4037 => x"c0",
          4038 => x"70",
          4039 => x"06",
          4040 => x"70",
          4041 => x"38",
          4042 => x"82",
          4043 => x"80",
          4044 => x"9e",
          4045 => x"81",
          4046 => x"51",
          4047 => x"80",
          4048 => x"81",
          4049 => x"d4",
          4050 => x"0b",
          4051 => x"90",
          4052 => x"c0",
          4053 => x"52",
          4054 => x"2e",
          4055 => x"52",
          4056 => x"ce",
          4057 => x"87",
          4058 => x"08",
          4059 => x"06",
          4060 => x"70",
          4061 => x"38",
          4062 => x"82",
          4063 => x"87",
          4064 => x"08",
          4065 => x"06",
          4066 => x"51",
          4067 => x"82",
          4068 => x"80",
          4069 => x"9e",
          4070 => x"84",
          4071 => x"52",
          4072 => x"2e",
          4073 => x"52",
          4074 => x"d1",
          4075 => x"9e",
          4076 => x"83",
          4077 => x"84",
          4078 => x"51",
          4079 => x"d2",
          4080 => x"87",
          4081 => x"08",
          4082 => x"51",
          4083 => x"80",
          4084 => x"81",
          4085 => x"d4",
          4086 => x"c0",
          4087 => x"70",
          4088 => x"51",
          4089 => x"d4",
          4090 => x"0d",
          4091 => x"0d",
          4092 => x"51",
          4093 => x"3f",
          4094 => x"33",
          4095 => x"2e",
          4096 => x"bd",
          4097 => x"93",
          4098 => x"be",
          4099 => x"af",
          4100 => x"d4",
          4101 => x"73",
          4102 => x"38",
          4103 => x"08",
          4104 => x"08",
          4105 => x"82",
          4106 => x"ff",
          4107 => x"82",
          4108 => x"54",
          4109 => x"94",
          4110 => x"98",
          4111 => x"9c",
          4112 => x"52",
          4113 => x"51",
          4114 => x"3f",
          4115 => x"33",
          4116 => x"2e",
          4117 => x"d4",
          4118 => x"d4",
          4119 => x"54",
          4120 => x"d0",
          4121 => x"f3",
          4122 => x"c9",
          4123 => x"80",
          4124 => x"82",
          4125 => x"82",
          4126 => x"11",
          4127 => x"be",
          4128 => x"92",
          4129 => x"d4",
          4130 => x"73",
          4131 => x"38",
          4132 => x"08",
          4133 => x"08",
          4134 => x"82",
          4135 => x"ff",
          4136 => x"82",
          4137 => x"54",
          4138 => x"8e",
          4139 => x"d0",
          4140 => x"bf",
          4141 => x"92",
          4142 => x"d4",
          4143 => x"73",
          4144 => x"38",
          4145 => x"33",
          4146 => x"c4",
          4147 => x"8b",
          4148 => x"d1",
          4149 => x"80",
          4150 => x"82",
          4151 => x"52",
          4152 => x"51",
          4153 => x"3f",
          4154 => x"33",
          4155 => x"2e",
          4156 => x"c0",
          4157 => x"ad",
          4158 => x"d4",
          4159 => x"73",
          4160 => x"38",
          4161 => x"51",
          4162 => x"3f",
          4163 => x"33",
          4164 => x"2e",
          4165 => x"c0",
          4166 => x"ad",
          4167 => x"d4",
          4168 => x"73",
          4169 => x"38",
          4170 => x"51",
          4171 => x"3f",
          4172 => x"33",
          4173 => x"2e",
          4174 => x"c0",
          4175 => x"ad",
          4176 => x"c0",
          4177 => x"ad",
          4178 => x"d4",
          4179 => x"82",
          4180 => x"ff",
          4181 => x"82",
          4182 => x"52",
          4183 => x"51",
          4184 => x"3f",
          4185 => x"08",
          4186 => x"9c",
          4187 => x"eb",
          4188 => x"c4",
          4189 => x"ee",
          4190 => x"b4",
          4191 => x"c1",
          4192 => x"90",
          4193 => x"d4",
          4194 => x"bd",
          4195 => x"75",
          4196 => x"3f",
          4197 => x"08",
          4198 => x"29",
          4199 => x"54",
          4200 => x"e4",
          4201 => x"c1",
          4202 => x"90",
          4203 => x"d4",
          4204 => x"73",
          4205 => x"38",
          4206 => x"08",
          4207 => x"c0",
          4208 => x"c4",
          4209 => x"d5",
          4210 => x"84",
          4211 => x"71",
          4212 => x"82",
          4213 => x"52",
          4214 => x"51",
          4215 => x"3f",
          4216 => x"33",
          4217 => x"2e",
          4218 => x"d4",
          4219 => x"bd",
          4220 => x"75",
          4221 => x"3f",
          4222 => x"08",
          4223 => x"29",
          4224 => x"54",
          4225 => x"e4",
          4226 => x"c2",
          4227 => x"8f",
          4228 => x"51",
          4229 => x"3f",
          4230 => x"04",
          4231 => x"02",
          4232 => x"ff",
          4233 => x"84",
          4234 => x"71",
          4235 => x"ad",
          4236 => x"71",
          4237 => x"c2",
          4238 => x"39",
          4239 => x"51",
          4240 => x"c3",
          4241 => x"39",
          4242 => x"51",
          4243 => x"c3",
          4244 => x"39",
          4245 => x"51",
          4246 => x"3f",
          4247 => x"04",
          4248 => x"0c",
          4249 => x"87",
          4250 => x"0c",
          4251 => x"d8",
          4252 => x"96",
          4253 => x"fd",
          4254 => x"98",
          4255 => x"2c",
          4256 => x"70",
          4257 => x"10",
          4258 => x"2b",
          4259 => x"54",
          4260 => x"0b",
          4261 => x"12",
          4262 => x"71",
          4263 => x"38",
          4264 => x"11",
          4265 => x"84",
          4266 => x"33",
          4267 => x"52",
          4268 => x"2e",
          4269 => x"83",
          4270 => x"72",
          4271 => x"0c",
          4272 => x"04",
          4273 => x"79",
          4274 => x"a3",
          4275 => x"33",
          4276 => x"72",
          4277 => x"38",
          4278 => x"08",
          4279 => x"ff",
          4280 => x"82",
          4281 => x"52",
          4282 => x"ad",
          4283 => x"f1",
          4284 => x"88",
          4285 => x"bd",
          4286 => x"ff",
          4287 => x"74",
          4288 => x"ff",
          4289 => x"39",
          4290 => x"8d",
          4291 => x"74",
          4292 => x"0d",
          4293 => x"0d",
          4294 => x"05",
          4295 => x"02",
          4296 => x"05",
          4297 => x"b4",
          4298 => x"29",
          4299 => x"05",
          4300 => x"59",
          4301 => x"59",
          4302 => x"86",
          4303 => x"9a",
          4304 => x"d5",
          4305 => x"84",
          4306 => x"dc",
          4307 => x"70",
          4308 => x"5a",
          4309 => x"82",
          4310 => x"75",
          4311 => x"b4",
          4312 => x"29",
          4313 => x"05",
          4314 => x"56",
          4315 => x"2e",
          4316 => x"53",
          4317 => x"51",
          4318 => x"3f",
          4319 => x"33",
          4320 => x"74",
          4321 => x"34",
          4322 => x"06",
          4323 => x"27",
          4324 => x"0b",
          4325 => x"34",
          4326 => x"b6",
          4327 => x"b0",
          4328 => x"80",
          4329 => x"82",
          4330 => x"55",
          4331 => x"8c",
          4332 => x"54",
          4333 => x"52",
          4334 => x"ec",
          4335 => x"d5",
          4336 => x"8a",
          4337 => x"d4",
          4338 => x"b0",
          4339 => x"ef",
          4340 => x"3d",
          4341 => x"3d",
          4342 => x"dc",
          4343 => x"72",
          4344 => x"80",
          4345 => x"71",
          4346 => x"3f",
          4347 => x"ff",
          4348 => x"54",
          4349 => x"25",
          4350 => x"0b",
          4351 => x"34",
          4352 => x"08",
          4353 => x"2e",
          4354 => x"51",
          4355 => x"3f",
          4356 => x"08",
          4357 => x"3f",
          4358 => x"d5",
          4359 => x"3d",
          4360 => x"3d",
          4361 => x"80",
          4362 => x"b0",
          4363 => x"f5",
          4364 => x"d5",
          4365 => x"d3",
          4366 => x"b0",
          4367 => x"f8",
          4368 => x"70",
          4369 => x"9f",
          4370 => x"d5",
          4371 => x"2e",
          4372 => x"51",
          4373 => x"3f",
          4374 => x"08",
          4375 => x"82",
          4376 => x"25",
          4377 => x"d5",
          4378 => x"05",
          4379 => x"55",
          4380 => x"75",
          4381 => x"81",
          4382 => x"98",
          4383 => x"8a",
          4384 => x"ff",
          4385 => x"06",
          4386 => x"a6",
          4387 => x"d9",
          4388 => x"3d",
          4389 => x"08",
          4390 => x"70",
          4391 => x"52",
          4392 => x"08",
          4393 => x"f0",
          4394 => x"e4",
          4395 => x"38",
          4396 => x"d5",
          4397 => x"55",
          4398 => x"8b",
          4399 => x"56",
          4400 => x"3f",
          4401 => x"08",
          4402 => x"38",
          4403 => x"b2",
          4404 => x"d5",
          4405 => x"18",
          4406 => x"0b",
          4407 => x"08",
          4408 => x"82",
          4409 => x"ff",
          4410 => x"55",
          4411 => x"34",
          4412 => x"30",
          4413 => x"9f",
          4414 => x"55",
          4415 => x"85",
          4416 => x"ac",
          4417 => x"b0",
          4418 => x"08",
          4419 => x"f4",
          4420 => x"d5",
          4421 => x"2e",
          4422 => x"c6",
          4423 => x"89",
          4424 => x"77",
          4425 => x"06",
          4426 => x"52",
          4427 => x"b2",
          4428 => x"51",
          4429 => x"3f",
          4430 => x"54",
          4431 => x"08",
          4432 => x"58",
          4433 => x"e4",
          4434 => x"0d",
          4435 => x"0d",
          4436 => x"5c",
          4437 => x"57",
          4438 => x"73",
          4439 => x"81",
          4440 => x"78",
          4441 => x"56",
          4442 => x"98",
          4443 => x"70",
          4444 => x"33",
          4445 => x"73",
          4446 => x"81",
          4447 => x"75",
          4448 => x"38",
          4449 => x"88",
          4450 => x"b8",
          4451 => x"52",
          4452 => x"f4",
          4453 => x"e4",
          4454 => x"52",
          4455 => x"ff",
          4456 => x"82",
          4457 => x"80",
          4458 => x"15",
          4459 => x"81",
          4460 => x"74",
          4461 => x"38",
          4462 => x"e6",
          4463 => x"81",
          4464 => x"3d",
          4465 => x"f8",
          4466 => x"ae",
          4467 => x"e4",
          4468 => x"9a",
          4469 => x"53",
          4470 => x"51",
          4471 => x"82",
          4472 => x"81",
          4473 => x"74",
          4474 => x"54",
          4475 => x"14",
          4476 => x"06",
          4477 => x"74",
          4478 => x"38",
          4479 => x"82",
          4480 => x"8c",
          4481 => x"d3",
          4482 => x"3d",
          4483 => x"08",
          4484 => x"59",
          4485 => x"0b",
          4486 => x"82",
          4487 => x"82",
          4488 => x"55",
          4489 => x"cb",
          4490 => x"d5",
          4491 => x"55",
          4492 => x"81",
          4493 => x"2e",
          4494 => x"81",
          4495 => x"55",
          4496 => x"2e",
          4497 => x"a8",
          4498 => x"3f",
          4499 => x"08",
          4500 => x"0c",
          4501 => x"08",
          4502 => x"92",
          4503 => x"76",
          4504 => x"e4",
          4505 => x"de",
          4506 => x"d5",
          4507 => x"2e",
          4508 => x"c6",
          4509 => x"a2",
          4510 => x"f7",
          4511 => x"e4",
          4512 => x"d5",
          4513 => x"80",
          4514 => x"3d",
          4515 => x"81",
          4516 => x"82",
          4517 => x"56",
          4518 => x"08",
          4519 => x"81",
          4520 => x"38",
          4521 => x"08",
          4522 => x"dc",
          4523 => x"e4",
          4524 => x"0b",
          4525 => x"08",
          4526 => x"82",
          4527 => x"ff",
          4528 => x"55",
          4529 => x"34",
          4530 => x"81",
          4531 => x"75",
          4532 => x"3f",
          4533 => x"81",
          4534 => x"54",
          4535 => x"83",
          4536 => x"74",
          4537 => x"81",
          4538 => x"38",
          4539 => x"82",
          4540 => x"76",
          4541 => x"d5",
          4542 => x"2e",
          4543 => x"d6",
          4544 => x"5d",
          4545 => x"82",
          4546 => x"98",
          4547 => x"2c",
          4548 => x"ff",
          4549 => x"78",
          4550 => x"82",
          4551 => x"70",
          4552 => x"98",
          4553 => x"9c",
          4554 => x"2b",
          4555 => x"71",
          4556 => x"70",
          4557 => x"c3",
          4558 => x"08",
          4559 => x"51",
          4560 => x"59",
          4561 => x"5d",
          4562 => x"73",
          4563 => x"e9",
          4564 => x"27",
          4565 => x"81",
          4566 => x"81",
          4567 => x"70",
          4568 => x"55",
          4569 => x"80",
          4570 => x"53",
          4571 => x"51",
          4572 => x"82",
          4573 => x"81",
          4574 => x"73",
          4575 => x"38",
          4576 => x"9c",
          4577 => x"b1",
          4578 => x"80",
          4579 => x"80",
          4580 => x"98",
          4581 => x"ff",
          4582 => x"55",
          4583 => x"97",
          4584 => x"74",
          4585 => x"f5",
          4586 => x"d5",
          4587 => x"ff",
          4588 => x"cc",
          4589 => x"80",
          4590 => x"2e",
          4591 => x"81",
          4592 => x"82",
          4593 => x"74",
          4594 => x"98",
          4595 => x"9c",
          4596 => x"2b",
          4597 => x"70",
          4598 => x"82",
          4599 => x"a8",
          4600 => x"51",
          4601 => x"58",
          4602 => x"77",
          4603 => x"06",
          4604 => x"82",
          4605 => x"08",
          4606 => x"0b",
          4607 => x"34",
          4608 => x"ed",
          4609 => x"39",
          4610 => x"a0",
          4611 => x"ed",
          4612 => x"af",
          4613 => x"7d",
          4614 => x"73",
          4615 => x"e1",
          4616 => x"29",
          4617 => x"05",
          4618 => x"04",
          4619 => x"33",
          4620 => x"2e",
          4621 => x"82",
          4622 => x"55",
          4623 => x"ab",
          4624 => x"2b",
          4625 => x"51",
          4626 => x"24",
          4627 => x"1a",
          4628 => x"81",
          4629 => x"81",
          4630 => x"81",
          4631 => x"70",
          4632 => x"ed",
          4633 => x"51",
          4634 => x"82",
          4635 => x"81",
          4636 => x"74",
          4637 => x"34",
          4638 => x"ae",
          4639 => x"34",
          4640 => x"33",
          4641 => x"25",
          4642 => x"14",
          4643 => x"ed",
          4644 => x"ed",
          4645 => x"81",
          4646 => x"81",
          4647 => x"70",
          4648 => x"ed",
          4649 => x"51",
          4650 => x"77",
          4651 => x"82",
          4652 => x"52",
          4653 => x"33",
          4654 => x"a1",
          4655 => x"81",
          4656 => x"81",
          4657 => x"70",
          4658 => x"ed",
          4659 => x"51",
          4660 => x"24",
          4661 => x"ed",
          4662 => x"98",
          4663 => x"2c",
          4664 => x"33",
          4665 => x"56",
          4666 => x"fc",
          4667 => x"f1",
          4668 => x"88",
          4669 => x"bd",
          4670 => x"80",
          4671 => x"80",
          4672 => x"98",
          4673 => x"a4",
          4674 => x"55",
          4675 => x"de",
          4676 => x"39",
          4677 => x"80",
          4678 => x"34",
          4679 => x"53",
          4680 => x"b6",
          4681 => x"9c",
          4682 => x"39",
          4683 => x"33",
          4684 => x"06",
          4685 => x"80",
          4686 => x"38",
          4687 => x"33",
          4688 => x"73",
          4689 => x"34",
          4690 => x"73",
          4691 => x"34",
          4692 => x"08",
          4693 => x"ff",
          4694 => x"82",
          4695 => x"70",
          4696 => x"98",
          4697 => x"a4",
          4698 => x"56",
          4699 => x"25",
          4700 => x"1a",
          4701 => x"33",
          4702 => x"f1",
          4703 => x"73",
          4704 => x"a0",
          4705 => x"81",
          4706 => x"81",
          4707 => x"70",
          4708 => x"ed",
          4709 => x"51",
          4710 => x"24",
          4711 => x"f1",
          4712 => x"a0",
          4713 => x"8d",
          4714 => x"a8",
          4715 => x"2b",
          4716 => x"82",
          4717 => x"57",
          4718 => x"74",
          4719 => x"c1",
          4720 => x"c8",
          4721 => x"51",
          4722 => x"3f",
          4723 => x"0a",
          4724 => x"0a",
          4725 => x"2c",
          4726 => x"33",
          4727 => x"75",
          4728 => x"38",
          4729 => x"82",
          4730 => x"7a",
          4731 => x"74",
          4732 => x"c8",
          4733 => x"51",
          4734 => x"3f",
          4735 => x"52",
          4736 => x"c9",
          4737 => x"e4",
          4738 => x"06",
          4739 => x"38",
          4740 => x"33",
          4741 => x"2e",
          4742 => x"53",
          4743 => x"51",
          4744 => x"84",
          4745 => x"34",
          4746 => x"ed",
          4747 => x"0b",
          4748 => x"34",
          4749 => x"e4",
          4750 => x"0d",
          4751 => x"a8",
          4752 => x"80",
          4753 => x"38",
          4754 => x"08",
          4755 => x"ff",
          4756 => x"82",
          4757 => x"ff",
          4758 => x"82",
          4759 => x"73",
          4760 => x"54",
          4761 => x"ed",
          4762 => x"ed",
          4763 => x"55",
          4764 => x"f9",
          4765 => x"14",
          4766 => x"ed",
          4767 => x"98",
          4768 => x"2c",
          4769 => x"06",
          4770 => x"74",
          4771 => x"38",
          4772 => x"81",
          4773 => x"34",
          4774 => x"08",
          4775 => x"51",
          4776 => x"3f",
          4777 => x"0a",
          4778 => x"0a",
          4779 => x"2c",
          4780 => x"33",
          4781 => x"75",
          4782 => x"38",
          4783 => x"08",
          4784 => x"ff",
          4785 => x"82",
          4786 => x"70",
          4787 => x"98",
          4788 => x"a4",
          4789 => x"56",
          4790 => x"24",
          4791 => x"82",
          4792 => x"52",
          4793 => x"9d",
          4794 => x"81",
          4795 => x"81",
          4796 => x"70",
          4797 => x"ed",
          4798 => x"51",
          4799 => x"25",
          4800 => x"fd",
          4801 => x"a8",
          4802 => x"ff",
          4803 => x"a4",
          4804 => x"54",
          4805 => x"f7",
          4806 => x"f1",
          4807 => x"81",
          4808 => x"82",
          4809 => x"74",
          4810 => x"52",
          4811 => x"85",
          4812 => x"a8",
          4813 => x"ff",
          4814 => x"a4",
          4815 => x"54",
          4816 => x"d6",
          4817 => x"39",
          4818 => x"53",
          4819 => x"b6",
          4820 => x"f0",
          4821 => x"82",
          4822 => x"80",
          4823 => x"a4",
          4824 => x"39",
          4825 => x"82",
          4826 => x"55",
          4827 => x"a6",
          4828 => x"ff",
          4829 => x"82",
          4830 => x"82",
          4831 => x"82",
          4832 => x"81",
          4833 => x"05",
          4834 => x"79",
          4835 => x"d8",
          4836 => x"81",
          4837 => x"84",
          4838 => x"dc",
          4839 => x"08",
          4840 => x"80",
          4841 => x"74",
          4842 => x"dc",
          4843 => x"e4",
          4844 => x"a4",
          4845 => x"e4",
          4846 => x"06",
          4847 => x"74",
          4848 => x"ff",
          4849 => x"ff",
          4850 => x"fa",
          4851 => x"55",
          4852 => x"f6",
          4853 => x"51",
          4854 => x"3f",
          4855 => x"93",
          4856 => x"06",
          4857 => x"d4",
          4858 => x"74",
          4859 => x"38",
          4860 => x"a4",
          4861 => x"d5",
          4862 => x"ed",
          4863 => x"d5",
          4864 => x"ff",
          4865 => x"53",
          4866 => x"51",
          4867 => x"3f",
          4868 => x"7a",
          4869 => x"d4",
          4870 => x"08",
          4871 => x"80",
          4872 => x"74",
          4873 => x"e0",
          4874 => x"e4",
          4875 => x"a4",
          4876 => x"e4",
          4877 => x"06",
          4878 => x"74",
          4879 => x"ff",
          4880 => x"81",
          4881 => x"81",
          4882 => x"89",
          4883 => x"ed",
          4884 => x"7a",
          4885 => x"a8",
          4886 => x"a4",
          4887 => x"51",
          4888 => x"f5",
          4889 => x"ed",
          4890 => x"81",
          4891 => x"ed",
          4892 => x"56",
          4893 => x"27",
          4894 => x"82",
          4895 => x"52",
          4896 => x"73",
          4897 => x"34",
          4898 => x"33",
          4899 => x"9a",
          4900 => x"ed",
          4901 => x"a8",
          4902 => x"80",
          4903 => x"38",
          4904 => x"08",
          4905 => x"ff",
          4906 => x"82",
          4907 => x"ff",
          4908 => x"82",
          4909 => x"f4",
          4910 => x"3d",
          4911 => x"f4",
          4912 => x"d4",
          4913 => x"0b",
          4914 => x"23",
          4915 => x"53",
          4916 => x"fa",
          4917 => x"aa",
          4918 => x"d5",
          4919 => x"80",
          4920 => x"34",
          4921 => x"81",
          4922 => x"d5",
          4923 => x"77",
          4924 => x"76",
          4925 => x"82",
          4926 => x"54",
          4927 => x"34",
          4928 => x"34",
          4929 => x"08",
          4930 => x"22",
          4931 => x"80",
          4932 => x"83",
          4933 => x"70",
          4934 => x"51",
          4935 => x"88",
          4936 => x"89",
          4937 => x"d5",
          4938 => x"88",
          4939 => x"d4",
          4940 => x"11",
          4941 => x"77",
          4942 => x"76",
          4943 => x"89",
          4944 => x"ff",
          4945 => x"52",
          4946 => x"72",
          4947 => x"fb",
          4948 => x"82",
          4949 => x"ff",
          4950 => x"51",
          4951 => x"d5",
          4952 => x"3d",
          4953 => x"3d",
          4954 => x"05",
          4955 => x"05",
          4956 => x"71",
          4957 => x"d4",
          4958 => x"2b",
          4959 => x"83",
          4960 => x"70",
          4961 => x"33",
          4962 => x"07",
          4963 => x"ae",
          4964 => x"81",
          4965 => x"07",
          4966 => x"53",
          4967 => x"54",
          4968 => x"53",
          4969 => x"77",
          4970 => x"18",
          4971 => x"d4",
          4972 => x"88",
          4973 => x"70",
          4974 => x"74",
          4975 => x"82",
          4976 => x"70",
          4977 => x"81",
          4978 => x"88",
          4979 => x"83",
          4980 => x"f8",
          4981 => x"56",
          4982 => x"73",
          4983 => x"06",
          4984 => x"54",
          4985 => x"82",
          4986 => x"81",
          4987 => x"72",
          4988 => x"82",
          4989 => x"16",
          4990 => x"34",
          4991 => x"34",
          4992 => x"04",
          4993 => x"82",
          4994 => x"02",
          4995 => x"05",
          4996 => x"2b",
          4997 => x"11",
          4998 => x"33",
          4999 => x"71",
          5000 => x"58",
          5001 => x"55",
          5002 => x"84",
          5003 => x"13",
          5004 => x"2b",
          5005 => x"2a",
          5006 => x"52",
          5007 => x"34",
          5008 => x"34",
          5009 => x"08",
          5010 => x"11",
          5011 => x"33",
          5012 => x"71",
          5013 => x"56",
          5014 => x"72",
          5015 => x"33",
          5016 => x"71",
          5017 => x"70",
          5018 => x"56",
          5019 => x"86",
          5020 => x"87",
          5021 => x"d5",
          5022 => x"70",
          5023 => x"33",
          5024 => x"07",
          5025 => x"ff",
          5026 => x"2a",
          5027 => x"53",
          5028 => x"34",
          5029 => x"34",
          5030 => x"04",
          5031 => x"02",
          5032 => x"82",
          5033 => x"71",
          5034 => x"11",
          5035 => x"12",
          5036 => x"2b",
          5037 => x"29",
          5038 => x"81",
          5039 => x"98",
          5040 => x"2b",
          5041 => x"53",
          5042 => x"56",
          5043 => x"71",
          5044 => x"f6",
          5045 => x"fe",
          5046 => x"d5",
          5047 => x"16",
          5048 => x"12",
          5049 => x"2b",
          5050 => x"07",
          5051 => x"33",
          5052 => x"71",
          5053 => x"70",
          5054 => x"ff",
          5055 => x"52",
          5056 => x"5a",
          5057 => x"05",
          5058 => x"54",
          5059 => x"13",
          5060 => x"13",
          5061 => x"d4",
          5062 => x"70",
          5063 => x"33",
          5064 => x"71",
          5065 => x"56",
          5066 => x"72",
          5067 => x"81",
          5068 => x"88",
          5069 => x"81",
          5070 => x"70",
          5071 => x"51",
          5072 => x"72",
          5073 => x"81",
          5074 => x"3d",
          5075 => x"3d",
          5076 => x"d4",
          5077 => x"05",
          5078 => x"70",
          5079 => x"11",
          5080 => x"83",
          5081 => x"8b",
          5082 => x"2b",
          5083 => x"59",
          5084 => x"73",
          5085 => x"81",
          5086 => x"88",
          5087 => x"8c",
          5088 => x"22",
          5089 => x"88",
          5090 => x"53",
          5091 => x"73",
          5092 => x"14",
          5093 => x"d4",
          5094 => x"70",
          5095 => x"33",
          5096 => x"71",
          5097 => x"56",
          5098 => x"72",
          5099 => x"33",
          5100 => x"71",
          5101 => x"70",
          5102 => x"55",
          5103 => x"82",
          5104 => x"83",
          5105 => x"d5",
          5106 => x"82",
          5107 => x"12",
          5108 => x"2b",
          5109 => x"e4",
          5110 => x"87",
          5111 => x"f7",
          5112 => x"82",
          5113 => x"31",
          5114 => x"83",
          5115 => x"70",
          5116 => x"fd",
          5117 => x"d5",
          5118 => x"83",
          5119 => x"82",
          5120 => x"12",
          5121 => x"2b",
          5122 => x"07",
          5123 => x"33",
          5124 => x"71",
          5125 => x"90",
          5126 => x"42",
          5127 => x"5b",
          5128 => x"54",
          5129 => x"8d",
          5130 => x"80",
          5131 => x"fe",
          5132 => x"84",
          5133 => x"33",
          5134 => x"71",
          5135 => x"83",
          5136 => x"11",
          5137 => x"53",
          5138 => x"55",
          5139 => x"34",
          5140 => x"06",
          5141 => x"14",
          5142 => x"d4",
          5143 => x"84",
          5144 => x"13",
          5145 => x"2b",
          5146 => x"2a",
          5147 => x"56",
          5148 => x"16",
          5149 => x"16",
          5150 => x"d4",
          5151 => x"80",
          5152 => x"34",
          5153 => x"14",
          5154 => x"d4",
          5155 => x"84",
          5156 => x"85",
          5157 => x"d5",
          5158 => x"70",
          5159 => x"33",
          5160 => x"07",
          5161 => x"80",
          5162 => x"2a",
          5163 => x"56",
          5164 => x"34",
          5165 => x"34",
          5166 => x"04",
          5167 => x"73",
          5168 => x"d4",
          5169 => x"f7",
          5170 => x"80",
          5171 => x"71",
          5172 => x"3f",
          5173 => x"04",
          5174 => x"80",
          5175 => x"f8",
          5176 => x"d5",
          5177 => x"ff",
          5178 => x"d5",
          5179 => x"11",
          5180 => x"33",
          5181 => x"07",
          5182 => x"56",
          5183 => x"ff",
          5184 => x"78",
          5185 => x"38",
          5186 => x"17",
          5187 => x"12",
          5188 => x"2b",
          5189 => x"ff",
          5190 => x"31",
          5191 => x"ff",
          5192 => x"27",
          5193 => x"56",
          5194 => x"79",
          5195 => x"73",
          5196 => x"38",
          5197 => x"5b",
          5198 => x"85",
          5199 => x"88",
          5200 => x"54",
          5201 => x"78",
          5202 => x"2e",
          5203 => x"79",
          5204 => x"76",
          5205 => x"d5",
          5206 => x"70",
          5207 => x"33",
          5208 => x"07",
          5209 => x"ff",
          5210 => x"5a",
          5211 => x"73",
          5212 => x"38",
          5213 => x"54",
          5214 => x"81",
          5215 => x"54",
          5216 => x"81",
          5217 => x"7a",
          5218 => x"06",
          5219 => x"51",
          5220 => x"81",
          5221 => x"80",
          5222 => x"52",
          5223 => x"c6",
          5224 => x"d4",
          5225 => x"86",
          5226 => x"12",
          5227 => x"2b",
          5228 => x"07",
          5229 => x"55",
          5230 => x"17",
          5231 => x"ff",
          5232 => x"2a",
          5233 => x"54",
          5234 => x"34",
          5235 => x"06",
          5236 => x"15",
          5237 => x"d4",
          5238 => x"2b",
          5239 => x"1e",
          5240 => x"87",
          5241 => x"88",
          5242 => x"88",
          5243 => x"5e",
          5244 => x"54",
          5245 => x"34",
          5246 => x"34",
          5247 => x"08",
          5248 => x"11",
          5249 => x"33",
          5250 => x"71",
          5251 => x"53",
          5252 => x"74",
          5253 => x"86",
          5254 => x"87",
          5255 => x"d5",
          5256 => x"16",
          5257 => x"11",
          5258 => x"33",
          5259 => x"07",
          5260 => x"53",
          5261 => x"56",
          5262 => x"16",
          5263 => x"16",
          5264 => x"d4",
          5265 => x"05",
          5266 => x"d5",
          5267 => x"3d",
          5268 => x"3d",
          5269 => x"82",
          5270 => x"84",
          5271 => x"3f",
          5272 => x"80",
          5273 => x"71",
          5274 => x"3f",
          5275 => x"08",
          5276 => x"d5",
          5277 => x"3d",
          5278 => x"3d",
          5279 => x"40",
          5280 => x"42",
          5281 => x"d4",
          5282 => x"09",
          5283 => x"38",
          5284 => x"7b",
          5285 => x"51",
          5286 => x"82",
          5287 => x"54",
          5288 => x"7e",
          5289 => x"51",
          5290 => x"7e",
          5291 => x"39",
          5292 => x"8f",
          5293 => x"e4",
          5294 => x"ff",
          5295 => x"d4",
          5296 => x"31",
          5297 => x"83",
          5298 => x"70",
          5299 => x"11",
          5300 => x"12",
          5301 => x"2b",
          5302 => x"31",
          5303 => x"ff",
          5304 => x"29",
          5305 => x"88",
          5306 => x"33",
          5307 => x"71",
          5308 => x"70",
          5309 => x"44",
          5310 => x"41",
          5311 => x"5b",
          5312 => x"5b",
          5313 => x"25",
          5314 => x"81",
          5315 => x"75",
          5316 => x"ff",
          5317 => x"54",
          5318 => x"83",
          5319 => x"88",
          5320 => x"88",
          5321 => x"33",
          5322 => x"71",
          5323 => x"90",
          5324 => x"47",
          5325 => x"54",
          5326 => x"8b",
          5327 => x"31",
          5328 => x"ff",
          5329 => x"77",
          5330 => x"fe",
          5331 => x"54",
          5332 => x"09",
          5333 => x"38",
          5334 => x"c0",
          5335 => x"ff",
          5336 => x"81",
          5337 => x"8e",
          5338 => x"24",
          5339 => x"51",
          5340 => x"81",
          5341 => x"18",
          5342 => x"24",
          5343 => x"79",
          5344 => x"33",
          5345 => x"71",
          5346 => x"53",
          5347 => x"f4",
          5348 => x"78",
          5349 => x"3f",
          5350 => x"08",
          5351 => x"06",
          5352 => x"53",
          5353 => x"82",
          5354 => x"11",
          5355 => x"55",
          5356 => x"ea",
          5357 => x"d4",
          5358 => x"05",
          5359 => x"ff",
          5360 => x"81",
          5361 => x"15",
          5362 => x"24",
          5363 => x"78",
          5364 => x"3f",
          5365 => x"08",
          5366 => x"33",
          5367 => x"71",
          5368 => x"53",
          5369 => x"9c",
          5370 => x"78",
          5371 => x"3f",
          5372 => x"08",
          5373 => x"06",
          5374 => x"53",
          5375 => x"82",
          5376 => x"11",
          5377 => x"55",
          5378 => x"92",
          5379 => x"d4",
          5380 => x"05",
          5381 => x"19",
          5382 => x"83",
          5383 => x"58",
          5384 => x"7f",
          5385 => x"b0",
          5386 => x"e4",
          5387 => x"d5",
          5388 => x"2e",
          5389 => x"53",
          5390 => x"d5",
          5391 => x"ff",
          5392 => x"73",
          5393 => x"3f",
          5394 => x"78",
          5395 => x"80",
          5396 => x"78",
          5397 => x"3f",
          5398 => x"2b",
          5399 => x"08",
          5400 => x"51",
          5401 => x"7b",
          5402 => x"d5",
          5403 => x"3d",
          5404 => x"3d",
          5405 => x"29",
          5406 => x"fb",
          5407 => x"d5",
          5408 => x"82",
          5409 => x"80",
          5410 => x"73",
          5411 => x"82",
          5412 => x"51",
          5413 => x"3f",
          5414 => x"e4",
          5415 => x"0d",
          5416 => x"0d",
          5417 => x"33",
          5418 => x"70",
          5419 => x"38",
          5420 => x"11",
          5421 => x"82",
          5422 => x"83",
          5423 => x"fc",
          5424 => x"9b",
          5425 => x"84",
          5426 => x"33",
          5427 => x"51",
          5428 => x"80",
          5429 => x"84",
          5430 => x"92",
          5431 => x"51",
          5432 => x"80",
          5433 => x"81",
          5434 => x"72",
          5435 => x"92",
          5436 => x"81",
          5437 => x"0b",
          5438 => x"8c",
          5439 => x"71",
          5440 => x"06",
          5441 => x"80",
          5442 => x"87",
          5443 => x"08",
          5444 => x"38",
          5445 => x"80",
          5446 => x"71",
          5447 => x"c0",
          5448 => x"51",
          5449 => x"87",
          5450 => x"d5",
          5451 => x"82",
          5452 => x"33",
          5453 => x"d5",
          5454 => x"3d",
          5455 => x"3d",
          5456 => x"64",
          5457 => x"bf",
          5458 => x"40",
          5459 => x"74",
          5460 => x"cd",
          5461 => x"e4",
          5462 => x"7a",
          5463 => x"81",
          5464 => x"72",
          5465 => x"87",
          5466 => x"11",
          5467 => x"8c",
          5468 => x"92",
          5469 => x"5a",
          5470 => x"58",
          5471 => x"c0",
          5472 => x"76",
          5473 => x"76",
          5474 => x"70",
          5475 => x"81",
          5476 => x"54",
          5477 => x"8e",
          5478 => x"52",
          5479 => x"81",
          5480 => x"81",
          5481 => x"74",
          5482 => x"53",
          5483 => x"83",
          5484 => x"78",
          5485 => x"8f",
          5486 => x"2e",
          5487 => x"c0",
          5488 => x"52",
          5489 => x"87",
          5490 => x"08",
          5491 => x"2e",
          5492 => x"84",
          5493 => x"38",
          5494 => x"87",
          5495 => x"15",
          5496 => x"70",
          5497 => x"52",
          5498 => x"ff",
          5499 => x"39",
          5500 => x"81",
          5501 => x"ff",
          5502 => x"57",
          5503 => x"90",
          5504 => x"80",
          5505 => x"71",
          5506 => x"78",
          5507 => x"38",
          5508 => x"80",
          5509 => x"80",
          5510 => x"81",
          5511 => x"72",
          5512 => x"0c",
          5513 => x"04",
          5514 => x"60",
          5515 => x"8c",
          5516 => x"33",
          5517 => x"5b",
          5518 => x"74",
          5519 => x"e1",
          5520 => x"e4",
          5521 => x"79",
          5522 => x"78",
          5523 => x"06",
          5524 => x"77",
          5525 => x"87",
          5526 => x"11",
          5527 => x"8c",
          5528 => x"92",
          5529 => x"59",
          5530 => x"85",
          5531 => x"98",
          5532 => x"7d",
          5533 => x"0c",
          5534 => x"08",
          5535 => x"70",
          5536 => x"53",
          5537 => x"2e",
          5538 => x"70",
          5539 => x"33",
          5540 => x"18",
          5541 => x"2a",
          5542 => x"51",
          5543 => x"2e",
          5544 => x"c0",
          5545 => x"52",
          5546 => x"87",
          5547 => x"08",
          5548 => x"2e",
          5549 => x"84",
          5550 => x"38",
          5551 => x"87",
          5552 => x"15",
          5553 => x"70",
          5554 => x"52",
          5555 => x"ff",
          5556 => x"39",
          5557 => x"81",
          5558 => x"80",
          5559 => x"52",
          5560 => x"90",
          5561 => x"80",
          5562 => x"71",
          5563 => x"7a",
          5564 => x"38",
          5565 => x"80",
          5566 => x"80",
          5567 => x"81",
          5568 => x"72",
          5569 => x"0c",
          5570 => x"04",
          5571 => x"7a",
          5572 => x"a3",
          5573 => x"88",
          5574 => x"33",
          5575 => x"56",
          5576 => x"3f",
          5577 => x"08",
          5578 => x"83",
          5579 => x"fe",
          5580 => x"87",
          5581 => x"0c",
          5582 => x"76",
          5583 => x"38",
          5584 => x"93",
          5585 => x"2b",
          5586 => x"8c",
          5587 => x"71",
          5588 => x"38",
          5589 => x"71",
          5590 => x"c6",
          5591 => x"39",
          5592 => x"81",
          5593 => x"06",
          5594 => x"71",
          5595 => x"38",
          5596 => x"8c",
          5597 => x"e8",
          5598 => x"98",
          5599 => x"71",
          5600 => x"73",
          5601 => x"92",
          5602 => x"72",
          5603 => x"06",
          5604 => x"f7",
          5605 => x"80",
          5606 => x"88",
          5607 => x"0c",
          5608 => x"80",
          5609 => x"56",
          5610 => x"56",
          5611 => x"82",
          5612 => x"88",
          5613 => x"fe",
          5614 => x"81",
          5615 => x"33",
          5616 => x"07",
          5617 => x"0c",
          5618 => x"3d",
          5619 => x"3d",
          5620 => x"11",
          5621 => x"33",
          5622 => x"71",
          5623 => x"81",
          5624 => x"72",
          5625 => x"75",
          5626 => x"82",
          5627 => x"52",
          5628 => x"54",
          5629 => x"0d",
          5630 => x"0d",
          5631 => x"05",
          5632 => x"52",
          5633 => x"70",
          5634 => x"34",
          5635 => x"51",
          5636 => x"83",
          5637 => x"ff",
          5638 => x"75",
          5639 => x"72",
          5640 => x"54",
          5641 => x"2a",
          5642 => x"70",
          5643 => x"34",
          5644 => x"51",
          5645 => x"81",
          5646 => x"70",
          5647 => x"70",
          5648 => x"3d",
          5649 => x"3d",
          5650 => x"77",
          5651 => x"70",
          5652 => x"38",
          5653 => x"05",
          5654 => x"70",
          5655 => x"34",
          5656 => x"eb",
          5657 => x"0d",
          5658 => x"0d",
          5659 => x"54",
          5660 => x"72",
          5661 => x"54",
          5662 => x"51",
          5663 => x"84",
          5664 => x"fc",
          5665 => x"77",
          5666 => x"53",
          5667 => x"05",
          5668 => x"70",
          5669 => x"33",
          5670 => x"ff",
          5671 => x"52",
          5672 => x"2e",
          5673 => x"80",
          5674 => x"71",
          5675 => x"0c",
          5676 => x"04",
          5677 => x"74",
          5678 => x"89",
          5679 => x"2e",
          5680 => x"11",
          5681 => x"52",
          5682 => x"70",
          5683 => x"e4",
          5684 => x"0d",
          5685 => x"82",
          5686 => x"04",
          5687 => x"77",
          5688 => x"70",
          5689 => x"33",
          5690 => x"55",
          5691 => x"ff",
          5692 => x"e4",
          5693 => x"72",
          5694 => x"38",
          5695 => x"72",
          5696 => x"a2",
          5697 => x"e4",
          5698 => x"ff",
          5699 => x"80",
          5700 => x"73",
          5701 => x"55",
          5702 => x"e4",
          5703 => x"0d",
          5704 => x"0d",
          5705 => x"0b",
          5706 => x"56",
          5707 => x"2e",
          5708 => x"81",
          5709 => x"08",
          5710 => x"70",
          5711 => x"33",
          5712 => x"e4",
          5713 => x"e4",
          5714 => x"09",
          5715 => x"38",
          5716 => x"08",
          5717 => x"b4",
          5718 => x"a8",
          5719 => x"a0",
          5720 => x"56",
          5721 => x"27",
          5722 => x"16",
          5723 => x"82",
          5724 => x"06",
          5725 => x"54",
          5726 => x"78",
          5727 => x"33",
          5728 => x"3f",
          5729 => x"5a",
          5730 => x"e4",
          5731 => x"0d",
          5732 => x"0d",
          5733 => x"56",
          5734 => x"b4",
          5735 => x"af",
          5736 => x"fe",
          5737 => x"d5",
          5738 => x"82",
          5739 => x"9f",
          5740 => x"74",
          5741 => x"52",
          5742 => x"51",
          5743 => x"82",
          5744 => x"80",
          5745 => x"ff",
          5746 => x"74",
          5747 => x"76",
          5748 => x"0c",
          5749 => x"04",
          5750 => x"7a",
          5751 => x"fe",
          5752 => x"d5",
          5753 => x"82",
          5754 => x"81",
          5755 => x"33",
          5756 => x"2e",
          5757 => x"80",
          5758 => x"17",
          5759 => x"81",
          5760 => x"06",
          5761 => x"84",
          5762 => x"d5",
          5763 => x"b8",
          5764 => x"56",
          5765 => x"82",
          5766 => x"84",
          5767 => x"fb",
          5768 => x"8b",
          5769 => x"52",
          5770 => x"eb",
          5771 => x"85",
          5772 => x"84",
          5773 => x"fb",
          5774 => x"17",
          5775 => x"a0",
          5776 => x"d3",
          5777 => x"08",
          5778 => x"17",
          5779 => x"3f",
          5780 => x"81",
          5781 => x"19",
          5782 => x"53",
          5783 => x"17",
          5784 => x"c4",
          5785 => x"18",
          5786 => x"80",
          5787 => x"33",
          5788 => x"3f",
          5789 => x"08",
          5790 => x"38",
          5791 => x"82",
          5792 => x"8a",
          5793 => x"fb",
          5794 => x"fe",
          5795 => x"08",
          5796 => x"56",
          5797 => x"74",
          5798 => x"38",
          5799 => x"75",
          5800 => x"16",
          5801 => x"53",
          5802 => x"e4",
          5803 => x"0d",
          5804 => x"0d",
          5805 => x"08",
          5806 => x"81",
          5807 => x"df",
          5808 => x"15",
          5809 => x"d7",
          5810 => x"33",
          5811 => x"82",
          5812 => x"38",
          5813 => x"89",
          5814 => x"2e",
          5815 => x"bf",
          5816 => x"2e",
          5817 => x"81",
          5818 => x"81",
          5819 => x"89",
          5820 => x"08",
          5821 => x"52",
          5822 => x"3f",
          5823 => x"08",
          5824 => x"74",
          5825 => x"14",
          5826 => x"81",
          5827 => x"2a",
          5828 => x"05",
          5829 => x"57",
          5830 => x"f5",
          5831 => x"e4",
          5832 => x"38",
          5833 => x"06",
          5834 => x"33",
          5835 => x"78",
          5836 => x"06",
          5837 => x"5c",
          5838 => x"53",
          5839 => x"38",
          5840 => x"06",
          5841 => x"39",
          5842 => x"a8",
          5843 => x"52",
          5844 => x"bd",
          5845 => x"e4",
          5846 => x"38",
          5847 => x"fe",
          5848 => x"b8",
          5849 => x"cf",
          5850 => x"e4",
          5851 => x"ff",
          5852 => x"39",
          5853 => x"a8",
          5854 => x"52",
          5855 => x"91",
          5856 => x"e4",
          5857 => x"76",
          5858 => x"fc",
          5859 => x"b8",
          5860 => x"ba",
          5861 => x"e4",
          5862 => x"06",
          5863 => x"81",
          5864 => x"d5",
          5865 => x"3d",
          5866 => x"3d",
          5867 => x"7e",
          5868 => x"82",
          5869 => x"27",
          5870 => x"76",
          5871 => x"27",
          5872 => x"75",
          5873 => x"79",
          5874 => x"38",
          5875 => x"89",
          5876 => x"2e",
          5877 => x"80",
          5878 => x"2e",
          5879 => x"81",
          5880 => x"81",
          5881 => x"89",
          5882 => x"08",
          5883 => x"52",
          5884 => x"3f",
          5885 => x"08",
          5886 => x"e4",
          5887 => x"38",
          5888 => x"06",
          5889 => x"81",
          5890 => x"06",
          5891 => x"77",
          5892 => x"2e",
          5893 => x"84",
          5894 => x"06",
          5895 => x"06",
          5896 => x"53",
          5897 => x"81",
          5898 => x"34",
          5899 => x"a8",
          5900 => x"52",
          5901 => x"d9",
          5902 => x"e4",
          5903 => x"d5",
          5904 => x"94",
          5905 => x"ff",
          5906 => x"05",
          5907 => x"54",
          5908 => x"38",
          5909 => x"74",
          5910 => x"06",
          5911 => x"07",
          5912 => x"74",
          5913 => x"39",
          5914 => x"a8",
          5915 => x"52",
          5916 => x"9d",
          5917 => x"e4",
          5918 => x"d5",
          5919 => x"d8",
          5920 => x"ff",
          5921 => x"76",
          5922 => x"06",
          5923 => x"05",
          5924 => x"3f",
          5925 => x"87",
          5926 => x"08",
          5927 => x"51",
          5928 => x"82",
          5929 => x"59",
          5930 => x"08",
          5931 => x"f0",
          5932 => x"82",
          5933 => x"06",
          5934 => x"05",
          5935 => x"54",
          5936 => x"3f",
          5937 => x"08",
          5938 => x"74",
          5939 => x"51",
          5940 => x"81",
          5941 => x"34",
          5942 => x"e4",
          5943 => x"0d",
          5944 => x"0d",
          5945 => x"72",
          5946 => x"56",
          5947 => x"27",
          5948 => x"9c",
          5949 => x"9d",
          5950 => x"2e",
          5951 => x"53",
          5952 => x"51",
          5953 => x"82",
          5954 => x"54",
          5955 => x"08",
          5956 => x"93",
          5957 => x"80",
          5958 => x"54",
          5959 => x"82",
          5960 => x"54",
          5961 => x"74",
          5962 => x"fb",
          5963 => x"d5",
          5964 => x"82",
          5965 => x"80",
          5966 => x"38",
          5967 => x"08",
          5968 => x"38",
          5969 => x"08",
          5970 => x"38",
          5971 => x"52",
          5972 => x"d6",
          5973 => x"e4",
          5974 => x"9c",
          5975 => x"11",
          5976 => x"57",
          5977 => x"74",
          5978 => x"81",
          5979 => x"0c",
          5980 => x"81",
          5981 => x"84",
          5982 => x"55",
          5983 => x"ff",
          5984 => x"54",
          5985 => x"e4",
          5986 => x"0d",
          5987 => x"0d",
          5988 => x"08",
          5989 => x"79",
          5990 => x"17",
          5991 => x"80",
          5992 => x"9c",
          5993 => x"26",
          5994 => x"58",
          5995 => x"52",
          5996 => x"fd",
          5997 => x"74",
          5998 => x"08",
          5999 => x"38",
          6000 => x"08",
          6001 => x"e4",
          6002 => x"82",
          6003 => x"17",
          6004 => x"e4",
          6005 => x"c7",
          6006 => x"94",
          6007 => x"56",
          6008 => x"2e",
          6009 => x"77",
          6010 => x"81",
          6011 => x"38",
          6012 => x"9c",
          6013 => x"26",
          6014 => x"56",
          6015 => x"51",
          6016 => x"80",
          6017 => x"e4",
          6018 => x"09",
          6019 => x"38",
          6020 => x"08",
          6021 => x"e4",
          6022 => x"30",
          6023 => x"80",
          6024 => x"07",
          6025 => x"08",
          6026 => x"55",
          6027 => x"ef",
          6028 => x"e4",
          6029 => x"95",
          6030 => x"08",
          6031 => x"27",
          6032 => x"9c",
          6033 => x"89",
          6034 => x"85",
          6035 => x"db",
          6036 => x"81",
          6037 => x"17",
          6038 => x"89",
          6039 => x"75",
          6040 => x"ac",
          6041 => x"7a",
          6042 => x"3f",
          6043 => x"08",
          6044 => x"38",
          6045 => x"d5",
          6046 => x"2e",
          6047 => x"86",
          6048 => x"e4",
          6049 => x"d5",
          6050 => x"70",
          6051 => x"07",
          6052 => x"7c",
          6053 => x"55",
          6054 => x"f8",
          6055 => x"2e",
          6056 => x"ff",
          6057 => x"55",
          6058 => x"ff",
          6059 => x"76",
          6060 => x"3f",
          6061 => x"08",
          6062 => x"08",
          6063 => x"d5",
          6064 => x"80",
          6065 => x"55",
          6066 => x"94",
          6067 => x"2e",
          6068 => x"53",
          6069 => x"51",
          6070 => x"82",
          6071 => x"55",
          6072 => x"75",
          6073 => x"9c",
          6074 => x"05",
          6075 => x"56",
          6076 => x"26",
          6077 => x"15",
          6078 => x"84",
          6079 => x"07",
          6080 => x"18",
          6081 => x"ff",
          6082 => x"2e",
          6083 => x"39",
          6084 => x"39",
          6085 => x"08",
          6086 => x"81",
          6087 => x"74",
          6088 => x"0c",
          6089 => x"04",
          6090 => x"7a",
          6091 => x"f3",
          6092 => x"d5",
          6093 => x"81",
          6094 => x"e4",
          6095 => x"38",
          6096 => x"51",
          6097 => x"82",
          6098 => x"82",
          6099 => x"b4",
          6100 => x"84",
          6101 => x"52",
          6102 => x"52",
          6103 => x"3f",
          6104 => x"39",
          6105 => x"8a",
          6106 => x"75",
          6107 => x"38",
          6108 => x"19",
          6109 => x"81",
          6110 => x"ed",
          6111 => x"d5",
          6112 => x"2e",
          6113 => x"15",
          6114 => x"70",
          6115 => x"07",
          6116 => x"53",
          6117 => x"75",
          6118 => x"0c",
          6119 => x"04",
          6120 => x"7a",
          6121 => x"58",
          6122 => x"f0",
          6123 => x"80",
          6124 => x"9f",
          6125 => x"80",
          6126 => x"90",
          6127 => x"17",
          6128 => x"aa",
          6129 => x"53",
          6130 => x"88",
          6131 => x"08",
          6132 => x"38",
          6133 => x"53",
          6134 => x"17",
          6135 => x"72",
          6136 => x"fe",
          6137 => x"08",
          6138 => x"80",
          6139 => x"16",
          6140 => x"2b",
          6141 => x"75",
          6142 => x"73",
          6143 => x"f5",
          6144 => x"d5",
          6145 => x"82",
          6146 => x"ff",
          6147 => x"81",
          6148 => x"e4",
          6149 => x"38",
          6150 => x"82",
          6151 => x"26",
          6152 => x"58",
          6153 => x"73",
          6154 => x"39",
          6155 => x"51",
          6156 => x"82",
          6157 => x"98",
          6158 => x"94",
          6159 => x"17",
          6160 => x"58",
          6161 => x"9a",
          6162 => x"81",
          6163 => x"74",
          6164 => x"98",
          6165 => x"83",
          6166 => x"b8",
          6167 => x"0c",
          6168 => x"82",
          6169 => x"8a",
          6170 => x"f8",
          6171 => x"70",
          6172 => x"08",
          6173 => x"57",
          6174 => x"0a",
          6175 => x"38",
          6176 => x"15",
          6177 => x"08",
          6178 => x"72",
          6179 => x"cb",
          6180 => x"ff",
          6181 => x"81",
          6182 => x"13",
          6183 => x"94",
          6184 => x"74",
          6185 => x"85",
          6186 => x"22",
          6187 => x"73",
          6188 => x"38",
          6189 => x"8a",
          6190 => x"05",
          6191 => x"06",
          6192 => x"8a",
          6193 => x"73",
          6194 => x"3f",
          6195 => x"08",
          6196 => x"81",
          6197 => x"e4",
          6198 => x"ff",
          6199 => x"82",
          6200 => x"ff",
          6201 => x"38",
          6202 => x"82",
          6203 => x"26",
          6204 => x"7b",
          6205 => x"98",
          6206 => x"55",
          6207 => x"94",
          6208 => x"73",
          6209 => x"3f",
          6210 => x"08",
          6211 => x"82",
          6212 => x"80",
          6213 => x"38",
          6214 => x"d5",
          6215 => x"2e",
          6216 => x"55",
          6217 => x"08",
          6218 => x"38",
          6219 => x"08",
          6220 => x"fb",
          6221 => x"d5",
          6222 => x"38",
          6223 => x"0c",
          6224 => x"51",
          6225 => x"82",
          6226 => x"98",
          6227 => x"90",
          6228 => x"16",
          6229 => x"15",
          6230 => x"74",
          6231 => x"0c",
          6232 => x"04",
          6233 => x"7b",
          6234 => x"5b",
          6235 => x"52",
          6236 => x"ac",
          6237 => x"e4",
          6238 => x"d5",
          6239 => x"ec",
          6240 => x"e4",
          6241 => x"17",
          6242 => x"51",
          6243 => x"82",
          6244 => x"54",
          6245 => x"08",
          6246 => x"82",
          6247 => x"9c",
          6248 => x"33",
          6249 => x"72",
          6250 => x"09",
          6251 => x"38",
          6252 => x"d5",
          6253 => x"72",
          6254 => x"55",
          6255 => x"53",
          6256 => x"8e",
          6257 => x"56",
          6258 => x"09",
          6259 => x"38",
          6260 => x"d5",
          6261 => x"81",
          6262 => x"fd",
          6263 => x"d5",
          6264 => x"82",
          6265 => x"80",
          6266 => x"38",
          6267 => x"09",
          6268 => x"38",
          6269 => x"82",
          6270 => x"8b",
          6271 => x"fd",
          6272 => x"9a",
          6273 => x"eb",
          6274 => x"d5",
          6275 => x"ff",
          6276 => x"70",
          6277 => x"53",
          6278 => x"09",
          6279 => x"38",
          6280 => x"eb",
          6281 => x"d5",
          6282 => x"2b",
          6283 => x"72",
          6284 => x"0c",
          6285 => x"04",
          6286 => x"77",
          6287 => x"ff",
          6288 => x"9a",
          6289 => x"55",
          6290 => x"76",
          6291 => x"53",
          6292 => x"09",
          6293 => x"38",
          6294 => x"52",
          6295 => x"eb",
          6296 => x"3d",
          6297 => x"3d",
          6298 => x"80",
          6299 => x"70",
          6300 => x"81",
          6301 => x"74",
          6302 => x"56",
          6303 => x"70",
          6304 => x"ff",
          6305 => x"51",
          6306 => x"38",
          6307 => x"e4",
          6308 => x"0d",
          6309 => x"0d",
          6310 => x"59",
          6311 => x"5f",
          6312 => x"70",
          6313 => x"19",
          6314 => x"83",
          6315 => x"19",
          6316 => x"51",
          6317 => x"82",
          6318 => x"5b",
          6319 => x"08",
          6320 => x"9c",
          6321 => x"33",
          6322 => x"86",
          6323 => x"82",
          6324 => x"15",
          6325 => x"70",
          6326 => x"58",
          6327 => x"1a",
          6328 => x"e4",
          6329 => x"81",
          6330 => x"81",
          6331 => x"81",
          6332 => x"e4",
          6333 => x"ae",
          6334 => x"06",
          6335 => x"53",
          6336 => x"53",
          6337 => x"82",
          6338 => x"77",
          6339 => x"56",
          6340 => x"09",
          6341 => x"38",
          6342 => x"7f",
          6343 => x"81",
          6344 => x"ef",
          6345 => x"2e",
          6346 => x"81",
          6347 => x"86",
          6348 => x"06",
          6349 => x"80",
          6350 => x"8d",
          6351 => x"81",
          6352 => x"90",
          6353 => x"1d",
          6354 => x"5d",
          6355 => x"09",
          6356 => x"9c",
          6357 => x"33",
          6358 => x"2e",
          6359 => x"81",
          6360 => x"1e",
          6361 => x"52",
          6362 => x"3f",
          6363 => x"08",
          6364 => x"06",
          6365 => x"f8",
          6366 => x"70",
          6367 => x"8d",
          6368 => x"51",
          6369 => x"58",
          6370 => x"e4",
          6371 => x"05",
          6372 => x"3f",
          6373 => x"08",
          6374 => x"06",
          6375 => x"2e",
          6376 => x"81",
          6377 => x"c8",
          6378 => x"1a",
          6379 => x"75",
          6380 => x"14",
          6381 => x"75",
          6382 => x"2e",
          6383 => x"b0",
          6384 => x"57",
          6385 => x"c1",
          6386 => x"70",
          6387 => x"81",
          6388 => x"55",
          6389 => x"8e",
          6390 => x"fe",
          6391 => x"73",
          6392 => x"80",
          6393 => x"1c",
          6394 => x"06",
          6395 => x"39",
          6396 => x"72",
          6397 => x"7b",
          6398 => x"51",
          6399 => x"82",
          6400 => x"81",
          6401 => x"72",
          6402 => x"38",
          6403 => x"1a",
          6404 => x"80",
          6405 => x"f8",
          6406 => x"d5",
          6407 => x"82",
          6408 => x"89",
          6409 => x"08",
          6410 => x"86",
          6411 => x"98",
          6412 => x"82",
          6413 => x"90",
          6414 => x"f2",
          6415 => x"70",
          6416 => x"80",
          6417 => x"f6",
          6418 => x"d5",
          6419 => x"82",
          6420 => x"83",
          6421 => x"ff",
          6422 => x"ff",
          6423 => x"0c",
          6424 => x"52",
          6425 => x"a9",
          6426 => x"e4",
          6427 => x"d5",
          6428 => x"85",
          6429 => x"08",
          6430 => x"57",
          6431 => x"84",
          6432 => x"39",
          6433 => x"bf",
          6434 => x"ff",
          6435 => x"73",
          6436 => x"75",
          6437 => x"82",
          6438 => x"83",
          6439 => x"06",
          6440 => x"8f",
          6441 => x"73",
          6442 => x"74",
          6443 => x"81",
          6444 => x"38",
          6445 => x"70",
          6446 => x"81",
          6447 => x"55",
          6448 => x"38",
          6449 => x"70",
          6450 => x"54",
          6451 => x"92",
          6452 => x"33",
          6453 => x"06",
          6454 => x"08",
          6455 => x"58",
          6456 => x"7c",
          6457 => x"06",
          6458 => x"8d",
          6459 => x"7d",
          6460 => x"81",
          6461 => x"38",
          6462 => x"9a",
          6463 => x"e5",
          6464 => x"d5",
          6465 => x"ff",
          6466 => x"74",
          6467 => x"76",
          6468 => x"06",
          6469 => x"05",
          6470 => x"75",
          6471 => x"c7",
          6472 => x"77",
          6473 => x"8f",
          6474 => x"e4",
          6475 => x"ff",
          6476 => x"80",
          6477 => x"77",
          6478 => x"80",
          6479 => x"51",
          6480 => x"3f",
          6481 => x"08",
          6482 => x"70",
          6483 => x"81",
          6484 => x"80",
          6485 => x"74",
          6486 => x"08",
          6487 => x"06",
          6488 => x"75",
          6489 => x"75",
          6490 => x"2e",
          6491 => x"b3",
          6492 => x"5b",
          6493 => x"ff",
          6494 => x"33",
          6495 => x"70",
          6496 => x"55",
          6497 => x"2e",
          6498 => x"80",
          6499 => x"77",
          6500 => x"22",
          6501 => x"8b",
          6502 => x"70",
          6503 => x"51",
          6504 => x"81",
          6505 => x"5c",
          6506 => x"93",
          6507 => x"f9",
          6508 => x"d5",
          6509 => x"ff",
          6510 => x"7e",
          6511 => x"ab",
          6512 => x"06",
          6513 => x"38",
          6514 => x"19",
          6515 => x"08",
          6516 => x"3f",
          6517 => x"08",
          6518 => x"38",
          6519 => x"ff",
          6520 => x"0c",
          6521 => x"51",
          6522 => x"82",
          6523 => x"58",
          6524 => x"08",
          6525 => x"e8",
          6526 => x"d5",
          6527 => x"3d",
          6528 => x"3d",
          6529 => x"08",
          6530 => x"81",
          6531 => x"5d",
          6532 => x"73",
          6533 => x"73",
          6534 => x"70",
          6535 => x"5d",
          6536 => x"8d",
          6537 => x"70",
          6538 => x"22",
          6539 => x"f0",
          6540 => x"a0",
          6541 => x"92",
          6542 => x"5f",
          6543 => x"3f",
          6544 => x"05",
          6545 => x"54",
          6546 => x"82",
          6547 => x"c0",
          6548 => x"34",
          6549 => x"1c",
          6550 => x"58",
          6551 => x"52",
          6552 => x"e2",
          6553 => x"27",
          6554 => x"7a",
          6555 => x"70",
          6556 => x"06",
          6557 => x"80",
          6558 => x"74",
          6559 => x"06",
          6560 => x"55",
          6561 => x"81",
          6562 => x"07",
          6563 => x"71",
          6564 => x"81",
          6565 => x"56",
          6566 => x"2e",
          6567 => x"84",
          6568 => x"56",
          6569 => x"76",
          6570 => x"38",
          6571 => x"55",
          6572 => x"05",
          6573 => x"57",
          6574 => x"bf",
          6575 => x"74",
          6576 => x"87",
          6577 => x"76",
          6578 => x"ff",
          6579 => x"2a",
          6580 => x"74",
          6581 => x"3d",
          6582 => x"54",
          6583 => x"34",
          6584 => x"b5",
          6585 => x"54",
          6586 => x"ad",
          6587 => x"70",
          6588 => x"e3",
          6589 => x"d5",
          6590 => x"2e",
          6591 => x"17",
          6592 => x"2e",
          6593 => x"15",
          6594 => x"55",
          6595 => x"89",
          6596 => x"70",
          6597 => x"d0",
          6598 => x"77",
          6599 => x"54",
          6600 => x"16",
          6601 => x"56",
          6602 => x"8a",
          6603 => x"81",
          6604 => x"58",
          6605 => x"78",
          6606 => x"27",
          6607 => x"51",
          6608 => x"82",
          6609 => x"8b",
          6610 => x"5b",
          6611 => x"27",
          6612 => x"87",
          6613 => x"e4",
          6614 => x"38",
          6615 => x"08",
          6616 => x"e4",
          6617 => x"09",
          6618 => x"df",
          6619 => x"cb",
          6620 => x"1b",
          6621 => x"cb",
          6622 => x"81",
          6623 => x"06",
          6624 => x"81",
          6625 => x"2e",
          6626 => x"52",
          6627 => x"fe",
          6628 => x"82",
          6629 => x"19",
          6630 => x"79",
          6631 => x"3f",
          6632 => x"08",
          6633 => x"e4",
          6634 => x"38",
          6635 => x"78",
          6636 => x"d4",
          6637 => x"2b",
          6638 => x"71",
          6639 => x"79",
          6640 => x"3f",
          6641 => x"08",
          6642 => x"e4",
          6643 => x"38",
          6644 => x"f5",
          6645 => x"d5",
          6646 => x"ff",
          6647 => x"1a",
          6648 => x"51",
          6649 => x"82",
          6650 => x"57",
          6651 => x"08",
          6652 => x"8c",
          6653 => x"1b",
          6654 => x"ff",
          6655 => x"5b",
          6656 => x"34",
          6657 => x"17",
          6658 => x"e4",
          6659 => x"34",
          6660 => x"08",
          6661 => x"51",
          6662 => x"77",
          6663 => x"05",
          6664 => x"73",
          6665 => x"2e",
          6666 => x"10",
          6667 => x"81",
          6668 => x"54",
          6669 => x"c7",
          6670 => x"76",
          6671 => x"b9",
          6672 => x"38",
          6673 => x"54",
          6674 => x"8c",
          6675 => x"38",
          6676 => x"ff",
          6677 => x"74",
          6678 => x"22",
          6679 => x"86",
          6680 => x"c0",
          6681 => x"76",
          6682 => x"83",
          6683 => x"52",
          6684 => x"f7",
          6685 => x"e4",
          6686 => x"d5",
          6687 => x"c9",
          6688 => x"59",
          6689 => x"38",
          6690 => x"52",
          6691 => x"81",
          6692 => x"e4",
          6693 => x"d5",
          6694 => x"38",
          6695 => x"d5",
          6696 => x"9c",
          6697 => x"df",
          6698 => x"53",
          6699 => x"9c",
          6700 => x"df",
          6701 => x"1a",
          6702 => x"33",
          6703 => x"55",
          6704 => x"34",
          6705 => x"1d",
          6706 => x"74",
          6707 => x"0c",
          6708 => x"04",
          6709 => x"78",
          6710 => x"12",
          6711 => x"08",
          6712 => x"55",
          6713 => x"94",
          6714 => x"74",
          6715 => x"3f",
          6716 => x"08",
          6717 => x"e4",
          6718 => x"38",
          6719 => x"52",
          6720 => x"8d",
          6721 => x"e4",
          6722 => x"d5",
          6723 => x"38",
          6724 => x"53",
          6725 => x"81",
          6726 => x"34",
          6727 => x"77",
          6728 => x"82",
          6729 => x"52",
          6730 => x"bf",
          6731 => x"e4",
          6732 => x"d5",
          6733 => x"2e",
          6734 => x"84",
          6735 => x"06",
          6736 => x"54",
          6737 => x"e4",
          6738 => x"0d",
          6739 => x"0d",
          6740 => x"08",
          6741 => x"80",
          6742 => x"34",
          6743 => x"80",
          6744 => x"38",
          6745 => x"ff",
          6746 => x"38",
          6747 => x"7f",
          6748 => x"70",
          6749 => x"5b",
          6750 => x"77",
          6751 => x"38",
          6752 => x"70",
          6753 => x"5b",
          6754 => x"97",
          6755 => x"80",
          6756 => x"ff",
          6757 => x"53",
          6758 => x"26",
          6759 => x"5b",
          6760 => x"76",
          6761 => x"81",
          6762 => x"58",
          6763 => x"b5",
          6764 => x"2b",
          6765 => x"80",
          6766 => x"82",
          6767 => x"83",
          6768 => x"55",
          6769 => x"27",
          6770 => x"76",
          6771 => x"74",
          6772 => x"72",
          6773 => x"97",
          6774 => x"55",
          6775 => x"30",
          6776 => x"78",
          6777 => x"72",
          6778 => x"52",
          6779 => x"80",
          6780 => x"80",
          6781 => x"74",
          6782 => x"55",
          6783 => x"80",
          6784 => x"08",
          6785 => x"70",
          6786 => x"54",
          6787 => x"38",
          6788 => x"80",
          6789 => x"79",
          6790 => x"53",
          6791 => x"05",
          6792 => x"82",
          6793 => x"70",
          6794 => x"5a",
          6795 => x"08",
          6796 => x"81",
          6797 => x"53",
          6798 => x"b7",
          6799 => x"2e",
          6800 => x"84",
          6801 => x"55",
          6802 => x"70",
          6803 => x"07",
          6804 => x"54",
          6805 => x"26",
          6806 => x"80",
          6807 => x"ae",
          6808 => x"05",
          6809 => x"17",
          6810 => x"70",
          6811 => x"34",
          6812 => x"8a",
          6813 => x"b5",
          6814 => x"88",
          6815 => x"0b",
          6816 => x"96",
          6817 => x"72",
          6818 => x"76",
          6819 => x"0b",
          6820 => x"81",
          6821 => x"39",
          6822 => x"1a",
          6823 => x"57",
          6824 => x"80",
          6825 => x"18",
          6826 => x"56",
          6827 => x"bf",
          6828 => x"72",
          6829 => x"38",
          6830 => x"8c",
          6831 => x"53",
          6832 => x"87",
          6833 => x"2a",
          6834 => x"72",
          6835 => x"72",
          6836 => x"72",
          6837 => x"38",
          6838 => x"83",
          6839 => x"56",
          6840 => x"70",
          6841 => x"34",
          6842 => x"15",
          6843 => x"33",
          6844 => x"59",
          6845 => x"38",
          6846 => x"05",
          6847 => x"82",
          6848 => x"1c",
          6849 => x"33",
          6850 => x"85",
          6851 => x"19",
          6852 => x"08",
          6853 => x"33",
          6854 => x"9c",
          6855 => x"11",
          6856 => x"aa",
          6857 => x"e4",
          6858 => x"96",
          6859 => x"87",
          6860 => x"e4",
          6861 => x"23",
          6862 => x"d8",
          6863 => x"d5",
          6864 => x"19",
          6865 => x"0d",
          6866 => x"0d",
          6867 => x"41",
          6868 => x"70",
          6869 => x"55",
          6870 => x"83",
          6871 => x"73",
          6872 => x"92",
          6873 => x"2e",
          6874 => x"98",
          6875 => x"1f",
          6876 => x"81",
          6877 => x"64",
          6878 => x"56",
          6879 => x"2e",
          6880 => x"83",
          6881 => x"73",
          6882 => x"70",
          6883 => x"25",
          6884 => x"51",
          6885 => x"38",
          6886 => x"0c",
          6887 => x"51",
          6888 => x"26",
          6889 => x"80",
          6890 => x"34",
          6891 => x"51",
          6892 => x"82",
          6893 => x"56",
          6894 => x"63",
          6895 => x"8c",
          6896 => x"54",
          6897 => x"3d",
          6898 => x"da",
          6899 => x"d5",
          6900 => x"2e",
          6901 => x"83",
          6902 => x"82",
          6903 => x"27",
          6904 => x"10",
          6905 => x"e4",
          6906 => x"55",
          6907 => x"23",
          6908 => x"82",
          6909 => x"83",
          6910 => x"70",
          6911 => x"30",
          6912 => x"71",
          6913 => x"51",
          6914 => x"73",
          6915 => x"80",
          6916 => x"38",
          6917 => x"26",
          6918 => x"52",
          6919 => x"51",
          6920 => x"82",
          6921 => x"81",
          6922 => x"81",
          6923 => x"d7",
          6924 => x"1a",
          6925 => x"23",
          6926 => x"ff",
          6927 => x"15",
          6928 => x"70",
          6929 => x"57",
          6930 => x"09",
          6931 => x"38",
          6932 => x"80",
          6933 => x"30",
          6934 => x"79",
          6935 => x"54",
          6936 => x"74",
          6937 => x"27",
          6938 => x"78",
          6939 => x"81",
          6940 => x"79",
          6941 => x"ae",
          6942 => x"80",
          6943 => x"82",
          6944 => x"06",
          6945 => x"82",
          6946 => x"73",
          6947 => x"81",
          6948 => x"38",
          6949 => x"73",
          6950 => x"81",
          6951 => x"78",
          6952 => x"80",
          6953 => x"0b",
          6954 => x"58",
          6955 => x"78",
          6956 => x"a0",
          6957 => x"70",
          6958 => x"34",
          6959 => x"8a",
          6960 => x"38",
          6961 => x"54",
          6962 => x"34",
          6963 => x"78",
          6964 => x"38",
          6965 => x"fe",
          6966 => x"22",
          6967 => x"72",
          6968 => x"30",
          6969 => x"51",
          6970 => x"56",
          6971 => x"2e",
          6972 => x"87",
          6973 => x"59",
          6974 => x"78",
          6975 => x"55",
          6976 => x"23",
          6977 => x"86",
          6978 => x"39",
          6979 => x"57",
          6980 => x"80",
          6981 => x"83",
          6982 => x"56",
          6983 => x"a0",
          6984 => x"06",
          6985 => x"1d",
          6986 => x"70",
          6987 => x"5d",
          6988 => x"f2",
          6989 => x"38",
          6990 => x"ff",
          6991 => x"ae",
          6992 => x"06",
          6993 => x"83",
          6994 => x"80",
          6995 => x"79",
          6996 => x"70",
          6997 => x"73",
          6998 => x"38",
          6999 => x"fe",
          7000 => x"19",
          7001 => x"2e",
          7002 => x"15",
          7003 => x"55",
          7004 => x"09",
          7005 => x"38",
          7006 => x"52",
          7007 => x"d5",
          7008 => x"70",
          7009 => x"5f",
          7010 => x"70",
          7011 => x"5f",
          7012 => x"80",
          7013 => x"38",
          7014 => x"96",
          7015 => x"32",
          7016 => x"80",
          7017 => x"54",
          7018 => x"8c",
          7019 => x"2e",
          7020 => x"83",
          7021 => x"39",
          7022 => x"5b",
          7023 => x"83",
          7024 => x"7c",
          7025 => x"30",
          7026 => x"80",
          7027 => x"07",
          7028 => x"55",
          7029 => x"a6",
          7030 => x"2e",
          7031 => x"7c",
          7032 => x"38",
          7033 => x"57",
          7034 => x"81",
          7035 => x"5d",
          7036 => x"7c",
          7037 => x"fc",
          7038 => x"ff",
          7039 => x"ff",
          7040 => x"38",
          7041 => x"57",
          7042 => x"75",
          7043 => x"ae",
          7044 => x"e4",
          7045 => x"ff",
          7046 => x"2a",
          7047 => x"51",
          7048 => x"80",
          7049 => x"75",
          7050 => x"82",
          7051 => x"33",
          7052 => x"ff",
          7053 => x"38",
          7054 => x"73",
          7055 => x"38",
          7056 => x"7f",
          7057 => x"c0",
          7058 => x"a0",
          7059 => x"2a",
          7060 => x"75",
          7061 => x"58",
          7062 => x"75",
          7063 => x"38",
          7064 => x"c7",
          7065 => x"cc",
          7066 => x"e4",
          7067 => x"8a",
          7068 => x"77",
          7069 => x"56",
          7070 => x"bf",
          7071 => x"99",
          7072 => x"7b",
          7073 => x"ff",
          7074 => x"73",
          7075 => x"38",
          7076 => x"e0",
          7077 => x"ff",
          7078 => x"55",
          7079 => x"a0",
          7080 => x"74",
          7081 => x"58",
          7082 => x"a0",
          7083 => x"73",
          7084 => x"09",
          7085 => x"38",
          7086 => x"1f",
          7087 => x"2e",
          7088 => x"88",
          7089 => x"2b",
          7090 => x"5c",
          7091 => x"54",
          7092 => x"8d",
          7093 => x"06",
          7094 => x"2e",
          7095 => x"85",
          7096 => x"07",
          7097 => x"2a",
          7098 => x"51",
          7099 => x"38",
          7100 => x"54",
          7101 => x"85",
          7102 => x"07",
          7103 => x"2a",
          7104 => x"51",
          7105 => x"2e",
          7106 => x"88",
          7107 => x"ab",
          7108 => x"51",
          7109 => x"82",
          7110 => x"ab",
          7111 => x"56",
          7112 => x"08",
          7113 => x"38",
          7114 => x"08",
          7115 => x"81",
          7116 => x"38",
          7117 => x"70",
          7118 => x"82",
          7119 => x"54",
          7120 => x"96",
          7121 => x"06",
          7122 => x"2e",
          7123 => x"ff",
          7124 => x"1f",
          7125 => x"80",
          7126 => x"81",
          7127 => x"bb",
          7128 => x"b7",
          7129 => x"2a",
          7130 => x"51",
          7131 => x"38",
          7132 => x"70",
          7133 => x"81",
          7134 => x"55",
          7135 => x"e1",
          7136 => x"08",
          7137 => x"60",
          7138 => x"52",
          7139 => x"ef",
          7140 => x"e4",
          7141 => x"0c",
          7142 => x"75",
          7143 => x"0c",
          7144 => x"04",
          7145 => x"7c",
          7146 => x"08",
          7147 => x"55",
          7148 => x"59",
          7149 => x"81",
          7150 => x"70",
          7151 => x"33",
          7152 => x"52",
          7153 => x"2e",
          7154 => x"ee",
          7155 => x"2e",
          7156 => x"81",
          7157 => x"33",
          7158 => x"81",
          7159 => x"52",
          7160 => x"26",
          7161 => x"14",
          7162 => x"06",
          7163 => x"52",
          7164 => x"80",
          7165 => x"0b",
          7166 => x"59",
          7167 => x"7a",
          7168 => x"70",
          7169 => x"33",
          7170 => x"05",
          7171 => x"9f",
          7172 => x"53",
          7173 => x"89",
          7174 => x"70",
          7175 => x"54",
          7176 => x"12",
          7177 => x"26",
          7178 => x"12",
          7179 => x"06",
          7180 => x"30",
          7181 => x"51",
          7182 => x"2e",
          7183 => x"85",
          7184 => x"be",
          7185 => x"74",
          7186 => x"30",
          7187 => x"9f",
          7188 => x"2a",
          7189 => x"54",
          7190 => x"2e",
          7191 => x"15",
          7192 => x"55",
          7193 => x"ff",
          7194 => x"39",
          7195 => x"86",
          7196 => x"7c",
          7197 => x"51",
          7198 => x"ed",
          7199 => x"70",
          7200 => x"0c",
          7201 => x"04",
          7202 => x"78",
          7203 => x"83",
          7204 => x"0b",
          7205 => x"79",
          7206 => x"d1",
          7207 => x"55",
          7208 => x"08",
          7209 => x"84",
          7210 => x"ce",
          7211 => x"d5",
          7212 => x"ff",
          7213 => x"83",
          7214 => x"d4",
          7215 => x"81",
          7216 => x"38",
          7217 => x"17",
          7218 => x"74",
          7219 => x"09",
          7220 => x"38",
          7221 => x"81",
          7222 => x"30",
          7223 => x"79",
          7224 => x"54",
          7225 => x"74",
          7226 => x"09",
          7227 => x"38",
          7228 => x"c7",
          7229 => x"ee",
          7230 => x"87",
          7231 => x"e4",
          7232 => x"d5",
          7233 => x"2e",
          7234 => x"53",
          7235 => x"52",
          7236 => x"51",
          7237 => x"82",
          7238 => x"55",
          7239 => x"08",
          7240 => x"38",
          7241 => x"82",
          7242 => x"88",
          7243 => x"f2",
          7244 => x"02",
          7245 => x"cb",
          7246 => x"55",
          7247 => x"60",
          7248 => x"3f",
          7249 => x"08",
          7250 => x"80",
          7251 => x"e4",
          7252 => x"c7",
          7253 => x"e4",
          7254 => x"82",
          7255 => x"70",
          7256 => x"8c",
          7257 => x"2e",
          7258 => x"73",
          7259 => x"81",
          7260 => x"33",
          7261 => x"80",
          7262 => x"81",
          7263 => x"c6",
          7264 => x"d5",
          7265 => x"ff",
          7266 => x"06",
          7267 => x"98",
          7268 => x"2e",
          7269 => x"74",
          7270 => x"81",
          7271 => x"8a",
          7272 => x"f7",
          7273 => x"39",
          7274 => x"77",
          7275 => x"d5",
          7276 => x"81",
          7277 => x"52",
          7278 => x"51",
          7279 => x"82",
          7280 => x"81",
          7281 => x"81",
          7282 => x"83",
          7283 => x"cb",
          7284 => x"2e",
          7285 => x"82",
          7286 => x"06",
          7287 => x"56",
          7288 => x"38",
          7289 => x"74",
          7290 => x"9c",
          7291 => x"e4",
          7292 => x"06",
          7293 => x"2e",
          7294 => x"81",
          7295 => x"38",
          7296 => x"19",
          7297 => x"7b",
          7298 => x"38",
          7299 => x"56",
          7300 => x"83",
          7301 => x"70",
          7302 => x"80",
          7303 => x"83",
          7304 => x"cb",
          7305 => x"d5",
          7306 => x"76",
          7307 => x"05",
          7308 => x"16",
          7309 => x"56",
          7310 => x"d7",
          7311 => x"82",
          7312 => x"33",
          7313 => x"9f",
          7314 => x"31",
          7315 => x"84",
          7316 => x"05",
          7317 => x"55",
          7318 => x"08",
          7319 => x"7a",
          7320 => x"38",
          7321 => x"51",
          7322 => x"82",
          7323 => x"81",
          7324 => x"80",
          7325 => x"d9",
          7326 => x"58",
          7327 => x"09",
          7328 => x"38",
          7329 => x"77",
          7330 => x"77",
          7331 => x"38",
          7332 => x"16",
          7333 => x"76",
          7334 => x"81",
          7335 => x"2e",
          7336 => x"8d",
          7337 => x"26",
          7338 => x"80",
          7339 => x"ca",
          7340 => x"d5",
          7341 => x"ff",
          7342 => x"72",
          7343 => x"09",
          7344 => x"d7",
          7345 => x"14",
          7346 => x"3f",
          7347 => x"08",
          7348 => x"06",
          7349 => x"38",
          7350 => x"51",
          7351 => x"82",
          7352 => x"58",
          7353 => x"0c",
          7354 => x"33",
          7355 => x"80",
          7356 => x"ff",
          7357 => x"ff",
          7358 => x"55",
          7359 => x"81",
          7360 => x"38",
          7361 => x"06",
          7362 => x"80",
          7363 => x"52",
          7364 => x"8a",
          7365 => x"80",
          7366 => x"ff",
          7367 => x"53",
          7368 => x"86",
          7369 => x"83",
          7370 => x"c9",
          7371 => x"87",
          7372 => x"e4",
          7373 => x"d5",
          7374 => x"15",
          7375 => x"06",
          7376 => x"76",
          7377 => x"80",
          7378 => x"c8",
          7379 => x"d5",
          7380 => x"ff",
          7381 => x"74",
          7382 => x"d8",
          7383 => x"ee",
          7384 => x"e4",
          7385 => x"c6",
          7386 => x"cb",
          7387 => x"e4",
          7388 => x"ff",
          7389 => x"56",
          7390 => x"83",
          7391 => x"14",
          7392 => x"71",
          7393 => x"5a",
          7394 => x"26",
          7395 => x"8a",
          7396 => x"74",
          7397 => x"fe",
          7398 => x"82",
          7399 => x"55",
          7400 => x"08",
          7401 => x"f3",
          7402 => x"e4",
          7403 => x"ff",
          7404 => x"83",
          7405 => x"74",
          7406 => x"26",
          7407 => x"57",
          7408 => x"26",
          7409 => x"57",
          7410 => x"56",
          7411 => x"82",
          7412 => x"15",
          7413 => x"0c",
          7414 => x"0c",
          7415 => x"a8",
          7416 => x"1d",
          7417 => x"54",
          7418 => x"2e",
          7419 => x"af",
          7420 => x"14",
          7421 => x"3f",
          7422 => x"08",
          7423 => x"06",
          7424 => x"72",
          7425 => x"79",
          7426 => x"80",
          7427 => x"c7",
          7428 => x"d5",
          7429 => x"15",
          7430 => x"2b",
          7431 => x"8d",
          7432 => x"2e",
          7433 => x"77",
          7434 => x"0c",
          7435 => x"76",
          7436 => x"38",
          7437 => x"70",
          7438 => x"81",
          7439 => x"53",
          7440 => x"89",
          7441 => x"56",
          7442 => x"08",
          7443 => x"38",
          7444 => x"15",
          7445 => x"90",
          7446 => x"80",
          7447 => x"34",
          7448 => x"09",
          7449 => x"92",
          7450 => x"14",
          7451 => x"3f",
          7452 => x"08",
          7453 => x"06",
          7454 => x"2e",
          7455 => x"80",
          7456 => x"1b",
          7457 => x"ca",
          7458 => x"d5",
          7459 => x"ea",
          7460 => x"e4",
          7461 => x"34",
          7462 => x"51",
          7463 => x"82",
          7464 => x"83",
          7465 => x"53",
          7466 => x"d5",
          7467 => x"06",
          7468 => x"b8",
          7469 => x"96",
          7470 => x"e4",
          7471 => x"85",
          7472 => x"09",
          7473 => x"38",
          7474 => x"51",
          7475 => x"82",
          7476 => x"86",
          7477 => x"f2",
          7478 => x"06",
          7479 => x"a0",
          7480 => x"ea",
          7481 => x"e4",
          7482 => x"0c",
          7483 => x"51",
          7484 => x"82",
          7485 => x"90",
          7486 => x"74",
          7487 => x"bc",
          7488 => x"53",
          7489 => x"bc",
          7490 => x"15",
          7491 => x"c4",
          7492 => x"0c",
          7493 => x"15",
          7494 => x"75",
          7495 => x"0c",
          7496 => x"04",
          7497 => x"77",
          7498 => x"73",
          7499 => x"38",
          7500 => x"72",
          7501 => x"38",
          7502 => x"71",
          7503 => x"38",
          7504 => x"84",
          7505 => x"52",
          7506 => x"09",
          7507 => x"38",
          7508 => x"51",
          7509 => x"3f",
          7510 => x"08",
          7511 => x"71",
          7512 => x"74",
          7513 => x"83",
          7514 => x"78",
          7515 => x"52",
          7516 => x"e4",
          7517 => x"0d",
          7518 => x"0d",
          7519 => x"33",
          7520 => x"3d",
          7521 => x"56",
          7522 => x"8b",
          7523 => x"82",
          7524 => x"24",
          7525 => x"d5",
          7526 => x"29",
          7527 => x"05",
          7528 => x"55",
          7529 => x"84",
          7530 => x"34",
          7531 => x"80",
          7532 => x"80",
          7533 => x"75",
          7534 => x"75",
          7535 => x"38",
          7536 => x"3d",
          7537 => x"05",
          7538 => x"3f",
          7539 => x"08",
          7540 => x"d5",
          7541 => x"3d",
          7542 => x"3d",
          7543 => x"84",
          7544 => x"05",
          7545 => x"89",
          7546 => x"2e",
          7547 => x"77",
          7548 => x"54",
          7549 => x"05",
          7550 => x"84",
          7551 => x"f6",
          7552 => x"d5",
          7553 => x"82",
          7554 => x"84",
          7555 => x"5c",
          7556 => x"3d",
          7557 => x"ea",
          7558 => x"d5",
          7559 => x"82",
          7560 => x"92",
          7561 => x"d7",
          7562 => x"98",
          7563 => x"73",
          7564 => x"38",
          7565 => x"9c",
          7566 => x"80",
          7567 => x"38",
          7568 => x"95",
          7569 => x"2e",
          7570 => x"aa",
          7571 => x"df",
          7572 => x"d5",
          7573 => x"9e",
          7574 => x"05",
          7575 => x"54",
          7576 => x"38",
          7577 => x"70",
          7578 => x"54",
          7579 => x"8e",
          7580 => x"83",
          7581 => x"88",
          7582 => x"83",
          7583 => x"83",
          7584 => x"06",
          7585 => x"80",
          7586 => x"38",
          7587 => x"51",
          7588 => x"82",
          7589 => x"56",
          7590 => x"0a",
          7591 => x"05",
          7592 => x"3f",
          7593 => x"0b",
          7594 => x"80",
          7595 => x"7a",
          7596 => x"3f",
          7597 => x"9c",
          7598 => x"db",
          7599 => x"81",
          7600 => x"34",
          7601 => x"80",
          7602 => x"b4",
          7603 => x"54",
          7604 => x"52",
          7605 => x"05",
          7606 => x"3f",
          7607 => x"08",
          7608 => x"e4",
          7609 => x"38",
          7610 => x"82",
          7611 => x"b2",
          7612 => x"84",
          7613 => x"06",
          7614 => x"73",
          7615 => x"38",
          7616 => x"ad",
          7617 => x"2a",
          7618 => x"51",
          7619 => x"2e",
          7620 => x"81",
          7621 => x"80",
          7622 => x"87",
          7623 => x"39",
          7624 => x"51",
          7625 => x"82",
          7626 => x"7b",
          7627 => x"12",
          7628 => x"82",
          7629 => x"81",
          7630 => x"83",
          7631 => x"06",
          7632 => x"80",
          7633 => x"77",
          7634 => x"58",
          7635 => x"08",
          7636 => x"63",
          7637 => x"63",
          7638 => x"57",
          7639 => x"82",
          7640 => x"82",
          7641 => x"88",
          7642 => x"9c",
          7643 => x"c0",
          7644 => x"d5",
          7645 => x"d5",
          7646 => x"1b",
          7647 => x"0c",
          7648 => x"22",
          7649 => x"77",
          7650 => x"80",
          7651 => x"34",
          7652 => x"1a",
          7653 => x"94",
          7654 => x"85",
          7655 => x"06",
          7656 => x"80",
          7657 => x"38",
          7658 => x"08",
          7659 => x"84",
          7660 => x"e4",
          7661 => x"0c",
          7662 => x"70",
          7663 => x"52",
          7664 => x"39",
          7665 => x"51",
          7666 => x"82",
          7667 => x"57",
          7668 => x"08",
          7669 => x"38",
          7670 => x"d5",
          7671 => x"2e",
          7672 => x"83",
          7673 => x"75",
          7674 => x"74",
          7675 => x"07",
          7676 => x"54",
          7677 => x"8a",
          7678 => x"75",
          7679 => x"73",
          7680 => x"98",
          7681 => x"a9",
          7682 => x"ff",
          7683 => x"80",
          7684 => x"76",
          7685 => x"c4",
          7686 => x"d5",
          7687 => x"38",
          7688 => x"39",
          7689 => x"82",
          7690 => x"05",
          7691 => x"84",
          7692 => x"0c",
          7693 => x"82",
          7694 => x"98",
          7695 => x"f2",
          7696 => x"63",
          7697 => x"40",
          7698 => x"7e",
          7699 => x"fc",
          7700 => x"51",
          7701 => x"82",
          7702 => x"55",
          7703 => x"08",
          7704 => x"19",
          7705 => x"80",
          7706 => x"74",
          7707 => x"39",
          7708 => x"81",
          7709 => x"56",
          7710 => x"82",
          7711 => x"39",
          7712 => x"1a",
          7713 => x"82",
          7714 => x"0b",
          7715 => x"81",
          7716 => x"39",
          7717 => x"94",
          7718 => x"55",
          7719 => x"83",
          7720 => x"7b",
          7721 => x"8c",
          7722 => x"08",
          7723 => x"06",
          7724 => x"81",
          7725 => x"8a",
          7726 => x"05",
          7727 => x"06",
          7728 => x"a8",
          7729 => x"38",
          7730 => x"55",
          7731 => x"19",
          7732 => x"51",
          7733 => x"82",
          7734 => x"55",
          7735 => x"ff",
          7736 => x"ff",
          7737 => x"38",
          7738 => x"0c",
          7739 => x"52",
          7740 => x"93",
          7741 => x"e4",
          7742 => x"ff",
          7743 => x"d5",
          7744 => x"7c",
          7745 => x"57",
          7746 => x"80",
          7747 => x"1a",
          7748 => x"22",
          7749 => x"75",
          7750 => x"38",
          7751 => x"58",
          7752 => x"53",
          7753 => x"1b",
          7754 => x"b8",
          7755 => x"d5",
          7756 => x"d6",
          7757 => x"11",
          7758 => x"74",
          7759 => x"38",
          7760 => x"77",
          7761 => x"78",
          7762 => x"84",
          7763 => x"16",
          7764 => x"08",
          7765 => x"2b",
          7766 => x"ff",
          7767 => x"77",
          7768 => x"ba",
          7769 => x"1a",
          7770 => x"08",
          7771 => x"84",
          7772 => x"57",
          7773 => x"27",
          7774 => x"56",
          7775 => x"52",
          7776 => x"8d",
          7777 => x"e4",
          7778 => x"38",
          7779 => x"19",
          7780 => x"06",
          7781 => x"52",
          7782 => x"bd",
          7783 => x"76",
          7784 => x"17",
          7785 => x"1e",
          7786 => x"18",
          7787 => x"5e",
          7788 => x"39",
          7789 => x"82",
          7790 => x"90",
          7791 => x"f2",
          7792 => x"63",
          7793 => x"40",
          7794 => x"7e",
          7795 => x"fc",
          7796 => x"51",
          7797 => x"82",
          7798 => x"55",
          7799 => x"08",
          7800 => x"18",
          7801 => x"80",
          7802 => x"74",
          7803 => x"39",
          7804 => x"70",
          7805 => x"81",
          7806 => x"56",
          7807 => x"80",
          7808 => x"38",
          7809 => x"0b",
          7810 => x"82",
          7811 => x"39",
          7812 => x"19",
          7813 => x"83",
          7814 => x"18",
          7815 => x"56",
          7816 => x"27",
          7817 => x"09",
          7818 => x"2e",
          7819 => x"94",
          7820 => x"83",
          7821 => x"56",
          7822 => x"38",
          7823 => x"22",
          7824 => x"89",
          7825 => x"55",
          7826 => x"75",
          7827 => x"18",
          7828 => x"9c",
          7829 => x"85",
          7830 => x"08",
          7831 => x"c6",
          7832 => x"d5",
          7833 => x"82",
          7834 => x"80",
          7835 => x"38",
          7836 => x"ff",
          7837 => x"ff",
          7838 => x"38",
          7839 => x"0c",
          7840 => x"85",
          7841 => x"19",
          7842 => x"b4",
          7843 => x"19",
          7844 => x"81",
          7845 => x"74",
          7846 => x"85",
          7847 => x"e4",
          7848 => x"38",
          7849 => x"52",
          7850 => x"bf",
          7851 => x"d5",
          7852 => x"2e",
          7853 => x"82",
          7854 => x"1b",
          7855 => x"5a",
          7856 => x"2e",
          7857 => x"78",
          7858 => x"11",
          7859 => x"55",
          7860 => x"85",
          7861 => x"31",
          7862 => x"76",
          7863 => x"81",
          7864 => x"ff",
          7865 => x"82",
          7866 => x"fe",
          7867 => x"b4",
          7868 => x"31",
          7869 => x"79",
          7870 => x"84",
          7871 => x"16",
          7872 => x"89",
          7873 => x"52",
          7874 => x"ff",
          7875 => x"7e",
          7876 => x"83",
          7877 => x"89",
          7878 => x"de",
          7879 => x"08",
          7880 => x"26",
          7881 => x"51",
          7882 => x"3f",
          7883 => x"08",
          7884 => x"7e",
          7885 => x"0c",
          7886 => x"19",
          7887 => x"08",
          7888 => x"84",
          7889 => x"57",
          7890 => x"27",
          7891 => x"56",
          7892 => x"52",
          7893 => x"bc",
          7894 => x"d5",
          7895 => x"b0",
          7896 => x"7c",
          7897 => x"08",
          7898 => x"1f",
          7899 => x"ff",
          7900 => x"7e",
          7901 => x"83",
          7902 => x"76",
          7903 => x"17",
          7904 => x"1e",
          7905 => x"18",
          7906 => x"0c",
          7907 => x"58",
          7908 => x"74",
          7909 => x"38",
          7910 => x"8c",
          7911 => x"89",
          7912 => x"33",
          7913 => x"55",
          7914 => x"34",
          7915 => x"82",
          7916 => x"90",
          7917 => x"f8",
          7918 => x"8b",
          7919 => x"53",
          7920 => x"f2",
          7921 => x"d5",
          7922 => x"82",
          7923 => x"81",
          7924 => x"16",
          7925 => x"2a",
          7926 => x"51",
          7927 => x"80",
          7928 => x"38",
          7929 => x"52",
          7930 => x"bb",
          7931 => x"d5",
          7932 => x"82",
          7933 => x"80",
          7934 => x"16",
          7935 => x"33",
          7936 => x"55",
          7937 => x"34",
          7938 => x"53",
          7939 => x"08",
          7940 => x"3f",
          7941 => x"52",
          7942 => x"ff",
          7943 => x"82",
          7944 => x"52",
          7945 => x"ff",
          7946 => x"76",
          7947 => x"51",
          7948 => x"3f",
          7949 => x"0b",
          7950 => x"78",
          7951 => x"98",
          7952 => x"e4",
          7953 => x"33",
          7954 => x"55",
          7955 => x"17",
          7956 => x"d5",
          7957 => x"3d",
          7958 => x"3d",
          7959 => x"52",
          7960 => x"3f",
          7961 => x"08",
          7962 => x"e4",
          7963 => x"86",
          7964 => x"52",
          7965 => x"ac",
          7966 => x"e4",
          7967 => x"d5",
          7968 => x"38",
          7969 => x"08",
          7970 => x"82",
          7971 => x"86",
          7972 => x"ff",
          7973 => x"3d",
          7974 => x"3f",
          7975 => x"0b",
          7976 => x"08",
          7977 => x"82",
          7978 => x"82",
          7979 => x"80",
          7980 => x"d5",
          7981 => x"3d",
          7982 => x"3d",
          7983 => x"94",
          7984 => x"52",
          7985 => x"e8",
          7986 => x"d5",
          7987 => x"82",
          7988 => x"80",
          7989 => x"58",
          7990 => x"3d",
          7991 => x"dc",
          7992 => x"d5",
          7993 => x"82",
          7994 => x"bc",
          7995 => x"c7",
          7996 => x"98",
          7997 => x"73",
          7998 => x"38",
          7999 => x"12",
          8000 => x"39",
          8001 => x"33",
          8002 => x"70",
          8003 => x"55",
          8004 => x"2e",
          8005 => x"7f",
          8006 => x"54",
          8007 => x"82",
          8008 => x"98",
          8009 => x"39",
          8010 => x"08",
          8011 => x"81",
          8012 => x"85",
          8013 => x"d5",
          8014 => x"3d",
          8015 => x"a3",
          8016 => x"e1",
          8017 => x"e1",
          8018 => x"5b",
          8019 => x"80",
          8020 => x"3d",
          8021 => x"52",
          8022 => x"51",
          8023 => x"82",
          8024 => x"57",
          8025 => x"08",
          8026 => x"7b",
          8027 => x"0c",
          8028 => x"11",
          8029 => x"3d",
          8030 => x"80",
          8031 => x"54",
          8032 => x"82",
          8033 => x"52",
          8034 => x"70",
          8035 => x"90",
          8036 => x"e4",
          8037 => x"d5",
          8038 => x"ef",
          8039 => x"3d",
          8040 => x"51",
          8041 => x"3f",
          8042 => x"08",
          8043 => x"e4",
          8044 => x"38",
          8045 => x"08",
          8046 => x"c8",
          8047 => x"d5",
          8048 => x"d6",
          8049 => x"52",
          8050 => x"d4",
          8051 => x"e4",
          8052 => x"d5",
          8053 => x"b3",
          8054 => x"74",
          8055 => x"3f",
          8056 => x"08",
          8057 => x"e4",
          8058 => x"80",
          8059 => x"52",
          8060 => x"8b",
          8061 => x"d5",
          8062 => x"a6",
          8063 => x"74",
          8064 => x"3f",
          8065 => x"08",
          8066 => x"e4",
          8067 => x"c9",
          8068 => x"2e",
          8069 => x"86",
          8070 => x"81",
          8071 => x"81",
          8072 => x"df",
          8073 => x"05",
          8074 => x"d6",
          8075 => x"93",
          8076 => x"82",
          8077 => x"56",
          8078 => x"80",
          8079 => x"02",
          8080 => x"55",
          8081 => x"16",
          8082 => x"56",
          8083 => x"38",
          8084 => x"73",
          8085 => x"99",
          8086 => x"2e",
          8087 => x"16",
          8088 => x"ff",
          8089 => x"3d",
          8090 => x"18",
          8091 => x"58",
          8092 => x"33",
          8093 => x"eb",
          8094 => x"80",
          8095 => x"11",
          8096 => x"74",
          8097 => x"39",
          8098 => x"09",
          8099 => x"38",
          8100 => x"e1",
          8101 => x"55",
          8102 => x"34",
          8103 => x"ed",
          8104 => x"84",
          8105 => x"d4",
          8106 => x"70",
          8107 => x"56",
          8108 => x"76",
          8109 => x"81",
          8110 => x"70",
          8111 => x"56",
          8112 => x"82",
          8113 => x"78",
          8114 => x"80",
          8115 => x"27",
          8116 => x"19",
          8117 => x"7a",
          8118 => x"5c",
          8119 => x"55",
          8120 => x"7a",
          8121 => x"5c",
          8122 => x"2e",
          8123 => x"85",
          8124 => x"97",
          8125 => x"3d",
          8126 => x"19",
          8127 => x"33",
          8128 => x"05",
          8129 => x"78",
          8130 => x"80",
          8131 => x"82",
          8132 => x"80",
          8133 => x"04",
          8134 => x"7b",
          8135 => x"fc",
          8136 => x"53",
          8137 => x"fc",
          8138 => x"e4",
          8139 => x"d5",
          8140 => x"fe",
          8141 => x"33",
          8142 => x"f6",
          8143 => x"08",
          8144 => x"27",
          8145 => x"15",
          8146 => x"2a",
          8147 => x"51",
          8148 => x"83",
          8149 => x"94",
          8150 => x"80",
          8151 => x"0c",
          8152 => x"2e",
          8153 => x"79",
          8154 => x"70",
          8155 => x"51",
          8156 => x"2e",
          8157 => x"52",
          8158 => x"fe",
          8159 => x"82",
          8160 => x"ff",
          8161 => x"70",
          8162 => x"fe",
          8163 => x"82",
          8164 => x"73",
          8165 => x"76",
          8166 => x"06",
          8167 => x"0c",
          8168 => x"98",
          8169 => x"58",
          8170 => x"39",
          8171 => x"54",
          8172 => x"73",
          8173 => x"ff",
          8174 => x"82",
          8175 => x"54",
          8176 => x"08",
          8177 => x"9d",
          8178 => x"e4",
          8179 => x"81",
          8180 => x"d5",
          8181 => x"16",
          8182 => x"16",
          8183 => x"2e",
          8184 => x"76",
          8185 => x"de",
          8186 => x"31",
          8187 => x"18",
          8188 => x"90",
          8189 => x"81",
          8190 => x"06",
          8191 => x"56",
          8192 => x"9b",
          8193 => x"74",
          8194 => x"81",
          8195 => x"e4",
          8196 => x"d5",
          8197 => x"38",
          8198 => x"08",
          8199 => x"73",
          8200 => x"ff",
          8201 => x"82",
          8202 => x"54",
          8203 => x"bf",
          8204 => x"27",
          8205 => x"53",
          8206 => x"08",
          8207 => x"73",
          8208 => x"ff",
          8209 => x"15",
          8210 => x"16",
          8211 => x"ff",
          8212 => x"80",
          8213 => x"73",
          8214 => x"ff",
          8215 => x"82",
          8216 => x"94",
          8217 => x"91",
          8218 => x"53",
          8219 => x"81",
          8220 => x"34",
          8221 => x"39",
          8222 => x"82",
          8223 => x"05",
          8224 => x"08",
          8225 => x"08",
          8226 => x"38",
          8227 => x"0c",
          8228 => x"80",
          8229 => x"72",
          8230 => x"73",
          8231 => x"53",
          8232 => x"8c",
          8233 => x"16",
          8234 => x"38",
          8235 => x"0c",
          8236 => x"82",
          8237 => x"8b",
          8238 => x"f9",
          8239 => x"56",
          8240 => x"80",
          8241 => x"38",
          8242 => x"3d",
          8243 => x"8a",
          8244 => x"51",
          8245 => x"82",
          8246 => x"55",
          8247 => x"08",
          8248 => x"77",
          8249 => x"52",
          8250 => x"dd",
          8251 => x"e4",
          8252 => x"d5",
          8253 => x"c4",
          8254 => x"33",
          8255 => x"55",
          8256 => x"24",
          8257 => x"16",
          8258 => x"2a",
          8259 => x"51",
          8260 => x"80",
          8261 => x"9c",
          8262 => x"77",
          8263 => x"3f",
          8264 => x"08",
          8265 => x"77",
          8266 => x"22",
          8267 => x"74",
          8268 => x"ff",
          8269 => x"82",
          8270 => x"55",
          8271 => x"09",
          8272 => x"38",
          8273 => x"39",
          8274 => x"84",
          8275 => x"0c",
          8276 => x"82",
          8277 => x"89",
          8278 => x"fc",
          8279 => x"87",
          8280 => x"53",
          8281 => x"e7",
          8282 => x"d5",
          8283 => x"38",
          8284 => x"08",
          8285 => x"3d",
          8286 => x"3d",
          8287 => x"89",
          8288 => x"54",
          8289 => x"54",
          8290 => x"82",
          8291 => x"53",
          8292 => x"08",
          8293 => x"74",
          8294 => x"d5",
          8295 => x"73",
          8296 => x"fc",
          8297 => x"e4",
          8298 => x"cb",
          8299 => x"e4",
          8300 => x"51",
          8301 => x"82",
          8302 => x"53",
          8303 => x"08",
          8304 => x"81",
          8305 => x"80",
          8306 => x"82",
          8307 => x"a7",
          8308 => x"73",
          8309 => x"3f",
          8310 => x"51",
          8311 => x"3f",
          8312 => x"08",
          8313 => x"30",
          8314 => x"9f",
          8315 => x"d5",
          8316 => x"51",
          8317 => x"72",
          8318 => x"0c",
          8319 => x"04",
          8320 => x"66",
          8321 => x"89",
          8322 => x"97",
          8323 => x"de",
          8324 => x"d5",
          8325 => x"82",
          8326 => x"b2",
          8327 => x"75",
          8328 => x"3f",
          8329 => x"08",
          8330 => x"e4",
          8331 => x"02",
          8332 => x"33",
          8333 => x"55",
          8334 => x"25",
          8335 => x"55",
          8336 => x"80",
          8337 => x"76",
          8338 => x"ce",
          8339 => x"82",
          8340 => x"95",
          8341 => x"f0",
          8342 => x"65",
          8343 => x"53",
          8344 => x"05",
          8345 => x"51",
          8346 => x"82",
          8347 => x"5b",
          8348 => x"08",
          8349 => x"7c",
          8350 => x"08",
          8351 => x"fe",
          8352 => x"08",
          8353 => x"55",
          8354 => x"91",
          8355 => x"0c",
          8356 => x"81",
          8357 => x"39",
          8358 => x"c9",
          8359 => x"e4",
          8360 => x"55",
          8361 => x"2e",
          8362 => x"80",
          8363 => x"75",
          8364 => x"52",
          8365 => x"05",
          8366 => x"f5",
          8367 => x"e4",
          8368 => x"cf",
          8369 => x"e4",
          8370 => x"cc",
          8371 => x"e4",
          8372 => x"82",
          8373 => x"07",
          8374 => x"05",
          8375 => x"53",
          8376 => x"9c",
          8377 => x"26",
          8378 => x"f9",
          8379 => x"08",
          8380 => x"08",
          8381 => x"98",
          8382 => x"81",
          8383 => x"58",
          8384 => x"3f",
          8385 => x"08",
          8386 => x"e4",
          8387 => x"38",
          8388 => x"77",
          8389 => x"5d",
          8390 => x"74",
          8391 => x"81",
          8392 => x"b8",
          8393 => x"a9",
          8394 => x"d5",
          8395 => x"ff",
          8396 => x"30",
          8397 => x"1b",
          8398 => x"5b",
          8399 => x"39",
          8400 => x"ff",
          8401 => x"82",
          8402 => x"f0",
          8403 => x"30",
          8404 => x"1b",
          8405 => x"5b",
          8406 => x"83",
          8407 => x"58",
          8408 => x"92",
          8409 => x"0c",
          8410 => x"12",
          8411 => x"33",
          8412 => x"54",
          8413 => x"34",
          8414 => x"e4",
          8415 => x"0d",
          8416 => x"0d",
          8417 => x"fc",
          8418 => x"52",
          8419 => x"3f",
          8420 => x"08",
          8421 => x"e4",
          8422 => x"38",
          8423 => x"56",
          8424 => x"38",
          8425 => x"70",
          8426 => x"81",
          8427 => x"55",
          8428 => x"80",
          8429 => x"38",
          8430 => x"54",
          8431 => x"08",
          8432 => x"38",
          8433 => x"82",
          8434 => x"53",
          8435 => x"52",
          8436 => x"b2",
          8437 => x"d5",
          8438 => x"88",
          8439 => x"80",
          8440 => x"17",
          8441 => x"51",
          8442 => x"3f",
          8443 => x"08",
          8444 => x"81",
          8445 => x"81",
          8446 => x"e4",
          8447 => x"09",
          8448 => x"38",
          8449 => x"39",
          8450 => x"77",
          8451 => x"e4",
          8452 => x"08",
          8453 => x"98",
          8454 => x"82",
          8455 => x"52",
          8456 => x"b1",
          8457 => x"d5",
          8458 => x"94",
          8459 => x"18",
          8460 => x"33",
          8461 => x"54",
          8462 => x"34",
          8463 => x"85",
          8464 => x"18",
          8465 => x"74",
          8466 => x"0c",
          8467 => x"04",
          8468 => x"82",
          8469 => x"ff",
          8470 => x"a3",
          8471 => x"cf",
          8472 => x"e4",
          8473 => x"d5",
          8474 => x"f9",
          8475 => x"a3",
          8476 => x"96",
          8477 => x"58",
          8478 => x"82",
          8479 => x"55",
          8480 => x"08",
          8481 => x"02",
          8482 => x"33",
          8483 => x"70",
          8484 => x"55",
          8485 => x"73",
          8486 => x"75",
          8487 => x"80",
          8488 => x"c1",
          8489 => x"da",
          8490 => x"81",
          8491 => x"87",
          8492 => x"b1",
          8493 => x"78",
          8494 => x"c3",
          8495 => x"e4",
          8496 => x"2a",
          8497 => x"51",
          8498 => x"80",
          8499 => x"38",
          8500 => x"d5",
          8501 => x"15",
          8502 => x"89",
          8503 => x"82",
          8504 => x"5c",
          8505 => x"3d",
          8506 => x"ff",
          8507 => x"82",
          8508 => x"55",
          8509 => x"08",
          8510 => x"82",
          8511 => x"52",
          8512 => x"bb",
          8513 => x"d5",
          8514 => x"82",
          8515 => x"86",
          8516 => x"80",
          8517 => x"d5",
          8518 => x"2e",
          8519 => x"d5",
          8520 => x"c1",
          8521 => x"c7",
          8522 => x"d5",
          8523 => x"d5",
          8524 => x"70",
          8525 => x"08",
          8526 => x"51",
          8527 => x"80",
          8528 => x"73",
          8529 => x"38",
          8530 => x"52",
          8531 => x"af",
          8532 => x"d5",
          8533 => x"74",
          8534 => x"51",
          8535 => x"3f",
          8536 => x"08",
          8537 => x"d5",
          8538 => x"3d",
          8539 => x"3d",
          8540 => x"9a",
          8541 => x"05",
          8542 => x"51",
          8543 => x"82",
          8544 => x"54",
          8545 => x"08",
          8546 => x"78",
          8547 => x"8e",
          8548 => x"58",
          8549 => x"82",
          8550 => x"54",
          8551 => x"08",
          8552 => x"54",
          8553 => x"82",
          8554 => x"84",
          8555 => x"06",
          8556 => x"02",
          8557 => x"33",
          8558 => x"81",
          8559 => x"86",
          8560 => x"fd",
          8561 => x"74",
          8562 => x"70",
          8563 => x"af",
          8564 => x"d5",
          8565 => x"55",
          8566 => x"e4",
          8567 => x"87",
          8568 => x"e4",
          8569 => x"09",
          8570 => x"38",
          8571 => x"d5",
          8572 => x"2e",
          8573 => x"86",
          8574 => x"81",
          8575 => x"81",
          8576 => x"d5",
          8577 => x"78",
          8578 => x"9c",
          8579 => x"e4",
          8580 => x"d5",
          8581 => x"9f",
          8582 => x"a0",
          8583 => x"51",
          8584 => x"3f",
          8585 => x"0b",
          8586 => x"78",
          8587 => x"80",
          8588 => x"82",
          8589 => x"52",
          8590 => x"51",
          8591 => x"3f",
          8592 => x"b8",
          8593 => x"ff",
          8594 => x"a0",
          8595 => x"11",
          8596 => x"05",
          8597 => x"ee",
          8598 => x"ae",
          8599 => x"15",
          8600 => x"78",
          8601 => x"53",
          8602 => x"cc",
          8603 => x"81",
          8604 => x"34",
          8605 => x"bf",
          8606 => x"d5",
          8607 => x"82",
          8608 => x"b3",
          8609 => x"b2",
          8610 => x"96",
          8611 => x"a3",
          8612 => x"53",
          8613 => x"51",
          8614 => x"3f",
          8615 => x"0b",
          8616 => x"78",
          8617 => x"83",
          8618 => x"51",
          8619 => x"3f",
          8620 => x"08",
          8621 => x"80",
          8622 => x"76",
          8623 => x"a1",
          8624 => x"d5",
          8625 => x"3d",
          8626 => x"3d",
          8627 => x"84",
          8628 => x"d0",
          8629 => x"aa",
          8630 => x"05",
          8631 => x"51",
          8632 => x"82",
          8633 => x"55",
          8634 => x"08",
          8635 => x"78",
          8636 => x"08",
          8637 => x"70",
          8638 => x"cd",
          8639 => x"e4",
          8640 => x"d5",
          8641 => x"be",
          8642 => x"9f",
          8643 => x"a0",
          8644 => x"55",
          8645 => x"38",
          8646 => x"3d",
          8647 => x"3d",
          8648 => x"51",
          8649 => x"3f",
          8650 => x"52",
          8651 => x"52",
          8652 => x"92",
          8653 => x"08",
          8654 => x"c8",
          8655 => x"d5",
          8656 => x"82",
          8657 => x"97",
          8658 => x"3d",
          8659 => x"81",
          8660 => x"65",
          8661 => x"2e",
          8662 => x"55",
          8663 => x"82",
          8664 => x"84",
          8665 => x"06",
          8666 => x"73",
          8667 => x"92",
          8668 => x"e4",
          8669 => x"d5",
          8670 => x"ca",
          8671 => x"93",
          8672 => x"ff",
          8673 => x"8d",
          8674 => x"a1",
          8675 => x"af",
          8676 => x"17",
          8677 => x"33",
          8678 => x"70",
          8679 => x"55",
          8680 => x"38",
          8681 => x"54",
          8682 => x"34",
          8683 => x"0b",
          8684 => x"8b",
          8685 => x"84",
          8686 => x"06",
          8687 => x"73",
          8688 => x"e7",
          8689 => x"2e",
          8690 => x"75",
          8691 => x"ff",
          8692 => x"82",
          8693 => x"52",
          8694 => x"a5",
          8695 => x"55",
          8696 => x"08",
          8697 => x"de",
          8698 => x"e4",
          8699 => x"51",
          8700 => x"3f",
          8701 => x"08",
          8702 => x"11",
          8703 => x"82",
          8704 => x"80",
          8705 => x"16",
          8706 => x"ae",
          8707 => x"06",
          8708 => x"53",
          8709 => x"51",
          8710 => x"3f",
          8711 => x"0b",
          8712 => x"87",
          8713 => x"e4",
          8714 => x"77",
          8715 => x"3f",
          8716 => x"08",
          8717 => x"e4",
          8718 => x"78",
          8719 => x"98",
          8720 => x"e4",
          8721 => x"82",
          8722 => x"aa",
          8723 => x"ec",
          8724 => x"80",
          8725 => x"02",
          8726 => x"e3",
          8727 => x"57",
          8728 => x"3d",
          8729 => x"97",
          8730 => x"c3",
          8731 => x"e4",
          8732 => x"d5",
          8733 => x"cf",
          8734 => x"66",
          8735 => x"d0",
          8736 => x"c5",
          8737 => x"e4",
          8738 => x"d5",
          8739 => x"38",
          8740 => x"05",
          8741 => x"06",
          8742 => x"73",
          8743 => x"a7",
          8744 => x"09",
          8745 => x"71",
          8746 => x"06",
          8747 => x"55",
          8748 => x"15",
          8749 => x"81",
          8750 => x"34",
          8751 => x"a2",
          8752 => x"d5",
          8753 => x"74",
          8754 => x"0c",
          8755 => x"04",
          8756 => x"65",
          8757 => x"94",
          8758 => x"52",
          8759 => x"d0",
          8760 => x"d5",
          8761 => x"82",
          8762 => x"80",
          8763 => x"58",
          8764 => x"3d",
          8765 => x"c4",
          8766 => x"d5",
          8767 => x"82",
          8768 => x"b4",
          8769 => x"c7",
          8770 => x"a0",
          8771 => x"55",
          8772 => x"84",
          8773 => x"17",
          8774 => x"2b",
          8775 => x"96",
          8776 => x"9d",
          8777 => x"54",
          8778 => x"15",
          8779 => x"ff",
          8780 => x"82",
          8781 => x"55",
          8782 => x"e4",
          8783 => x"0d",
          8784 => x"0d",
          8785 => x"5a",
          8786 => x"3d",
          8787 => x"9a",
          8788 => x"db",
          8789 => x"e4",
          8790 => x"e4",
          8791 => x"82",
          8792 => x"07",
          8793 => x"55",
          8794 => x"2e",
          8795 => x"81",
          8796 => x"55",
          8797 => x"2e",
          8798 => x"7b",
          8799 => x"80",
          8800 => x"70",
          8801 => x"ac",
          8802 => x"d5",
          8803 => x"82",
          8804 => x"80",
          8805 => x"52",
          8806 => x"b1",
          8807 => x"d5",
          8808 => x"82",
          8809 => x"bf",
          8810 => x"e4",
          8811 => x"e4",
          8812 => x"59",
          8813 => x"81",
          8814 => x"56",
          8815 => x"33",
          8816 => x"16",
          8817 => x"27",
          8818 => x"56",
          8819 => x"80",
          8820 => x"80",
          8821 => x"ff",
          8822 => x"70",
          8823 => x"56",
          8824 => x"e8",
          8825 => x"76",
          8826 => x"81",
          8827 => x"80",
          8828 => x"57",
          8829 => x"78",
          8830 => x"51",
          8831 => x"2e",
          8832 => x"73",
          8833 => x"38",
          8834 => x"08",
          8835 => x"9f",
          8836 => x"d5",
          8837 => x"82",
          8838 => x"a7",
          8839 => x"33",
          8840 => x"c3",
          8841 => x"2e",
          8842 => x"e4",
          8843 => x"2e",
          8844 => x"56",
          8845 => x"05",
          8846 => x"92",
          8847 => x"e4",
          8848 => x"76",
          8849 => x"0c",
          8850 => x"04",
          8851 => x"82",
          8852 => x"ff",
          8853 => x"9d",
          8854 => x"d3",
          8855 => x"e4",
          8856 => x"e4",
          8857 => x"82",
          8858 => x"82",
          8859 => x"53",
          8860 => x"3d",
          8861 => x"ff",
          8862 => x"73",
          8863 => x"51",
          8864 => x"74",
          8865 => x"38",
          8866 => x"3d",
          8867 => x"cc",
          8868 => x"e4",
          8869 => x"ff",
          8870 => x"38",
          8871 => x"08",
          8872 => x"3f",
          8873 => x"82",
          8874 => x"51",
          8875 => x"82",
          8876 => x"83",
          8877 => x"55",
          8878 => x"a3",
          8879 => x"82",
          8880 => x"ff",
          8881 => x"82",
          8882 => x"93",
          8883 => x"75",
          8884 => x"75",
          8885 => x"38",
          8886 => x"76",
          8887 => x"86",
          8888 => x"39",
          8889 => x"27",
          8890 => x"88",
          8891 => x"77",
          8892 => x"59",
          8893 => x"56",
          8894 => x"81",
          8895 => x"81",
          8896 => x"33",
          8897 => x"73",
          8898 => x"fe",
          8899 => x"33",
          8900 => x"73",
          8901 => x"81",
          8902 => x"80",
          8903 => x"02",
          8904 => x"75",
          8905 => x"51",
          8906 => x"2e",
          8907 => x"87",
          8908 => x"56",
          8909 => x"78",
          8910 => x"80",
          8911 => x"70",
          8912 => x"a8",
          8913 => x"d5",
          8914 => x"82",
          8915 => x"80",
          8916 => x"52",
          8917 => x"ae",
          8918 => x"d5",
          8919 => x"82",
          8920 => x"8d",
          8921 => x"c4",
          8922 => x"e5",
          8923 => x"c6",
          8924 => x"e4",
          8925 => x"09",
          8926 => x"cc",
          8927 => x"75",
          8928 => x"c4",
          8929 => x"74",
          8930 => x"d8",
          8931 => x"e4",
          8932 => x"d5",
          8933 => x"38",
          8934 => x"d5",
          8935 => x"66",
          8936 => x"c5",
          8937 => x"88",
          8938 => x"34",
          8939 => x"52",
          8940 => x"99",
          8941 => x"54",
          8942 => x"15",
          8943 => x"ff",
          8944 => x"82",
          8945 => x"54",
          8946 => x"82",
          8947 => x"9c",
          8948 => x"f2",
          8949 => x"62",
          8950 => x"80",
          8951 => x"93",
          8952 => x"55",
          8953 => x"5e",
          8954 => x"3f",
          8955 => x"08",
          8956 => x"e4",
          8957 => x"38",
          8958 => x"58",
          8959 => x"38",
          8960 => x"97",
          8961 => x"08",
          8962 => x"38",
          8963 => x"70",
          8964 => x"81",
          8965 => x"55",
          8966 => x"87",
          8967 => x"39",
          8968 => x"90",
          8969 => x"82",
          8970 => x"8a",
          8971 => x"89",
          8972 => x"7f",
          8973 => x"56",
          8974 => x"3f",
          8975 => x"06",
          8976 => x"72",
          8977 => x"82",
          8978 => x"05",
          8979 => x"7c",
          8980 => x"55",
          8981 => x"27",
          8982 => x"16",
          8983 => x"83",
          8984 => x"76",
          8985 => x"80",
          8986 => x"79",
          8987 => x"c1",
          8988 => x"7f",
          8989 => x"14",
          8990 => x"83",
          8991 => x"82",
          8992 => x"81",
          8993 => x"38",
          8994 => x"08",
          8995 => x"95",
          8996 => x"e4",
          8997 => x"81",
          8998 => x"7b",
          8999 => x"06",
          9000 => x"39",
          9001 => x"56",
          9002 => x"09",
          9003 => x"b9",
          9004 => x"80",
          9005 => x"80",
          9006 => x"78",
          9007 => x"7a",
          9008 => x"38",
          9009 => x"73",
          9010 => x"81",
          9011 => x"ff",
          9012 => x"74",
          9013 => x"ff",
          9014 => x"82",
          9015 => x"58",
          9016 => x"08",
          9017 => x"74",
          9018 => x"16",
          9019 => x"73",
          9020 => x"39",
          9021 => x"7e",
          9022 => x"0c",
          9023 => x"2e",
          9024 => x"88",
          9025 => x"8c",
          9026 => x"1a",
          9027 => x"07",
          9028 => x"1b",
          9029 => x"08",
          9030 => x"16",
          9031 => x"75",
          9032 => x"38",
          9033 => x"94",
          9034 => x"15",
          9035 => x"54",
          9036 => x"34",
          9037 => x"82",
          9038 => x"90",
          9039 => x"e8",
          9040 => x"6e",
          9041 => x"80",
          9042 => x"9e",
          9043 => x"5c",
          9044 => x"3f",
          9045 => x"0b",
          9046 => x"08",
          9047 => x"38",
          9048 => x"08",
          9049 => x"ed",
          9050 => x"08",
          9051 => x"80",
          9052 => x"80",
          9053 => x"d5",
          9054 => x"d5",
          9055 => x"82",
          9056 => x"33",
          9057 => x"12",
          9058 => x"55",
          9059 => x"51",
          9060 => x"3f",
          9061 => x"08",
          9062 => x"70",
          9063 => x"57",
          9064 => x"8c",
          9065 => x"82",
          9066 => x"06",
          9067 => x"56",
          9068 => x"38",
          9069 => x"05",
          9070 => x"7f",
          9071 => x"cc",
          9072 => x"e4",
          9073 => x"68",
          9074 => x"2e",
          9075 => x"82",
          9076 => x"8b",
          9077 => x"75",
          9078 => x"80",
          9079 => x"81",
          9080 => x"2e",
          9081 => x"80",
          9082 => x"38",
          9083 => x"0a",
          9084 => x"ff",
          9085 => x"55",
          9086 => x"86",
          9087 => x"8b",
          9088 => x"89",
          9089 => x"2a",
          9090 => x"77",
          9091 => x"59",
          9092 => x"81",
          9093 => x"70",
          9094 => x"07",
          9095 => x"56",
          9096 => x"38",
          9097 => x"80",
          9098 => x"54",
          9099 => x"52",
          9100 => x"8e",
          9101 => x"56",
          9102 => x"08",
          9103 => x"83",
          9104 => x"ff",
          9105 => x"82",
          9106 => x"83",
          9107 => x"55",
          9108 => x"82",
          9109 => x"09",
          9110 => x"a3",
          9111 => x"29",
          9112 => x"11",
          9113 => x"74",
          9114 => x"93",
          9115 => x"17",
          9116 => x"da",
          9117 => x"e4",
          9118 => x"18",
          9119 => x"92",
          9120 => x"d5",
          9121 => x"b7",
          9122 => x"f8",
          9123 => x"52",
          9124 => x"90",
          9125 => x"56",
          9126 => x"08",
          9127 => x"62",
          9128 => x"77",
          9129 => x"e4",
          9130 => x"55",
          9131 => x"bf",
          9132 => x"8e",
          9133 => x"26",
          9134 => x"74",
          9135 => x"8e",
          9136 => x"68",
          9137 => x"38",
          9138 => x"81",
          9139 => x"af",
          9140 => x"2a",
          9141 => x"56",
          9142 => x"2e",
          9143 => x"87",
          9144 => x"82",
          9145 => x"38",
          9146 => x"55",
          9147 => x"83",
          9148 => x"81",
          9149 => x"56",
          9150 => x"80",
          9151 => x"38",
          9152 => x"83",
          9153 => x"06",
          9154 => x"78",
          9155 => x"91",
          9156 => x"0b",
          9157 => x"22",
          9158 => x"80",
          9159 => x"74",
          9160 => x"38",
          9161 => x"56",
          9162 => x"17",
          9163 => x"57",
          9164 => x"2e",
          9165 => x"75",
          9166 => x"79",
          9167 => x"fe",
          9168 => x"82",
          9169 => x"84",
          9170 => x"05",
          9171 => x"5e",
          9172 => x"80",
          9173 => x"e4",
          9174 => x"8a",
          9175 => x"fd",
          9176 => x"75",
          9177 => x"38",
          9178 => x"78",
          9179 => x"8c",
          9180 => x"0b",
          9181 => x"22",
          9182 => x"80",
          9183 => x"74",
          9184 => x"38",
          9185 => x"56",
          9186 => x"17",
          9187 => x"57",
          9188 => x"2e",
          9189 => x"75",
          9190 => x"79",
          9191 => x"fe",
          9192 => x"82",
          9193 => x"10",
          9194 => x"82",
          9195 => x"9f",
          9196 => x"38",
          9197 => x"d5",
          9198 => x"82",
          9199 => x"05",
          9200 => x"2a",
          9201 => x"56",
          9202 => x"17",
          9203 => x"81",
          9204 => x"7b",
          9205 => x"67",
          9206 => x"12",
          9207 => x"30",
          9208 => x"74",
          9209 => x"59",
          9210 => x"7d",
          9211 => x"81",
          9212 => x"76",
          9213 => x"42",
          9214 => x"76",
          9215 => x"90",
          9216 => x"60",
          9217 => x"51",
          9218 => x"26",
          9219 => x"75",
          9220 => x"31",
          9221 => x"67",
          9222 => x"fe",
          9223 => x"82",
          9224 => x"58",
          9225 => x"09",
          9226 => x"38",
          9227 => x"08",
          9228 => x"26",
          9229 => x"78",
          9230 => x"79",
          9231 => x"78",
          9232 => x"87",
          9233 => x"82",
          9234 => x"06",
          9235 => x"83",
          9236 => x"82",
          9237 => x"27",
          9238 => x"8f",
          9239 => x"55",
          9240 => x"26",
          9241 => x"59",
          9242 => x"63",
          9243 => x"74",
          9244 => x"38",
          9245 => x"88",
          9246 => x"e4",
          9247 => x"26",
          9248 => x"86",
          9249 => x"1a",
          9250 => x"79",
          9251 => x"38",
          9252 => x"80",
          9253 => x"2e",
          9254 => x"83",
          9255 => x"9f",
          9256 => x"8b",
          9257 => x"06",
          9258 => x"74",
          9259 => x"84",
          9260 => x"52",
          9261 => x"8f",
          9262 => x"53",
          9263 => x"52",
          9264 => x"8f",
          9265 => x"80",
          9266 => x"51",
          9267 => x"3f",
          9268 => x"34",
          9269 => x"ff",
          9270 => x"1b",
          9271 => x"99",
          9272 => x"90",
          9273 => x"83",
          9274 => x"70",
          9275 => x"80",
          9276 => x"55",
          9277 => x"ff",
          9278 => x"67",
          9279 => x"ff",
          9280 => x"38",
          9281 => x"ff",
          9282 => x"1b",
          9283 => x"e9",
          9284 => x"74",
          9285 => x"51",
          9286 => x"3f",
          9287 => x"1c",
          9288 => x"98",
          9289 => x"8d",
          9290 => x"ff",
          9291 => x"51",
          9292 => x"3f",
          9293 => x"1b",
          9294 => x"db",
          9295 => x"2e",
          9296 => x"80",
          9297 => x"88",
          9298 => x"80",
          9299 => x"ff",
          9300 => x"7c",
          9301 => x"51",
          9302 => x"3f",
          9303 => x"1b",
          9304 => x"b3",
          9305 => x"b0",
          9306 => x"8d",
          9307 => x"52",
          9308 => x"ff",
          9309 => x"ff",
          9310 => x"c0",
          9311 => x"0b",
          9312 => x"34",
          9313 => x"c7",
          9314 => x"c7",
          9315 => x"39",
          9316 => x"0a",
          9317 => x"51",
          9318 => x"3f",
          9319 => x"ff",
          9320 => x"1b",
          9321 => x"d1",
          9322 => x"0b",
          9323 => x"a9",
          9324 => x"34",
          9325 => x"c7",
          9326 => x"1b",
          9327 => x"86",
          9328 => x"d5",
          9329 => x"1b",
          9330 => x"ff",
          9331 => x"81",
          9332 => x"7a",
          9333 => x"ff",
          9334 => x"81",
          9335 => x"e4",
          9336 => x"38",
          9337 => x"09",
          9338 => x"ec",
          9339 => x"86",
          9340 => x"52",
          9341 => x"88",
          9342 => x"80",
          9343 => x"7a",
          9344 => x"e5",
          9345 => x"85",
          9346 => x"7a",
          9347 => x"87",
          9348 => x"85",
          9349 => x"83",
          9350 => x"ff",
          9351 => x"ff",
          9352 => x"e8",
          9353 => x"8b",
          9354 => x"52",
          9355 => x"51",
          9356 => x"3f",
          9357 => x"52",
          9358 => x"8b",
          9359 => x"54",
          9360 => x"7a",
          9361 => x"ff",
          9362 => x"75",
          9363 => x"53",
          9364 => x"51",
          9365 => x"3f",
          9366 => x"52",
          9367 => x"8c",
          9368 => x"56",
          9369 => x"83",
          9370 => x"06",
          9371 => x"52",
          9372 => x"8b",
          9373 => x"52",
          9374 => x"ff",
          9375 => x"f0",
          9376 => x"1b",
          9377 => x"87",
          9378 => x"55",
          9379 => x"83",
          9380 => x"74",
          9381 => x"ff",
          9382 => x"7c",
          9383 => x"74",
          9384 => x"38",
          9385 => x"54",
          9386 => x"52",
          9387 => x"86",
          9388 => x"d5",
          9389 => x"be",
          9390 => x"53",
          9391 => x"08",
          9392 => x"ff",
          9393 => x"76",
          9394 => x"31",
          9395 => x"cd",
          9396 => x"58",
          9397 => x"ff",
          9398 => x"55",
          9399 => x"83",
          9400 => x"61",
          9401 => x"26",
          9402 => x"57",
          9403 => x"53",
          9404 => x"51",
          9405 => x"3f",
          9406 => x"08",
          9407 => x"76",
          9408 => x"31",
          9409 => x"db",
          9410 => x"7d",
          9411 => x"38",
          9412 => x"83",
          9413 => x"8a",
          9414 => x"7d",
          9415 => x"38",
          9416 => x"80",
          9417 => x"81",
          9418 => x"7a",
          9419 => x"ff",
          9420 => x"81",
          9421 => x"e4",
          9422 => x"38",
          9423 => x"1b",
          9424 => x"b2",
          9425 => x"54",
          9426 => x"08",
          9427 => x"7f",
          9428 => x"d4",
          9429 => x"39",
          9430 => x"81",
          9431 => x"80",
          9432 => x"80",
          9433 => x"7a",
          9434 => x"fd",
          9435 => x"d5",
          9436 => x"ff",
          9437 => x"83",
          9438 => x"77",
          9439 => x"0b",
          9440 => x"81",
          9441 => x"34",
          9442 => x"34",
          9443 => x"34",
          9444 => x"80",
          9445 => x"75",
          9446 => x"95",
          9447 => x"85",
          9448 => x"d5",
          9449 => x"2a",
          9450 => x"75",
          9451 => x"82",
          9452 => x"87",
          9453 => x"52",
          9454 => x"51",
          9455 => x"3f",
          9456 => x"ca",
          9457 => x"88",
          9458 => x"54",
          9459 => x"52",
          9460 => x"84",
          9461 => x"56",
          9462 => x"08",
          9463 => x"53",
          9464 => x"51",
          9465 => x"3f",
          9466 => x"d5",
          9467 => x"38",
          9468 => x"56",
          9469 => x"56",
          9470 => x"d5",
          9471 => x"75",
          9472 => x"0c",
          9473 => x"04",
          9474 => x"7d",
          9475 => x"80",
          9476 => x"05",
          9477 => x"76",
          9478 => x"38",
          9479 => x"11",
          9480 => x"53",
          9481 => x"79",
          9482 => x"3f",
          9483 => x"09",
          9484 => x"38",
          9485 => x"55",
          9486 => x"db",
          9487 => x"70",
          9488 => x"34",
          9489 => x"74",
          9490 => x"81",
          9491 => x"80",
          9492 => x"55",
          9493 => x"76",
          9494 => x"d5",
          9495 => x"3d",
          9496 => x"3d",
          9497 => x"84",
          9498 => x"33",
          9499 => x"8a",
          9500 => x"06",
          9501 => x"52",
          9502 => x"3f",
          9503 => x"56",
          9504 => x"be",
          9505 => x"08",
          9506 => x"05",
          9507 => x"75",
          9508 => x"56",
          9509 => x"a1",
          9510 => x"fc",
          9511 => x"53",
          9512 => x"76",
          9513 => x"97",
          9514 => x"32",
          9515 => x"72",
          9516 => x"70",
          9517 => x"56",
          9518 => x"18",
          9519 => x"88",
          9520 => x"3d",
          9521 => x"3d",
          9522 => x"11",
          9523 => x"80",
          9524 => x"38",
          9525 => x"05",
          9526 => x"8c",
          9527 => x"08",
          9528 => x"3f",
          9529 => x"08",
          9530 => x"16",
          9531 => x"09",
          9532 => x"38",
          9533 => x"55",
          9534 => x"55",
          9535 => x"e4",
          9536 => x"0d",
          9537 => x"0d",
          9538 => x"cc",
          9539 => x"73",
          9540 => x"d5",
          9541 => x"0c",
          9542 => x"04",
          9543 => x"02",
          9544 => x"33",
          9545 => x"3d",
          9546 => x"54",
          9547 => x"52",
          9548 => x"ae",
          9549 => x"ff",
          9550 => x"3d",
          9551 => x"3d",
          9552 => x"84",
          9553 => x"22",
          9554 => x"52",
          9555 => x"26",
          9556 => x"83",
          9557 => x"52",
          9558 => x"83",
          9559 => x"27",
          9560 => x"b5",
          9561 => x"06",
          9562 => x"80",
          9563 => x"82",
          9564 => x"51",
          9565 => x"9c",
          9566 => x"70",
          9567 => x"06",
          9568 => x"80",
          9569 => x"38",
          9570 => x"c9",
          9571 => x"22",
          9572 => x"39",
          9573 => x"70",
          9574 => x"53",
          9575 => x"d5",
          9576 => x"3d",
          9577 => x"3d",
          9578 => x"05",
          9579 => x"05",
          9580 => x"53",
          9581 => x"70",
          9582 => x"85",
          9583 => x"9a",
          9584 => x"b5",
          9585 => x"06",
          9586 => x"81",
          9587 => x"38",
          9588 => x"c7",
          9589 => x"22",
          9590 => x"82",
          9591 => x"84",
          9592 => x"fb",
          9593 => x"51",
          9594 => x"ff",
          9595 => x"38",
          9596 => x"ff",
          9597 => x"a8",
          9598 => x"ff",
          9599 => x"38",
          9600 => x"56",
          9601 => x"05",
          9602 => x"30",
          9603 => x"72",
          9604 => x"51",
          9605 => x"80",
          9606 => x"70",
          9607 => x"22",
          9608 => x"71",
          9609 => x"70",
          9610 => x"55",
          9611 => x"25",
          9612 => x"73",
          9613 => x"dc",
          9614 => x"29",
          9615 => x"05",
          9616 => x"04",
          9617 => x"10",
          9618 => x"22",
          9619 => x"80",
          9620 => x"75",
          9621 => x"72",
          9622 => x"51",
          9623 => x"12",
          9624 => x"e0",
          9625 => x"39",
          9626 => x"95",
          9627 => x"51",
          9628 => x"12",
          9629 => x"ff",
          9630 => x"85",
          9631 => x"12",
          9632 => x"ff",
          9633 => x"8c",
          9634 => x"f8",
          9635 => x"16",
          9636 => x"39",
          9637 => x"82",
          9638 => x"87",
          9639 => x"00",
          9640 => x"ff",
          9641 => x"ff",
          9642 => x"ff",
          9643 => x"00",
          9644 => x"00",
          9645 => x"00",
          9646 => x"00",
          9647 => x"00",
          9648 => x"00",
          9649 => x"00",
          9650 => x"00",
          9651 => x"00",
          9652 => x"00",
          9653 => x"00",
          9654 => x"00",
          9655 => x"00",
          9656 => x"00",
          9657 => x"00",
          9658 => x"00",
          9659 => x"00",
          9660 => x"00",
          9661 => x"00",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"00",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"00",
          9683 => x"00",
          9684 => x"00",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"00",
          9787 => x"00",
          9788 => x"64",
          9789 => x"74",
          9790 => x"64",
          9791 => x"74",
          9792 => x"66",
          9793 => x"74",
          9794 => x"66",
          9795 => x"64",
          9796 => x"66",
          9797 => x"63",
          9798 => x"6d",
          9799 => x"61",
          9800 => x"6d",
          9801 => x"79",
          9802 => x"6d",
          9803 => x"66",
          9804 => x"6d",
          9805 => x"70",
          9806 => x"6d",
          9807 => x"6d",
          9808 => x"6d",
          9809 => x"68",
          9810 => x"68",
          9811 => x"68",
          9812 => x"68",
          9813 => x"63",
          9814 => x"00",
          9815 => x"6a",
          9816 => x"72",
          9817 => x"61",
          9818 => x"72",
          9819 => x"74",
          9820 => x"69",
          9821 => x"00",
          9822 => x"74",
          9823 => x"00",
          9824 => x"74",
          9825 => x"69",
          9826 => x"6d",
          9827 => x"69",
          9828 => x"6b",
          9829 => x"00",
          9830 => x"65",
          9831 => x"44",
          9832 => x"20",
          9833 => x"6f",
          9834 => x"49",
          9835 => x"72",
          9836 => x"20",
          9837 => x"6f",
          9838 => x"44",
          9839 => x"20",
          9840 => x"20",
          9841 => x"64",
          9842 => x"4e",
          9843 => x"69",
          9844 => x"66",
          9845 => x"64",
          9846 => x"4e",
          9847 => x"61",
          9848 => x"66",
          9849 => x"64",
          9850 => x"49",
          9851 => x"6c",
          9852 => x"66",
          9853 => x"6e",
          9854 => x"2e",
          9855 => x"41",
          9856 => x"73",
          9857 => x"65",
          9858 => x"64",
          9859 => x"46",
          9860 => x"20",
          9861 => x"65",
          9862 => x"20",
          9863 => x"73",
          9864 => x"00",
          9865 => x"46",
          9866 => x"20",
          9867 => x"64",
          9868 => x"69",
          9869 => x"6c",
          9870 => x"00",
          9871 => x"53",
          9872 => x"73",
          9873 => x"69",
          9874 => x"70",
          9875 => x"65",
          9876 => x"64",
          9877 => x"44",
          9878 => x"65",
          9879 => x"6d",
          9880 => x"20",
          9881 => x"69",
          9882 => x"6c",
          9883 => x"00",
          9884 => x"44",
          9885 => x"20",
          9886 => x"20",
          9887 => x"62",
          9888 => x"2e",
          9889 => x"4e",
          9890 => x"6f",
          9891 => x"74",
          9892 => x"65",
          9893 => x"6c",
          9894 => x"73",
          9895 => x"20",
          9896 => x"6e",
          9897 => x"6e",
          9898 => x"73",
          9899 => x"46",
          9900 => x"61",
          9901 => x"62",
          9902 => x"65",
          9903 => x"54",
          9904 => x"6f",
          9905 => x"20",
          9906 => x"72",
          9907 => x"6f",
          9908 => x"61",
          9909 => x"6c",
          9910 => x"2e",
          9911 => x"46",
          9912 => x"20",
          9913 => x"6c",
          9914 => x"65",
          9915 => x"49",
          9916 => x"66",
          9917 => x"69",
          9918 => x"20",
          9919 => x"6f",
          9920 => x"00",
          9921 => x"54",
          9922 => x"6d",
          9923 => x"20",
          9924 => x"6e",
          9925 => x"6c",
          9926 => x"00",
          9927 => x"50",
          9928 => x"6d",
          9929 => x"72",
          9930 => x"6e",
          9931 => x"72",
          9932 => x"2e",
          9933 => x"53",
          9934 => x"65",
          9935 => x"00",
          9936 => x"55",
          9937 => x"6f",
          9938 => x"65",
          9939 => x"72",
          9940 => x"0a",
          9941 => x"20",
          9942 => x"65",
          9943 => x"73",
          9944 => x"20",
          9945 => x"20",
          9946 => x"65",
          9947 => x"65",
          9948 => x"00",
          9949 => x"72",
          9950 => x"00",
          9951 => x"25",
          9952 => x"58",
          9953 => x"3a",
          9954 => x"25",
          9955 => x"00",
          9956 => x"20",
          9957 => x"20",
          9958 => x"00",
          9959 => x"25",
          9960 => x"00",
          9961 => x"20",
          9962 => x"20",
          9963 => x"7c",
          9964 => x"7a",
          9965 => x"0a",
          9966 => x"25",
          9967 => x"00",
          9968 => x"31",
          9969 => x"32",
          9970 => x"32",
          9971 => x"76",
          9972 => x"62",
          9973 => x"20",
          9974 => x"2c",
          9975 => x"76",
          9976 => x"32",
          9977 => x"25",
          9978 => x"73",
          9979 => x"0a",
          9980 => x"5a",
          9981 => x"49",
          9982 => x"72",
          9983 => x"74",
          9984 => x"6e",
          9985 => x"72",
          9986 => x"54",
          9987 => x"72",
          9988 => x"74",
          9989 => x"75",
          9990 => x"50",
          9991 => x"69",
          9992 => x"72",
          9993 => x"74",
          9994 => x"49",
          9995 => x"4c",
          9996 => x"20",
          9997 => x"65",
          9998 => x"70",
          9999 => x"49",
         10000 => x"4c",
         10001 => x"20",
         10002 => x"65",
         10003 => x"70",
         10004 => x"55",
         10005 => x"30",
         10006 => x"20",
         10007 => x"65",
         10008 => x"70",
         10009 => x"55",
         10010 => x"30",
         10011 => x"20",
         10012 => x"65",
         10013 => x"70",
         10014 => x"55",
         10015 => x"31",
         10016 => x"20",
         10017 => x"65",
         10018 => x"70",
         10019 => x"55",
         10020 => x"31",
         10021 => x"20",
         10022 => x"65",
         10023 => x"70",
         10024 => x"53",
         10025 => x"69",
         10026 => x"75",
         10027 => x"69",
         10028 => x"2e",
         10029 => x"45",
         10030 => x"6c",
         10031 => x"20",
         10032 => x"65",
         10033 => x"2e",
         10034 => x"61",
         10035 => x"65",
         10036 => x"2e",
         10037 => x"00",
         10038 => x"7a",
         10039 => x"7a",
         10040 => x"68",
         10041 => x"30",
         10042 => x"46",
         10043 => x"65",
         10044 => x"6f",
         10045 => x"69",
         10046 => x"6c",
         10047 => x"20",
         10048 => x"63",
         10049 => x"20",
         10050 => x"70",
         10051 => x"73",
         10052 => x"6e",
         10053 => x"6d",
         10054 => x"61",
         10055 => x"2e",
         10056 => x"2a",
         10057 => x"43",
         10058 => x"72",
         10059 => x"2e",
         10060 => x"00",
         10061 => x"43",
         10062 => x"69",
         10063 => x"2e",
         10064 => x"43",
         10065 => x"61",
         10066 => x"67",
         10067 => x"00",
         10068 => x"25",
         10069 => x"78",
         10070 => x"38",
         10071 => x"3e",
         10072 => x"6c",
         10073 => x"30",
         10074 => x"0a",
         10075 => x"44",
         10076 => x"20",
         10077 => x"6f",
         10078 => x"0a",
         10079 => x"70",
         10080 => x"65",
         10081 => x"25",
         10082 => x"58",
         10083 => x"32",
         10084 => x"3f",
         10085 => x"25",
         10086 => x"58",
         10087 => x"34",
         10088 => x"25",
         10089 => x"58",
         10090 => x"38",
         10091 => x"00",
         10092 => x"45",
         10093 => x"75",
         10094 => x"67",
         10095 => x"64",
         10096 => x"20",
         10097 => x"6c",
         10098 => x"2e",
         10099 => x"43",
         10100 => x"69",
         10101 => x"63",
         10102 => x"20",
         10103 => x"30",
         10104 => x"20",
         10105 => x"0a",
         10106 => x"43",
         10107 => x"20",
         10108 => x"75",
         10109 => x"64",
         10110 => x"64",
         10111 => x"25",
         10112 => x"0a",
         10113 => x"52",
         10114 => x"61",
         10115 => x"6e",
         10116 => x"70",
         10117 => x"63",
         10118 => x"6f",
         10119 => x"2e",
         10120 => x"43",
         10121 => x"20",
         10122 => x"6f",
         10123 => x"6e",
         10124 => x"2e",
         10125 => x"5a",
         10126 => x"62",
         10127 => x"25",
         10128 => x"25",
         10129 => x"73",
         10130 => x"00",
         10131 => x"25",
         10132 => x"25",
         10133 => x"73",
         10134 => x"25",
         10135 => x"25",
         10136 => x"42",
         10137 => x"63",
         10138 => x"61",
         10139 => x"00",
         10140 => x"4d",
         10141 => x"72",
         10142 => x"78",
         10143 => x"73",
         10144 => x"2c",
         10145 => x"6e",
         10146 => x"20",
         10147 => x"63",
         10148 => x"20",
         10149 => x"6d",
         10150 => x"2e",
         10151 => x"52",
         10152 => x"69",
         10153 => x"2e",
         10154 => x"45",
         10155 => x"6c",
         10156 => x"20",
         10157 => x"65",
         10158 => x"70",
         10159 => x"2e",
         10160 => x"25",
         10161 => x"64",
         10162 => x"20",
         10163 => x"25",
         10164 => x"64",
         10165 => x"25",
         10166 => x"53",
         10167 => x"43",
         10168 => x"69",
         10169 => x"61",
         10170 => x"6e",
         10171 => x"20",
         10172 => x"6f",
         10173 => x"6f",
         10174 => x"6f",
         10175 => x"67",
         10176 => x"3a",
         10177 => x"76",
         10178 => x"73",
         10179 => x"70",
         10180 => x"65",
         10181 => x"64",
         10182 => x"20",
         10183 => x"57",
         10184 => x"44",
         10185 => x"20",
         10186 => x"30",
         10187 => x"25",
         10188 => x"29",
         10189 => x"20",
         10190 => x"53",
         10191 => x"4d",
         10192 => x"20",
         10193 => x"30",
         10194 => x"25",
         10195 => x"29",
         10196 => x"20",
         10197 => x"49",
         10198 => x"20",
         10199 => x"4d",
         10200 => x"30",
         10201 => x"25",
         10202 => x"29",
         10203 => x"20",
         10204 => x"42",
         10205 => x"20",
         10206 => x"20",
         10207 => x"30",
         10208 => x"25",
         10209 => x"29",
         10210 => x"20",
         10211 => x"52",
         10212 => x"20",
         10213 => x"20",
         10214 => x"30",
         10215 => x"25",
         10216 => x"29",
         10217 => x"20",
         10218 => x"53",
         10219 => x"41",
         10220 => x"20",
         10221 => x"65",
         10222 => x"65",
         10223 => x"25",
         10224 => x"29",
         10225 => x"20",
         10226 => x"54",
         10227 => x"52",
         10228 => x"20",
         10229 => x"69",
         10230 => x"73",
         10231 => x"25",
         10232 => x"29",
         10233 => x"20",
         10234 => x"49",
         10235 => x"20",
         10236 => x"4c",
         10237 => x"68",
         10238 => x"65",
         10239 => x"25",
         10240 => x"29",
         10241 => x"20",
         10242 => x"57",
         10243 => x"42",
         10244 => x"20",
         10245 => x"00",
         10246 => x"20",
         10247 => x"57",
         10248 => x"32",
         10249 => x"20",
         10250 => x"49",
         10251 => x"4c",
         10252 => x"20",
         10253 => x"50",
         10254 => x"20",
         10255 => x"53",
         10256 => x"41",
         10257 => x"65",
         10258 => x"73",
         10259 => x"20",
         10260 => x"43",
         10261 => x"52",
         10262 => x"74",
         10263 => x"63",
         10264 => x"20",
         10265 => x"72",
         10266 => x"20",
         10267 => x"30",
         10268 => x"00",
         10269 => x"20",
         10270 => x"43",
         10271 => x"4d",
         10272 => x"72",
         10273 => x"74",
         10274 => x"20",
         10275 => x"72",
         10276 => x"20",
         10277 => x"30",
         10278 => x"00",
         10279 => x"20",
         10280 => x"53",
         10281 => x"6b",
         10282 => x"61",
         10283 => x"41",
         10284 => x"65",
         10285 => x"20",
         10286 => x"20",
         10287 => x"30",
         10288 => x"00",
         10289 => x"4d",
         10290 => x"3a",
         10291 => x"20",
         10292 => x"5a",
         10293 => x"49",
         10294 => x"20",
         10295 => x"20",
         10296 => x"20",
         10297 => x"20",
         10298 => x"20",
         10299 => x"30",
         10300 => x"00",
         10301 => x"20",
         10302 => x"53",
         10303 => x"65",
         10304 => x"6c",
         10305 => x"20",
         10306 => x"71",
         10307 => x"20",
         10308 => x"20",
         10309 => x"64",
         10310 => x"34",
         10311 => x"7a",
         10312 => x"20",
         10313 => x"53",
         10314 => x"4d",
         10315 => x"6f",
         10316 => x"46",
         10317 => x"20",
         10318 => x"20",
         10319 => x"20",
         10320 => x"64",
         10321 => x"34",
         10322 => x"7a",
         10323 => x"20",
         10324 => x"57",
         10325 => x"62",
         10326 => x"20",
         10327 => x"41",
         10328 => x"6c",
         10329 => x"20",
         10330 => x"71",
         10331 => x"64",
         10332 => x"34",
         10333 => x"7a",
         10334 => x"53",
         10335 => x"6c",
         10336 => x"4d",
         10337 => x"75",
         10338 => x"46",
         10339 => x"00",
         10340 => x"45",
         10341 => x"45",
         10342 => x"00",
         10343 => x"55",
         10344 => x"6f",
         10345 => x"00",
         10346 => x"01",
         10347 => x"00",
         10348 => x"00",
         10349 => x"01",
         10350 => x"00",
         10351 => x"00",
         10352 => x"01",
         10353 => x"00",
         10354 => x"00",
         10355 => x"01",
         10356 => x"00",
         10357 => x"00",
         10358 => x"01",
         10359 => x"00",
         10360 => x"00",
         10361 => x"01",
         10362 => x"00",
         10363 => x"00",
         10364 => x"01",
         10365 => x"00",
         10366 => x"00",
         10367 => x"01",
         10368 => x"00",
         10369 => x"00",
         10370 => x"01",
         10371 => x"00",
         10372 => x"00",
         10373 => x"01",
         10374 => x"00",
         10375 => x"00",
         10376 => x"01",
         10377 => x"00",
         10378 => x"00",
         10379 => x"04",
         10380 => x"00",
         10381 => x"00",
         10382 => x"04",
         10383 => x"00",
         10384 => x"00",
         10385 => x"04",
         10386 => x"00",
         10387 => x"00",
         10388 => x"03",
         10389 => x"00",
         10390 => x"00",
         10391 => x"04",
         10392 => x"00",
         10393 => x"00",
         10394 => x"04",
         10395 => x"00",
         10396 => x"00",
         10397 => x"04",
         10398 => x"00",
         10399 => x"00",
         10400 => x"03",
         10401 => x"00",
         10402 => x"00",
         10403 => x"03",
         10404 => x"00",
         10405 => x"00",
         10406 => x"03",
         10407 => x"00",
         10408 => x"00",
         10409 => x"03",
         10410 => x"00",
         10411 => x"1b",
         10412 => x"1b",
         10413 => x"1b",
         10414 => x"1b",
         10415 => x"1b",
         10416 => x"1b",
         10417 => x"1b",
         10418 => x"1b",
         10419 => x"1b",
         10420 => x"1b",
         10421 => x"1b",
         10422 => x"10",
         10423 => x"0e",
         10424 => x"0d",
         10425 => x"0b",
         10426 => x"08",
         10427 => x"06",
         10428 => x"05",
         10429 => x"04",
         10430 => x"03",
         10431 => x"02",
         10432 => x"01",
         10433 => x"68",
         10434 => x"6f",
         10435 => x"68",
         10436 => x"00",
         10437 => x"21",
         10438 => x"25",
         10439 => x"75",
         10440 => x"73",
         10441 => x"46",
         10442 => x"65",
         10443 => x"6f",
         10444 => x"73",
         10445 => x"74",
         10446 => x"68",
         10447 => x"6f",
         10448 => x"66",
         10449 => x"20",
         10450 => x"45",
         10451 => x"00",
         10452 => x"43",
         10453 => x"6f",
         10454 => x"70",
         10455 => x"63",
         10456 => x"74",
         10457 => x"69",
         10458 => x"72",
         10459 => x"69",
         10460 => x"20",
         10461 => x"61",
         10462 => x"6e",
         10463 => x"53",
         10464 => x"22",
         10465 => x"3e",
         10466 => x"00",
         10467 => x"2b",
         10468 => x"5b",
         10469 => x"46",
         10470 => x"46",
         10471 => x"32",
         10472 => x"eb",
         10473 => x"53",
         10474 => x"35",
         10475 => x"4e",
         10476 => x"41",
         10477 => x"20",
         10478 => x"41",
         10479 => x"20",
         10480 => x"4e",
         10481 => x"41",
         10482 => x"20",
         10483 => x"41",
         10484 => x"20",
         10485 => x"00",
         10486 => x"00",
         10487 => x"00",
         10488 => x"00",
         10489 => x"01",
         10490 => x"09",
         10491 => x"14",
         10492 => x"1e",
         10493 => x"80",
         10494 => x"8e",
         10495 => x"45",
         10496 => x"49",
         10497 => x"90",
         10498 => x"99",
         10499 => x"59",
         10500 => x"9c",
         10501 => x"41",
         10502 => x"a5",
         10503 => x"a8",
         10504 => x"ac",
         10505 => x"b0",
         10506 => x"b4",
         10507 => x"b8",
         10508 => x"bc",
         10509 => x"c0",
         10510 => x"c4",
         10511 => x"c8",
         10512 => x"cc",
         10513 => x"d0",
         10514 => x"d4",
         10515 => x"d8",
         10516 => x"dc",
         10517 => x"e0",
         10518 => x"e4",
         10519 => x"e8",
         10520 => x"ec",
         10521 => x"f0",
         10522 => x"f4",
         10523 => x"f8",
         10524 => x"fc",
         10525 => x"2b",
         10526 => x"3d",
         10527 => x"5c",
         10528 => x"3c",
         10529 => x"7f",
         10530 => x"00",
         10531 => x"00",
         10532 => x"01",
         10533 => x"00",
         10534 => x"00",
         10535 => x"00",
         10536 => x"00",
         10537 => x"00",
         10538 => x"00",
         10539 => x"00",
         10540 => x"00",
         10541 => x"00",
         10542 => x"00",
         10543 => x"00",
         10544 => x"00",
         10545 => x"00",
         10546 => x"00",
         10547 => x"00",
         10548 => x"00",
         10549 => x"00",
         10550 => x"00",
         10551 => x"00",
         10552 => x"00",
         10553 => x"20",
         10554 => x"00",
         10555 => x"00",
         10556 => x"00",
         10557 => x"00",
         10558 => x"00",
         10559 => x"00",
         10560 => x"00",
         10561 => x"00",
         10562 => x"25",
         10563 => x"25",
         10564 => x"25",
         10565 => x"25",
         10566 => x"25",
         10567 => x"25",
         10568 => x"25",
         10569 => x"25",
         10570 => x"25",
         10571 => x"25",
         10572 => x"25",
         10573 => x"25",
         10574 => x"25",
         10575 => x"25",
         10576 => x"25",
         10577 => x"25",
         10578 => x"25",
         10579 => x"25",
         10580 => x"25",
         10581 => x"25",
         10582 => x"25",
         10583 => x"25",
         10584 => x"25",
         10585 => x"25",
         10586 => x"03",
         10587 => x"03",
         10588 => x"03",
         10589 => x"00",
         10590 => x"03",
         10591 => x"03",
         10592 => x"22",
         10593 => x"03",
         10594 => x"22",
         10595 => x"22",
         10596 => x"23",
         10597 => x"00",
         10598 => x"00",
         10599 => x"00",
         10600 => x"20",
         10601 => x"25",
         10602 => x"00",
         10603 => x"00",
         10604 => x"00",
         10605 => x"00",
         10606 => x"01",
         10607 => x"01",
         10608 => x"01",
         10609 => x"01",
         10610 => x"01",
         10611 => x"01",
         10612 => x"00",
         10613 => x"01",
         10614 => x"01",
         10615 => x"01",
         10616 => x"01",
         10617 => x"01",
         10618 => x"01",
         10619 => x"01",
         10620 => x"01",
         10621 => x"01",
         10622 => x"01",
         10623 => x"01",
         10624 => x"01",
         10625 => x"01",
         10626 => x"01",
         10627 => x"01",
         10628 => x"01",
         10629 => x"01",
         10630 => x"01",
         10631 => x"01",
         10632 => x"01",
         10633 => x"01",
         10634 => x"01",
         10635 => x"01",
         10636 => x"01",
         10637 => x"01",
         10638 => x"01",
         10639 => x"01",
         10640 => x"01",
         10641 => x"01",
         10642 => x"01",
         10643 => x"01",
         10644 => x"01",
         10645 => x"01",
         10646 => x"01",
         10647 => x"01",
         10648 => x"01",
         10649 => x"01",
         10650 => x"01",
         10651 => x"01",
         10652 => x"01",
         10653 => x"01",
         10654 => x"01",
         10655 => x"00",
         10656 => x"01",
         10657 => x"01",
         10658 => x"02",
         10659 => x"02",
         10660 => x"2c",
         10661 => x"02",
         10662 => x"2c",
         10663 => x"02",
         10664 => x"02",
         10665 => x"01",
         10666 => x"00",
         10667 => x"01",
         10668 => x"01",
         10669 => x"02",
         10670 => x"02",
         10671 => x"02",
         10672 => x"02",
         10673 => x"01",
         10674 => x"02",
         10675 => x"02",
         10676 => x"02",
         10677 => x"01",
         10678 => x"02",
         10679 => x"02",
         10680 => x"02",
         10681 => x"02",
         10682 => x"01",
         10683 => x"02",
         10684 => x"02",
         10685 => x"02",
         10686 => x"02",
         10687 => x"02",
         10688 => x"02",
         10689 => x"01",
         10690 => x"02",
         10691 => x"02",
         10692 => x"02",
         10693 => x"01",
         10694 => x"01",
         10695 => x"02",
         10696 => x"02",
         10697 => x"02",
         10698 => x"01",
         10699 => x"00",
         10700 => x"03",
         10701 => x"03",
         10702 => x"03",
         10703 => x"03",
         10704 => x"03",
         10705 => x"03",
         10706 => x"03",
         10707 => x"03",
         10708 => x"03",
         10709 => x"03",
         10710 => x"03",
         10711 => x"01",
         10712 => x"00",
         10713 => x"03",
         10714 => x"03",
         10715 => x"03",
         10716 => x"03",
         10717 => x"03",
         10718 => x"03",
         10719 => x"07",
         10720 => x"01",
         10721 => x"01",
         10722 => x"01",
         10723 => x"00",
         10724 => x"04",
         10725 => x"05",
         10726 => x"00",
         10727 => x"1d",
         10728 => x"2c",
         10729 => x"01",
         10730 => x"01",
         10731 => x"06",
         10732 => x"06",
         10733 => x"06",
         10734 => x"06",
         10735 => x"06",
         10736 => x"00",
         10737 => x"1f",
         10738 => x"1f",
         10739 => x"1f",
         10740 => x"1f",
         10741 => x"1f",
         10742 => x"1f",
         10743 => x"1f",
         10744 => x"1f",
         10745 => x"1f",
         10746 => x"1f",
         10747 => x"1f",
         10748 => x"1f",
         10749 => x"1f",
         10750 => x"1f",
         10751 => x"1f",
         10752 => x"1f",
         10753 => x"1f",
         10754 => x"1f",
         10755 => x"1f",
         10756 => x"1f",
         10757 => x"06",
         10758 => x"06",
         10759 => x"00",
         10760 => x"1f",
         10761 => x"1f",
         10762 => x"00",
         10763 => x"21",
         10764 => x"21",
         10765 => x"21",
         10766 => x"05",
         10767 => x"04",
         10768 => x"01",
         10769 => x"01",
         10770 => x"01",
         10771 => x"01",
         10772 => x"08",
         10773 => x"03",
         10774 => x"00",
         10775 => x"00",
         10776 => x"01",
         10777 => x"00",
         10778 => x"00",
         10779 => x"00",
         10780 => x"01",
         10781 => x"00",
         10782 => x"00",
         10783 => x"00",
         10784 => x"01",
         10785 => x"00",
         10786 => x"00",
         10787 => x"00",
         10788 => x"01",
         10789 => x"00",
         10790 => x"00",
         10791 => x"00",
         10792 => x"01",
         10793 => x"00",
         10794 => x"00",
         10795 => x"00",
         10796 => x"01",
         10797 => x"00",
         10798 => x"00",
         10799 => x"00",
         10800 => x"01",
         10801 => x"00",
         10802 => x"00",
         10803 => x"00",
         10804 => x"01",
         10805 => x"00",
         10806 => x"00",
         10807 => x"00",
         10808 => x"01",
         10809 => x"00",
         10810 => x"00",
         10811 => x"00",
         10812 => x"01",
         10813 => x"00",
         10814 => x"00",
         10815 => x"00",
         10816 => x"01",
         10817 => x"00",
         10818 => x"00",
         10819 => x"00",
         10820 => x"01",
         10821 => x"00",
         10822 => x"00",
         10823 => x"00",
         10824 => x"01",
         10825 => x"00",
         10826 => x"00",
         10827 => x"00",
         10828 => x"01",
         10829 => x"00",
         10830 => x"00",
         10831 => x"00",
         10832 => x"01",
         10833 => x"00",
         10834 => x"00",
         10835 => x"00",
         10836 => x"01",
         10837 => x"00",
         10838 => x"00",
         10839 => x"00",
         10840 => x"01",
         10841 => x"00",
         10842 => x"00",
         10843 => x"00",
         10844 => x"01",
         10845 => x"00",
         10846 => x"00",
         10847 => x"00",
         10848 => x"01",
         10849 => x"00",
         10850 => x"00",
         10851 => x"00",
         10852 => x"01",
         10853 => x"00",
         10854 => x"00",
         10855 => x"00",
         10856 => x"01",
         10857 => x"00",
         10858 => x"00",
         10859 => x"00",
         10860 => x"01",
         10861 => x"00",
         10862 => x"00",
         10863 => x"00",
         10864 => x"01",
         10865 => x"00",
         10866 => x"00",
         10867 => x"00",
         10868 => x"01",
         10869 => x"00",
         10870 => x"00",
         10871 => x"00",
         10872 => x"01",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"01",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"01",
         10889 => x"01",
         10890 => x"00",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"05",
         10895 => x"05",
         10896 => x"05",
         10897 => x"00",
         10898 => x"01",
         10899 => x"01",
         10900 => x"01",
         10901 => x"01",
         10902 => x"00",
         10903 => x"00",
         10904 => x"00",
         10905 => x"00",
         10906 => x"00",
         10907 => x"00",
         10908 => x"00",
         10909 => x"00",
         10910 => x"00",
         10911 => x"00",
         10912 => x"00",
         10913 => x"00",
         10914 => x"00",
         10915 => x"00",
         10916 => x"00",
         10917 => x"00",
         10918 => x"00",
         10919 => x"00",
         10920 => x"00",
         10921 => x"00",
         10922 => x"00",
         10923 => x"00",
         10924 => x"00",
         10925 => x"00",
         10926 => x"00",
         10927 => x"01",
         10928 => x"00",
         10929 => x"01",
         10930 => x"00",
         10931 => x"02",
         10932 => x"00",
         10933 => x"00",
         10934 => x"00",
         10935 => x"00",
         10936 => x"01",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"ad",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"f0",
           193 => x"f0",
           194 => x"f0",
           195 => x"08",
           196 => x"0c",
           197 => x"84",
           198 => x"af",
           199 => x"80",
           200 => x"ad",
           201 => x"90",
           202 => x"2d",
           203 => x"04",
           204 => x"2d",
           205 => x"04",
           206 => x"2d",
           207 => x"04",
           208 => x"82",
           209 => x"82",
           210 => x"d5",
           211 => x"d5",
           212 => x"f0",
           213 => x"f0",
           214 => x"f0",
           215 => x"f0",
           216 => x"f0",
           217 => x"f0",
           218 => x"f0",
           219 => x"f0",
           220 => x"f0",
           221 => x"f0",
           222 => x"f0",
           223 => x"f0",
           224 => x"f0",
           225 => x"f0",
           226 => x"f0",
           227 => x"f0",
           228 => x"f0",
           229 => x"f0",
           230 => x"f0",
           231 => x"f0",
           232 => x"f0",
           233 => x"f0",
           234 => x"f0",
           235 => x"f0",
           236 => x"f0",
           237 => x"f0",
           238 => x"f0",
           239 => x"f0",
           240 => x"f0",
           241 => x"f0",
           242 => x"f0",
           243 => x"f0",
           244 => x"f0",
           245 => x"f0",
           246 => x"f0",
           247 => x"f0",
           248 => x"f0",
           249 => x"f0",
           250 => x"f0",
           251 => x"f0",
           252 => x"f0",
           253 => x"f0",
           254 => x"f0",
           255 => x"f0",
           256 => x"f0",
           257 => x"f0",
           258 => x"f0",
           259 => x"f0",
           260 => x"f0",
           261 => x"f0",
           262 => x"f0",
           263 => x"f0",
           264 => x"f0",
           265 => x"f0",
           266 => x"f0",
           267 => x"f0",
           268 => x"f0",
           269 => x"f0",
           270 => x"f0",
           271 => x"f0",
           272 => x"f0",
           273 => x"f0",
           274 => x"f0",
           275 => x"f0",
           276 => x"f0",
           277 => x"f0",
           278 => x"f0",
           279 => x"f0",
           280 => x"f0",
           281 => x"f0",
           282 => x"f0",
           283 => x"f0",
           284 => x"f0",
           285 => x"f0",
           286 => x"f0",
           287 => x"f0",
           288 => x"f0",
           289 => x"f0",
           290 => x"f0",
           291 => x"f0",
           292 => x"f0",
           293 => x"f0",
           294 => x"f0",
           295 => x"f0",
           296 => x"f0",
           297 => x"f0",
           298 => x"f0",
           299 => x"00",
           300 => x"10",
           301 => x"10",
           302 => x"10",
           303 => x"10",
           304 => x"ff",
           305 => x"83",
           306 => x"fc",
           307 => x"80",
           308 => x"06",
           309 => x"0a",
           310 => x"51",
           311 => x"d0",
           312 => x"05",
           313 => x"04",
           314 => x"00",
           315 => x"f0",
           316 => x"08",
           317 => x"fc",
           318 => x"05",
           319 => x"05",
           320 => x"54",
           321 => x"70",
           322 => x"82",
           323 => x"82",
           324 => x"0d",
           325 => x"f0",
           326 => x"3d",
           327 => x"08",
           328 => x"81",
           329 => x"38",
           330 => x"05",
           331 => x"0b",
           332 => x"81",
           333 => x"05",
           334 => x"8c",
           335 => x"08",
           336 => x"88",
           337 => x"05",
           338 => x"08",
           339 => x"82",
           340 => x"80",
           341 => x"05",
           342 => x"e4",
           343 => x"05",
           344 => x"05",
           345 => x"38",
           346 => x"05",
           347 => x"08",
           348 => x"f8",
           349 => x"82",
           350 => x"05",
           351 => x"82",
           352 => x"05",
           353 => x"ff",
           354 => x"05",
           355 => x"f0",
           356 => x"f0",
           357 => x"f0",
           358 => x"0c",
           359 => x"04",
           360 => x"f0",
           361 => x"d5",
           362 => x"f0",
           363 => x"08",
           364 => x"d5",
           365 => x"f0",
           366 => x"08",
           367 => x"fc",
           368 => x"8c",
           369 => x"e0",
           370 => x"3f",
           371 => x"f0",
           372 => x"08",
           373 => x"88",
           374 => x"34",
           375 => x"70",
           376 => x"0d",
           377 => x"f0",
           378 => x"3d",
           379 => x"70",
           380 => x"82",
           381 => x"82",
           382 => x"82",
           383 => x"54",
           384 => x"82",
           385 => x"d5",
           386 => x"d5",
           387 => x"82",
           388 => x"08",
           389 => x"0d",
           390 => x"05",
           391 => x"08",
           392 => x"d5",
           393 => x"33",
           394 => x"81",
           395 => x"80",
           396 => x"f0",
           397 => x"82",
           398 => x"72",
           399 => x"f8",
           400 => x"72",
           401 => x"f0",
           402 => x"d5",
           403 => x"f0",
           404 => x"51",
           405 => x"82",
           406 => x"af",
           407 => x"f0",
           408 => x"26",
           409 => x"f8",
           410 => x"81",
           411 => x"08",
           412 => x"98",
           413 => x"82",
           414 => x"83",
           415 => x"51",
           416 => x"38",
           417 => x"70",
           418 => x"d5",
           419 => x"39",
           420 => x"70",
           421 => x"83",
           422 => x"51",
           423 => x"f0",
           424 => x"08",
           425 => x"08",
           426 => x"51",
           427 => x"e8",
           428 => x"05",
           429 => x"51",
           430 => x"80",
           431 => x"05",
           432 => x"22",
           433 => x"51",
           434 => x"f0",
           435 => x"70",
           436 => x"2c",
           437 => x"d5",
           438 => x"39",
           439 => x"70",
           440 => x"53",
           441 => x"f0",
           442 => x"70",
           443 => x"38",
           444 => x"05",
           445 => x"33",
           446 => x"05",
           447 => x"05",
           448 => x"82",
           449 => x"82",
           450 => x"51",
           451 => x"f0",
           452 => x"51",
           453 => x"05",
           454 => x"22",
           455 => x"d5",
           456 => x"39",
           457 => x"70",
           458 => x"d5",
           459 => x"39",
           460 => x"70",
           461 => x"d5",
           462 => x"39",
           463 => x"70",
           464 => x"f0",
           465 => x"d5",
           466 => x"39",
           467 => x"70",
           468 => x"f0",
           469 => x"bf",
           470 => x"34",
           471 => x"ff",
           472 => x"08",
           473 => x"d5",
           474 => x"39",
           475 => x"82",
           476 => x"05",
           477 => x"70",
           478 => x"08",
           479 => x"ec",
           480 => x"82",
           481 => x"ef",
           482 => x"08",
           483 => x"84",
           484 => x"0c",
           485 => x"05",
           486 => x"22",
           487 => x"51",
           488 => x"82",
           489 => x"98",
           490 => x"d5",
           491 => x"a4",
           492 => x"72",
           493 => x"99",
           494 => x"08",
           495 => x"08",
           496 => x"05",
           497 => x"22",
           498 => x"22",
           499 => x"d5",
           500 => x"39",
           501 => x"82",
           502 => x"05",
           503 => x"70",
           504 => x"0c",
           505 => x"70",
           506 => x"51",
           507 => x"d5",
           508 => x"2b",
           509 => x"f0",
           510 => x"ec",
           511 => x"82",
           512 => x"39",
           513 => x"51",
           514 => x"53",
           515 => x"23",
           516 => x"53",
           517 => x"73",
           518 => x"f0",
           519 => x"82",
           520 => x"82",
           521 => x"72",
           522 => x"08",
           523 => x"90",
           524 => x"08",
           525 => x"f0",
           526 => x"82",
           527 => x"d5",
           528 => x"82",
           529 => x"08",
           530 => x"53",
           531 => x"82",
           532 => x"d5",
           533 => x"a4",
           534 => x"22",
           535 => x"d5",
           536 => x"f0",
           537 => x"f0",
           538 => x"08",
           539 => x"51",
           540 => x"05",
           541 => x"d5",
           542 => x"82",
           543 => x"80",
           544 => x"f0",
           545 => x"82",
           546 => x"0b",
           547 => x"82",
           548 => x"82",
           549 => x"72",
           550 => x"08",
           551 => x"90",
           552 => x"08",
           553 => x"f0",
           554 => x"82",
           555 => x"d5",
           556 => x"82",
           557 => x"08",
           558 => x"53",
           559 => x"82",
           560 => x"d5",
           561 => x"06",
           562 => x"e4",
           563 => x"d5",
           564 => x"f0",
           565 => x"08",
           566 => x"fc",
           567 => x"54",
           568 => x"08",
           569 => x"08",
           570 => x"d4",
           571 => x"05",
           572 => x"27",
           573 => x"05",
           574 => x"f0",
           575 => x"11",
           576 => x"08",
           577 => x"f0",
           578 => x"b0",
           579 => x"08",
           580 => x"d4",
           581 => x"d0",
           582 => x"08",
           583 => x"f0",
           584 => x"08",
           585 => x"f0",
           586 => x"d6",
           587 => x"d5",
           588 => x"d5",
           589 => x"84",
           590 => x"08",
           591 => x"55",
           592 => x"53",
           593 => x"34",
           594 => x"70",
           595 => x"94",
           596 => x"22",
           597 => x"f0",
           598 => x"08",
           599 => x"81",
           600 => x"80",
           601 => x"05",
           602 => x"08",
           603 => x"cc",
           604 => x"08",
           605 => x"f4",
           606 => x"09",
           607 => x"08",
           608 => x"82",
           609 => x"39",
           610 => x"ff",
           611 => x"c8",
           612 => x"05",
           613 => x"23",
           614 => x"70",
           615 => x"53",
           616 => x"d5",
           617 => x"2b",
           618 => x"fc",
           619 => x"74",
           620 => x"e4",
           621 => x"72",
           622 => x"9d",
           623 => x"33",
           624 => x"33",
           625 => x"d5",
           626 => x"f0",
           627 => x"70",
           628 => x"2e",
           629 => x"05",
           630 => x"70",
           631 => x"51",
           632 => x"08",
           633 => x"53",
           634 => x"23",
           635 => x"05",
           636 => x"70",
           637 => x"51",
           638 => x"08",
           639 => x"53",
           640 => x"23",
           641 => x"70",
           642 => x"38",
           643 => x"ff",
           644 => x"08",
           645 => x"90",
           646 => x"38",
           647 => x"52",
           648 => x"82",
           649 => x"81",
           650 => x"72",
           651 => x"08",
           652 => x"ca",
           653 => x"08",
           654 => x"81",
           655 => x"90",
           656 => x"08",
           657 => x"39",
           658 => x"70",
           659 => x"53",
           660 => x"f0",
           661 => x"8a",
           662 => x"05",
           663 => x"51",
           664 => x"82",
           665 => x"b0",
           666 => x"08",
           667 => x"09",
           668 => x"08",
           669 => x"08",
           670 => x"82",
           671 => x"88",
           672 => x"72",
           673 => x"08",
           674 => x"72",
           675 => x"73",
           676 => x"80",
           677 => x"08",
           678 => x"fa",
           679 => x"e4",
           680 => x"06",
           681 => x"38",
           682 => x"ff",
           683 => x"08",
           684 => x"98",
           685 => x"38",
           686 => x"52",
           687 => x"82",
           688 => x"87",
           689 => x"72",
           690 => x"05",
           691 => x"d5",
           692 => x"2b",
           693 => x"25",
           694 => x"05",
           695 => x"d2",
           696 => x"33",
           697 => x"06",
           698 => x"05",
           699 => x"05",
           700 => x"39",
           701 => x"53",
           702 => x"80",
           703 => x"05",
           704 => x"d5",
           705 => x"ff",
           706 => x"2e",
           707 => x"88",
           708 => x"fc",
           709 => x"f0",
           710 => x"d5",
           711 => x"f2",
           712 => x"08",
           713 => x"2e",
           714 => x"d5",
           715 => x"51",
           716 => x"05",
           717 => x"72",
           718 => x"82",
           719 => x"82",
           720 => x"33",
           721 => x"f0",
           722 => x"d5",
           723 => x"39",
           724 => x"82",
           725 => x"f0",
           726 => x"f0",
           727 => x"d5",
           728 => x"f0",
           729 => x"53",
           730 => x"f0",
           731 => x"70",
           732 => x"2e",
           733 => x"ec",
           734 => x"82",
           735 => x"90",
           736 => x"73",
           737 => x"88",
           738 => x"3f",
           739 => x"05",
           740 => x"05",
           741 => x"82",
           742 => x"b7",
           743 => x"33",
           744 => x"a8",
           745 => x"e4",
           746 => x"08",
           747 => x"f0",
           748 => x"d5",
           749 => x"39",
           750 => x"52",
           751 => x"51",
           752 => x"d5",
           753 => x"08",
           754 => x"0c",
           755 => x"05",
           756 => x"0d",
           757 => x"f0",
           758 => x"3d",
           759 => x"d5",
           760 => x"d5",
           761 => x"dd",
           762 => x"d5",
           763 => x"d5",
           764 => x"02",
           765 => x"80",
           766 => x"0c",
           767 => x"70",
           768 => x"06",
           769 => x"2e",
           770 => x"08",
           771 => x"d5",
           772 => x"33",
           773 => x"81",
           774 => x"0c",
           775 => x"05",
           776 => x"80",
           777 => x"82",
           778 => x"08",
           779 => x"51",
           780 => x"53",
           781 => x"0b",
           782 => x"ff",
           783 => x"f1",
           784 => x"13",
           785 => x"08",
           786 => x"0b",
           787 => x"82",
           788 => x"82",
           789 => x"82",
           790 => x"d5",
           791 => x"f0",
           792 => x"82",
           793 => x"0b",
           794 => x"82",
           795 => x"11",
           796 => x"70",
           797 => x"72",
           798 => x"d5",
           799 => x"39",
           800 => x"53",
           801 => x"05",
           802 => x"88",
           803 => x"08",
           804 => x"53",
           805 => x"f0",
           806 => x"08",
           807 => x"08",
           808 => x"51",
           809 => x"53",
           810 => x"0b",
           811 => x"ff",
           812 => x"05",
           813 => x"05",
           814 => x"05",
           815 => x"0d",
           816 => x"f0",
           817 => x"3d",
           818 => x"d5",
           819 => x"3f",
           820 => x"e4",
           821 => x"f0",
           822 => x"82",
           823 => x"d5",
           824 => x"33",
           825 => x"81",
           826 => x"80",
           827 => x"f0",
           828 => x"82",
           829 => x"11",
           830 => x"51",
           831 => x"db",
           832 => x"08",
           833 => x"54",
           834 => x"25",
           835 => x"05",
           836 => x"08",
           837 => x"72",
           838 => x"0c",
           839 => x"8c",
           840 => x"82",
           841 => x"82",
           842 => x"53",
           843 => x"8c",
           844 => x"05",
           845 => x"05",
           846 => x"12",
           847 => x"d5",
           848 => x"d5",
           849 => x"08",
           850 => x"f0",
           851 => x"f0",
           852 => x"39",
           853 => x"05",
           854 => x"08",
           855 => x"82",
           856 => x"08",
           857 => x"0d",
           858 => x"85",
           859 => x"06",
           860 => x"8d",
           861 => x"f8",
           862 => x"f0",
           863 => x"70",
           864 => x"51",
           865 => x"82",
           866 => x"d5",
           867 => x"85",
           868 => x"52",
           869 => x"08",
           870 => x"05",
           871 => x"88",
           872 => x"d5",
           873 => x"52",
           874 => x"88",
           875 => x"2a",
           876 => x"71",
           877 => x"f0",
           878 => x"33",
           879 => x"51",
           880 => x"08",
           881 => x"05",
           882 => x"08",
           883 => x"07",
           884 => x"0b",
           885 => x"81",
           886 => x"05",
           887 => x"52",
           888 => x"88",
           889 => x"05",
           890 => x"71",
           891 => x"d5",
           892 => x"d5",
           893 => x"80",
           894 => x"05",
           895 => x"0c",
           896 => x"85",
           897 => x"05",
           898 => x"05",
           899 => x"38",
           900 => x"90",
           901 => x"ec",
           902 => x"08",
           903 => x"82",
           904 => x"d5",
           905 => x"d5",
           906 => x"34",
           907 => x"05",
           908 => x"88",
           909 => x"8c",
           910 => x"05",
           911 => x"d5",
           912 => x"52",
           913 => x"82",
           914 => x"d5",
           915 => x"02",
           916 => x"82",
           917 => x"d5",
           918 => x"f0",
           919 => x"08",
           920 => x"90",
           921 => x"82",
           922 => x"d5",
           923 => x"ac",
           924 => x"08",
           925 => x"05",
           926 => x"08",
           927 => x"f0",
           928 => x"08",
           929 => x"08",
           930 => x"f8",
           931 => x"05",
           932 => x"05",
           933 => x"08",
           934 => x"05",
           935 => x"08",
           936 => x"05",
           937 => x"08",
           938 => x"f0",
           939 => x"d5",
           940 => x"f0",
           941 => x"d5",
           942 => x"f0",
           943 => x"08",
           944 => x"71",
           945 => x"08",
           946 => x"f0",
           947 => x"08",
           948 => x"f0",
           949 => x"08",
           950 => x"82",
           951 => x"70",
           952 => x"08",
           953 => x"05",
           954 => x"08",
           955 => x"f0",
           956 => x"d5",
           957 => x"39",
           958 => x"70",
           959 => x"0d",
           960 => x"f0",
           961 => x"3d",
           962 => x"08",
           963 => x"82",
           964 => x"71",
           965 => x"08",
           966 => x"05",
           967 => x"70",
           968 => x"d5",
           969 => x"82",
           970 => x"d5",
           971 => x"f0",
           972 => x"d5",
           973 => x"d5",
           974 => x"02",
           975 => x"82",
           976 => x"d5",
           977 => x"f0",
           978 => x"82",
           979 => x"05",
           980 => x"82",
           981 => x"51",
           982 => x"fc",
           983 => x"08",
           984 => x"51",
           985 => x"39",
           986 => x"70",
           987 => x"0d",
           988 => x"f0",
           989 => x"3d",
           990 => x"08",
           991 => x"82",
           992 => x"d5",
           993 => x"f0",
           994 => x"e5",
           995 => x"08",
           996 => x"05",
           997 => x"08",
           998 => x"05",
           999 => x"08",
          1000 => x"08",
          1001 => x"d5",
          1002 => x"82",
          1003 => x"d5",
          1004 => x"71",
          1005 => x"05",
          1006 => x"fc",
          1007 => x"f0",
          1008 => x"e4",
          1009 => x"f0",
          1010 => x"82",
          1011 => x"d5",
          1012 => x"81",
          1013 => x"05",
          1014 => x"08",
          1015 => x"f0",
          1016 => x"08",
          1017 => x"ff",
          1018 => x"2e",
          1019 => x"f0",
          1020 => x"82",
          1021 => x"05",
          1022 => x"70",
          1023 => x"38",
          1024 => x"05",
          1025 => x"08",
          1026 => x"f0",
          1027 => x"08",
          1028 => x"ff",
          1029 => x"05",
          1030 => x"d5",
          1031 => x"52",
          1032 => x"d5",
          1033 => x"39",
          1034 => x"ff",
          1035 => x"0c",
          1036 => x"70",
          1037 => x"0b",
          1038 => x"ae",
          1039 => x"08",
          1040 => x"05",
          1041 => x"82",
          1042 => x"55",
          1043 => x"82",
          1044 => x"d5",
          1045 => x"e4",
          1046 => x"0c",
          1047 => x"d5",
          1048 => x"f0",
          1049 => x"f0",
          1050 => x"3f",
          1051 => x"f0",
          1052 => x"08",
          1053 => x"51",
          1054 => x"e4",
          1055 => x"05",
          1056 => x"05",
          1057 => x"f0",
          1058 => x"d5",
          1059 => x"f0",
          1060 => x"74",
          1061 => x"08",
          1062 => x"08",
          1063 => x"08",
          1064 => x"08",
          1065 => x"0c",
          1066 => x"08",
          1067 => x"82",
          1068 => x"08",
          1069 => x"0d",
          1070 => x"82",
          1071 => x"d5",
          1072 => x"80",
          1073 => x"0c",
          1074 => x"f8",
          1075 => x"f0",
          1076 => x"d5",
          1077 => x"ff",
          1078 => x"38",
          1079 => x"ff",
          1080 => x"0c",
          1081 => x"ff",
          1082 => x"d5",
          1083 => x"82",
          1084 => x"d5",
          1085 => x"f0",
          1086 => x"d5",
          1087 => x"d5",
          1088 => x"e4",
          1089 => x"0c",
          1090 => x"d5",
          1091 => x"f0",
          1092 => x"08",
          1093 => x"90",
          1094 => x"82",
          1095 => x"05",
          1096 => x"82",
          1097 => x"05",
          1098 => x"82",
          1099 => x"2e",
          1100 => x"05",
          1101 => x"fc",
          1102 => x"82",
          1103 => x"05",
          1104 => x"ff",
          1105 => x"05",
          1106 => x"84",
          1107 => x"82",
          1108 => x"0c",
          1109 => x"f0",
          1110 => x"08",
          1111 => x"82",
          1112 => x"82",
          1113 => x"0b",
          1114 => x"82",
          1115 => x"38",
          1116 => x"05",
          1117 => x"08",
          1118 => x"82",
          1119 => x"25",
          1120 => x"05",
          1121 => x"05",
          1122 => x"f0",
          1123 => x"05",
          1124 => x"f0",
          1125 => x"08",
          1126 => x"fc",
          1127 => x"08",
          1128 => x"08",
          1129 => x"82",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"82",
          1134 => x"d5",
          1135 => x"d5",
          1136 => x"d5",
          1137 => x"02",
          1138 => x"80",
          1139 => x"0c",
          1140 => x"80",
          1141 => x"88",
          1142 => x"88",
          1143 => x"08",
          1144 => x"8c",
          1145 => x"d5",
          1146 => x"d5",
          1147 => x"82",
          1148 => x"82",
          1149 => x"81",
          1150 => x"82",
          1151 => x"82",
          1152 => x"2e",
          1153 => x"05",
          1154 => x"05",
          1155 => x"08",
          1156 => x"3d",
          1157 => x"d5",
          1158 => x"fd",
          1159 => x"08",
          1160 => x"08",
          1161 => x"82",
          1162 => x"0c",
          1163 => x"0c",
          1164 => x"d5",
          1165 => x"82",
          1166 => x"82",
          1167 => x"93",
          1168 => x"d5",
          1169 => x"d5",
          1170 => x"02",
          1171 => x"81",
          1172 => x"0c",
          1173 => x"05",
          1174 => x"08",
          1175 => x"27",
          1176 => x"05",
          1177 => x"82",
          1178 => x"a2",
          1179 => x"08",
          1180 => x"0c",
          1181 => x"10",
          1182 => x"ff",
          1183 => x"05",
          1184 => x"d5",
          1185 => x"f0",
          1186 => x"82",
          1187 => x"d5",
          1188 => x"d5",
          1189 => x"f0",
          1190 => x"08",
          1191 => x"08",
          1192 => x"fc",
          1193 => x"08",
          1194 => x"8c",
          1195 => x"08",
          1196 => x"d5",
          1197 => x"93",
          1198 => x"08",
          1199 => x"0c",
          1200 => x"f8",
          1201 => x"f4",
          1202 => x"f4",
          1203 => x"3d",
          1204 => x"d5",
          1205 => x"f7",
          1206 => x"08",
          1207 => x"8c",
          1208 => x"d5",
          1209 => x"51",
          1210 => x"f0",
          1211 => x"06",
          1212 => x"91",
          1213 => x"08",
          1214 => x"ce",
          1215 => x"33",
          1216 => x"a4",
          1217 => x"f0",
          1218 => x"05",
          1219 => x"70",
          1220 => x"f0",
          1221 => x"08",
          1222 => x"09",
          1223 => x"f0",
          1224 => x"05",
          1225 => x"33",
          1226 => x"82",
          1227 => x"d5",
          1228 => x"f0",
          1229 => x"b6",
          1230 => x"08",
          1231 => x"39",
          1232 => x"05",
          1233 => x"08",
          1234 => x"08",
          1235 => x"08",
          1236 => x"0b",
          1237 => x"82",
          1238 => x"08",
          1239 => x"53",
          1240 => x"05",
          1241 => x"08",
          1242 => x"8d",
          1243 => x"ec",
          1244 => x"f0",
          1245 => x"27",
          1246 => x"05",
          1247 => x"8d",
          1248 => x"ec",
          1249 => x"82",
          1250 => x"39",
          1251 => x"53",
          1252 => x"f0",
          1253 => x"26",
          1254 => x"d5",
          1255 => x"39",
          1256 => x"05",
          1257 => x"fc",
          1258 => x"05",
          1259 => x"38",
          1260 => x"53",
          1261 => x"d5",
          1262 => x"51",
          1263 => x"05",
          1264 => x"33",
          1265 => x"f0",
          1266 => x"08",
          1267 => x"ad",
          1268 => x"33",
          1269 => x"f0",
          1270 => x"08",
          1271 => x"8d",
          1272 => x"ec",
          1273 => x"f0",
          1274 => x"08",
          1275 => x"26",
          1276 => x"08",
          1277 => x"d5",
          1278 => x"d5",
          1279 => x"d5",
          1280 => x"82",
          1281 => x"d5",
          1282 => x"81",
          1283 => x"52",
          1284 => x"08",
          1285 => x"d5",
          1286 => x"80",
          1287 => x"fc",
          1288 => x"fc",
          1289 => x"05",
          1290 => x"08",
          1291 => x"f0",
          1292 => x"08",
          1293 => x"8b",
          1294 => x"82",
          1295 => x"0c",
          1296 => x"f0",
          1297 => x"08",
          1298 => x"82",
          1299 => x"08",
          1300 => x"d5",
          1301 => x"ff",
          1302 => x"06",
          1303 => x"05",
          1304 => x"53",
          1305 => x"05",
          1306 => x"06",
          1307 => x"08",
          1308 => x"88",
          1309 => x"0c",
          1310 => x"d5",
          1311 => x"f0",
          1312 => x"2e",
          1313 => x"d5",
          1314 => x"81",
          1315 => x"72",
          1316 => x"34",
          1317 => x"82",
          1318 => x"d5",
          1319 => x"2e",
          1320 => x"05",
          1321 => x"cd",
          1322 => x"f4",
          1323 => x"05",
          1324 => x"70",
          1325 => x"f0",
          1326 => x"82",
          1327 => x"34",
          1328 => x"70",
          1329 => x"51",
          1330 => x"f8",
          1331 => x"f0",
          1332 => x"26",
          1333 => x"08",
          1334 => x"d5",
          1335 => x"73",
          1336 => x"f8",
          1337 => x"38",
          1338 => x"08",
          1339 => x"0b",
          1340 => x"b2",
          1341 => x"33",
          1342 => x"d5",
          1343 => x"b9",
          1344 => x"82",
          1345 => x"a5",
          1346 => x"f4",
          1347 => x"08",
          1348 => x"f8",
          1349 => x"cf",
          1350 => x"33",
          1351 => x"82",
          1352 => x"11",
          1353 => x"f8",
          1354 => x"05",
          1355 => x"d5",
          1356 => x"f0",
          1357 => x"27",
          1358 => x"05",
          1359 => x"d5",
          1360 => x"f0",
          1361 => x"26",
          1362 => x"08",
          1363 => x"d5",
          1364 => x"f0",
          1365 => x"74",
          1366 => x"f0",
          1367 => x"82",
          1368 => x"82",
          1369 => x"82",
          1370 => x"12",
          1371 => x"82",
          1372 => x"08",
          1373 => x"51",
          1374 => x"f0",
          1375 => x"82",
          1376 => x"72",
          1377 => x"08",
          1378 => x"08",
          1379 => x"8c",
          1380 => x"05",
          1381 => x"d5",
          1382 => x"f0",
          1383 => x"0c",
          1384 => x"04",
          1385 => x"56",
          1386 => x"38",
          1387 => x"16",
          1388 => x"54",
          1389 => x"38",
          1390 => x"76",
          1391 => x"08",
          1392 => x"e4",
          1393 => x"53",
          1394 => x"82",
          1395 => x"33",
          1396 => x"81",
          1397 => x"99",
          1398 => x"82",
          1399 => x"ff",
          1400 => x"81",
          1401 => x"ac",
          1402 => x"9c",
          1403 => x"51",
          1404 => x"80",
          1405 => x"eb",
          1406 => x"39",
          1407 => x"82",
          1408 => x"b4",
          1409 => x"a4",
          1410 => x"51",
          1411 => x"bb",
          1412 => x"82",
          1413 => x"ac",
          1414 => x"a3",
          1415 => x"82",
          1416 => x"84",
          1417 => x"8b",
          1418 => x"82",
          1419 => x"3d",
          1420 => x"56",
          1421 => x"74",
          1422 => x"39",
          1423 => x"3f",
          1424 => x"ef",
          1425 => x"79",
          1426 => x"ff",
          1427 => x"ec",
          1428 => x"e3",
          1429 => x"30",
          1430 => x"59",
          1431 => x"83",
          1432 => x"81",
          1433 => x"81",
          1434 => x"3d",
          1435 => x"82",
          1436 => x"08",
          1437 => x"c0",
          1438 => x"59",
          1439 => x"53",
          1440 => x"3f",
          1441 => x"e4",
          1442 => x"2e",
          1443 => x"59",
          1444 => x"81",
          1445 => x"07",
          1446 => x"72",
          1447 => x"2e",
          1448 => x"c0",
          1449 => x"92",
          1450 => x"0c",
          1451 => x"7c",
          1452 => x"59",
          1453 => x"51",
          1454 => x"a8",
          1455 => x"81",
          1456 => x"c4",
          1457 => x"e4",
          1458 => x"82",
          1459 => x"04",
          1460 => x"0d",
          1461 => x"02",
          1462 => x"73",
          1463 => x"5e",
          1464 => x"ff",
          1465 => x"ff",
          1466 => x"27",
          1467 => x"38",
          1468 => x"39",
          1469 => x"38",
          1470 => x"ff",
          1471 => x"94",
          1472 => x"55",
          1473 => x"7a",
          1474 => x"b6",
          1475 => x"39",
          1476 => x"3f",
          1477 => x"53",
          1478 => x"52",
          1479 => x"3f",
          1480 => x"b7",
          1481 => x"c8",
          1482 => x"fe",
          1483 => x"b6",
          1484 => x"80",
          1485 => x"53",
          1486 => x"81",
          1487 => x"38",
          1488 => x"ff",
          1489 => x"38",
          1490 => x"f1",
          1491 => x"82",
          1492 => x"8a",
          1493 => x"82",
          1494 => x"18",
          1495 => x"82",
          1496 => x"2c",
          1497 => x"06",
          1498 => x"e4",
          1499 => x"a0",
          1500 => x"30",
          1501 => x"51",
          1502 => x"73",
          1503 => x"81",
          1504 => x"7c",
          1505 => x"38",
          1506 => x"8f",
          1507 => x"9b",
          1508 => x"b7",
          1509 => x"82",
          1510 => x"82",
          1511 => x"82",
          1512 => x"51",
          1513 => x"84",
          1514 => x"04",
          1515 => x"08",
          1516 => x"cd",
          1517 => x"3f",
          1518 => x"2a",
          1519 => x"2e",
          1520 => x"82",
          1521 => x"51",
          1522 => x"81",
          1523 => x"38",
          1524 => x"98",
          1525 => x"85",
          1526 => x"51",
          1527 => x"51",
          1528 => x"99",
          1529 => x"72",
          1530 => x"71",
          1531 => x"d5",
          1532 => x"3f",
          1533 => x"2a",
          1534 => x"2e",
          1535 => x"82",
          1536 => x"51",
          1537 => x"81",
          1538 => x"38",
          1539 => x"e4",
          1540 => x"8d",
          1541 => x"51",
          1542 => x"51",
          1543 => x"98",
          1544 => x"72",
          1545 => x"71",
          1546 => x"dd",
          1547 => x"3f",
          1548 => x"3f",
          1549 => x"77",
          1550 => x"55",
          1551 => x"91",
          1552 => x"54",
          1553 => x"c8",
          1554 => x"bf",
          1555 => x"82",
          1556 => x"71",
          1557 => x"82",
          1558 => x"d8",
          1559 => x"06",
          1560 => x"52",
          1561 => x"d5",
          1562 => x"d5",
          1563 => x"39",
          1564 => x"3f",
          1565 => x"34",
          1566 => x"73",
          1567 => x"82",
          1568 => x"a9",
          1569 => x"0c",
          1570 => x"80",
          1571 => x"f0",
          1572 => x"c7",
          1573 => x"ff",
          1574 => x"06",
          1575 => x"82",
          1576 => x"3f",
          1577 => x"51",
          1578 => x"08",
          1579 => x"51",
          1580 => x"82",
          1581 => x"97",
          1582 => x"79",
          1583 => x"84",
          1584 => x"e4",
          1585 => x"59",
          1586 => x"78",
          1587 => x"2e",
          1588 => x"38",
          1589 => x"bc",
          1590 => x"78",
          1591 => x"80",
          1592 => x"2e",
          1593 => x"80",
          1594 => x"f9",
          1595 => x"88",
          1596 => x"a3",
          1597 => x"2e",
          1598 => x"8b",
          1599 => x"38",
          1600 => x"89",
          1601 => x"ff",
          1602 => x"ec",
          1603 => x"2e",
          1604 => x"11",
          1605 => x"3f",
          1606 => x"af",
          1607 => x"ff",
          1608 => x"d5",
          1609 => x"08",
          1610 => x"80",
          1611 => x"27",
          1612 => x"70",
          1613 => x"f5",
          1614 => x"80",
          1615 => x"f7",
          1616 => x"fd",
          1617 => x"53",
          1618 => x"82",
          1619 => x"38",
          1620 => x"84",
          1621 => x"e4",
          1622 => x"ba",
          1623 => x"5a",
          1624 => x"59",
          1625 => x"34",
          1626 => x"3d",
          1627 => x"51",
          1628 => x"80",
          1629 => x"fc",
          1630 => x"ff",
          1631 => x"fc",
          1632 => x"53",
          1633 => x"82",
          1634 => x"38",
          1635 => x"3f",
          1636 => x"62",
          1637 => x"78",
          1638 => x"54",
          1639 => x"d0",
          1640 => x"63",
          1641 => x"51",
          1642 => x"3d",
          1643 => x"51",
          1644 => x"80",
          1645 => x"78",
          1646 => x"08",
          1647 => x"33",
          1648 => x"d4",
          1649 => x"ca",
          1650 => x"82",
          1651 => x"d4",
          1652 => x"38",
          1653 => x"82",
          1654 => x"88",
          1655 => x"39",
          1656 => x"45",
          1657 => x"84",
          1658 => x"e4",
          1659 => x"33",
          1660 => x"d4",
          1661 => x"d4",
          1662 => x"38",
          1663 => x"82",
          1664 => x"88",
          1665 => x"39",
          1666 => x"2e",
          1667 => x"99",
          1668 => x"80",
          1669 => x"44",
          1670 => x"05",
          1671 => x"ff",
          1672 => x"d5",
          1673 => x"63",
          1674 => x"81",
          1675 => x"72",
          1676 => x"51",
          1677 => x"7a",
          1678 => x"ba",
          1679 => x"64",
          1680 => x"f2",
          1681 => x"b1",
          1682 => x"ff",
          1683 => x"d5",
          1684 => x"b5",
          1685 => x"05",
          1686 => x"08",
          1687 => x"80",
          1688 => x"05",
          1689 => x"ff",
          1690 => x"d5",
          1691 => x"64",
          1692 => x"51",
          1693 => x"08",
          1694 => x"aa",
          1695 => x"78",
          1696 => x"27",
          1697 => x"53",
          1698 => x"82",
          1699 => x"64",
          1700 => x"34",
          1701 => x"82",
          1702 => x"a7",
          1703 => x"ff",
          1704 => x"d5",
          1705 => x"b5",
          1706 => x"05",
          1707 => x"08",
          1708 => x"80",
          1709 => x"5b",
          1710 => x"11",
          1711 => x"3f",
          1712 => x"df",
          1713 => x"bb",
          1714 => x"f1",
          1715 => x"51",
          1716 => x"33",
          1717 => x"78",
          1718 => x"42",
          1719 => x"53",
          1720 => x"82",
          1721 => x"61",
          1722 => x"70",
          1723 => x"a9",
          1724 => x"3f",
          1725 => x"11",
          1726 => x"3f",
          1727 => x"e7",
          1728 => x"ff",
          1729 => x"d5",
          1730 => x"61",
          1731 => x"b5",
          1732 => x"05",
          1733 => x"08",
          1734 => x"08",
          1735 => x"a7",
          1736 => x"80",
          1737 => x"3f",
          1738 => x"2e",
          1739 => x"38",
          1740 => x"84",
          1741 => x"e4",
          1742 => x"71",
          1743 => x"b5",
          1744 => x"3f",
          1745 => x"11",
          1746 => x"3f",
          1747 => x"c7",
          1748 => x"ff",
          1749 => x"b5",
          1750 => x"05",
          1751 => x"08",
          1752 => x"82",
          1753 => x"64",
          1754 => x"80",
          1755 => x"08",
          1756 => x"f0",
          1757 => x"51",
          1758 => x"f4",
          1759 => x"e3",
          1760 => x"e2",
          1761 => x"59",
          1762 => x"f8",
          1763 => x"d5",
          1764 => x"80",
          1765 => x"08",
          1766 => x"83",
          1767 => x"7f",
          1768 => x"d2",
          1769 => x"b5",
          1770 => x"81",
          1771 => x"b2",
          1772 => x"81",
          1773 => x"83",
          1774 => x"bc",
          1775 => x"54",
          1776 => x"3d",
          1777 => x"3f",
          1778 => x"b0",
          1779 => x"7b",
          1780 => x"82",
          1781 => x"05",
          1782 => x"7b",
          1783 => x"b5",
          1784 => x"f8",
          1785 => x"94",
          1786 => x"84",
          1787 => x"b5",
          1788 => x"3f",
          1789 => x"08",
          1790 => x"25",
          1791 => x"83",
          1792 => x"06",
          1793 => x"1b",
          1794 => x"fe",
          1795 => x"32",
          1796 => x"2e",
          1797 => x"e0",
          1798 => x"b1",
          1799 => x"f0",
          1800 => x"39",
          1801 => x"94",
          1802 => x"54",
          1803 => x"d7",
          1804 => x"2b",
          1805 => x"52",
          1806 => x"d5",
          1807 => x"94",
          1808 => x"80",
          1809 => x"d5",
          1810 => x"53",
          1811 => x"8e",
          1812 => x"75",
          1813 => x"94",
          1814 => x"c0",
          1815 => x"80",
          1816 => x"99",
          1817 => x"0b",
          1818 => x"72",
          1819 => x"be",
          1820 => x"51",
          1821 => x"51",
          1822 => x"51",
          1823 => x"3f",
          1824 => x"0d",
          1825 => x"52",
          1826 => x"81",
          1827 => x"52",
          1828 => x"d5",
          1829 => x"3d",
          1830 => x"73",
          1831 => x"38",
          1832 => x"81",
          1833 => x"39",
          1834 => x"81",
          1835 => x"54",
          1836 => x"06",
          1837 => x"80",
          1838 => x"83",
          1839 => x"38",
          1840 => x"52",
          1841 => x"2e",
          1842 => x"84",
          1843 => x"52",
          1844 => x"83",
          1845 => x"30",
          1846 => x"51",
          1847 => x"70",
          1848 => x"72",
          1849 => x"3d",
          1850 => x"72",
          1851 => x"fc",
          1852 => x"82",
          1853 => x"83",
          1854 => x"0c",
          1855 => x"76",
          1856 => x"81",
          1857 => x"83",
          1858 => x"70",
          1859 => x"33",
          1860 => x"fe",
          1861 => x"70",
          1862 => x"33",
          1863 => x"e6",
          1864 => x"74",
          1865 => x"13",
          1866 => x"26",
          1867 => x"98",
          1868 => x"bc",
          1869 => x"b8",
          1870 => x"b4",
          1871 => x"b0",
          1872 => x"ac",
          1873 => x"a8",
          1874 => x"73",
          1875 => x"87",
          1876 => x"82",
          1877 => x"f3",
          1878 => x"9c",
          1879 => x"bc",
          1880 => x"98",
          1881 => x"87",
          1882 => x"1c",
          1883 => x"79",
          1884 => x"08",
          1885 => x"98",
          1886 => x"87",
          1887 => x"1c",
          1888 => x"79",
          1889 => x"83",
          1890 => x"ff",
          1891 => x"1b",
          1892 => x"1b",
          1893 => x"83",
          1894 => x"51",
          1895 => x"04",
          1896 => x"82",
          1897 => x"58",
          1898 => x"75",
          1899 => x"94",
          1900 => x"81",
          1901 => x"8c",
          1902 => x"51",
          1903 => x"70",
          1904 => x"8d",
          1905 => x"51",
          1906 => x"ff",
          1907 => x"70",
          1908 => x"90",
          1909 => x"e4",
          1910 => x"0d",
          1911 => x"9f",
          1912 => x"fc",
          1913 => x"0d",
          1914 => x"2e",
          1915 => x"8d",
          1916 => x"70",
          1917 => x"94",
          1918 => x"87",
          1919 => x"96",
          1920 => x"72",
          1921 => x"70",
          1922 => x"74",
          1923 => x"72",
          1924 => x"70",
          1925 => x"38",
          1926 => x"94",
          1927 => x"87",
          1928 => x"80",
          1929 => x"0d",
          1930 => x"74",
          1931 => x"57",
          1932 => x"81",
          1933 => x"33",
          1934 => x"58",
          1935 => x"2e",
          1936 => x"70",
          1937 => x"53",
          1938 => x"71",
          1939 => x"70",
          1940 => x"06",
          1941 => x"71",
          1942 => x"70",
          1943 => x"51",
          1944 => x"2e",
          1945 => x"77",
          1946 => x"81",
          1947 => x"86",
          1948 => x"3d",
          1949 => x"fc",
          1950 => x"87",
          1951 => x"86",
          1952 => x"08",
          1953 => x"51",
          1954 => x"81",
          1955 => x"52",
          1956 => x"94",
          1957 => x"06",
          1958 => x"0d",
          1959 => x"08",
          1960 => x"04",
          1961 => x"70",
          1962 => x"94",
          1963 => x"87",
          1964 => x"82",
          1965 => x"ff",
          1966 => x"81",
          1967 => x"52",
          1968 => x"94",
          1969 => x"70",
          1970 => x"d5",
          1971 => x"3d",
          1972 => x"9c",
          1973 => x"2e",
          1974 => x"08",
          1975 => x"a8",
          1976 => x"9e",
          1977 => x"c0",
          1978 => x"87",
          1979 => x"0c",
          1980 => x"94",
          1981 => x"d4",
          1982 => x"82",
          1983 => x"08",
          1984 => x"b8",
          1985 => x"9e",
          1986 => x"c0",
          1987 => x"87",
          1988 => x"0c",
          1989 => x"82",
          1990 => x"08",
          1991 => x"88",
          1992 => x"9e",
          1993 => x"0b",
          1994 => x"c0",
          1995 => x"06",
          1996 => x"38",
          1997 => x"80",
          1998 => x"88",
          1999 => x"80",
          2000 => x"d4",
          2001 => x"90",
          2002 => x"52",
          2003 => x"52",
          2004 => x"87",
          2005 => x"80",
          2006 => x"83",
          2007 => x"34",
          2008 => x"70",
          2009 => x"70",
          2010 => x"82",
          2011 => x"9e",
          2012 => x"51",
          2013 => x"81",
          2014 => x"0b",
          2015 => x"80",
          2016 => x"2e",
          2017 => x"cb",
          2018 => x"08",
          2019 => x"52",
          2020 => x"71",
          2021 => x"c0",
          2022 => x"06",
          2023 => x"38",
          2024 => x"80",
          2025 => x"80",
          2026 => x"80",
          2027 => x"d4",
          2028 => x"90",
          2029 => x"52",
          2030 => x"71",
          2031 => x"90",
          2032 => x"2a",
          2033 => x"34",
          2034 => x"70",
          2035 => x"80",
          2036 => x"d4",
          2037 => x"70",
          2038 => x"51",
          2039 => x"0b",
          2040 => x"06",
          2041 => x"38",
          2042 => x"87",
          2043 => x"51",
          2044 => x"3d",
          2045 => x"d8",
          2046 => x"c4",
          2047 => x"82",
          2048 => x"82",
          2049 => x"82",
          2050 => x"94",
          2051 => x"a4",
          2052 => x"51",
          2053 => x"33",
          2054 => x"d4",
          2055 => x"54",
          2056 => x"90",
          2057 => x"80",
          2058 => x"82",
          2059 => x"be",
          2060 => x"d4",
          2061 => x"38",
          2062 => x"08",
          2063 => x"ff",
          2064 => x"54",
          2065 => x"90",
          2066 => x"52",
          2067 => x"3f",
          2068 => x"2e",
          2069 => x"82",
          2070 => x"82",
          2071 => x"8e",
          2072 => x"bf",
          2073 => x"d4",
          2074 => x"38",
          2075 => x"e4",
          2076 => x"c5",
          2077 => x"82",
          2078 => x"82",
          2079 => x"89",
          2080 => x"db",
          2081 => x"80",
          2082 => x"ff",
          2083 => x"54",
          2084 => x"b0",
          2085 => x"ce",
          2086 => x"82",
          2087 => x"82",
          2088 => x"82",
          2089 => x"51",
          2090 => x"08",
          2091 => x"f8",
          2092 => x"c1",
          2093 => x"c1",
          2094 => x"d4",
          2095 => x"ff",
          2096 => x"56",
          2097 => x"9e",
          2098 => x"c0",
          2099 => x"d5",
          2100 => x"ff",
          2101 => x"54",
          2102 => x"bc",
          2103 => x"51",
          2104 => x"bd",
          2105 => x"54",
          2106 => x"a0",
          2107 => x"c6",
          2108 => x"82",
          2109 => x"52",
          2110 => x"e4",
          2111 => x"31",
          2112 => x"82",
          2113 => x"8a",
          2114 => x"0d",
          2115 => x"33",
          2116 => x"38",
          2117 => x"52",
          2118 => x"9d",
          2119 => x"82",
          2120 => x"90",
          2121 => x"85",
          2122 => x"80",
          2123 => x"80",
          2124 => x"84",
          2125 => x"c0",
          2126 => x"76",
          2127 => x"2b",
          2128 => x"82",
          2129 => x"80",
          2130 => x"53",
          2131 => x"a4",
          2132 => x"05",
          2133 => x"72",
          2134 => x"53",
          2135 => x"0d",
          2136 => x"05",
          2137 => x"54",
          2138 => x"c8",
          2139 => x"3f",
          2140 => x"ff",
          2141 => x"52",
          2142 => x"33",
          2143 => x"81",
          2144 => x"ff",
          2145 => x"3d",
          2146 => x"84",
          2147 => x"bb",
          2148 => x"84",
          2149 => x"51",
          2150 => x"2e",
          2151 => x"82",
          2152 => x"d4",
          2153 => x"56",
          2154 => x"08",
          2155 => x"84",
          2156 => x"51",
          2157 => x"75",
          2158 => x"ed",
          2159 => x"55",
          2160 => x"ff",
          2161 => x"80",
          2162 => x"2e",
          2163 => x"75",
          2164 => x"33",
          2165 => x"05",
          2166 => x"80",
          2167 => x"52",
          2168 => x"d5",
          2169 => x"8c",
          2170 => x"d4",
          2171 => x"71",
          2172 => x"d1",
          2173 => x"14",
          2174 => x"80",
          2175 => x"b0",
          2176 => x"71",
          2177 => x"b0",
          2178 => x"82",
          2179 => x"dc",
          2180 => x"d5",
          2181 => x"82",
          2182 => x"d5",
          2183 => x"3d",
          2184 => x"82",
          2185 => x"75",
          2186 => x"e4",
          2187 => x"08",
          2188 => x"ff",
          2189 => x"34",
          2190 => x"c6",
          2191 => x"74",
          2192 => x"38",
          2193 => x"aa",
          2194 => x"81",
          2195 => x"b0",
          2196 => x"d5",
          2197 => x"82",
          2198 => x"52",
          2199 => x"c5",
          2200 => x"a5",
          2201 => x"82",
          2202 => x"80",
          2203 => x"38",
          2204 => x"17",
          2205 => x"70",
          2206 => x"55",
          2207 => x"ff",
          2208 => x"11",
          2209 => x"82",
          2210 => x"82",
          2211 => x"78",
          2212 => x"75",
          2213 => x"79",
          2214 => x"08",
          2215 => x"80",
          2216 => x"3d",
          2217 => x"71",
          2218 => x"58",
          2219 => x"38",
          2220 => x"27",
          2221 => x"71",
          2222 => x"09",
          2223 => x"ea",
          2224 => x"d5",
          2225 => x"b0",
          2226 => x"79",
          2227 => x"3f",
          2228 => x"84",
          2229 => x"38",
          2230 => x"fc",
          2231 => x"8c",
          2232 => x"c5",
          2233 => x"2e",
          2234 => x"77",
          2235 => x"08",
          2236 => x"74",
          2237 => x"ff",
          2238 => x"8b",
          2239 => x"0c",
          2240 => x"b0",
          2241 => x"08",
          2242 => x"34",
          2243 => x"08",
          2244 => x"82",
          2245 => x"38",
          2246 => x"38",
          2247 => x"80",
          2248 => x"87",
          2249 => x"b0",
          2250 => x"81",
          2251 => x"d5",
          2252 => x"82",
          2253 => x"82",
          2254 => x"80",
          2255 => x"82",
          2256 => x"90",
          2257 => x"3f",
          2258 => x"e4",
          2259 => x"d0",
          2260 => x"ae",
          2261 => x"80",
          2262 => x"38",
          2263 => x"17",
          2264 => x"74",
          2265 => x"c2",
          2266 => x"5c",
          2267 => x"5b",
          2268 => x"97",
          2269 => x"34",
          2270 => x"80",
          2271 => x"3d",
          2272 => x"08",
          2273 => x"78",
          2274 => x"06",
          2275 => x"70",
          2276 => x"98",
          2277 => x"05",
          2278 => x"70",
          2279 => x"51",
          2280 => x"56",
          2281 => x"74",
          2282 => x"29",
          2283 => x"51",
          2284 => x"76",
          2285 => x"3f",
          2286 => x"54",
          2287 => x"ed",
          2288 => x"81",
          2289 => x"70",
          2290 => x"51",
          2291 => x"53",
          2292 => x"82",
          2293 => x"73",
          2294 => x"80",
          2295 => x"74",
          2296 => x"70",
          2297 => x"98",
          2298 => x"70",
          2299 => x"5e",
          2300 => x"74",
          2301 => x"38",
          2302 => x"80",
          2303 => x"82",
          2304 => x"ed",
          2305 => x"78",
          2306 => x"54",
          2307 => x"84",
          2308 => x"08",
          2309 => x"7e",
          2310 => x"33",
          2311 => x"98",
          2312 => x"75",
          2313 => x"33",
          2314 => x"29",
          2315 => x"82",
          2316 => x"39",
          2317 => x"54",
          2318 => x"54",
          2319 => x"a4",
          2320 => x"81",
          2321 => x"82",
          2322 => x"29",
          2323 => x"82",
          2324 => x"74",
          2325 => x"08",
          2326 => x"ff",
          2327 => x"29",
          2328 => x"82",
          2329 => x"75",
          2330 => x"70",
          2331 => x"a4",
          2332 => x"25",
          2333 => x"52",
          2334 => x"81",
          2335 => x"70",
          2336 => x"51",
          2337 => x"ee",
          2338 => x"1b",
          2339 => x"82",
          2340 => x"fd",
          2341 => x"ff",
          2342 => x"c6",
          2343 => x"54",
          2344 => x"54",
          2345 => x"c8",
          2346 => x"3f",
          2347 => x"70",
          2348 => x"51",
          2349 => x"74",
          2350 => x"82",
          2351 => x"ff",
          2352 => x"29",
          2353 => x"82",
          2354 => x"75",
          2355 => x"52",
          2356 => x"ed",
          2357 => x"2c",
          2358 => x"57",
          2359 => x"f1",
          2360 => x"ea",
          2361 => x"80",
          2362 => x"a4",
          2363 => x"de",
          2364 => x"33",
          2365 => x"f1",
          2366 => x"ba",
          2367 => x"f6",
          2368 => x"ff",
          2369 => x"a4",
          2370 => x"81",
          2371 => x"3f",
          2372 => x"82",
          2373 => x"a4",
          2374 => x"3d",
          2375 => x"73",
          2376 => x"c8",
          2377 => x"3f",
          2378 => x"73",
          2379 => x"06",
          2380 => x"82",
          2381 => x"2e",
          2382 => x"82",
          2383 => x"98",
          2384 => x"55",
          2385 => x"54",
          2386 => x"c8",
          2387 => x"92",
          2388 => x"80",
          2389 => x"a4",
          2390 => x"d5",
          2391 => x"51",
          2392 => x"33",
          2393 => x"ed",
          2394 => x"74",
          2395 => x"08",
          2396 => x"74",
          2397 => x"05",
          2398 => x"58",
          2399 => x"f7",
          2400 => x"81",
          2401 => x"56",
          2402 => x"82",
          2403 => x"73",
          2404 => x"33",
          2405 => x"ed",
          2406 => x"ed",
          2407 => x"26",
          2408 => x"a8",
          2409 => x"ee",
          2410 => x"34",
          2411 => x"9e",
          2412 => x"08",
          2413 => x"51",
          2414 => x"08",
          2415 => x"08",
          2416 => x"52",
          2417 => x"5b",
          2418 => x"d4",
          2419 => x"74",
          2420 => x"a4",
          2421 => x"ed",
          2422 => x"ff",
          2423 => x"51",
          2424 => x"80",
          2425 => x"2e",
          2426 => x"ad",
          2427 => x"81",
          2428 => x"55",
          2429 => x"ff",
          2430 => x"82",
          2431 => x"81",
          2432 => x"79",
          2433 => x"39",
          2434 => x"70",
          2435 => x"38",
          2436 => x"d5",
          2437 => x"d5",
          2438 => x"53",
          2439 => x"3f",
          2440 => x"5b",
          2441 => x"74",
          2442 => x"ed",
          2443 => x"3f",
          2444 => x"70",
          2445 => x"59",
          2446 => x"38",
          2447 => x"54",
          2448 => x"70",
          2449 => x"f4",
          2450 => x"73",
          2451 => x"c8",
          2452 => x"3f",
          2453 => x"73",
          2454 => x"f9",
          2455 => x"d5",
          2456 => x"d0",
          2457 => x"84",
          2458 => x"82",
          2459 => x"74",
          2460 => x"82",
          2461 => x"34",
          2462 => x"08",
          2463 => x"15",
          2464 => x"d0",
          2465 => x"70",
          2466 => x"58",
          2467 => x"73",
          2468 => x"70",
          2469 => x"f8",
          2470 => x"34",
          2471 => x"04",
          2472 => x"84",
          2473 => x"2a",
          2474 => x"51",
          2475 => x"83",
          2476 => x"a6",
          2477 => x"22",
          2478 => x"83",
          2479 => x"11",
          2480 => x"2b",
          2481 => x"71",
          2482 => x"2a",
          2483 => x"57",
          2484 => x"81",
          2485 => x"75",
          2486 => x"34",
          2487 => x"08",
          2488 => x"71",
          2489 => x"ff",
          2490 => x"05",
          2491 => x"2a",
          2492 => x"72",
          2493 => x"34",
          2494 => x"76",
          2495 => x"0d",
          2496 => x"08",
          2497 => x"83",
          2498 => x"12",
          2499 => x"07",
          2500 => x"05",
          2501 => x"88",
          2502 => x"56",
          2503 => x"13",
          2504 => x"84",
          2505 => x"2b",
          2506 => x"52",
          2507 => x"33",
          2508 => x"54",
          2509 => x"73",
          2510 => x"13",
          2511 => x"2b",
          2512 => x"88",
          2513 => x"73",
          2514 => x"0d",
          2515 => x"22",
          2516 => x"71",
          2517 => x"88",
          2518 => x"33",
          2519 => x"90",
          2520 => x"5a",
          2521 => x"80",
          2522 => x"82",
          2523 => x"81",
          2524 => x"2b",
          2525 => x"33",
          2526 => x"8f",
          2527 => x"53",
          2528 => x"2a",
          2529 => x"83",
          2530 => x"16",
          2531 => x"2b",
          2532 => x"55",
          2533 => x"71",
          2534 => x"06",
          2535 => x"52",
          2536 => x"88",
          2537 => x"d5",
          2538 => x"22",
          2539 => x"33",
          2540 => x"83",
          2541 => x"52",
          2542 => x"71",
          2543 => x"05",
          2544 => x"51",
          2545 => x"81",
          2546 => x"15",
          2547 => x"2b",
          2548 => x"52",
          2549 => x"33",
          2550 => x"54",
          2551 => x"72",
          2552 => x"14",
          2553 => x"88",
          2554 => x"54",
          2555 => x"7b",
          2556 => x"70",
          2557 => x"53",
          2558 => x"76",
          2559 => x"83",
          2560 => x"2b",
          2561 => x"33",
          2562 => x"53",
          2563 => x"59",
          2564 => x"80",
          2565 => x"81",
          2566 => x"33",
          2567 => x"76",
          2568 => x"58",
          2569 => x"ff",
          2570 => x"d5",
          2571 => x"85",
          2572 => x"88",
          2573 => x"84",
          2574 => x"d5",
          2575 => x"14",
          2576 => x"d5",
          2577 => x"75",
          2578 => x"18",
          2579 => x"2b",
          2580 => x"88",
          2581 => x"74",
          2582 => x"0d",
          2583 => x"d5",
          2584 => x"71",
          2585 => x"8c",
          2586 => x"0d",
          2587 => x"82",
          2588 => x"82",
          2589 => x"12",
          2590 => x"59",
          2591 => x"75",
          2592 => x"29",
          2593 => x"88",
          2594 => x"79",
          2595 => x"7f",
          2596 => x"77",
          2597 => x"85",
          2598 => x"33",
          2599 => x"57",
          2600 => x"ff",
          2601 => x"80",
          2602 => x"11",
          2603 => x"2b",
          2604 => x"52",
          2605 => x"83",
          2606 => x"26",
          2607 => x"2e",
          2608 => x"81",
          2609 => x"3f",
          2610 => x"79",
          2611 => x"d5",
          2612 => x"87",
          2613 => x"2b",
          2614 => x"7a",
          2615 => x"88",
          2616 => x"15",
          2617 => x"85",
          2618 => x"83",
          2619 => x"33",
          2620 => x"70",
          2621 => x"56",
          2622 => x"19",
          2623 => x"84",
          2624 => x"2b",
          2625 => x"55",
          2626 => x"76",
          2627 => x"70",
          2628 => x"12",
          2629 => x"2a",
          2630 => x"84",
          2631 => x"d5",
          2632 => x"82",
          2633 => x"fe",
          2634 => x"08",
          2635 => x"71",
          2636 => x"ed",
          2637 => x"82",
          2638 => x"ee",
          2639 => x"70",
          2640 => x"2e",
          2641 => x"3f",
          2642 => x"3f",
          2643 => x"39",
          2644 => x"3f",
          2645 => x"f5",
          2646 => x"ff",
          2647 => x"71",
          2648 => x"06",
          2649 => x"81",
          2650 => x"75",
          2651 => x"88",
          2652 => x"70",
          2653 => x"07",
          2654 => x"48",
          2655 => x"56",
          2656 => x"76",
          2657 => x"83",
          2658 => x"33",
          2659 => x"70",
          2660 => x"33",
          2661 => x"53",
          2662 => x"25",
          2663 => x"ff",
          2664 => x"81",
          2665 => x"2e",
          2666 => x"f6",
          2667 => x"58",
          2668 => x"74",
          2669 => x"3f",
          2670 => x"75",
          2671 => x"11",
          2672 => x"07",
          2673 => x"52",
          2674 => x"e4",
          2675 => x"7c",
          2676 => x"08",
          2677 => x"91",
          2678 => x"84",
          2679 => x"5c",
          2680 => x"74",
          2681 => x"c9",
          2682 => x"11",
          2683 => x"07",
          2684 => x"52",
          2685 => x"e4",
          2686 => x"7c",
          2687 => x"08",
          2688 => x"91",
          2689 => x"84",
          2690 => x"73",
          2691 => x"7b",
          2692 => x"d5",
          2693 => x"80",
          2694 => x"82",
          2695 => x"3f",
          2696 => x"7a",
          2697 => x"52",
          2698 => x"83",
          2699 => x"05",
          2700 => x"82",
          2701 => x"fc",
          2702 => x"54",
          2703 => x"55",
          2704 => x"38",
          2705 => x"08",
          2706 => x"d5",
          2707 => x"3d",
          2708 => x"52",
          2709 => x"e0",
          2710 => x"0c",
          2711 => x"02",
          2712 => x"05",
          2713 => x"26",
          2714 => x"c0",
          2715 => x"74",
          2716 => x"73",
          2717 => x"51",
          2718 => x"98",
          2719 => x"82",
          2720 => x"38",
          2721 => x"ec",
          2722 => x"52",
          2723 => x"08",
          2724 => x"82",
          2725 => x"13",
          2726 => x"86",
          2727 => x"62",
          2728 => x"57",
          2729 => x"fe",
          2730 => x"06",
          2731 => x"71",
          2732 => x"80",
          2733 => x"c0",
          2734 => x"5a",
          2735 => x"0c",
          2736 => x"08",
          2737 => x"53",
          2738 => x"08",
          2739 => x"34",
          2740 => x"53",
          2741 => x"53",
          2742 => x"80",
          2743 => x"08",
          2744 => x"8c",
          2745 => x"78",
          2746 => x"0c",
          2747 => x"08",
          2748 => x"38",
          2749 => x"17",
          2750 => x"53",
          2751 => x"fc",
          2752 => x"7d",
          2753 => x"80",
          2754 => x"38",
          2755 => x"e4",
          2756 => x"0d",
          2757 => x"05",
          2758 => x"80",
          2759 => x"d5",
          2760 => x"71",
          2761 => x"38",
          2762 => x"80",
          2763 => x"c0",
          2764 => x"5a",
          2765 => x"76",
          2766 => x"75",
          2767 => x"51",
          2768 => x"7a",
          2769 => x"81",
          2770 => x"06",
          2771 => x"87",
          2772 => x"38",
          2773 => x"80",
          2774 => x"99",
          2775 => x"8c",
          2776 => x"51",
          2777 => x"8d",
          2778 => x"84",
          2779 => x"2e",
          2780 => x"52",
          2781 => x"f8",
          2782 => x"71",
          2783 => x"53",
          2784 => x"0d",
          2785 => x"05",
          2786 => x"05",
          2787 => x"fe",
          2788 => x"53",
          2789 => x"0b",
          2790 => x"71",
          2791 => x"24",
          2792 => x"92",
          2793 => x"8d",
          2794 => x"80",
          2795 => x"70",
          2796 => x"52",
          2797 => x"98",
          2798 => x"c0",
          2799 => x"81",
          2800 => x"53",
          2801 => x"71",
          2802 => x"39",
          2803 => x"81",
          2804 => x"84",
          2805 => x"0c",
          2806 => x"74",
          2807 => x"2b",
          2808 => x"84",
          2809 => x"83",
          2810 => x"2b",
          2811 => x"70",
          2812 => x"07",
          2813 => x"56",
          2814 => x"3d",
          2815 => x"22",
          2816 => x"54",
          2817 => x"34",
          2818 => x"73",
          2819 => x"05",
          2820 => x"72",
          2821 => x"2a",
          2822 => x"34",
          2823 => x"83",
          2824 => x"75",
          2825 => x"92",
          2826 => x"73",
          2827 => x"51",
          2828 => x"3d",
          2829 => x"72",
          2830 => x"11",
          2831 => x"04",
          2832 => x"56",
          2833 => x"74",
          2834 => x"31",
          2835 => x"80",
          2836 => x"38",
          2837 => x"0d",
          2838 => x"51",
          2839 => x"81",
          2840 => x"38",
          2841 => x"3d",
          2842 => x"0c",
          2843 => x"70",
          2844 => x"55",
          2845 => x"d5",
          2846 => x"98",
          2847 => x"f9",
          2848 => x"ff",
          2849 => x"38",
          2850 => x"d5",
          2851 => x"3d",
          2852 => x"33",
          2853 => x"38",
          2854 => x"16",
          2855 => x"f9",
          2856 => x"2e",
          2857 => x"e4",
          2858 => x"70",
          2859 => x"59",
          2860 => x"82",
          2861 => x"81",
          2862 => x"53",
          2863 => x"a5",
          2864 => x"d5",
          2865 => x"3d",
          2866 => x"74",
          2867 => x"51",
          2868 => x"57",
          2869 => x"54",
          2870 => x"33",
          2871 => x"08",
          2872 => x"57",
          2873 => x"e4",
          2874 => x"0d",
          2875 => x"82",
          2876 => x"08",
          2877 => x"83",
          2878 => x"84",
          2879 => x"81",
          2880 => x"82",
          2881 => x"52",
          2882 => x"52",
          2883 => x"84",
          2884 => x"fb",
          2885 => x"52",
          2886 => x"94",
          2887 => x"fb",
          2888 => x"a4",
          2889 => x"08",
          2890 => x"55",
          2891 => x"f7",
          2892 => x"53",
          2893 => x"99",
          2894 => x"83",
          2895 => x"0c",
          2896 => x"77",
          2897 => x"55",
          2898 => x"8d",
          2899 => x"b0",
          2900 => x"d5",
          2901 => x"3d",
          2902 => x"57",
          2903 => x"9c",
          2904 => x"74",
          2905 => x"f5",
          2906 => x"81",
          2907 => x"83",
          2908 => x"76",
          2909 => x"16",
          2910 => x"96",
          2911 => x"38",
          2912 => x"33",
          2913 => x"08",
          2914 => x"fc",
          2915 => x"fe",
          2916 => x"11",
          2917 => x"81",
          2918 => x"51",
          2919 => x"ff",
          2920 => x"2a",
          2921 => x"fc",
          2922 => x"c6",
          2923 => x"05",
          2924 => x"d5",
          2925 => x"ae",
          2926 => x"05",
          2927 => x"d5",
          2928 => x"83",
          2929 => x"f8",
          2930 => x"0a",
          2931 => x"82",
          2932 => x"f8",
          2933 => x"56",
          2934 => x"38",
          2935 => x"38",
          2936 => x"9d",
          2937 => x"81",
          2938 => x"83",
          2939 => x"76",
          2940 => x"18",
          2941 => x"9e",
          2942 => x"d5",
          2943 => x"ff",
          2944 => x"81",
          2945 => x"80",
          2946 => x"f0",
          2947 => x"51",
          2948 => x"17",
          2949 => x"05",
          2950 => x"d5",
          2951 => x"81",
          2952 => x"b8",
          2953 => x"8f",
          2954 => x"f0",
          2955 => x"72",
          2956 => x"2a",
          2957 => x"fa",
          2958 => x"82",
          2959 => x"83",
          2960 => x"fe",
          2961 => x"e6",
          2962 => x"17",
          2963 => x"3f",
          2964 => x"e4",
          2965 => x"77",
          2966 => x"b8",
          2967 => x"8b",
          2968 => x"06",
          2969 => x"3f",
          2970 => x"d5",
          2971 => x"3d",
          2972 => x"56",
          2973 => x"74",
          2974 => x"80",
          2975 => x"75",
          2976 => x"08",
          2977 => x"38",
          2978 => x"81",
          2979 => x"08",
          2980 => x"51",
          2981 => x"58",
          2982 => x"c7",
          2983 => x"d2",
          2984 => x"cf",
          2985 => x"fc",
          2986 => x"38",
          2987 => x"08",
          2988 => x"38",
          2989 => x"33",
          2990 => x"77",
          2991 => x"80",
          2992 => x"3d",
          2993 => x"71",
          2994 => x"90",
          2995 => x"38",
          2996 => x"81",
          2997 => x"f9",
          2998 => x"e4",
          2999 => x"e4",
          3000 => x"2e",
          3001 => x"d5",
          3002 => x"58",
          3003 => x"80",
          3004 => x"09",
          3005 => x"56",
          3006 => x"82",
          3007 => x"3f",
          3008 => x"2e",
          3009 => x"e4",
          3010 => x"70",
          3011 => x"7c",
          3012 => x"51",
          3013 => x"d5",
          3014 => x"17",
          3015 => x"73",
          3016 => x"58",
          3017 => x"56",
          3018 => x"26",
          3019 => x"81",
          3020 => x"c6",
          3021 => x"b8",
          3022 => x"81",
          3023 => x"d5",
          3024 => x"09",
          3025 => x"70",
          3026 => x"80",
          3027 => x"06",
          3028 => x"39",
          3029 => x"f7",
          3030 => x"e4",
          3031 => x"07",
          3032 => x"2e",
          3033 => x"75",
          3034 => x"3f",
          3035 => x"38",
          3036 => x"fe",
          3037 => x"74",
          3038 => x"0c",
          3039 => x"84",
          3040 => x"81",
          3041 => x"8c",
          3042 => x"39",
          3043 => x"e4",
          3044 => x"0d",
          3045 => x"82",
          3046 => x"d5",
          3047 => x"74",
          3048 => x"08",
          3049 => x"59",
          3050 => x"70",
          3051 => x"84",
          3052 => x"58",
          3053 => x"75",
          3054 => x"51",
          3055 => x"80",
          3056 => x"32",
          3057 => x"2a",
          3058 => x"e4",
          3059 => x"0d",
          3060 => x"74",
          3061 => x"74",
          3062 => x"74",
          3063 => x"73",
          3064 => x"27",
          3065 => x"9b",
          3066 => x"88",
          3067 => x"80",
          3068 => x"0c",
          3069 => x"89",
          3070 => x"38",
          3071 => x"82",
          3072 => x"08",
          3073 => x"d5",
          3074 => x"08",
          3075 => x"82",
          3076 => x"cb",
          3077 => x"3f",
          3078 => x"73",
          3079 => x"82",
          3080 => x"39",
          3081 => x"13",
          3082 => x"16",
          3083 => x"77",
          3084 => x"04",
          3085 => x"12",
          3086 => x"80",
          3087 => x"98",
          3088 => x"55",
          3089 => x"83",
          3090 => x"81",
          3091 => x"55",
          3092 => x"17",
          3093 => x"9b",
          3094 => x"ff",
          3095 => x"81",
          3096 => x"e6",
          3097 => x"55",
          3098 => x"80",
          3099 => x"08",
          3100 => x"08",
          3101 => x"38",
          3102 => x"84",
          3103 => x"52",
          3104 => x"e4",
          3105 => x"08",
          3106 => x"82",
          3107 => x"81",
          3108 => x"b0",
          3109 => x"51",
          3110 => x"a0",
          3111 => x"75",
          3112 => x"08",
          3113 => x"77",
          3114 => x"55",
          3115 => x"0d",
          3116 => x"08",
          3117 => x"fc",
          3118 => x"82",
          3119 => x"d5",
          3120 => x"78",
          3121 => x"08",
          3122 => x"38",
          3123 => x"70",
          3124 => x"2e",
          3125 => x"82",
          3126 => x"81",
          3127 => x"2e",
          3128 => x"2e",
          3129 => x"82",
          3130 => x"51",
          3131 => x"54",
          3132 => x"9b",
          3133 => x"83",
          3134 => x"0c",
          3135 => x"76",
          3136 => x"82",
          3137 => x"76",
          3138 => x"2e",
          3139 => x"51",
          3140 => x"90",
          3141 => x"e4",
          3142 => x"0d",
          3143 => x"54",
          3144 => x"3f",
          3145 => x"2e",
          3146 => x"2a",
          3147 => x"86",
          3148 => x"54",
          3149 => x"71",
          3150 => x"05",
          3151 => x"06",
          3152 => x"e4",
          3153 => x"3d",
          3154 => x"40",
          3155 => x"ff",
          3156 => x"2e",
          3157 => x"7d",
          3158 => x"08",
          3159 => x"38",
          3160 => x"73",
          3161 => x"8b",
          3162 => x"06",
          3163 => x"d5",
          3164 => x"09",
          3165 => x"d5",
          3166 => x"81",
          3167 => x"07",
          3168 => x"08",
          3169 => x"2e",
          3170 => x"75",
          3171 => x"81",
          3172 => x"06",
          3173 => x"81",
          3174 => x"38",
          3175 => x"70",
          3176 => x"5d",
          3177 => x"81",
          3178 => x"73",
          3179 => x"8c",
          3180 => x"cc",
          3181 => x"ff",
          3182 => x"33",
          3183 => x"05",
          3184 => x"c7",
          3185 => x"a4",
          3186 => x"ff",
          3187 => x"73",
          3188 => x"10",
          3189 => x"81",
          3190 => x"ff",
          3191 => x"17",
          3192 => x"33",
          3193 => x"54",
          3194 => x"81",
          3195 => x"53",
          3196 => x"ff",
          3197 => x"53",
          3198 => x"74",
          3199 => x"08",
          3200 => x"a7",
          3201 => x"39",
          3202 => x"82",
          3203 => x"08",
          3204 => x"38",
          3205 => x"7a",
          3206 => x"04",
          3207 => x"59",
          3208 => x"82",
          3209 => x"08",
          3210 => x"5c",
          3211 => x"08",
          3212 => x"d5",
          3213 => x"83",
          3214 => x"57",
          3215 => x"f6",
          3216 => x"81",
          3217 => x"34",
          3218 => x"74",
          3219 => x"74",
          3220 => x"38",
          3221 => x"f7",
          3222 => x"70",
          3223 => x"a1",
          3224 => x"51",
          3225 => x"17",
          3226 => x"1c",
          3227 => x"75",
          3228 => x"38",
          3229 => x"09",
          3230 => x"08",
          3231 => x"82",
          3232 => x"55",
          3233 => x"bf",
          3234 => x"81",
          3235 => x"33",
          3236 => x"d5",
          3237 => x"79",
          3238 => x"26",
          3239 => x"a0",
          3240 => x"1e",
          3241 => x"55",
          3242 => x"e4",
          3243 => x"38",
          3244 => x"ff",
          3245 => x"1b",
          3246 => x"76",
          3247 => x"51",
          3248 => x"73",
          3249 => x"70",
          3250 => x"1c",
          3251 => x"39",
          3252 => x"7b",
          3253 => x"82",
          3254 => x"73",
          3255 => x"81",
          3256 => x"a0",
          3257 => x"b0",
          3258 => x"9e",
          3259 => x"1a",
          3260 => x"3f",
          3261 => x"e4",
          3262 => x"82",
          3263 => x"ee",
          3264 => x"33",
          3265 => x"55",
          3266 => x"08",
          3267 => x"2e",
          3268 => x"70",
          3269 => x"53",
          3270 => x"53",
          3271 => x"cb",
          3272 => x"2e",
          3273 => x"1b",
          3274 => x"56",
          3275 => x"e3",
          3276 => x"38",
          3277 => x"ff",
          3278 => x"38",
          3279 => x"59",
          3280 => x"10",
          3281 => x"70",
          3282 => x"80",
          3283 => x"32",
          3284 => x"db",
          3285 => x"84",
          3286 => x"07",
          3287 => x"38",
          3288 => x"16",
          3289 => x"56",
          3290 => x"17",
          3291 => x"27",
          3292 => x"2e",
          3293 => x"54",
          3294 => x"80",
          3295 => x"74",
          3296 => x"15",
          3297 => x"19",
          3298 => x"3d",
          3299 => x"81",
          3300 => x"26",
          3301 => x"33",
          3302 => x"75",
          3303 => x"3f",
          3304 => x"1b",
          3305 => x"38",
          3306 => x"f0",
          3307 => x"d5",
          3308 => x"82",
          3309 => x"ab",
          3310 => x"70",
          3311 => x"5e",
          3312 => x"8d",
          3313 => x"3f",
          3314 => x"52",
          3315 => x"e4",
          3316 => x"9e",
          3317 => x"81",
          3318 => x"08",
          3319 => x"dd",
          3320 => x"d5",
          3321 => x"51",
          3322 => x"81",
          3323 => x"7b",
          3324 => x"08",
          3325 => x"38",
          3326 => x"81",
          3327 => x"17",
          3328 => x"d5",
          3329 => x"e4",
          3330 => x"3f",
          3331 => x"55",
          3332 => x"74",
          3333 => x"51",
          3334 => x"33",
          3335 => x"85",
          3336 => x"57",
          3337 => x"ff",
          3338 => x"70",
          3339 => x"80",
          3340 => x"0b",
          3341 => x"ef",
          3342 => x"82",
          3343 => x"19",
          3344 => x"08",
          3345 => x"d5",
          3346 => x"ae",
          3347 => x"52",
          3348 => x"8b",
          3349 => x"51",
          3350 => x"1b",
          3351 => x"16",
          3352 => x"55",
          3353 => x"0d",
          3354 => x"90",
          3355 => x"57",
          3356 => x"52",
          3357 => x"e4",
          3358 => x"c9",
          3359 => x"e1",
          3360 => x"82",
          3361 => x"08",
          3362 => x"17",
          3363 => x"38",
          3364 => x"ee",
          3365 => x"82",
          3366 => x"73",
          3367 => x"82",
          3368 => x"3d",
          3369 => x"71",
          3370 => x"19",
          3371 => x"e2",
          3372 => x"bb",
          3373 => x"08",
          3374 => x"72",
          3375 => x"14",
          3376 => x"7a",
          3377 => x"83",
          3378 => x"ff",
          3379 => x"39",
          3380 => x"31",
          3381 => x"90",
          3382 => x"3f",
          3383 => x"06",
          3384 => x"81",
          3385 => x"53",
          3386 => x"82",
          3387 => x"70",
          3388 => x"07",
          3389 => x"38",
          3390 => x"81",
          3391 => x"1d",
          3392 => x"54",
          3393 => x"70",
          3394 => x"51",
          3395 => x"0b",
          3396 => x"58",
          3397 => x"33",
          3398 => x"2e",
          3399 => x"06",
          3400 => x"32",
          3401 => x"51",
          3402 => x"72",
          3403 => x"81",
          3404 => x"76",
          3405 => x"57",
          3406 => x"17",
          3407 => x"34",
          3408 => x"38",
          3409 => x"34",
          3410 => x"89",
          3411 => x"2e",
          3412 => x"55",
          3413 => x"55",
          3414 => x"08",
          3415 => x"27",
          3416 => x"39",
          3417 => x"53",
          3418 => x"70",
          3419 => x"76",
          3420 => x"81",
          3421 => x"55",
          3422 => x"94",
          3423 => x"9c",
          3424 => x"72",
          3425 => x"1c",
          3426 => x"34",
          3427 => x"d9",
          3428 => x"0c",
          3429 => x"d5",
          3430 => x"51",
          3431 => x"84",
          3432 => x"3d",
          3433 => x"64",
          3434 => x"2e",
          3435 => x"2e",
          3436 => x"7f",
          3437 => x"39",
          3438 => x"56",
          3439 => x"06",
          3440 => x"32",
          3441 => x"51",
          3442 => x"1f",
          3443 => x"9f",
          3444 => x"1f",
          3445 => x"3f",
          3446 => x"39",
          3447 => x"5b",
          3448 => x"51",
          3449 => x"ff",
          3450 => x"0b",
          3451 => x"78",
          3452 => x"2a",
          3453 => x"59",
          3454 => x"06",
          3455 => x"27",
          3456 => x"56",
          3457 => x"ae",
          3458 => x"75",
          3459 => x"3f",
          3460 => x"78",
          3461 => x"10",
          3462 => x"59",
          3463 => x"61",
          3464 => x"2e",
          3465 => x"73",
          3466 => x"25",
          3467 => x"38",
          3468 => x"57",
          3469 => x"38",
          3470 => x"38",
          3471 => x"81",
          3472 => x"54",
          3473 => x"c1",
          3474 => x"09",
          3475 => x"54",
          3476 => x"56",
          3477 => x"38",
          3478 => x"57",
          3479 => x"e9",
          3480 => x"1f",
          3481 => x"a8",
          3482 => x"74",
          3483 => x"70",
          3484 => x"58",
          3485 => x"73",
          3486 => x"38",
          3487 => x"74",
          3488 => x"90",
          3489 => x"39",
          3490 => x"06",
          3491 => x"81",
          3492 => x"1b",
          3493 => x"2e",
          3494 => x"ff",
          3495 => x"81",
          3496 => x"78",
          3497 => x"05",
          3498 => x"9d",
          3499 => x"ff",
          3500 => x"fe",
          3501 => x"2e",
          3502 => x"a0",
          3503 => x"80",
          3504 => x"1a",
          3505 => x"75",
          3506 => x"2e",
          3507 => x"70",
          3508 => x"2e",
          3509 => x"76",
          3510 => x"73",
          3511 => x"5b",
          3512 => x"07",
          3513 => x"55",
          3514 => x"8b",
          3515 => x"8b",
          3516 => x"26",
          3517 => x"8b",
          3518 => x"5f",
          3519 => x"af",
          3520 => x"52",
          3521 => x"d5",
          3522 => x"87",
          3523 => x"73",
          3524 => x"06",
          3525 => x"81",
          3526 => x"54",
          3527 => x"07",
          3528 => x"18",
          3529 => x"73",
          3530 => x"39",
          3531 => x"82",
          3532 => x"d5",
          3533 => x"df",
          3534 => x"ff",
          3535 => x"38",
          3536 => x"54",
          3537 => x"07",
          3538 => x"58",
          3539 => x"75",
          3540 => x"39",
          3541 => x"2e",
          3542 => x"a0",
          3543 => x"06",
          3544 => x"06",
          3545 => x"2e",
          3546 => x"83",
          3547 => x"82",
          3548 => x"06",
          3549 => x"06",
          3550 => x"90",
          3551 => x"06",
          3552 => x"76",
          3553 => x"7d",
          3554 => x"08",
          3555 => x"e4",
          3556 => x"e4",
          3557 => x"e8",
          3558 => x"76",
          3559 => x"2e",
          3560 => x"80",
          3561 => x"ab",
          3562 => x"74",
          3563 => x"56",
          3564 => x"06",
          3565 => x"33",
          3566 => x"55",
          3567 => x"1e",
          3568 => x"05",
          3569 => x"d5",
          3570 => x"39",
          3571 => x"0d",
          3572 => x"7b",
          3573 => x"55",
          3574 => x"75",
          3575 => x"26",
          3576 => x"70",
          3577 => x"06",
          3578 => x"70",
          3579 => x"89",
          3580 => x"ff",
          3581 => x"2e",
          3582 => x"d4",
          3583 => x"76",
          3584 => x"81",
          3585 => x"53",
          3586 => x"13",
          3587 => x"9f",
          3588 => x"e0",
          3589 => x"72",
          3590 => x"72",
          3591 => x"ff",
          3592 => x"70",
          3593 => x"9f",
          3594 => x"80",
          3595 => x"59",
          3596 => x"8b",
          3597 => x"76",
          3598 => x"82",
          3599 => x"e4",
          3600 => x"0d",
          3601 => x"ff",
          3602 => x"51",
          3603 => x"e4",
          3604 => x"51",
          3605 => x"83",
          3606 => x"82",
          3607 => x"e3",
          3608 => x"57",
          3609 => x"83",
          3610 => x"70",
          3611 => x"51",
          3612 => x"2e",
          3613 => x"82",
          3614 => x"cf",
          3615 => x"82",
          3616 => x"85",
          3617 => x"16",
          3618 => x"08",
          3619 => x"83",
          3620 => x"0c",
          3621 => x"61",
          3622 => x"58",
          3623 => x"e1",
          3624 => x"56",
          3625 => x"87",
          3626 => x"29",
          3627 => x"53",
          3628 => x"38",
          3629 => x"74",
          3630 => x"38",
          3631 => x"82",
          3632 => x"81",
          3633 => x"80",
          3634 => x"70",
          3635 => x"86",
          3636 => x"34",
          3637 => x"33",
          3638 => x"33",
          3639 => x"08",
          3640 => x"55",
          3641 => x"80",
          3642 => x"81",
          3643 => x"b8",
          3644 => x"fd",
          3645 => x"ff",
          3646 => x"76",
          3647 => x"d9",
          3648 => x"90",
          3649 => x"56",
          3650 => x"72",
          3651 => x"51",
          3652 => x"57",
          3653 => x"ff",
          3654 => x"25",
          3655 => x"11",
          3656 => x"71",
          3657 => x"f0",
          3658 => x"74",
          3659 => x"90",
          3660 => x"3f",
          3661 => x"57",
          3662 => x"54",
          3663 => x"83",
          3664 => x"38",
          3665 => x"84",
          3666 => x"38",
          3667 => x"38",
          3668 => x"38",
          3669 => x"82",
          3670 => x"53",
          3671 => x"84",
          3672 => x"ec",
          3673 => x"ff",
          3674 => x"14",
          3675 => x"08",
          3676 => x"14",
          3677 => x"33",
          3678 => x"54",
          3679 => x"98",
          3680 => x"29",
          3681 => x"72",
          3682 => x"38",
          3683 => x"2e",
          3684 => x"80",
          3685 => x"d5",
          3686 => x"88",
          3687 => x"56",
          3688 => x"51",
          3689 => x"83",
          3690 => x"80",
          3691 => x"d5",
          3692 => x"c8",
          3693 => x"ff",
          3694 => x"2e",
          3695 => x"14",
          3696 => x"75",
          3697 => x"52",
          3698 => x"3f",
          3699 => x"e4",
          3700 => x"d5",
          3701 => x"26",
          3702 => x"f5",
          3703 => x"f5",
          3704 => x"8d",
          3705 => x"82",
          3706 => x"16",
          3707 => x"7a",
          3708 => x"83",
          3709 => x"e2",
          3710 => x"e4",
          3711 => x"56",
          3712 => x"38",
          3713 => x"82",
          3714 => x"82",
          3715 => x"80",
          3716 => x"15",
          3717 => x"8d",
          3718 => x"76",
          3719 => x"13",
          3720 => x"15",
          3721 => x"94",
          3722 => x"ff",
          3723 => x"2e",
          3724 => x"e8",
          3725 => x"e4",
          3726 => x"81",
          3727 => x"81",
          3728 => x"82",
          3729 => x"d5",
          3730 => x"14",
          3731 => x"08",
          3732 => x"d4",
          3733 => x"38",
          3734 => x"d5",
          3735 => x"2e",
          3736 => x"14",
          3737 => x"08",
          3738 => x"81",
          3739 => x"c5",
          3740 => x"15",
          3741 => x"3f",
          3742 => x"76",
          3743 => x"05",
          3744 => x"86",
          3745 => x"15",
          3746 => x"56",
          3747 => x"0d",
          3748 => x"55",
          3749 => x"53",
          3750 => x"52",
          3751 => x"22",
          3752 => x"2e",
          3753 => x"33",
          3754 => x"e4",
          3755 => x"71",
          3756 => x"53",
          3757 => x"d5",
          3758 => x"3d",
          3759 => x"89",
          3760 => x"3f",
          3761 => x"08",
          3762 => x"84",
          3763 => x"55",
          3764 => x"74",
          3765 => x"38",
          3766 => x"54",
          3767 => x"89",
          3768 => x"e4",
          3769 => x"82",
          3770 => x"ea",
          3771 => x"eb",
          3772 => x"80",
          3773 => x"70",
          3774 => x"3d",
          3775 => x"82",
          3776 => x"08",
          3777 => x"8c",
          3778 => x"82",
          3779 => x"08",
          3780 => x"70",
          3781 => x"83",
          3782 => x"73",
          3783 => x"2e",
          3784 => x"06",
          3785 => x"82",
          3786 => x"b2",
          3787 => x"b8",
          3788 => x"51",
          3789 => x"55",
          3790 => x"74",
          3791 => x"81",
          3792 => x"af",
          3793 => x"3f",
          3794 => x"b2",
          3795 => x"f4",
          3796 => x"34",
          3797 => x"85",
          3798 => x"c2",
          3799 => x"15",
          3800 => x"7a",
          3801 => x"75",
          3802 => x"86",
          3803 => x"d5",
          3804 => x"74",
          3805 => x"70",
          3806 => x"56",
          3807 => x"82",
          3808 => x"06",
          3809 => x"75",
          3810 => x"38",
          3811 => x"7a",
          3812 => x"08",
          3813 => x"55",
          3814 => x"77",
          3815 => x"73",
          3816 => x"07",
          3817 => x"0c",
          3818 => x"52",
          3819 => x"08",
          3820 => x"63",
          3821 => x"82",
          3822 => x"8c",
          3823 => x"17",
          3824 => x"34",
          3825 => x"9c",
          3826 => x"77",
          3827 => x"73",
          3828 => x"e4",
          3829 => x"d5",
          3830 => x"22",
          3831 => x"a8",
          3832 => x"3f",
          3833 => x"e4",
          3834 => x"82",
          3835 => x"06",
          3836 => x"56",
          3837 => x"51",
          3838 => x"70",
          3839 => x"76",
          3840 => x"83",
          3841 => x"38",
          3842 => x"82",
          3843 => x"8e",
          3844 => x"08",
          3845 => x"79",
          3846 => x"0c",
          3847 => x"60",
          3848 => x"80",
          3849 => x"78",
          3850 => x"08",
          3851 => x"91",
          3852 => x"38",
          3853 => x"33",
          3854 => x"2e",
          3855 => x"91",
          3856 => x"81",
          3857 => x"a3",
          3858 => x"31",
          3859 => x"5c",
          3860 => x"19",
          3861 => x"74",
          3862 => x"ff",
          3863 => x"79",
          3864 => x"08",
          3865 => x"78",
          3866 => x"08",
          3867 => x"74",
          3868 => x"1a",
          3869 => x"c3",
          3870 => x"2e",
          3871 => x"1a",
          3872 => x"2e",
          3873 => x"11",
          3874 => x"85",
          3875 => x"76",
          3876 => x"ff",
          3877 => x"fe",
          3878 => x"56",
          3879 => x"08",
          3880 => x"38",
          3881 => x"16",
          3882 => x"51",
          3883 => x"56",
          3884 => x"19",
          3885 => x"31",
          3886 => x"7b",
          3887 => x"c0",
          3888 => x"ff",
          3889 => x"ff",
          3890 => x"ff",
          3891 => x"08",
          3892 => x"08",
          3893 => x"f0",
          3894 => x"0c",
          3895 => x"60",
          3896 => x"80",
          3897 => x"77",
          3898 => x"08",
          3899 => x"91",
          3900 => x"38",
          3901 => x"33",
          3902 => x"56",
          3903 => x"ab",
          3904 => x"34",
          3905 => x"91",
          3906 => x"94",
          3907 => x"76",
          3908 => x"80",
          3909 => x"70",
          3910 => x"82",
          3911 => x"77",
          3912 => x"38",
          3913 => x"74",
          3914 => x"18",
          3915 => x"82",
          3916 => x"08",
          3917 => x"2e",
          3918 => x"95",
          3919 => x"08",
          3920 => x"55",
          3921 => x"09",
          3922 => x"bd",
          3923 => x"ed",
          3924 => x"ff",
          3925 => x"80",
          3926 => x"08",
          3927 => x"80",
          3928 => x"8a",
          3929 => x"27",
          3930 => x"54",
          3931 => x"51",
          3932 => x"08",
          3933 => x"78",
          3934 => x"38",
          3935 => x"31",
          3936 => x"51",
          3937 => x"0b",
          3938 => x"80",
          3939 => x"08",
          3940 => x"f6",
          3941 => x"38",
          3942 => x"9c",
          3943 => x"06",
          3944 => x"76",
          3945 => x"08",
          3946 => x"82",
          3947 => x"53",
          3948 => x"06",
          3949 => x"3f",
          3950 => x"7b",
          3951 => x"76",
          3952 => x"1c",
          3953 => x"5c",
          3954 => x"74",
          3955 => x"18",
          3956 => x"19",
          3957 => x"0c",
          3958 => x"7a",
          3959 => x"56",
          3960 => x"57",
          3961 => x"90",
          3962 => x"06",
          3963 => x"ee",
          3964 => x"ff",
          3965 => x"57",
          3966 => x"a4",
          3967 => x"55",
          3968 => x"08",
          3969 => x"a5",
          3970 => x"51",
          3971 => x"0a",
          3972 => x"3f",
          3973 => x"c6",
          3974 => x"34",
          3975 => x"d5",
          3976 => x"06",
          3977 => x"82",
          3978 => x"fc",
          3979 => x"d4",
          3980 => x"d5",
          3981 => x"05",
          3982 => x"d5",
          3983 => x"87",
          3984 => x"72",
          3985 => x"04",
          3986 => x"89",
          3987 => x"e4",
          3988 => x"08",
          3989 => x"82",
          3990 => x"ee",
          3991 => x"05",
          3992 => x"82",
          3993 => x"08",
          3994 => x"94",
          3995 => x"82",
          3996 => x"08",
          3997 => x"70",
          3998 => x"89",
          3999 => x"b2",
          4000 => x"2a",
          4001 => x"80",
          4002 => x"52",
          4003 => x"08",
          4004 => x"e4",
          4005 => x"38",
          4006 => x"94",
          4007 => x"80",
          4008 => x"5b",
          4009 => x"df",
          4010 => x"3d",
          4011 => x"08",
          4012 => x"38",
          4013 => x"98",
          4014 => x"58",
          4015 => x"2e",
          4016 => x"3d",
          4017 => x"d5",
          4018 => x"82",
          4019 => x"7b",
          4020 => x"e4",
          4021 => x"d8",
          4022 => x"51",
          4023 => x"80",
          4024 => x"c3",
          4025 => x"82",
          4026 => x"52",
          4027 => x"e4",
          4028 => x"38",
          4029 => x"c8",
          4030 => x"2e",
          4031 => x"e8",
          4032 => x"d5",
          4033 => x"84",
          4034 => x"57",
          4035 => x"80",
          4036 => x"51",
          4037 => x"11",
          4038 => x"73",
          4039 => x"05",
          4040 => x"56",
          4041 => x"54",
          4042 => x"80",
          4043 => x"55",
          4044 => x"ff",
          4045 => x"74",
          4046 => x"18",
          4047 => x"af",
          4048 => x"2e",
          4049 => x"80",
          4050 => x"74",
          4051 => x"70",
          4052 => x"08",
          4053 => x"73",
          4054 => x"1a",
          4055 => x"38",
          4056 => x"38",
          4057 => x"74",
          4058 => x"05",
          4059 => x"ba",
          4060 => x"ff",
          4061 => x"57",
          4062 => x"81",
          4063 => x"81",
          4064 => x"38",
          4065 => x"0c",
          4066 => x"0d",
          4067 => x"71",
          4068 => x"d5",
          4069 => x"82",
          4070 => x"82",
          4071 => x"76",
          4072 => x"81",
          4073 => x"72",
          4074 => x"54",
          4075 => x"78",
          4076 => x"22",
          4077 => x"78",
          4078 => x"51",
          4079 => x"08",
          4080 => x"53",
          4081 => x"08",
          4082 => x"75",
          4083 => x"31",
          4084 => x"b2",
          4085 => x"38",
          4086 => x"3f",
          4087 => x"e4",
          4088 => x"d5",
          4089 => x"82",
          4090 => x"98",
          4091 => x"38",
          4092 => x"77",
          4093 => x"0c",
          4094 => x"81",
          4095 => x"2e",
          4096 => x"bb",
          4097 => x"82",
          4098 => x"e4",
          4099 => x"51",
          4100 => x"08",
          4101 => x"74",
          4102 => x"14",
          4103 => x"0c",
          4104 => x"94",
          4105 => x"72",
          4106 => x"51",
          4107 => x"08",
          4108 => x"82",
          4109 => x"16",
          4110 => x"2a",
          4111 => x"15",
          4112 => x"90",
          4113 => x"33",
          4114 => x"34",
          4115 => x"2e",
          4116 => x"85",
          4117 => x"72",
          4118 => x"04",
          4119 => x"75",
          4120 => x"89",
          4121 => x"05",
          4122 => x"08",
          4123 => x"38",
          4124 => x"d4",
          4125 => x"82",
          4126 => x"16",
          4127 => x"74",
          4128 => x"84",
          4129 => x"73",
          4130 => x"52",
          4131 => x"e4",
          4132 => x"14",
          4133 => x"51",
          4134 => x"08",
          4135 => x"85",
          4136 => x"2e",
          4137 => x"73",
          4138 => x"04",
          4139 => x"05",
          4140 => x"82",
          4141 => x"e4",
          4142 => x"fb",
          4143 => x"05",
          4144 => x"3f",
          4145 => x"e4",
          4146 => x"82",
          4147 => x"bb",
          4148 => x"80",
          4149 => x"73",
          4150 => x"08",
          4151 => x"09",
          4152 => x"39",
          4153 => x"52",
          4154 => x"73",
          4155 => x"e4",
          4156 => x"07",
          4157 => x"06",
          4158 => x"e4",
          4159 => x"0d",
          4160 => x"53",
          4161 => x"82",
          4162 => x"08",
          4163 => x"a6",
          4164 => x"d5",
          4165 => x"05",
          4166 => x"80",
          4167 => x"76",
          4168 => x"51",
          4169 => x"0c",
          4170 => x"63",
          4171 => x"ec",
          4172 => x"3f",
          4173 => x"e4",
          4174 => x"73",
          4175 => x"13",
          4176 => x"26",
          4177 => x"39",
          4178 => x"81",
          4179 => x"33",
          4180 => x"06",
          4181 => x"76",
          4182 => x"af",
          4183 => x"2e",
          4184 => x"2e",
          4185 => x"70",
          4186 => x"7a",
          4187 => x"54",
          4188 => x"80",
          4189 => x"e4",
          4190 => x"52",
          4191 => x"8e",
          4192 => x"d5",
          4193 => x"33",
          4194 => x"54",
          4195 => x"38",
          4196 => x"82",
          4197 => x"70",
          4198 => x"59",
          4199 => x"51",
          4200 => x"08",
          4201 => x"25",
          4202 => x"75",
          4203 => x"ff",
          4204 => x"94",
          4205 => x"56",
          4206 => x"d5",
          4207 => x"3d",
          4208 => x"70",
          4209 => x"e4",
          4210 => x"aa",
          4211 => x"a2",
          4212 => x"70",
          4213 => x"73",
          4214 => x"08",
          4215 => x"82",
          4216 => x"08",
          4217 => x"ff",
          4218 => x"74",
          4219 => x"98",
          4220 => x"c6",
          4221 => x"09",
          4222 => x"d5",
          4223 => x"85",
          4224 => x"38",
          4225 => x"15",
          4226 => x"53",
          4227 => x"ff",
          4228 => x"56",
          4229 => x"17",
          4230 => x"18",
          4231 => x"91",
          4232 => x"e4",
          4233 => x"0d",
          4234 => x"52",
          4235 => x"d5",
          4236 => x"81",
          4237 => x"52",
          4238 => x"3f",
          4239 => x"e4",
          4240 => x"05",
          4241 => x"51",
          4242 => x"38",
          4243 => x"81",
          4244 => x"70",
          4245 => x"81",
          4246 => x"ba",
          4247 => x"84",
          4248 => x"73",
          4249 => x"82",
          4250 => x"81",
          4251 => x"08",
          4252 => x"54",
          4253 => x"08",
          4254 => x"38",
          4255 => x"ff",
          4256 => x"55",
          4257 => x"55",
          4258 => x"84",
          4259 => x"80",
          4260 => x"82",
          4261 => x"30",
          4262 => x"25",
          4263 => x"38",
          4264 => x"75",
          4265 => x"82",
          4266 => x"78",
          4267 => x"e4",
          4268 => x"a2",
          4269 => x"53",
          4270 => x"3d",
          4271 => x"08",
          4272 => x"38",
          4273 => x"52",
          4274 => x"08",
          4275 => x"88",
          4276 => x"08",
          4277 => x"38",
          4278 => x"2a",
          4279 => x"81",
          4280 => x"3d",
          4281 => x"82",
          4282 => x"d5",
          4283 => x"d5",
          4284 => x"83",
          4285 => x"ff",
          4286 => x"54",
          4287 => x"82",
          4288 => x"b2",
          4289 => x"82",
          4290 => x"53",
          4291 => x"c6",
          4292 => x"34",
          4293 => x"34",
          4294 => x"19",
          4295 => x"78",
          4296 => x"3f",
          4297 => x"d8",
          4298 => x"54",
          4299 => x"53",
          4300 => x"b7",
          4301 => x"15",
          4302 => x"82",
          4303 => x"08",
          4304 => x"64",
          4305 => x"75",
          4306 => x"9d",
          4307 => x"34",
          4308 => x"78",
          4309 => x"e4",
          4310 => x"52",
          4311 => x"82",
          4312 => x"d8",
          4313 => x"d1",
          4314 => x"fc",
          4315 => x"3f",
          4316 => x"e4",
          4317 => x"3d",
          4318 => x"c8",
          4319 => x"82",
          4320 => x"81",
          4321 => x"86",
          4322 => x"a5",
          4323 => x"05",
          4324 => x"77",
          4325 => x"a2",
          4326 => x"51",
          4327 => x"55",
          4328 => x"a1",
          4329 => x"38",
          4330 => x"88",
          4331 => x"08",
          4332 => x"38",
          4333 => x"d5",
          4334 => x"81",
          4335 => x"3d",
          4336 => x"ff",
          4337 => x"8b",
          4338 => x"2a",
          4339 => x"89",
          4340 => x"17",
          4341 => x"34",
          4342 => x"81",
          4343 => x"80",
          4344 => x"38",
          4345 => x"3f",
          4346 => x"ff",
          4347 => x"e4",
          4348 => x"d5",
          4349 => x"9e",
          4350 => x"d8",
          4351 => x"08",
          4352 => x"73",
          4353 => x"63",
          4354 => x"9d",
          4355 => x"34",
          4356 => x"38",
          4357 => x"e4",
          4358 => x"38",
          4359 => x"d5",
          4360 => x"0c",
          4361 => x"02",
          4362 => x"80",
          4363 => x"96",
          4364 => x"d1",
          4365 => x"82",
          4366 => x"5a",
          4367 => x"c5",
          4368 => x"82",
          4369 => x"cf",
          4370 => x"55",
          4371 => x"71",
          4372 => x"74",
          4373 => x"8b",
          4374 => x"15",
          4375 => x"82",
          4376 => x"e4",
          4377 => x"0d",
          4378 => x"05",
          4379 => x"82",
          4380 => x"08",
          4381 => x"94",
          4382 => x"82",
          4383 => x"08",
          4384 => x"81",
          4385 => x"38",
          4386 => x"90",
          4387 => x"ff",
          4388 => x"83",
          4389 => x"3f",
          4390 => x"d5",
          4391 => x"3d",
          4392 => x"99",
          4393 => x"cf",
          4394 => x"d5",
          4395 => x"08",
          4396 => x"80",
          4397 => x"06",
          4398 => x"38",
          4399 => x"3d",
          4400 => x"82",
          4401 => x"08",
          4402 => x"ff",
          4403 => x"57",
          4404 => x"d5",
          4405 => x"5b",
          4406 => x"18",
          4407 => x"81",
          4408 => x"8b",
          4409 => x"75",
          4410 => x"1b",
          4411 => x"2e",
          4412 => x"09",
          4413 => x"80",
          4414 => x"25",
          4415 => x"38",
          4416 => x"11",
          4417 => x"82",
          4418 => x"08",
          4419 => x"80",
          4420 => x"80",
          4421 => x"a7",
          4422 => x"9b",
          4423 => x"0c",
          4424 => x"0d",
          4425 => x"3d",
          4426 => x"cd",
          4427 => x"d5",
          4428 => x"08",
          4429 => x"8a",
          4430 => x"3f",
          4431 => x"9f",
          4432 => x"9d",
          4433 => x"d5",
          4434 => x"c4",
          4435 => x"c0",
          4436 => x"08",
          4437 => x"08",
          4438 => x"2e",
          4439 => x"51",
          4440 => x"08",
          4441 => x"38",
          4442 => x"8a",
          4443 => x"e7",
          4444 => x"74",
          4445 => x"05",
          4446 => x"70",
          4447 => x"70",
          4448 => x"fe",
          4449 => x"55",
          4450 => x"75",
          4451 => x"55",
          4452 => x"a0",
          4453 => x"16",
          4454 => x"42",
          4455 => x"ff",
          4456 => x"54",
          4457 => x"81",
          4458 => x"82",
          4459 => x"08",
          4460 => x"54",
          4461 => x"d5",
          4462 => x"80",
          4463 => x"80",
          4464 => x"ab",
          4465 => x"82",
          4466 => x"82",
          4467 => x"99",
          4468 => x"15",
          4469 => x"ff",
          4470 => x"83",
          4471 => x"3f",
          4472 => x"74",
          4473 => x"04",
          4474 => x"05",
          4475 => x"05",
          4476 => x"b9",
          4477 => x"d5",
          4478 => x"33",
          4479 => x"2e",
          4480 => x"90",
          4481 => x"70",
          4482 => x"38",
          4483 => x"82",
          4484 => x"7e",
          4485 => x"55",
          4486 => x"f6",
          4487 => x"70",
          4488 => x"08",
          4489 => x"5d",
          4490 => x"9c",
          4491 => x"57",
          4492 => x"52",
          4493 => x"15",
          4494 => x"26",
          4495 => x"08",
          4496 => x"e4",
          4497 => x"d5",
          4498 => x"75",
          4499 => x"93",
          4500 => x"2e",
          4501 => x"58",
          4502 => x"38",
          4503 => x"b4",
          4504 => x"09",
          4505 => x"53",
          4506 => x"3f",
          4507 => x"e4",
          4508 => x"ff",
          4509 => x"84",
          4510 => x"12",
          4511 => x"78",
          4512 => x"90",
          4513 => x"90",
          4514 => x"94",
          4515 => x"91",
          4516 => x"84",
          4517 => x"16",
          4518 => x"0c",
          4519 => x"6c",
          4520 => x"33",
          4521 => x"d1",
          4522 => x"e4",
          4523 => x"e4",
          4524 => x"70",
          4525 => x"38",
          4526 => x"82",
          4527 => x"11",
          4528 => x"41",
          4529 => x"ac",
          4530 => x"06",
          4531 => x"74",
          4532 => x"81",
          4533 => x"cc",
          4534 => x"52",
          4535 => x"d5",
          4536 => x"80",
          4537 => x"26",
          4538 => x"74",
          4539 => x"80",
          4540 => x"92",
          4541 => x"38",
          4542 => x"2e",
          4543 => x"78",
          4544 => x"2b",
          4545 => x"38",
          4546 => x"77",
          4547 => x"dc",
          4548 => x"81",
          4549 => x"ff",
          4550 => x"e4",
          4551 => x"51",
          4552 => x"08",
          4553 => x"74",
          4554 => x"8b",
          4555 => x"b2",
          4556 => x"8b",
          4557 => x"92",
          4558 => x"ba",
          4559 => x"82",
          4560 => x"3d",
          4561 => x"ff",
          4562 => x"e4",
          4563 => x"70",
          4564 => x"51",
          4565 => x"55",
          4566 => x"38",
          4567 => x"ff",
          4568 => x"78",
          4569 => x"81",
          4570 => x"80",
          4571 => x"74",
          4572 => x"06",
          4573 => x"62",
          4574 => x"74",
          4575 => x"7d",
          4576 => x"38",
          4577 => x"81",
          4578 => x"74",
          4579 => x"98",
          4580 => x"82",
          4581 => x"80",
          4582 => x"38",
          4583 => x"3f",
          4584 => x"87",
          4585 => x"5c",
          4586 => x"80",
          4587 => x"0a",
          4588 => x"39",
          4589 => x"81",
          4590 => x"74",
          4591 => x"98",
          4592 => x"82",
          4593 => x"80",
          4594 => x"38",
          4595 => x"3f",
          4596 => x"57",
          4597 => x"96",
          4598 => x"10",
          4599 => x"72",
          4600 => x"ff",
          4601 => x"46",
          4602 => x"70",
          4603 => x"06",
          4604 => x"41",
          4605 => x"38",
          4606 => x"39",
          4607 => x"70",
          4608 => x"76",
          4609 => x"7d",
          4610 => x"55",
          4611 => x"08",
          4612 => x"9b",
          4613 => x"f5",
          4614 => x"38",
          4615 => x"38",
          4616 => x"81",
          4617 => x"0b",
          4618 => x"78",
          4619 => x"c0",
          4620 => x"39",
          4621 => x"8f",
          4622 => x"d5",
          4623 => x"78",
          4624 => x"80",
          4625 => x"39",
          4626 => x"06",
          4627 => x"27",
          4628 => x"56",
          4629 => x"80",
          4630 => x"8b",
          4631 => x"ff",
          4632 => x"1b",
          4633 => x"1c",
          4634 => x"8e",
          4635 => x"0b",
          4636 => x"30",
          4637 => x"51",
          4638 => x"3f",
          4639 => x"90",
          4640 => x"93",
          4641 => x"39",
          4642 => x"fc",
          4643 => x"52",
          4644 => x"81",
          4645 => x"c6",
          4646 => x"8d",
          4647 => x"06",
          4648 => x"52",
          4649 => x"3f",
          4650 => x"bc",
          4651 => x"8d",
          4652 => x"ff",
          4653 => x"51",
          4654 => x"80",
          4655 => x"1c",
          4656 => x"80",
          4657 => x"b2",
          4658 => x"fc",
          4659 => x"96",
          4660 => x"80",
          4661 => x"1c",
          4662 => x"ab",
          4663 => x"d4",
          4664 => x"59",
          4665 => x"53",
          4666 => x"3f",
          4667 => x"9c",
          4668 => x"80",
          4669 => x"7a",
          4670 => x"84",
          4671 => x"8c",
          4672 => x"52",
          4673 => x"8a",
          4674 => x"51",
          4675 => x"83",
          4676 => x"82",
          4677 => x"e4",
          4678 => x"ff",
          4679 => x"53",
          4680 => x"3f",
          4681 => x"7f",
          4682 => x"80",
          4683 => x"60",
          4684 => x"81",
          4685 => x"ff",
          4686 => x"51",
          4687 => x"88",
          4688 => x"f8",
          4689 => x"55",
          4690 => x"3f",
          4691 => x"83",
          4692 => x"7a",
          4693 => x"82",
          4694 => x"80",
          4695 => x"51",
          4696 => x"78",
          4697 => x"18",
          4698 => x"79",
          4699 => x"55",
          4700 => x"74",
          4701 => x"7f",
          4702 => x"e4",
          4703 => x"78",
          4704 => x"57",
          4705 => x"67",
          4706 => x"57",
          4707 => x"64",
          4708 => x"53",
          4709 => x"3f",
          4710 => x"c4",
          4711 => x"83",
          4712 => x"e4",
          4713 => x"85",
          4714 => x"2a",
          4715 => x"84",
          4716 => x"89",
          4717 => x"51",
          4718 => x"55",
          4719 => x"34",
          4720 => x"16",
          4721 => x"56",
          4722 => x"a1",
          4723 => x"82",
          4724 => x"56",
          4725 => x"08",
          4726 => x"1b",
          4727 => x"83",
          4728 => x"81",
          4729 => x"ff",
          4730 => x"e4",
          4731 => x"7f",
          4732 => x"82",
          4733 => x"8e",
          4734 => x"82",
          4735 => x"e4",
          4736 => x"0d",
          4737 => x"ff",
          4738 => x"b4",
          4739 => x"81",
          4740 => x"94",
          4741 => x"9c",
          4742 => x"2e",
          4743 => x"58",
          4744 => x"09",
          4745 => x"78",
          4746 => x"82",
          4747 => x"f7",
          4748 => x"05",
          4749 => x"81",
          4750 => x"e7",
          4751 => x"24",
          4752 => x"8c",
          4753 => x"16",
          4754 => x"3d",
          4755 => x"52",
          4756 => x"76",
          4757 => x"2a",
          4758 => x"84",
          4759 => x"8b",
          4760 => x"84",
          4761 => x"a7",
          4762 => x"53",
          4763 => x"dc",
          4764 => x"84",
          4765 => x"87",
          4766 => x"ff",
          4767 => x"3d",
          4768 => x"80",
          4769 => x"86",
          4770 => x"0d",
          4771 => x"05",
          4772 => x"54",
          4773 => x"fe",
          4774 => x"98",
          4775 => x"02",
          4776 => x"80",
          4777 => x"72",
          4778 => x"39",
          4779 => x"83",
          4780 => x"70",
          4781 => x"22",
          4782 => x"12",
          4783 => x"71",
          4784 => x"82",
          4785 => x"e1",
          4786 => x"06",
          4787 => x"85",
          4788 => x"92",
          4789 => x"22",
          4790 => x"26",
          4791 => x"83",
          4792 => x"70",
          4793 => x"82",
          4794 => x"72",
          4795 => x"04",
          4796 => x"ff",
          4797 => x"ff",
          4798 => x"9f",
          4799 => x"9c",
          4800 => x"70",
          4801 => x"07",
          4802 => x"75",
          4803 => x"2a",
          4804 => x"52",
          4805 => x"38",
          4806 => x"84",
          4807 => x"08",
          4808 => x"70",
          4809 => x"71",
          4810 => x"51",
          4811 => x"39",
          4812 => x"51",
          4813 => x"88",
          4814 => x"51",
          4815 => x"83",
          4816 => x"fe",
          4817 => x"f1",
          4818 => x"0c",
          4819 => x"ff",
          4820 => x"ff",
          4821 => x"51",
          4822 => x"dc",
          4823 => x"ea",
          4824 => x"f8",
          4825 => x"06",
          4826 => x"14",
          4827 => x"21",
          4828 => x"2d",
          4829 => x"39",
          4830 => x"45",
          4831 => x"33",
          4832 => x"3f",
          4833 => x"4b",
          4834 => x"29",
          4835 => x"92",
          4836 => x"fe",
          4837 => x"63",
          4838 => x"db",
          4839 => x"e4",
          4840 => x"3a",
          4841 => x"02",
          4842 => x"fe",
          4843 => x"db",
          4844 => x"92",
          4845 => x"4f",
          4846 => x"60",
          4847 => x"6a",
          4848 => x"74",
          4849 => x"31",
          4850 => x"1a",
          4851 => x"1a",
          4852 => x"1a",
          4853 => x"1a",
          4854 => x"1a",
          4855 => x"1a",
          4856 => x"78",
          4857 => x"1a",
          4858 => x"1a",
          4859 => x"1a",
          4860 => x"1a",
          4861 => x"1a",
          4862 => x"1a",
          4863 => x"1a",
          4864 => x"1a",
          4865 => x"1a",
          4866 => x"1a",
          4867 => x"1a",
          4868 => x"1a",
          4869 => x"1a",
          4870 => x"1a",
          4871 => x"1a",
          4872 => x"1a",
          4873 => x"1a",
          4874 => x"1a",
          4875 => x"1a",
          4876 => x"1a",
          4877 => x"16",
          4878 => x"1a",
          4879 => x"1a",
          4880 => x"1a",
          4881 => x"1a",
          4882 => x"1a",
          4883 => x"3f",
          4884 => x"af",
          4885 => x"1a",
          4886 => x"1a",
          4887 => x"98",
          4888 => x"1a",
          4889 => x"f7",
          4890 => x"1a",
          4891 => x"1a",
          4892 => x"1a",
          4893 => x"16",
          4894 => x"00",
          4895 => x"00",
          4896 => x"00",
          4897 => x"00",
          4898 => x"00",
          4899 => x"00",
          4900 => x"00",
          4901 => x"00",
          4902 => x"00",
          4903 => x"00",
          4904 => x"00",
          4905 => x"00",
          4906 => x"6c",
          4907 => x"00",
          4908 => x"00",
          4909 => x"00",
          4910 => x"00",
          4911 => x"00",
          4912 => x"00",
          4913 => x"00",
          4914 => x"00",
          4915 => x"6b",
          4916 => x"00",
          4917 => x"6c",
          4918 => x"00",
          4919 => x"74",
          4920 => x"00",
          4921 => x"20",
          4922 => x"00",
          4923 => x"20",
          4924 => x"00",
          4925 => x"20",
          4926 => x"65",
          4927 => x"65",
          4928 => x"65",
          4929 => x"65",
          4930 => x"79",
          4931 => x"2e",
          4932 => x"65",
          4933 => x"20",
          4934 => x"2e",
          4935 => x"69",
          4936 => x"20",
          4937 => x"65",
          4938 => x"76",
          4939 => x"72",
          4940 => x"61",
          4941 => x"00",
          4942 => x"74",
          4943 => x"64",
          4944 => x"63",
          4945 => x"6c",
          4946 => x"79",
          4947 => x"75",
          4948 => x"69",
          4949 => x"6d",
          4950 => x"74",
          4951 => x"65",
          4952 => x"65",
          4953 => x"63",
          4954 => x"64",
          4955 => x"65",
          4956 => x"6b",
          4957 => x"75",
          4958 => x"74",
          4959 => x"2e",
          4960 => x"20",
          4961 => x"65",
          4962 => x"2e",
          4963 => x"61",
          4964 => x"69",
          4965 => x"74",
          4966 => x"63",
          4967 => x"00",
          4968 => x"20",
          4969 => x"00",
          4970 => x"74",
          4971 => x"74",
          4972 => x"74",
          4973 => x"0a",
          4974 => x"64",
          4975 => x"6c",
          4976 => x"00",
          4977 => x"00",
          4978 => x"20",
          4979 => x"58",
          4980 => x"00",
          4981 => x"00",
          4982 => x"20",
          4983 => x"00",
          4984 => x"30",
          4985 => x"31",
          4986 => x"55",
          4987 => x"30",
          4988 => x"25",
          4989 => x"00",
          4990 => x"65",
          4991 => x"61",
          4992 => x"00",
          4993 => x"6e",
          4994 => x"00",
          4995 => x"65",
          4996 => x"00",
          4997 => x"44",
          4998 => x"75",
          4999 => x"54",
          5000 => x"74",
          5001 => x"00",
          5002 => x"58",
          5003 => x"75",
          5004 => x"54",
          5005 => x"74",
          5006 => x"00",
          5007 => x"58",
          5008 => x"75",
          5009 => x"54",
          5010 => x"74",
          5011 => x"00",
          5012 => x"20",
          5013 => x"72",
          5014 => x"62",
          5015 => x"6d",
          5016 => x"00",
          5017 => x"63",
          5018 => x"00",
          5019 => x"2e",
          5020 => x"00",
          5021 => x"74",
          5022 => x"61",
          5023 => x"20",
          5024 => x"20",
          5025 => x"69",
          5026 => x"75",
          5027 => x"00",
          5028 => x"61",
          5029 => x"2e",
          5030 => x"79",
          5031 => x"00",
          5032 => x"6e",
          5033 => x"00",
          5034 => x"30",
          5035 => x"38",
          5036 => x"29",
          5037 => x"70",
          5038 => x"00",
          5039 => x"74",
          5040 => x"6c",
          5041 => x"00",
          5042 => x"6c",
          5043 => x"00",
          5044 => x"30",
          5045 => x"00",
          5046 => x"6e",
          5047 => x"40",
          5048 => x"2e",
          5049 => x"6c",
          5050 => x"65",
          5051 => x"78",
          5052 => x"00",
          5053 => x"74",
          5054 => x"6f",
          5055 => x"2e",
          5056 => x"74",
          5057 => x"61",
          5058 => x"69",
          5059 => x"00",
          5060 => x"62",
          5061 => x"2e",
          5062 => x"00",
          5063 => x"5c",
          5064 => x"73",
          5065 => x"5c",
          5066 => x"00",
          5067 => x"00",
          5068 => x"6d",
          5069 => x"00",
          5070 => x"65",
          5071 => x"64",
          5072 => x"74",
          5073 => x"73",
          5074 => x"64",
          5075 => x"6e",
          5076 => x"00",
          5077 => x"67",
          5078 => x"75",
          5079 => x"00",
          5080 => x"64",
          5081 => x"25",
          5082 => x"00",
          5083 => x"66",
          5084 => x"6f",
          5085 => x"72",
          5086 => x"63",
          5087 => x"00",
          5088 => x"65",
          5089 => x"6d",
          5090 => x"00",
          5091 => x"53",
          5092 => x"25",
          5093 => x"58",
          5094 => x"20",
          5095 => x"20",
          5096 => x"3a",
          5097 => x"00",
          5098 => x"4e",
          5099 => x"25",
          5100 => x"58",
          5101 => x"20",
          5102 => x"20",
          5103 => x"3a",
          5104 => x"00",
          5105 => x"20",
          5106 => x"25",
          5107 => x"58",
          5108 => x"20",
          5109 => x"20",
          5110 => x"63",
          5111 => x"64",
          5112 => x"20",
          5113 => x"20",
          5114 => x"72",
          5115 => x"64",
          5116 => x"20",
          5117 => x"52",
          5118 => x"6e",
          5119 => x"64",
          5120 => x"20",
          5121 => x"45",
          5122 => x"00",
          5123 => x"49",
          5124 => x"20",
          5125 => x"00",
          5126 => x"00",
          5127 => x"00",
          5128 => x"65",
          5129 => x"20",
          5130 => x"65",
          5131 => x"72",
          5132 => x"73",
          5133 => x"0a",
          5134 => x"20",
          5135 => x"6f",
          5136 => x"74",
          5137 => x"73",
          5138 => x"0a",
          5139 => x"20",
          5140 => x"74",
          5141 => x"72",
          5142 => x"20",
          5143 => x"0a",
          5144 => x"63",
          5145 => x"20",
          5146 => x"20",
          5147 => x"20",
          5148 => x"20",
          5149 => x"0a",
          5150 => x"20",
          5151 => x"43",
          5152 => x"65",
          5153 => x"20",
          5154 => x"30",
          5155 => x"00",
          5156 => x"41",
          5157 => x"20",
          5158 => x"20",
          5159 => x"25",
          5160 => x"48",
          5161 => x"20",
          5162 => x"65",
          5163 => x"43",
          5164 => x"65",
          5165 => x"30",
          5166 => x"00",
          5167 => x"00",
          5168 => x"00",
          5169 => x"00",
          5170 => x"6d",
          5171 => x"6e",
          5172 => x"00",
          5173 => x"02",
          5174 => x"00",
          5175 => x"f8",
          5176 => x"04",
          5177 => x"00",
          5178 => x"f0",
          5179 => x"06",
          5180 => x"00",
          5181 => x"e8",
          5182 => x"01",
          5183 => x"00",
          5184 => x"e0",
          5185 => x"0b",
          5186 => x"00",
          5187 => x"d8",
          5188 => x"0a",
          5189 => x"00",
          5190 => x"d0",
          5191 => x"0c",
          5192 => x"00",
          5193 => x"c8",
          5194 => x"0f",
          5195 => x"00",
          5196 => x"c0",
          5197 => x"10",
          5198 => x"00",
          5199 => x"b8",
          5200 => x"12",
          5201 => x"00",
          5202 => x"b0",
          5203 => x"14",
          5204 => x"00",
          5205 => x"00",
          5206 => x"00",
          5207 => x"7e",
          5208 => x"7e",
          5209 => x"7e",
          5210 => x"7e",
          5211 => x"00",
          5212 => x"00",
          5213 => x"00",
          5214 => x"00",
          5215 => x"00",
          5216 => x"74",
          5217 => x"74",
          5218 => x"00",
          5219 => x"25",
          5220 => x"6c",
          5221 => x"65",
          5222 => x"20",
          5223 => x"20",
          5224 => x"20",
          5225 => x"00",
          5226 => x"6f",
          5227 => x"61",
          5228 => x"6f",
          5229 => x"2c",
          5230 => x"69",
          5231 => x"00",
          5232 => x"7f",
          5233 => x"3d",
          5234 => x"00",
          5235 => x"00",
          5236 => x"53",
          5237 => x"4e",
          5238 => x"46",
          5239 => x"00",
          5240 => x"20",
          5241 => x"20",
          5242 => x"7c",
          5243 => x"00",
          5244 => x"07",
          5245 => x"1c",
          5246 => x"41",
          5247 => x"49",
          5248 => x"4f",
          5249 => x"9b",
          5250 => x"55",
          5251 => x"ab",
          5252 => x"b3",
          5253 => x"bb",
          5254 => x"c3",
          5255 => x"cb",
          5256 => x"d3",
          5257 => x"db",
          5258 => x"e3",
          5259 => x"eb",
          5260 => x"f3",
          5261 => x"fb",
          5262 => x"3b",
          5263 => x"3a",
          5264 => x"00",
          5265 => x"40",
          5266 => x"00",
          5267 => x"08",
          5268 => x"00",
          5269 => x"e2",
          5270 => x"e7",
          5271 => x"ef",
          5272 => x"c5",
          5273 => x"f4",
          5274 => x"f9",
          5275 => x"a2",
          5276 => x"92",
          5277 => x"fa",
          5278 => x"ba",
          5279 => x"bd",
          5280 => x"bb",
          5281 => x"02",
          5282 => x"56",
          5283 => x"57",
          5284 => x"10",
          5285 => x"1c",
          5286 => x"5f",
          5287 => x"66",
          5288 => x"67",
          5289 => x"59",
          5290 => x"6b",
          5291 => x"88",
          5292 => x"80",
          5293 => x"c0",
          5294 => x"c4",
          5295 => x"b4",
          5296 => x"29",
          5297 => x"64",
          5298 => x"48",
          5299 => x"1a",
          5300 => x"a0",
          5301 => x"17",
          5302 => x"01",
          5303 => x"32",
          5304 => x"4a",
          5305 => x"80",
          5306 => x"82",
          5307 => x"86",
          5308 => x"8a",
          5309 => x"8e",
          5310 => x"91",
          5311 => x"96",
          5312 => x"3d",
          5313 => x"20",
          5314 => x"a2",
          5315 => x"a6",
          5316 => x"aa",
          5317 => x"ae",
          5318 => x"b2",
          5319 => x"b5",
          5320 => x"ba",
          5321 => x"be",
          5322 => x"c2",
          5323 => x"c4",
          5324 => x"ca",
          5325 => x"10",
          5326 => x"de",
          5327 => x"f1",
          5328 => x"28",
          5329 => x"09",
          5330 => x"3d",
          5331 => x"41",
          5332 => x"53",
          5333 => x"55",
          5334 => x"8f",
          5335 => x"5d",
          5336 => x"61",
          5337 => x"65",
          5338 => x"96",
          5339 => x"6d",
          5340 => x"71",
          5341 => x"9f",
          5342 => x"79",
          5343 => x"64",
          5344 => x"81",
          5345 => x"85",
          5346 => x"44",
          5347 => x"8d",
          5348 => x"91",
          5349 => x"fd",
          5350 => x"04",
          5351 => x"8a",
          5352 => x"02",
          5353 => x"08",
          5354 => x"8e",
          5355 => x"f2",
          5356 => x"f4",
          5357 => x"f7",
          5358 => x"30",
          5359 => x"60",
          5360 => x"c1",
          5361 => x"c0",
          5362 => x"26",
          5363 => x"01",
          5364 => x"a0",
          5365 => x"10",
          5366 => x"30",
          5367 => x"51",
          5368 => x"5b",
          5369 => x"5f",
          5370 => x"0e",
          5371 => x"c9",
          5372 => x"db",
          5373 => x"eb",
          5374 => x"08",
          5375 => x"08",
          5376 => x"b9",
          5377 => x"01",
          5378 => x"e0",
          5379 => x"ec",
          5380 => x"4e",
          5381 => x"10",
          5382 => x"d0",
          5383 => x"60",
          5384 => x"75",
          5385 => x"00",
          5386 => x"00",
          5387 => x"f0",
          5388 => x"00",
          5389 => x"f8",
          5390 => x"00",
          5391 => x"00",
          5392 => x"00",
          5393 => x"08",
          5394 => x"00",
          5395 => x"10",
          5396 => x"00",
          5397 => x"18",
          5398 => x"00",
          5399 => x"20",
          5400 => x"00",
          5401 => x"28",
          5402 => x"00",
          5403 => x"30",
          5404 => x"00",
          5405 => x"38",
          5406 => x"00",
          5407 => x"3c",
          5408 => x"00",
          5409 => x"40",
          5410 => x"00",
          5411 => x"44",
          5412 => x"00",
          5413 => x"48",
          5414 => x"00",
          5415 => x"4c",
          5416 => x"00",
          5417 => x"50",
          5418 => x"00",
          5419 => x"54",
          5420 => x"00",
          5421 => x"5c",
          5422 => x"00",
          5423 => x"60",
          5424 => x"00",
          5425 => x"68",
          5426 => x"00",
          5427 => x"70",
          5428 => x"00",
          5429 => x"78",
          5430 => x"00",
          5431 => x"80",
          5432 => x"00",
          5433 => x"88",
          5434 => x"00",
          5435 => x"90",
          5436 => x"00",
          5437 => x"98",
          5438 => x"00",
          5439 => x"00",
          5440 => x"ff",
          5441 => x"ff",
          5442 => x"ff",
          5443 => x"00",
          5444 => x"ff",
          5445 => x"00",
          5446 => x"00",
          5447 => x"00",
          5448 => x"00",
          5449 => x"01",
          5450 => x"00",
          5451 => x"00",
          5452 => x"00",
          5453 => x"00",
          5454 => x"00",
          5455 => x"00",
          5456 => x"00",
          5457 => x"00",
          5458 => x"00",
          5459 => x"00",
          5460 => x"00",
          5461 => x"00",
          5462 => x"00",
          5463 => x"00",
          5464 => x"00",
          5465 => x"00",
          5466 => x"00",
          5467 => x"04",
          5468 => x"04",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"82",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a4",
           135 => x"0b",
           136 => x"0b",
           137 => x"e0",
           138 => x"0b",
           139 => x"0b",
           140 => x"9e",
           141 => x"0b",
           142 => x"0b",
           143 => x"dd",
           144 => x"0b",
           145 => x"0b",
           146 => x"9d",
           147 => x"0b",
           148 => x"0b",
           149 => x"dd",
           150 => x"0b",
           151 => x"0b",
           152 => x"9d",
           153 => x"0b",
           154 => x"0b",
           155 => x"dd",
           156 => x"0b",
           157 => x"0b",
           158 => x"9d",
           159 => x"0b",
           160 => x"0b",
           161 => x"dd",
           162 => x"0b",
           163 => x"0b",
           164 => x"9d",
           165 => x"0b",
           166 => x"0b",
           167 => x"dd",
           168 => x"0b",
           169 => x"0b",
           170 => x"9d",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"d5",
           193 => x"d5",
           194 => x"d5",
           195 => x"f0",
           196 => x"f0",
           197 => x"08",
           198 => x"0c",
           199 => x"84",
           200 => x"94",
           201 => x"80",
           202 => x"c2",
           203 => x"90",
           204 => x"f7",
           205 => x"90",
           206 => x"a6",
           207 => x"90",
           208 => x"2d",
           209 => x"04",
           210 => x"82",
           211 => x"82",
           212 => x"d5",
           213 => x"d5",
           214 => x"d5",
           215 => x"d5",
           216 => x"d5",
           217 => x"d5",
           218 => x"d5",
           219 => x"d5",
           220 => x"d5",
           221 => x"d5",
           222 => x"d5",
           223 => x"d5",
           224 => x"d5",
           225 => x"d5",
           226 => x"d5",
           227 => x"d5",
           228 => x"d5",
           229 => x"d5",
           230 => x"d5",
           231 => x"d5",
           232 => x"d5",
           233 => x"d5",
           234 => x"d5",
           235 => x"d5",
           236 => x"d5",
           237 => x"d5",
           238 => x"d5",
           239 => x"d5",
           240 => x"d5",
           241 => x"d5",
           242 => x"d5",
           243 => x"d5",
           244 => x"d5",
           245 => x"d5",
           246 => x"d5",
           247 => x"d5",
           248 => x"d5",
           249 => x"d5",
           250 => x"d5",
           251 => x"d5",
           252 => x"d5",
           253 => x"d5",
           254 => x"d5",
           255 => x"d5",
           256 => x"d5",
           257 => x"d5",
           258 => x"d5",
           259 => x"d5",
           260 => x"d5",
           261 => x"d5",
           262 => x"d5",
           263 => x"d5",
           264 => x"d5",
           265 => x"d5",
           266 => x"d5",
           267 => x"d5",
           268 => x"d5",
           269 => x"d5",
           270 => x"d5",
           271 => x"d5",
           272 => x"d5",
           273 => x"d5",
           274 => x"d5",
           275 => x"d5",
           276 => x"d5",
           277 => x"d5",
           278 => x"d5",
           279 => x"d5",
           280 => x"d5",
           281 => x"d5",
           282 => x"d5",
           283 => x"d5",
           284 => x"d5",
           285 => x"d5",
           286 => x"d5",
           287 => x"d5",
           288 => x"d5",
           289 => x"d5",
           290 => x"d5",
           291 => x"d5",
           292 => x"d5",
           293 => x"d5",
           294 => x"d5",
           295 => x"d5",
           296 => x"d5",
           297 => x"d5",
           298 => x"d5",
           299 => x"04",
           300 => x"10",
           301 => x"10",
           302 => x"10",
           303 => x"10",
           304 => x"81",
           305 => x"05",
           306 => x"72",
           307 => x"72",
           308 => x"72",
           309 => x"10",
           310 => x"53",
           311 => x"f1",
           312 => x"84",
           313 => x"bc",
           314 => x"04",
           315 => x"d5",
           316 => x"f0",
           317 => x"08",
           318 => x"fc",
           319 => x"88",
           320 => x"52",
           321 => x"08",
           322 => x"0c",
           323 => x"70",
           324 => x"3d",
           325 => x"d5",
           326 => x"fb",
           327 => x"05",
           328 => x"70",
           329 => x"8f",
           330 => x"8c",
           331 => x"80",
           332 => x"0c",
           333 => x"8c",
           334 => x"08",
           335 => x"f0",
           336 => x"08",
           337 => x"fc",
           338 => x"05",
           339 => x"0b",
           340 => x"25",
           341 => x"90",
           342 => x"d5",
           343 => x"f8",
           344 => x"f8",
           345 => x"8d",
           346 => x"f4",
           347 => x"f0",
           348 => x"08",
           349 => x"34",
           350 => x"ff",
           351 => x"0c",
           352 => x"81",
           353 => x"0c",
           354 => x"fc",
           355 => x"d5",
           356 => x"d5",
           357 => x"d5",
           358 => x"e4",
           359 => x"0c",
           360 => x"d5",
           361 => x"82",
           362 => x"d5",
           363 => x"f0",
           364 => x"82",
           365 => x"d5",
           366 => x"f0",
           367 => x"08",
           368 => x"08",
           369 => x"08",
           370 => x"8d",
           371 => x"d5",
           372 => x"f0",
           373 => x"08",
           374 => x"74",
           375 => x"08",
           376 => x"3d",
           377 => x"d5",
           378 => x"fb",
           379 => x"05",
           380 => x"0c",
           381 => x"54",
           382 => x"53",
           383 => x"52",
           384 => x"70",
           385 => x"82",
           386 => x"82",
           387 => x"0d",
           388 => x"f0",
           389 => x"3d",
           390 => x"e4",
           391 => x"05",
           392 => x"82",
           393 => x"11",
           394 => x"70",
           395 => x"72",
           396 => x"d5",
           397 => x"39",
           398 => x"53",
           399 => x"08",
           400 => x"53",
           401 => x"d5",
           402 => x"82",
           403 => x"d5",
           404 => x"06",
           405 => x"38",
           406 => x"53",
           407 => x"d5",
           408 => x"b9",
           409 => x"08",
           410 => x"09",
           411 => x"f0",
           412 => x"70",
           413 => x"38",
           414 => x"70",
           415 => x"06",
           416 => x"99",
           417 => x"22",
           418 => x"82",
           419 => x"d0",
           420 => x"33",
           421 => x"70",
           422 => x"51",
           423 => x"d5",
           424 => x"f0",
           425 => x"f0",
           426 => x"11",
           427 => x"08",
           428 => x"e8",
           429 => x"2c",
           430 => x"38",
           431 => x"e8",
           432 => x"05",
           433 => x"51",
           434 => x"d5",
           435 => x"2b",
           436 => x"88",
           437 => x"82",
           438 => x"b8",
           439 => x"22",
           440 => x"51",
           441 => x"d5",
           442 => x"2b",
           443 => x"8a",
           444 => x"e8",
           445 => x"05",
           446 => x"c4",
           447 => x"c4",
           448 => x"38",
           449 => x"70",
           450 => x"08",
           451 => x"d5",
           452 => x"07",
           453 => x"e4",
           454 => x"05",
           455 => x"82",
           456 => x"a8",
           457 => x"22",
           458 => x"82",
           459 => x"90",
           460 => x"22",
           461 => x"82",
           462 => x"f8",
           463 => x"22",
           464 => x"d5",
           465 => x"82",
           466 => x"d8",
           467 => x"22",
           468 => x"d5",
           469 => x"39",
           470 => x"05",
           471 => x"22",
           472 => x"f0",
           473 => x"82",
           474 => x"a8",
           475 => x"08",
           476 => x"84",
           477 => x"0c",
           478 => x"f0",
           479 => x"08",
           480 => x"72",
           481 => x"8c",
           482 => x"05",
           483 => x"08",
           484 => x"05",
           485 => x"fc",
           486 => x"05",
           487 => x"51",
           488 => x"38",
           489 => x"70",
           490 => x"82",
           491 => x"53",
           492 => x"53",
           493 => x"23",
           494 => x"05",
           495 => x"e4",
           496 => x"f4",
           497 => x"05",
           498 => x"05",
           499 => x"82",
           500 => x"d8",
           501 => x"08",
           502 => x"84",
           503 => x"0c",
           504 => x"05",
           505 => x"22",
           506 => x"51",
           507 => x"82",
           508 => x"98",
           509 => x"d5",
           510 => x"a2",
           511 => x"72",
           512 => x"99",
           513 => x"08",
           514 => x"08",
           515 => x"05",
           516 => x"22",
           517 => x"22",
           518 => x"d5",
           519 => x"39",
           520 => x"70",
           521 => x"53",
           522 => x"f0",
           523 => x"08",
           524 => x"f0",
           525 => x"d5",
           526 => x"39",
           527 => x"82",
           528 => x"05",
           529 => x"70",
           530 => x"0c",
           531 => x"08",
           532 => x"82",
           533 => x"25",
           534 => x"05",
           535 => x"82",
           536 => x"d5",
           537 => x"d5",
           538 => x"f0",
           539 => x"06",
           540 => x"e4",
           541 => x"82",
           542 => x"39",
           543 => x"70",
           544 => x"d5",
           545 => x"0b",
           546 => x"90",
           547 => x"23",
           548 => x"70",
           549 => x"53",
           550 => x"f0",
           551 => x"08",
           552 => x"f0",
           553 => x"d5",
           554 => x"39",
           555 => x"82",
           556 => x"05",
           557 => x"70",
           558 => x"0c",
           559 => x"08",
           560 => x"82",
           561 => x"cf",
           562 => x"08",
           563 => x"82",
           564 => x"d5",
           565 => x"f0",
           566 => x"08",
           567 => x"56",
           568 => x"e4",
           569 => x"f0",
           570 => x"08",
           571 => x"f0",
           572 => x"73",
           573 => x"f0",
           574 => x"d5",
           575 => x"df",
           576 => x"f0",
           577 => x"d5",
           578 => x"33",
           579 => x"f0",
           580 => x"08",
           581 => x"08",
           582 => x"f0",
           583 => x"d5",
           584 => x"f0",
           585 => x"d5",
           586 => x"a3",
           587 => x"82",
           588 => x"82",
           589 => x"2e",
           590 => x"f0",
           591 => x"54",
           592 => x"51",
           593 => x"05",
           594 => x"22",
           595 => x"2e",
           596 => x"05",
           597 => x"d5",
           598 => x"f0",
           599 => x"70",
           600 => x"2e",
           601 => x"ec",
           602 => x"f0",
           603 => x"08",
           604 => x"f0",
           605 => x"08",
           606 => x"2e",
           607 => x"f0",
           608 => x"72",
           609 => x"93",
           610 => x"08",
           611 => x"08",
           612 => x"c8",
           613 => x"05",
           614 => x"22",
           615 => x"51",
           616 => x"82",
           617 => x"98",
           618 => x"08",
           619 => x"72",
           620 => x"08",
           621 => x"53",
           622 => x"23",
           623 => x"05",
           624 => x"05",
           625 => x"82",
           626 => x"d5",
           627 => x"2a",
           628 => x"80",
           629 => x"e8",
           630 => x"2b",
           631 => x"51",
           632 => x"f0",
           633 => x"51",
           634 => x"05",
           635 => x"fc",
           636 => x"2b",
           637 => x"51",
           638 => x"f0",
           639 => x"51",
           640 => x"05",
           641 => x"22",
           642 => x"b0",
           643 => x"22",
           644 => x"f0",
           645 => x"70",
           646 => x"90",
           647 => x"08",
           648 => x"39",
           649 => x"70",
           650 => x"53",
           651 => x"f0",
           652 => x"8a",
           653 => x"f0",
           654 => x"70",
           655 => x"2e",
           656 => x"05",
           657 => x"a3",
           658 => x"22",
           659 => x"51",
           660 => x"d5",
           661 => x"51",
           662 => x"e4",
           663 => x"06",
           664 => x"38",
           665 => x"52",
           666 => x"f0",
           667 => x"2e",
           668 => x"f0",
           669 => x"f0",
           670 => x"3f",
           671 => x"70",
           672 => x"53",
           673 => x"f0",
           674 => x"54",
           675 => x"23",
           676 => x"53",
           677 => x"f0",
           678 => x"88",
           679 => x"08",
           680 => x"81",
           681 => x"b0",
           682 => x"33",
           683 => x"f0",
           684 => x"70",
           685 => x"90",
           686 => x"08",
           687 => x"39",
           688 => x"70",
           689 => x"53",
           690 => x"ec",
           691 => x"82",
           692 => x"90",
           693 => x"73",
           694 => x"88",
           695 => x"3f",
           696 => x"05",
           697 => x"81",
           698 => x"88",
           699 => x"fc",
           700 => x"ee",
           701 => x"33",
           702 => x"06",
           703 => x"f4",
           704 => x"82",
           705 => x"83",
           706 => x"ff",
           707 => x"08",
           708 => x"08",
           709 => x"d5",
           710 => x"82",
           711 => x"86",
           712 => x"f0",
           713 => x"d3",
           714 => x"82",
           715 => x"11",
           716 => x"f4",
           717 => x"53",
           718 => x"38",
           719 => x"52",
           720 => x"70",
           721 => x"d5",
           722 => x"82",
           723 => x"b7",
           724 => x"08",
           725 => x"d5",
           726 => x"d5",
           727 => x"82",
           728 => x"d5",
           729 => x"52",
           730 => x"d5",
           731 => x"2a",
           732 => x"80",
           733 => x"08",
           734 => x"72",
           735 => x"73",
           736 => x"80",
           737 => x"08",
           738 => x"9b",
           739 => x"88",
           740 => x"f8",
           741 => x"0b",
           742 => x"ea",
           743 => x"05",
           744 => x"06",
           745 => x"08",
           746 => x"f0",
           747 => x"d5",
           748 => x"82",
           749 => x"80",
           750 => x"08",
           751 => x"33",
           752 => x"82",
           753 => x"11",
           754 => x"05",
           755 => x"e0",
           756 => x"3d",
           757 => x"d5",
           758 => x"fd",
           759 => x"82",
           760 => x"82",
           761 => x"e4",
           762 => x"82",
           763 => x"82",
           764 => x"08",
           765 => x"0d",
           766 => x"05",
           767 => x"33",
           768 => x"81",
           769 => x"80",
           770 => x"f0",
           771 => x"82",
           772 => x"72",
           773 => x"08",
           774 => x"05",
           775 => x"fc",
           776 => x"72",
           777 => x"08",
           778 => x"f0",
           779 => x"08",
           780 => x"08",
           781 => x"ff",
           782 => x"0c",
           783 => x"82",
           784 => x"90",
           785 => x"e4",
           786 => x"ff",
           787 => x"0c",
           788 => x"70",
           789 => x"53",
           790 => x"82",
           791 => x"d5",
           792 => x"02",
           793 => x"80",
           794 => x"0c",
           795 => x"85",
           796 => x"32",
           797 => x"53",
           798 => x"82",
           799 => x"f3",
           800 => x"08",
           801 => x"88",
           802 => x"08",
           803 => x"f0",
           804 => x"06",
           805 => x"d5",
           806 => x"f0",
           807 => x"f0",
           808 => x"08",
           809 => x"08",
           810 => x"ff",
           811 => x"0c",
           812 => x"f8",
           813 => x"f4",
           814 => x"f4",
           815 => x"3d",
           816 => x"d5",
           817 => x"fe",
           818 => x"82",
           819 => x"93",
           820 => x"d5",
           821 => x"d5",
           822 => x"02",
           823 => x"82",
           824 => x"11",
           825 => x"70",
           826 => x"72",
           827 => x"d5",
           828 => x"39",
           829 => x"85",
           830 => x"06",
           831 => x"80",
           832 => x"05",
           833 => x"08",
           834 => x"08",
           835 => x"8c",
           836 => x"f0",
           837 => x"54",
           838 => x"74",
           839 => x"08",
           840 => x"0c",
           841 => x"70",
           842 => x"51",
           843 => x"08",
           844 => x"8c",
           845 => x"88",
           846 => x"90",
           847 => x"82",
           848 => x"82",
           849 => x"11",
           850 => x"d5",
           851 => x"d5",
           852 => x"8a",
           853 => x"fc",
           854 => x"05",
           855 => x"0d",
           856 => x"f0",
           857 => x"3d",
           858 => x"08",
           859 => x"81",
           860 => x"2e",
           861 => x"08",
           862 => x"d5",
           863 => x"33",
           864 => x"51",
           865 => x"38",
           866 => x"82",
           867 => x"53",
           868 => x"51",
           869 => x"f0",
           870 => x"81",
           871 => x"08",
           872 => x"82",
           873 => x"51",
           874 => x"08",
           875 => x"82",
           876 => x"52",
           877 => x"d5",
           878 => x"70",
           879 => x"0c",
           880 => x"05",
           881 => x"88",
           882 => x"05",
           883 => x"a0",
           884 => x"ff",
           885 => x"0c",
           886 => x"88",
           887 => x"0c",
           888 => x"08",
           889 => x"88",
           890 => x"52",
           891 => x"82",
           892 => x"82",
           893 => x"25",
           894 => x"88",
           895 => x"05",
           896 => x"08",
           897 => x"f0",
           898 => x"fc",
           899 => x"95",
           900 => x"08",
           901 => x"08",
           902 => x"f0",
           903 => x"71",
           904 => x"82",
           905 => x"82",
           906 => x"13",
           907 => x"f8",
           908 => x"08",
           909 => x"05",
           910 => x"fc",
           911 => x"82",
           912 => x"51",
           913 => x"08",
           914 => x"82",
           915 => x"08",
           916 => x"0d",
           917 => x"82",
           918 => x"d5",
           919 => x"f0",
           920 => x"08",
           921 => x"38",
           922 => x"82",
           923 => x"81",
           924 => x"05",
           925 => x"08",
           926 => x"05",
           927 => x"d5",
           928 => x"f0",
           929 => x"f0",
           930 => x"08",
           931 => x"90",
           932 => x"f8",
           933 => x"05",
           934 => x"90",
           935 => x"05",
           936 => x"90",
           937 => x"05",
           938 => x"d5",
           939 => x"82",
           940 => x"d5",
           941 => x"82",
           942 => x"d5",
           943 => x"f0",
           944 => x"33",
           945 => x"f0",
           946 => x"d5",
           947 => x"f0",
           948 => x"d5",
           949 => x"f0",
           950 => x"38",
           951 => x"51",
           952 => x"05",
           953 => x"f8",
           954 => x"05",
           955 => x"d5",
           956 => x"82",
           957 => x"ad",
           958 => x"08",
           959 => x"3d",
           960 => x"d5",
           961 => x"fe",
           962 => x"05",
           963 => x"0c",
           964 => x"52",
           965 => x"05",
           966 => x"fc",
           967 => x"51",
           968 => x"82",
           969 => x"05",
           970 => x"82",
           971 => x"d5",
           972 => x"82",
           973 => x"82",
           974 => x"08",
           975 => x"0d",
           976 => x"82",
           977 => x"d5",
           978 => x"33",
           979 => x"81",
           980 => x"0c",
           981 => x"53",
           982 => x"08",
           983 => x"f0",
           984 => x"06",
           985 => x"be",
           986 => x"08",
           987 => x"3d",
           988 => x"d5",
           989 => x"fd",
           990 => x"05",
           991 => x"0c",
           992 => x"82",
           993 => x"d5",
           994 => x"80",
           995 => x"05",
           996 => x"90",
           997 => x"05",
           998 => x"90",
           999 => x"05",
          1000 => x"f0",
          1001 => x"82",
          1002 => x"05",
          1003 => x"82",
          1004 => x"52",
          1005 => x"fc",
          1006 => x"08",
          1007 => x"d5",
          1008 => x"d5",
          1009 => x"d5",
          1010 => x"02",
          1011 => x"82",
          1012 => x"2e",
          1013 => x"8c",
          1014 => x"f0",
          1015 => x"d5",
          1016 => x"f0",
          1017 => x"81",
          1018 => x"71",
          1019 => x"d5",
          1020 => x"33",
          1021 => x"81",
          1022 => x"0c",
          1023 => x"8d",
          1024 => x"fc",
          1025 => x"f0",
          1026 => x"d5",
          1027 => x"f0",
          1028 => x"38",
          1029 => x"90",
          1030 => x"82",
          1031 => x"33",
          1032 => x"82",
          1033 => x"d7",
          1034 => x"08",
          1035 => x"05",
          1036 => x"08",
          1037 => x"81",
          1038 => x"0c",
          1039 => x"05",
          1040 => x"8c",
          1041 => x"70",
          1042 => x"53",
          1043 => x"0b",
          1044 => x"82",
          1045 => x"d5",
          1046 => x"f0",
          1047 => x"82",
          1048 => x"d5",
          1049 => x"d5",
          1050 => x"8d",
          1051 => x"d5",
          1052 => x"f0",
          1053 => x"53",
          1054 => x"d5",
          1055 => x"fc",
          1056 => x"fc",
          1057 => x"d5",
          1058 => x"82",
          1059 => x"d5",
          1060 => x"80",
          1061 => x"05",
          1062 => x"05",
          1063 => x"05",
          1064 => x"e4",
          1065 => x"05",
          1066 => x"05",
          1067 => x"0d",
          1068 => x"f0",
          1069 => x"3d",
          1070 => x"08",
          1071 => x"82",
          1072 => x"38",
          1073 => x"05",
          1074 => x"08",
          1075 => x"d5",
          1076 => x"82",
          1077 => x"81",
          1078 => x"9f",
          1079 => x"08",
          1080 => x"05",
          1081 => x"08",
          1082 => x"82",
          1083 => x"05",
          1084 => x"82",
          1085 => x"d5",
          1086 => x"82",
          1087 => x"82",
          1088 => x"d5",
          1089 => x"f0",
          1090 => x"82",
          1091 => x"d5",
          1092 => x"f0",
          1093 => x"08",
          1094 => x"38",
          1095 => x"81",
          1096 => x"0c",
          1097 => x"ff",
          1098 => x"0c",
          1099 => x"80",
          1100 => x"8c",
          1101 => x"08",
          1102 => x"34",
          1103 => x"81",
          1104 => x"0c",
          1105 => x"88",
          1106 => x"51",
          1107 => x"04",
          1108 => x"f0",
          1109 => x"d5",
          1110 => x"f0",
          1111 => x"38",
          1112 => x"30",
          1113 => x"80",
          1114 => x"0c",
          1115 => x"8a",
          1116 => x"f4",
          1117 => x"05",
          1118 => x"0c",
          1119 => x"80",
          1120 => x"8c",
          1121 => x"8c",
          1122 => x"08",
          1123 => x"fc",
          1124 => x"d5",
          1125 => x"f0",
          1126 => x"08",
          1127 => x"f0",
          1128 => x"f0",
          1129 => x"3f",
          1130 => x"f0",
          1131 => x"f0",
          1132 => x"38",
          1133 => x"30",
          1134 => x"82",
          1135 => x"82",
          1136 => x"82",
          1137 => x"08",
          1138 => x"0d",
          1139 => x"05",
          1140 => x"08",
          1141 => x"08",
          1142 => x"08",
          1143 => x"f0",
          1144 => x"08",
          1145 => x"82",
          1146 => x"82",
          1147 => x"53",
          1148 => x"52",
          1149 => x"51",
          1150 => x"70",
          1151 => x"54",
          1152 => x"80",
          1153 => x"f8",
          1154 => x"f8",
          1155 => x"05",
          1156 => x"87",
          1157 => x"82",
          1158 => x"0c",
          1159 => x"f0",
          1160 => x"f0",
          1161 => x"3f",
          1162 => x"e4",
          1163 => x"f0",
          1164 => x"82",
          1165 => x"53",
          1166 => x"52",
          1167 => x"51",
          1168 => x"82",
          1169 => x"82",
          1170 => x"08",
          1171 => x"0d",
          1172 => x"05",
          1173 => x"f8",
          1174 => x"05",
          1175 => x"08",
          1176 => x"fc",
          1177 => x"0b",
          1178 => x"24",
          1179 => x"05",
          1180 => x"05",
          1181 => x"08",
          1182 => x"0c",
          1183 => x"fc",
          1184 => x"82",
          1185 => x"d5",
          1186 => x"38",
          1187 => x"82",
          1188 => x"82",
          1189 => x"d5",
          1190 => x"f0",
          1191 => x"f0",
          1192 => x"08",
          1193 => x"f0",
          1194 => x"08",
          1195 => x"f0",
          1196 => x"82",
          1197 => x"2e",
          1198 => x"05",
          1199 => x"05",
          1200 => x"08",
          1201 => x"08",
          1202 => x"08",
          1203 => x"85",
          1204 => x"82",
          1205 => x"0c",
          1206 => x"f0",
          1207 => x"08",
          1208 => x"82",
          1209 => x"08",
          1210 => x"d5",
          1211 => x"ff",
          1212 => x"06",
          1213 => x"05",
          1214 => x"53",
          1215 => x"05",
          1216 => x"06",
          1217 => x"08",
          1218 => x"88",
          1219 => x"0c",
          1220 => x"d5",
          1221 => x"f0",
          1222 => x"2e",
          1223 => x"d5",
          1224 => x"81",
          1225 => x"72",
          1226 => x"34",
          1227 => x"82",
          1228 => x"d5",
          1229 => x"2e",
          1230 => x"05",
          1231 => x"cd",
          1232 => x"f4",
          1233 => x"05",
          1234 => x"70",
          1235 => x"f0",
          1236 => x"82",
          1237 => x"34",
          1238 => x"70",
          1239 => x"51",
          1240 => x"f8",
          1241 => x"f0",
          1242 => x"26",
          1243 => x"08",
          1244 => x"d5",
          1245 => x"73",
          1246 => x"f8",
          1247 => x"38",
          1248 => x"08",
          1249 => x"0b",
          1250 => x"b2",
          1251 => x"33",
          1252 => x"d5",
          1253 => x"b9",
          1254 => x"82",
          1255 => x"a5",
          1256 => x"f4",
          1257 => x"08",
          1258 => x"f8",
          1259 => x"cf",
          1260 => x"33",
          1261 => x"82",
          1262 => x"11",
          1263 => x"f8",
          1264 => x"05",
          1265 => x"d5",
          1266 => x"f0",
          1267 => x"27",
          1268 => x"05",
          1269 => x"d5",
          1270 => x"f0",
          1271 => x"26",
          1272 => x"08",
          1273 => x"d5",
          1274 => x"f0",
          1275 => x"74",
          1276 => x"f0",
          1277 => x"82",
          1278 => x"82",
          1279 => x"82",
          1280 => x"12",
          1281 => x"82",
          1282 => x"08",
          1283 => x"51",
          1284 => x"f0",
          1285 => x"82",
          1286 => x"72",
          1287 => x"08",
          1288 => x"08",
          1289 => x"8c",
          1290 => x"05",
          1291 => x"d5",
          1292 => x"f0",
          1293 => x"0c",
          1294 => x"04",
          1295 => x"f0",
          1296 => x"d5",
          1297 => x"f0",
          1298 => x"0c",
          1299 => x"70",
          1300 => x"82",
          1301 => x"81",
          1302 => x"81",
          1303 => x"88",
          1304 => x"0c",
          1305 => x"f8",
          1306 => x"81",
          1307 => x"f0",
          1308 => x"08",
          1309 => x"71",
          1310 => x"82",
          1311 => x"d5",
          1312 => x"b0",
          1313 => x"82",
          1314 => x"08",
          1315 => x"53",
          1316 => x"05",
          1317 => x"33",
          1318 => x"82",
          1319 => x"e2",
          1320 => x"e8",
          1321 => x"80",
          1322 => x"08",
          1323 => x"88",
          1324 => x"0c",
          1325 => x"d5",
          1326 => x"39",
          1327 => x"05",
          1328 => x"08",
          1329 => x"08",
          1330 => x"08",
          1331 => x"d5",
          1332 => x"a0",
          1333 => x"f0",
          1334 => x"82",
          1335 => x"af",
          1336 => x"08",
          1337 => x"83",
          1338 => x"f0",
          1339 => x"88",
          1340 => x"34",
          1341 => x"05",
          1342 => x"82",
          1343 => x"72",
          1344 => x"0b",
          1345 => x"82",
          1346 => x"08",
          1347 => x"f0",
          1348 => x"08",
          1349 => x"81",
          1350 => x"05",
          1351 => x"38",
          1352 => x"e0",
          1353 => x"08",
          1354 => x"f8",
          1355 => x"82",
          1356 => x"d5",
          1357 => x"73",
          1358 => x"f8",
          1359 => x"82",
          1360 => x"d5",
          1361 => x"89",
          1362 => x"f0",
          1363 => x"82",
          1364 => x"d5",
          1365 => x"72",
          1366 => x"d5",
          1367 => x"39",
          1368 => x"70",
          1369 => x"29",
          1370 => x"70",
          1371 => x"0c",
          1372 => x"70",
          1373 => x"51",
          1374 => x"d5",
          1375 => x"39",
          1376 => x"53",
          1377 => x"f0",
          1378 => x"f0",
          1379 => x"08",
          1380 => x"fc",
          1381 => x"82",
          1382 => x"d5",
          1383 => x"e4",
          1384 => x"0c",
          1385 => x"70",
          1386 => x"df",
          1387 => x"85",
          1388 => x"33",
          1389 => x"86",
          1390 => x"57",
          1391 => x"70",
          1392 => x"d5",
          1393 => x"75",
          1394 => x"3f",
          1395 => x"16",
          1396 => x"38",
          1397 => x"54",
          1398 => x"73",
          1399 => x"04",
          1400 => x"26",
          1401 => x"ad",
          1402 => x"b3",
          1403 => x"a8",
          1404 => x"51",
          1405 => x"80",
          1406 => x"e4",
          1407 => x"39",
          1408 => x"82",
          1409 => x"b4",
          1410 => x"bc",
          1411 => x"51",
          1412 => x"39",
          1413 => x"b5",
          1414 => x"51",
          1415 => x"39",
          1416 => x"b6",
          1417 => x"51",
          1418 => x"39",
          1419 => x"83",
          1420 => x"79",
          1421 => x"38",
          1422 => x"90",
          1423 => x"af",
          1424 => x"51",
          1425 => x"54",
          1426 => x"51",
          1427 => x"04",
          1428 => x"80",
          1429 => x"78",
          1430 => x"57",
          1431 => x"26",
          1432 => x"70",
          1433 => x"74",
          1434 => x"8c",
          1435 => x"3f",
          1436 => x"e4",
          1437 => x"87",
          1438 => x"08",
          1439 => x"80",
          1440 => x"b5",
          1441 => x"d5",
          1442 => x"80",
          1443 => x"59",
          1444 => x"51",
          1445 => x"78",
          1446 => x"2a",
          1447 => x"80",
          1448 => x"87",
          1449 => x"fe",
          1450 => x"e4",
          1451 => x"0d",
          1452 => x"58",
          1453 => x"7a",
          1454 => x"08",
          1455 => x"76",
          1456 => x"f1",
          1457 => x"d5",
          1458 => x"2d",
          1459 => x"78",
          1460 => x"3d",
          1461 => x"63",
          1462 => x"73",
          1463 => x"5e",
          1464 => x"51",
          1465 => x"51",
          1466 => x"79",
          1467 => x"89",
          1468 => x"c6",
          1469 => x"8e",
          1470 => x"51",
          1471 => x"b7",
          1472 => x"15",
          1473 => x"72",
          1474 => x"82",
          1475 => x"89",
          1476 => x"b1",
          1477 => x"18",
          1478 => x"33",
          1479 => x"99",
          1480 => x"ff",
          1481 => x"f1",
          1482 => x"3f",
          1483 => x"ff",
          1484 => x"27",
          1485 => x"55",
          1486 => x"38",
          1487 => x"83",
          1488 => x"81",
          1489 => x"90",
          1490 => x"82",
          1491 => x"39",
          1492 => x"d6",
          1493 => x"39",
          1494 => x"78",
          1495 => x"3f",
          1496 => x"98",
          1497 => x"81",
          1498 => x"d5",
          1499 => x"70",
          1500 => x"70",
          1501 => x"06",
          1502 => x"80",
          1503 => x"09",
          1504 => x"39",
          1505 => x"b2",
          1506 => x"0c",
          1507 => x"02",
          1508 => x"82",
          1509 => x"3f",
          1510 => x"3f",
          1511 => x"53",
          1512 => x"d4",
          1513 => x"2e",
          1514 => x"0d",
          1515 => x"80",
          1516 => x"98",
          1517 => x"e2",
          1518 => x"81",
          1519 => x"80",
          1520 => x"3f",
          1521 => x"80",
          1522 => x"70",
          1523 => x"92",
          1524 => x"b8",
          1525 => x"98",
          1526 => x"06",
          1527 => x"81",
          1528 => x"51",
          1529 => x"3f",
          1530 => x"52",
          1531 => x"97",
          1532 => x"ea",
          1533 => x"85",
          1534 => x"80",
          1535 => x"3f",
          1536 => x"80",
          1537 => x"70",
          1538 => x"92",
          1539 => x"b8",
          1540 => x"97",
          1541 => x"06",
          1542 => x"81",
          1543 => x"51",
          1544 => x"3f",
          1545 => x"52",
          1546 => x"96",
          1547 => x"f2",
          1548 => x"83",
          1549 => x"0d",
          1550 => x"70",
          1551 => x"e3",
          1552 => x"33",
          1553 => x"b9",
          1554 => x"8a",
          1555 => x"70",
          1556 => x"82",
          1557 => x"0b",
          1558 => x"d0",
          1559 => x"81",
          1560 => x"74",
          1561 => x"82",
          1562 => x"82",
          1563 => x"91",
          1564 => x"f0",
          1565 => x"d8",
          1566 => x"54",
          1567 => x"38",
          1568 => x"51",
          1569 => x"e4",
          1570 => x"0d",
          1571 => x"ec",
          1572 => x"80",
          1573 => x"81",
          1574 => x"81",
          1575 => x"53",
          1576 => x"9e",
          1577 => x"90",
          1578 => x"e4",
          1579 => x"e8",
          1580 => x"5e",
          1581 => x"3f",
          1582 => x"52",
          1583 => x"ff",
          1584 => x"d5",
          1585 => x"51",
          1586 => x"38",
          1587 => x"bd",
          1588 => x"90",
          1589 => x"78",
          1590 => x"39",
          1591 => x"78",
          1592 => x"bf",
          1593 => x"78",
          1594 => x"80",
          1595 => x"2e",
          1596 => x"89",
          1597 => x"83",
          1598 => x"24",
          1599 => x"ed",
          1600 => x"2e",
          1601 => x"3d",
          1602 => x"51",
          1603 => x"80",
          1604 => x"fc",
          1605 => x"c8",
          1606 => x"fe",
          1607 => x"53",
          1608 => x"82",
          1609 => x"e4",
          1610 => x"af",
          1611 => x"7b",
          1612 => x"7a",
          1613 => x"26",
          1614 => x"ff",
          1615 => x"eb",
          1616 => x"2e",
          1617 => x"11",
          1618 => x"3f",
          1619 => x"c8",
          1620 => x"ff",
          1621 => x"d5",
          1622 => x"82",
          1623 => x"64",
          1624 => x"62",
          1625 => x"79",
          1626 => x"b5",
          1627 => x"05",
          1628 => x"08",
          1629 => x"fe",
          1630 => x"ea",
          1631 => x"2e",
          1632 => x"11",
          1633 => x"3f",
          1634 => x"d0",
          1635 => x"b9",
          1636 => x"38",
          1637 => x"5b",
          1638 => x"7a",
          1639 => x"ba",
          1640 => x"1a",
          1641 => x"8a",
          1642 => x"b5",
          1643 => x"05",
          1644 => x"08",
          1645 => x"59",
          1646 => x"80",
          1647 => x"c9",
          1648 => x"82",
          1649 => x"d4",
          1650 => x"38",
          1651 => x"82",
          1652 => x"88",
          1653 => x"39",
          1654 => x"2e",
          1655 => x"89",
          1656 => x"05",
          1657 => x"ff",
          1658 => x"d5",
          1659 => x"c8",
          1660 => x"82",
          1661 => x"82",
          1662 => x"88",
          1663 => x"39",
          1664 => x"2e",
          1665 => x"aa",
          1666 => x"80",
          1667 => x"44",
          1668 => x"78",
          1669 => x"08",
          1670 => x"88",
          1671 => x"53",
          1672 => x"82",
          1673 => x"80",
          1674 => x"38",
          1675 => x"70",
          1676 => x"51",
          1677 => x"38",
          1678 => x"82",
          1679 => x"55",
          1680 => x"51",
          1681 => x"87",
          1682 => x"53",
          1683 => x"82",
          1684 => x"38",
          1685 => x"84",
          1686 => x"e4",
          1687 => x"02",
          1688 => x"81",
          1689 => x"53",
          1690 => x"82",
          1691 => x"39",
          1692 => x"84",
          1693 => x"c4",
          1694 => x"ff",
          1695 => x"59",
          1696 => x"79",
          1697 => x"11",
          1698 => x"3f",
          1699 => x"38",
          1700 => x"79",
          1701 => x"39",
          1702 => x"ff",
          1703 => x"53",
          1704 => x"82",
          1705 => x"38",
          1706 => x"84",
          1707 => x"e4",
          1708 => x"02",
          1709 => x"05",
          1710 => x"f0",
          1711 => x"a7",
          1712 => x"f7",
          1713 => x"82",
          1714 => x"82",
          1715 => x"79",
          1716 => x"79",
          1717 => x"38",
          1718 => x"05",
          1719 => x"11",
          1720 => x"3f",
          1721 => x"38",
          1722 => x"79",
          1723 => x"ff",
          1724 => x"fc",
          1725 => x"f4",
          1726 => x"af",
          1727 => x"f6",
          1728 => x"53",
          1729 => x"82",
          1730 => x"61",
          1731 => x"42",
          1732 => x"84",
          1733 => x"e4",
          1734 => x"70",
          1735 => x"ff",
          1736 => x"53",
          1737 => x"de",
          1738 => x"ae",
          1739 => x"9b",
          1740 => x"ff",
          1741 => x"d5",
          1742 => x"61",
          1743 => x"ff",
          1744 => x"dc",
          1745 => x"80",
          1746 => x"e0",
          1747 => x"f5",
          1748 => x"51",
          1749 => x"04",
          1750 => x"84",
          1751 => x"e4",
          1752 => x"52",
          1753 => x"3f",
          1754 => x"08",
          1755 => x"e4",
          1756 => x"a5",
          1757 => x"84",
          1758 => x"3f",
          1759 => x"c1",
          1760 => x"91",
          1761 => x"33",
          1762 => x"80",
          1763 => x"82",
          1764 => x"08",
          1765 => x"e4",
          1766 => x"51",
          1767 => x"60",
          1768 => x"81",
          1769 => x"cd",
          1770 => x"26",
          1771 => x"2e",
          1772 => x"7a",
          1773 => x"7a",
          1774 => x"82",
          1775 => x"b8",
          1776 => x"b5",
          1777 => x"b1",
          1778 => x"ff",
          1779 => x"39",
          1780 => x"53",
          1781 => x"b0",
          1782 => x"39",
          1783 => x"52",
          1784 => x"a6",
          1785 => x"d6",
          1786 => x"54",
          1787 => x"52",
          1788 => x"f5",
          1789 => x"e4",
          1790 => x"80",
          1791 => x"7a",
          1792 => x"7a",
          1793 => x"81",
          1794 => x"7a",
          1795 => x"81",
          1796 => x"ff",
          1797 => x"bc",
          1798 => x"51",
          1799 => x"bc",
          1800 => x"a0",
          1801 => x"d6",
          1802 => x"08",
          1803 => x"51",
          1804 => x"90",
          1805 => x"80",
          1806 => x"82",
          1807 => x"c0",
          1808 => x"84",
          1809 => x"82",
          1810 => x"55",
          1811 => x"d7",
          1812 => x"07",
          1813 => x"c0",
          1814 => x"87",
          1815 => x"5a",
          1816 => x"05",
          1817 => x"c4",
          1818 => x"70",
          1819 => x"89",
          1820 => x"9c",
          1821 => x"a8",
          1822 => x"d8",
          1823 => x"9c",
          1824 => x"3d",
          1825 => x"2b",
          1826 => x"08",
          1827 => x"54",
          1828 => x"82",
          1829 => x"fc",
          1830 => x"80",
          1831 => x"8a",
          1832 => x"09",
          1833 => x"f1",
          1834 => x"09",
          1835 => x"81",
          1836 => x"81",
          1837 => x"52",
          1838 => x"2e",
          1839 => x"9d",
          1840 => x"12",
          1841 => x"a0",
          1842 => x"2e",
          1843 => x"33",
          1844 => x"06",
          1845 => x"70",
          1846 => x"51",
          1847 => x"72",
          1848 => x"0c",
          1849 => x"86",
          1850 => x"53",
          1851 => x"3d",
          1852 => x"3f",
          1853 => x"53",
          1854 => x"e4",
          1855 => x"0d",
          1856 => x"53",
          1857 => x"38",
          1858 => x"52",
          1859 => x"13",
          1860 => x"80",
          1861 => x"52",
          1862 => x"13",
          1863 => x"80",
          1864 => x"52",
          1865 => x"8a",
          1866 => x"e7",
          1867 => x"c0",
          1868 => x"98",
          1869 => x"98",
          1870 => x"98",
          1871 => x"98",
          1872 => x"98",
          1873 => x"98",
          1874 => x"0c",
          1875 => x"0b",
          1876 => x"71",
          1877 => x"04",
          1878 => x"98",
          1879 => x"98",
          1880 => x"c0",
          1881 => x"34",
          1882 => x"83",
          1883 => x"5a",
          1884 => x"ac",
          1885 => x"c0",
          1886 => x"34",
          1887 => x"88",
          1888 => x"5a",
          1889 => x"79",
          1890 => x"ff",
          1891 => x"85",
          1892 => x"83",
          1893 => x"7d",
          1894 => x"c0",
          1895 => x"0d",
          1896 => x"33",
          1897 => x"06",
          1898 => x"51",
          1899 => x"94",
          1900 => x"70",
          1901 => x"2e",
          1902 => x"06",
          1903 => x"32",
          1904 => x"2e",
          1905 => x"06",
          1906 => x"81",
          1907 => x"52",
          1908 => x"94",
          1909 => x"d5",
          1910 => x"3d",
          1911 => x"70",
          1912 => x"d3",
          1913 => x"3d",
          1914 => x"8a",
          1915 => x"52",
          1916 => x"33",
          1917 => x"c0",
          1918 => x"38",
          1919 => x"70",
          1920 => x"54",
          1921 => x"2a",
          1922 => x"38",
          1923 => x"53",
          1924 => x"2a",
          1925 => x"be",
          1926 => x"c0",
          1927 => x"38",
          1928 => x"0c",
          1929 => x"3d",
          1930 => x"80",
          1931 => x"53",
          1932 => x"71",
          1933 => x"fc",
          1934 => x"55",
          1935 => x"80",
          1936 => x"51",
          1937 => x"06",
          1938 => x"38",
          1939 => x"51",
          1940 => x"81",
          1941 => x"38",
          1942 => x"51",
          1943 => x"06",
          1944 => x"80",
          1945 => x"52",
          1946 => x"70",
          1947 => x"ff",
          1948 => x"89",
          1949 => x"d3",
          1950 => x"52",
          1951 => x"2e",
          1952 => x"70",
          1953 => x"51",
          1954 => x"71",
          1955 => x"80",
          1956 => x"c0",
          1957 => x"ff",
          1958 => x"3d",
          1959 => x"e4",
          1960 => x"0c",
          1961 => x"33",
          1962 => x"c0",
          1963 => x"38",
          1964 => x"70",
          1965 => x"51",
          1966 => x"72",
          1967 => x"80",
          1968 => x"c0",
          1969 => x"2b",
          1970 => x"82",
          1971 => x"ff",
          1972 => x"70",
          1973 => x"80",
          1974 => x"a4",
          1975 => x"9e",
          1976 => x"c0",
          1977 => x"87",
          1978 => x"0c",
          1979 => x"90",
          1980 => x"d4",
          1981 => x"82",
          1982 => x"08",
          1983 => x"b4",
          1984 => x"9e",
          1985 => x"c0",
          1986 => x"87",
          1987 => x"0c",
          1988 => x"b0",
          1989 => x"70",
          1990 => x"84",
          1991 => x"9e",
          1992 => x"c0",
          1993 => x"81",
          1994 => x"87",
          1995 => x"0a",
          1996 => x"83",
          1997 => x"34",
          1998 => x"70",
          1999 => x"70",
          2000 => x"82",
          2001 => x"9e",
          2002 => x"51",
          2003 => x"81",
          2004 => x"0b",
          2005 => x"80",
          2006 => x"2e",
          2007 => x"c8",
          2008 => x"08",
          2009 => x"52",
          2010 => x"71",
          2011 => x"c0",
          2012 => x"06",
          2013 => x"38",
          2014 => x"80",
          2015 => x"84",
          2016 => x"80",
          2017 => x"d4",
          2018 => x"90",
          2019 => x"52",
          2020 => x"52",
          2021 => x"87",
          2022 => x"80",
          2023 => x"83",
          2024 => x"34",
          2025 => x"70",
          2026 => x"70",
          2027 => x"82",
          2028 => x"9e",
          2029 => x"52",
          2030 => x"52",
          2031 => x"9e",
          2032 => x"8a",
          2033 => x"d0",
          2034 => x"08",
          2035 => x"70",
          2036 => x"82",
          2037 => x"08",
          2038 => x"51",
          2039 => x"80",
          2040 => x"88",
          2041 => x"83",
          2042 => x"34",
          2043 => x"06",
          2044 => x"83",
          2045 => x"bd",
          2046 => x"d4",
          2047 => x"38",
          2048 => x"3f",
          2049 => x"3f",
          2050 => x"2e",
          2051 => x"d4",
          2052 => x"98",
          2053 => x"cb",
          2054 => x"82",
          2055 => x"11",
          2056 => x"93",
          2057 => x"73",
          2058 => x"08",
          2059 => x"82",
          2060 => x"82",
          2061 => x"94",
          2062 => x"8c",
          2063 => x"51",
          2064 => x"33",
          2065 => x"d4",
          2066 => x"54",
          2067 => x"b9",
          2068 => x"80",
          2069 => x"52",
          2070 => x"3f",
          2071 => x"2e",
          2072 => x"82",
          2073 => x"82",
          2074 => x"8e",
          2075 => x"bf",
          2076 => x"d4",
          2077 => x"38",
          2078 => x"3f",
          2079 => x"2e",
          2080 => x"ad",
          2081 => x"73",
          2082 => x"51",
          2083 => x"33",
          2084 => x"c0",
          2085 => x"d4",
          2086 => x"38",
          2087 => x"3f",
          2088 => x"3f",
          2089 => x"cc",
          2090 => x"ac",
          2091 => x"90",
          2092 => x"82",
          2093 => x"82",
          2094 => x"82",
          2095 => x"51",
          2096 => x"08",
          2097 => x"c5",
          2098 => x"84",
          2099 => x"82",
          2100 => x"51",
          2101 => x"33",
          2102 => x"d4",
          2103 => x"75",
          2104 => x"08",
          2105 => x"54",
          2106 => x"c2",
          2107 => x"d4",
          2108 => x"38",
          2109 => x"c0",
          2110 => x"d5",
          2111 => x"71",
          2112 => x"52",
          2113 => x"3f",
          2114 => x"3d",
          2115 => x"05",
          2116 => x"aa",
          2117 => x"05",
          2118 => x"51",
          2119 => x"39",
          2120 => x"c3",
          2121 => x"51",
          2122 => x"8f",
          2123 => x"88",
          2124 => x"96",
          2125 => x"87",
          2126 => x"0d",
          2127 => x"98",
          2128 => x"70",
          2129 => x"51",
          2130 => x"55",
          2131 => x"c3",
          2132 => x"97",
          2133 => x"70",
          2134 => x"81",
          2135 => x"3d",
          2136 => x"84",
          2137 => x"56",
          2138 => x"f1",
          2139 => x"d3",
          2140 => x"51",
          2141 => x"08",
          2142 => x"73",
          2143 => x"72",
          2144 => x"51",
          2145 => x"87",
          2146 => x"02",
          2147 => x"05",
          2148 => x"70",
          2149 => x"08",
          2150 => x"80",
          2151 => x"3f",
          2152 => x"82",
          2153 => x"58",
          2154 => x"e4",
          2155 => x"70",
          2156 => x"08",
          2157 => x"38",
          2158 => x"b6",
          2159 => x"05",
          2160 => x"81",
          2161 => x"38",
          2162 => x"80",
          2163 => x"56",
          2164 => x"ac",
          2165 => x"fc",
          2166 => x"51",
          2167 => x"08",
          2168 => x"82",
          2169 => x"3f",
          2170 => x"82",
          2171 => x"52",
          2172 => x"99",
          2173 => x"84",
          2174 => x"38",
          2175 => x"d5",
          2176 => x"38",
          2177 => x"d5",
          2178 => x"0b",
          2179 => x"04",
          2180 => x"82",
          2181 => x"3f",
          2182 => x"82",
          2183 => x"88",
          2184 => x"3f",
          2185 => x"38",
          2186 => x"d5",
          2187 => x"e4",
          2188 => x"08",
          2189 => x"74",
          2190 => x"82",
          2191 => x"3f",
          2192 => x"af",
          2193 => x"0d",
          2194 => x"5a",
          2195 => x"d5",
          2196 => x"82",
          2197 => x"0b",
          2198 => x"f8",
          2199 => x"9e",
          2200 => x"2e",
          2201 => x"3f",
          2202 => x"55",
          2203 => x"8e",
          2204 => x"70",
          2205 => x"09",
          2206 => x"51",
          2207 => x"73",
          2208 => x"8c",
          2209 => x"3f",
          2210 => x"38",
          2211 => x"3f",
          2212 => x"38",
          2213 => x"3f",
          2214 => x"3d",
          2215 => x"34",
          2216 => x"a9",
          2217 => x"7e",
          2218 => x"5a",
          2219 => x"a2",
          2220 => x"76",
          2221 => x"70",
          2222 => x"2e",
          2223 => x"26",
          2224 => x"82",
          2225 => x"ff",
          2226 => x"53",
          2227 => x"f3",
          2228 => x"38",
          2229 => x"88",
          2230 => x"39",
          2231 => x"5a",
          2232 => x"51",
          2233 => x"80",
          2234 => x"52",
          2235 => x"e4",
          2236 => x"38",
          2237 => x"81",
          2238 => x"ff",
          2239 => x"e4",
          2240 => x"0d",
          2241 => x"3d",
          2242 => x"3d",
          2243 => x"b0",
          2244 => x"73",
          2245 => x"83",
          2246 => x"bc",
          2247 => x"73",
          2248 => x"98",
          2249 => x"d5",
          2250 => x"2e",
          2251 => x"82",
          2252 => x"3f",
          2253 => x"38",
          2254 => x"3f",
          2255 => x"5b",
          2256 => x"52",
          2257 => x"f6",
          2258 => x"d5",
          2259 => x"80",
          2260 => x"ff",
          2261 => x"55",
          2262 => x"a9",
          2263 => x"70",
          2264 => x"53",
          2265 => x"f8",
          2266 => x"06",
          2267 => x"80",
          2268 => x"ff",
          2269 => x"ac",
          2270 => x"08",
          2271 => x"8f",
          2272 => x"e4",
          2273 => x"59",
          2274 => x"ff",
          2275 => x"2b",
          2276 => x"70",
          2277 => x"2c",
          2278 => x"05",
          2279 => x"51",
          2280 => x"81",
          2281 => x"77",
          2282 => x"0a",
          2283 => x"2c",
          2284 => x"38",
          2285 => x"85",
          2286 => x"06",
          2287 => x"82",
          2288 => x"74",
          2289 => x"05",
          2290 => x"56",
          2291 => x"76",
          2292 => x"3f",
          2293 => x"54",
          2294 => x"75",
          2295 => x"55",
          2296 => x"2b",
          2297 => x"70",
          2298 => x"11",
          2299 => x"33",
          2300 => x"55",
          2301 => x"92",
          2302 => x"0c",
          2303 => x"0b",
          2304 => x"82",
          2305 => x"34",
          2306 => x"7e",
          2307 => x"73",
          2308 => x"73",
          2309 => x"73",
          2310 => x"a4",
          2311 => x"74",
          2312 => x"73",
          2313 => x"73",
          2314 => x"0a",
          2315 => x"2c",
          2316 => x"df",
          2317 => x"56",
          2318 => x"1a",
          2319 => x"ed",
          2320 => x"38",
          2321 => x"34",
          2322 => x"0a",
          2323 => x"2c",
          2324 => x"56",
          2325 => x"c8",
          2326 => x"54",
          2327 => x"0a",
          2328 => x"2c",
          2329 => x"73",
          2330 => x"33",
          2331 => x"ed",
          2332 => x"77",
          2333 => x"08",
          2334 => x"74",
          2335 => x"05",
          2336 => x"56",
          2337 => x"fb",
          2338 => x"81",
          2339 => x"52",
          2340 => x"81",
          2341 => x"81",
          2342 => x"fb",
          2343 => x"05",
          2344 => x"15",
          2345 => x"f1",
          2346 => x"db",
          2347 => x"2b",
          2348 => x"57",
          2349 => x"38",
          2350 => x"34",
          2351 => x"51",
          2352 => x"0a",
          2353 => x"2c",
          2354 => x"75",
          2355 => x"08",
          2356 => x"82",
          2357 => x"98",
          2358 => x"56",
          2359 => x"82",
          2360 => x"9f",
          2361 => x"81",
          2362 => x"ed",
          2363 => x"25",
          2364 => x"a4",
          2365 => x"82",
          2366 => x"9f",
          2367 => x"51",
          2368 => x"81",
          2369 => x"ed",
          2370 => x"38",
          2371 => x"f3",
          2372 => x"0b",
          2373 => x"ed",
          2374 => x"af",
          2375 => x"54",
          2376 => x"f1",
          2377 => x"e3",
          2378 => x"54",
          2379 => x"ff",
          2380 => x"33",
          2381 => x"75",
          2382 => x"73",
          2383 => x"70",
          2384 => x"51",
          2385 => x"1a",
          2386 => x"f1",
          2387 => x"9e",
          2388 => x"81",
          2389 => x"ed",
          2390 => x"24",
          2391 => x"a0",
          2392 => x"a8",
          2393 => x"82",
          2394 => x"74",
          2395 => x"c8",
          2396 => x"3f",
          2397 => x"0a",
          2398 => x"33",
          2399 => x"38",
          2400 => x"70",
          2401 => x"59",
          2402 => x"38",
          2403 => x"54",
          2404 => x"70",
          2405 => x"82",
          2406 => x"82",
          2407 => x"75",
          2408 => x"ed",
          2409 => x"51",
          2410 => x"a8",
          2411 => x"f7",
          2412 => x"a8",
          2413 => x"74",
          2414 => x"e4",
          2415 => x"e4",
          2416 => x"74",
          2417 => x"93",
          2418 => x"82",
          2419 => x"54",
          2420 => x"ff",
          2421 => x"82",
          2422 => x"81",
          2423 => x"79",
          2424 => x"54",
          2425 => x"80",
          2426 => x"a4",
          2427 => x"09",
          2428 => x"08",
          2429 => x"51",
          2430 => x"08",
          2431 => x"08",
          2432 => x"52",
          2433 => x"c3",
          2434 => x"05",
          2435 => x"ab",
          2436 => x"82",
          2437 => x"82",
          2438 => x"05",
          2439 => x"a6",
          2440 => x"06",
          2441 => x"34",
          2442 => x"82",
          2443 => x"e2",
          2444 => x"33",
          2445 => x"33",
          2446 => x"87",
          2447 => x"14",
          2448 => x"1a",
          2449 => x"3f",
          2450 => x"54",
          2451 => x"f1",
          2452 => x"8b",
          2453 => x"54",
          2454 => x"39",
          2455 => x"82",
          2456 => x"d5",
          2457 => x"52",
          2458 => x"3f",
          2459 => x"77",
          2460 => x"34",
          2461 => x"15",
          2462 => x"d4",
          2463 => x"87",
          2464 => x"d5",
          2465 => x"07",
          2466 => x"2a",
          2467 => x"34",
          2468 => x"22",
          2469 => x"05",
          2470 => x"15",
          2471 => x"0d",
          2472 => x"51",
          2473 => x"83",
          2474 => x"06",
          2475 => x"0c",
          2476 => x"02",
          2477 => x"05",
          2478 => x"71",
          2479 => x"73",
          2480 => x"88",
          2481 => x"22",
          2482 => x"88",
          2483 => x"5b",
          2484 => x"70",
          2485 => x"14",
          2486 => x"15",
          2487 => x"d4",
          2488 => x"33",
          2489 => x"8f",
          2490 => x"71",
          2491 => x"88",
          2492 => x"34",
          2493 => x"12",
          2494 => x"71",
          2495 => x"3d",
          2496 => x"d4",
          2497 => x"70",
          2498 => x"87",
          2499 => x"2b",
          2500 => x"72",
          2501 => x"71",
          2502 => x"56",
          2503 => x"85",
          2504 => x"14",
          2505 => x"8b",
          2506 => x"57",
          2507 => x"13",
          2508 => x"2a",
          2509 => x"34",
          2510 => x"08",
          2511 => x"88",
          2512 => x"70",
          2513 => x"71",
          2514 => x"3d",
          2515 => x"05",
          2516 => x"2b",
          2517 => x"71",
          2518 => x"70",
          2519 => x"71",
          2520 => x"52",
          2521 => x"25",
          2522 => x"3f",
          2523 => x"33",
          2524 => x"83",
          2525 => x"12",
          2526 => x"2b",
          2527 => x"51",
          2528 => x"88",
          2529 => x"73",
          2530 => x"70",
          2531 => x"8b",
          2532 => x"57",
          2533 => x"33",
          2534 => x"ff",
          2535 => x"58",
          2536 => x"34",
          2537 => x"82",
          2538 => x"05",
          2539 => x"11",
          2540 => x"71",
          2541 => x"56",
          2542 => x"33",
          2543 => x"a2",
          2544 => x"53",
          2545 => x"70",
          2546 => x"70",
          2547 => x"8b",
          2548 => x"57",
          2549 => x"13",
          2550 => x"2a",
          2551 => x"34",
          2552 => x"08",
          2553 => x"71",
          2554 => x"52",
          2555 => x"0d",
          2556 => x"2a",
          2557 => x"57",
          2558 => x"08",
          2559 => x"33",
          2560 => x"83",
          2561 => x"12",
          2562 => x"07",
          2563 => x"55",
          2564 => x"82",
          2565 => x"3f",
          2566 => x"15",
          2567 => x"07",
          2568 => x"55",
          2569 => x"81",
          2570 => x"82",
          2571 => x"33",
          2572 => x"70",
          2573 => x"72",
          2574 => x"82",
          2575 => x"86",
          2576 => x"82",
          2577 => x"34",
          2578 => x"08",
          2579 => x"88",
          2580 => x"70",
          2581 => x"74",
          2582 => x"3d",
          2583 => x"82",
          2584 => x"3f",
          2585 => x"fe",
          2586 => x"3d",
          2587 => x"3f",
          2588 => x"06",
          2589 => x"85",
          2590 => x"5f",
          2591 => x"59",
          2592 => x"88",
          2593 => x"71",
          2594 => x"06",
          2595 => x"70",
          2596 => x"55",
          2597 => x"2e",
          2598 => x"15",
          2599 => x"07",
          2600 => x"ff",
          2601 => x"56",
          2602 => x"08",
          2603 => x"88",
          2604 => x"51",
          2605 => x"2e",
          2606 => x"78",
          2607 => x"80",
          2608 => x"09",
          2609 => x"f2",
          2610 => x"53",
          2611 => x"82",
          2612 => x"33",
          2613 => x"83",
          2614 => x"05",
          2615 => x"70",
          2616 => x"84",
          2617 => x"76",
          2618 => x"75",
          2619 => x"11",
          2620 => x"07",
          2621 => x"5a",
          2622 => x"87",
          2623 => x"1c",
          2624 => x"8b",
          2625 => x"5a",
          2626 => x"34",
          2627 => x"08",
          2628 => x"85",
          2629 => x"88",
          2630 => x"73",
          2631 => x"82",
          2632 => x"73",
          2633 => x"04",
          2634 => x"d4",
          2635 => x"53",
          2636 => x"fc",
          2637 => x"72",
          2638 => x"04",
          2639 => x"80",
          2640 => x"60",
          2641 => x"a8",
          2642 => x"b8",
          2643 => x"c7",
          2644 => x"92",
          2645 => x"51",
          2646 => x"83",
          2647 => x"7d",
          2648 => x"ff",
          2649 => x"33",
          2650 => x"70",
          2651 => x"70",
          2652 => x"1a",
          2653 => x"2b",
          2654 => x"53",
          2655 => x"5c",
          2656 => x"38",
          2657 => x"70",
          2658 => x"16",
          2659 => x"07",
          2660 => x"12",
          2661 => x"07",
          2662 => x"80",
          2663 => x"83",
          2664 => x"27",
          2665 => x"7b",
          2666 => x"51",
          2667 => x"06",
          2668 => x"7a",
          2669 => x"aa",
          2670 => x"7a",
          2671 => x"82",
          2672 => x"2b",
          2673 => x"80",
          2674 => x"d5",
          2675 => x"54",
          2676 => x"d4",
          2677 => x"ff",
          2678 => x"14",
          2679 => x"59",
          2680 => x"7a",
          2681 => x"f5",
          2682 => x"82",
          2683 => x"2b",
          2684 => x"80",
          2685 => x"d5",
          2686 => x"54",
          2687 => x"d4",
          2688 => x"ff",
          2689 => x"14",
          2690 => x"5c",
          2691 => x"39",
          2692 => x"82",
          2693 => x"08",
          2694 => x"52",
          2695 => x"a6",
          2696 => x"58",
          2697 => x"7a",
          2698 => x"19",
          2699 => x"84",
          2700 => x"73",
          2701 => x"04",
          2702 => x"52",
          2703 => x"08",
          2704 => x"8e",
          2705 => x"e4",
          2706 => x"82",
          2707 => x"ff",
          2708 => x"81",
          2709 => x"d5",
          2710 => x"e4",
          2711 => x"0d",
          2712 => x"9f",
          2713 => x"81",
          2714 => x"87",
          2715 => x"54",
          2716 => x"54",
          2717 => x"11",
          2718 => x"c0",
          2719 => x"70",
          2720 => x"8a",
          2721 => x"70",
          2722 => x"06",
          2723 => x"8c",
          2724 => x"71",
          2725 => x"e0",
          2726 => x"0c",
          2727 => x"60",
          2728 => x"33",
          2729 => x"5a",
          2730 => x"81",
          2731 => x"38",
          2732 => x"92",
          2733 => x"87",
          2734 => x"57",
          2735 => x"8c",
          2736 => x"75",
          2737 => x"51",
          2738 => x"7b",
          2739 => x"5d",
          2740 => x"06",
          2741 => x"81",
          2742 => x"72",
          2743 => x"8c",
          2744 => x"98",
          2745 => x"38",
          2746 => x"76",
          2747 => x"72",
          2748 => x"f7",
          2749 => x"80",
          2750 => x"5a",
          2751 => x"73",
          2752 => x"38",
          2753 => x"fc",
          2754 => x"83",
          2755 => x"d5",
          2756 => x"3d",
          2757 => x"bf",
          2758 => x"59",
          2759 => x"82",
          2760 => x"52",
          2761 => x"b1",
          2762 => x"92",
          2763 => x"87",
          2764 => x"56",
          2765 => x"0c",
          2766 => x"58",
          2767 => x"06",
          2768 => x"38",
          2769 => x"0c",
          2770 => x"81",
          2771 => x"38",
          2772 => x"d0",
          2773 => x"71",
          2774 => x"2e",
          2775 => x"92",
          2776 => x"06",
          2777 => x"59",
          2778 => x"06",
          2779 => x"80",
          2780 => x"06",
          2781 => x"fe",
          2782 => x"52",
          2783 => x"71",
          2784 => x"3d",
          2785 => x"84",
          2786 => x"a7",
          2787 => x"fa",
          2788 => x"06",
          2789 => x"85",
          2790 => x"56",
          2791 => x"76",
          2792 => x"c0",
          2793 => x"2e",
          2794 => x"2e",
          2795 => x"08",
          2796 => x"51",
          2797 => x"c0",
          2798 => x"87",
          2799 => x"38",
          2800 => x"14",
          2801 => x"52",
          2802 => x"92",
          2803 => x"39",
          2804 => x"39",
          2805 => x"e4",
          2806 => x"0d",
          2807 => x"88",
          2808 => x"51",
          2809 => x"75",
          2810 => x"90",
          2811 => x"33",
          2812 => x"71",
          2813 => x"54",
          2814 => x"ff",
          2815 => x"05",
          2816 => x"05",
          2817 => x"72",
          2818 => x"0d",
          2819 => x"81",
          2820 => x"70",
          2821 => x"88",
          2822 => x"54",
          2823 => x"34",
          2824 => x"76",
          2825 => x"2e",
          2826 => x"33",
          2827 => x"11",
          2828 => x"fe",
          2829 => x"53",
          2830 => x"ff",
          2831 => x"0d",
          2832 => x"56",
          2833 => x"33",
          2834 => x"71",
          2835 => x"72",
          2836 => x"e2",
          2837 => x"3d",
          2838 => x"54",
          2839 => x"38",
          2840 => x"f3",
          2841 => x"84",
          2842 => x"e4",
          2843 => x"08",
          2844 => x"54",
          2845 => x"82",
          2846 => x"2e",
          2847 => x"80",
          2848 => x"83",
          2849 => x"86",
          2850 => x"82",
          2851 => x"f7",
          2852 => x"17",
          2853 => x"d6",
          2854 => x"b8",
          2855 => x"59",
          2856 => x"7a",
          2857 => x"d5",
          2858 => x"08",
          2859 => x"08",
          2860 => x"38",
          2861 => x"09",
          2862 => x"18",
          2863 => x"f9",
          2864 => x"82",
          2865 => x"fa",
          2866 => x"57",
          2867 => x"75",
          2868 => x"08",
          2869 => x"81",
          2870 => x"16",
          2871 => x"e4",
          2872 => x"81",
          2873 => x"d5",
          2874 => x"3d",
          2875 => x"3f",
          2876 => x"e4",
          2877 => x"74",
          2878 => x"38",
          2879 => x"09",
          2880 => x"53",
          2881 => x"70",
          2882 => x"d5",
          2883 => x"3f",
          2884 => x"51",
          2885 => x"f2",
          2886 => x"3f",
          2887 => x"51",
          2888 => x"84",
          2889 => x"17",
          2890 => x"79",
          2891 => x"51",
          2892 => x"80",
          2893 => x"f9",
          2894 => x"2e",
          2895 => x"e4",
          2896 => x"0d",
          2897 => x"05",
          2898 => x"27",
          2899 => x"29",
          2900 => x"82",
          2901 => x"f9",
          2902 => x"54",
          2903 => x"76",
          2904 => x"ff",
          2905 => x"80",
          2906 => x"72",
          2907 => x"72",
          2908 => x"39",
          2909 => x"a8",
          2910 => x"fd",
          2911 => x"9f",
          2912 => x"11",
          2913 => x"18",
          2914 => x"53",
          2915 => x"80",
          2916 => x"b8",
          2917 => x"79",
          2918 => x"58",
          2919 => x"9f",
          2920 => x"88",
          2921 => x"51",
          2922 => x"80",
          2923 => x"74",
          2924 => x"82",
          2925 => x"58",
          2926 => x"08",
          2927 => x"82",
          2928 => x"2b",
          2929 => x"51",
          2930 => x"f0",
          2931 => x"77",
          2932 => x"04",
          2933 => x"58",
          2934 => x"9e",
          2935 => x"96",
          2936 => x"81",
          2937 => x"72",
          2938 => x"72",
          2939 => x"39",
          2940 => x"a8",
          2941 => x"fb",
          2942 => x"82",
          2943 => x"83",
          2944 => x"78",
          2945 => x"76",
          2946 => x"9f",
          2947 => x"07",
          2948 => x"83",
          2949 => x"08",
          2950 => x"82",
          2951 => x"08",
          2952 => x"16",
          2953 => x"76",
          2954 => x"81",
          2955 => x"53",
          2956 => x"88",
          2957 => x"51",
          2958 => x"59",
          2959 => x"77",
          2960 => x"83",
          2961 => x"f6",
          2962 => x"a8",
          2963 => x"ef",
          2964 => x"d5",
          2965 => x"06",
          2966 => x"18",
          2967 => x"f6",
          2968 => x"0a",
          2969 => x"c5",
          2970 => x"82",
          2971 => x"f8",
          2972 => x"59",
          2973 => x"38",
          2974 => x"73",
          2975 => x"52",
          2976 => x"e4",
          2977 => x"f2",
          2978 => x"39",
          2979 => x"e4",
          2980 => x"78",
          2981 => x"08",
          2982 => x"80",
          2983 => x"2e",
          2984 => x"2e",
          2985 => x"51",
          2986 => x"c5",
          2987 => x"18",
          2988 => x"90",
          2989 => x"16",
          2990 => x"34",
          2991 => x"38",
          2992 => x"8a",
          2993 => x"7e",
          2994 => x"38",
          2995 => x"88",
          2996 => x"38",
          2997 => x"51",
          2998 => x"d5",
          2999 => x"d5",
          3000 => x"ff",
          3001 => x"82",
          3002 => x"79",
          3003 => x"73",
          3004 => x"2e",
          3005 => x"1a",
          3006 => x"38",
          3007 => x"af",
          3008 => x"81",
          3009 => x"d5",
          3010 => x"09",
          3011 => x"70",
          3012 => x"51",
          3013 => x"82",
          3014 => x"90",
          3015 => x"38",
          3016 => x"73",
          3017 => x"77",
          3018 => x"76",
          3019 => x"26",
          3020 => x"f8",
          3021 => x"2e",
          3022 => x"08",
          3023 => x"82",
          3024 => x"08",
          3025 => x"25",
          3026 => x"73",
          3027 => x"81",
          3028 => x"f5",
          3029 => x"f9",
          3030 => x"d5",
          3031 => x"08",
          3032 => x"80",
          3033 => x"38",
          3034 => x"d0",
          3035 => x"a5",
          3036 => x"08",
          3037 => x"74",
          3038 => x"18",
          3039 => x"73",
          3040 => x"74",
          3041 => x"55",
          3042 => x"85",
          3043 => x"d5",
          3044 => x"3d",
          3045 => x"3f",
          3046 => x"82",
          3047 => x"52",
          3048 => x"e4",
          3049 => x"0c",
          3050 => x"15",
          3051 => x"56",
          3052 => x"22",
          3053 => x"54",
          3054 => x"33",
          3055 => x"08",
          3056 => x"76",
          3057 => x"9f",
          3058 => x"d5",
          3059 => x"3d",
          3060 => x"57",
          3061 => x"38",
          3062 => x"38",
          3063 => x"54",
          3064 => x"73",
          3065 => x"73",
          3066 => x"0b",
          3067 => x"27",
          3068 => x"18",
          3069 => x"70",
          3070 => x"b2",
          3071 => x"3f",
          3072 => x"e4",
          3073 => x"82",
          3074 => x"16",
          3075 => x"38",
          3076 => x"55",
          3077 => x"d5",
          3078 => x"0c",
          3079 => x"53",
          3080 => x"85",
          3081 => x"2a",
          3082 => x"06",
          3083 => x"58",
          3084 => x"0d",
          3085 => x"90",
          3086 => x"f0",
          3087 => x"0b",
          3088 => x"84",
          3089 => x"76",
          3090 => x"38",
          3091 => x"08",
          3092 => x"88",
          3093 => x"81",
          3094 => x"22",
          3095 => x"72",
          3096 => x"f3",
          3097 => x"82",
          3098 => x"27",
          3099 => x"e4",
          3100 => x"16",
          3101 => x"ca",
          3102 => x"0c",
          3103 => x"08",
          3104 => x"d5",
          3105 => x"e4",
          3106 => x"55",
          3107 => x"38",
          3108 => x"2e",
          3109 => x"75",
          3110 => x"08",
          3111 => x"52",
          3112 => x"e4",
          3113 => x"0c",
          3114 => x"80",
          3115 => x"3d",
          3116 => x"71",
          3117 => x"51",
          3118 => x"54",
          3119 => x"82",
          3120 => x"52",
          3121 => x"e4",
          3122 => x"d2",
          3123 => x"08",
          3124 => x"e5",
          3125 => x"58",
          3126 => x"38",
          3127 => x"80",
          3128 => x"7a",
          3129 => x"39",
          3130 => x"76",
          3131 => x"08",
          3132 => x"ff",
          3133 => x"06",
          3134 => x"e4",
          3135 => x"0d",
          3136 => x"3f",
          3137 => x"06",
          3138 => x"83",
          3139 => x"14",
          3140 => x"08",
          3141 => x"d5",
          3142 => x"3d",
          3143 => x"06",
          3144 => x"af",
          3145 => x"83",
          3146 => x"90",
          3147 => x"3f",
          3148 => x"75",
          3149 => x"2a",
          3150 => x"81",
          3151 => x"ff",
          3152 => x"72",
          3153 => x"85",
          3154 => x"62",
          3155 => x"81",
          3156 => x"80",
          3157 => x"52",
          3158 => x"e4",
          3159 => x"eb",
          3160 => x"55",
          3161 => x"39",
          3162 => x"ff",
          3163 => x"82",
          3164 => x"2e",
          3165 => x"82",
          3166 => x"09",
          3167 => x"73",
          3168 => x"e4",
          3169 => x"88",
          3170 => x"56",
          3171 => x"5c",
          3172 => x"81",
          3173 => x"70",
          3174 => x"92",
          3175 => x"06",
          3176 => x"56",
          3177 => x"06",
          3178 => x"7c",
          3179 => x"38",
          3180 => x"e8",
          3181 => x"ff",
          3182 => x"74",
          3183 => x"f3",
          3184 => x"82",
          3185 => x"e8",
          3186 => x"ff",
          3187 => x"38",
          3188 => x"73",
          3189 => x"23",
          3190 => x"ff",
          3191 => x"81",
          3192 => x"74",
          3193 => x"51",
          3194 => x"73",
          3195 => x"1a",
          3196 => x"81",
          3197 => x"ff",
          3198 => x"38",
          3199 => x"e4",
          3200 => x"2e",
          3201 => x"a0",
          3202 => x"3f",
          3203 => x"e4",
          3204 => x"84",
          3205 => x"0c",
          3206 => x"0d",
          3207 => x"40",
          3208 => x"3f",
          3209 => x"e4",
          3210 => x"5f",
          3211 => x"19",
          3212 => x"82",
          3213 => x"08",
          3214 => x"33",
          3215 => x"82",
          3216 => x"70",
          3217 => x"1a",
          3218 => x"38",
          3219 => x"54",
          3220 => x"b2",
          3221 => x"81",
          3222 => x"2a",
          3223 => x"82",
          3224 => x"06",
          3225 => x"8d",
          3226 => x"90",
          3227 => x"5e",
          3228 => x"b9",
          3229 => x"2e",
          3230 => x"1f",
          3231 => x"3f",
          3232 => x"06",
          3233 => x"70",
          3234 => x"56",
          3235 => x"1b",
          3236 => x"82",
          3237 => x"56",
          3238 => x"fe",
          3239 => x"e1",
          3240 => x"10",
          3241 => x"59",
          3242 => x"d5",
          3243 => x"c1",
          3244 => x"ff",
          3245 => x"81",
          3246 => x"38",
          3247 => x"06",
          3248 => x"38",
          3249 => x"1d",
          3250 => x"ff",
          3251 => x"84",
          3252 => x"39",
          3253 => x"3f",
          3254 => x"54",
          3255 => x"33",
          3256 => x"53",
          3257 => x"e5",
          3258 => x"2e",
          3259 => x"ac",
          3260 => x"81",
          3261 => x"d5",
          3262 => x"77",
          3263 => x"04",
          3264 => x"12",
          3265 => x"86",
          3266 => x"1d",
          3267 => x"80",
          3268 => x"16",
          3269 => x"8c",
          3270 => x"70",
          3271 => x"80",
          3272 => x"80",
          3273 => x"ab",
          3274 => x"7b",
          3275 => x"51",
          3276 => x"c6",
          3277 => x"ff",
          3278 => x"b4",
          3279 => x"19",
          3280 => x"76",
          3281 => x"2a",
          3282 => x"73",
          3283 => x"a1",
          3284 => x"25",
          3285 => x"02",
          3286 => x"b0",
          3287 => x"84",
          3288 => x"ff",
          3289 => x"58",
          3290 => x"05",
          3291 => x"77",
          3292 => x"a0",
          3293 => x"52",
          3294 => x"08",
          3295 => x"74",
          3296 => x"81",
          3297 => x"74",
          3298 => x"94",
          3299 => x"15",
          3300 => x"87",
          3301 => x"70",
          3302 => x"87",
          3303 => x"f9",
          3304 => x"81",
          3305 => x"84",
          3306 => x"82",
          3307 => x"82",
          3308 => x"06",
          3309 => x"33",
          3310 => x"33",
          3311 => x"55",
          3312 => x"38",
          3313 => x"9f",
          3314 => x"78",
          3315 => x"d5",
          3316 => x"82",
          3317 => x"2e",
          3318 => x"1b",
          3319 => x"ef",
          3320 => x"82",
          3321 => x"1a",
          3322 => x"08",
          3323 => x"52",
          3324 => x"e4",
          3325 => x"d7",
          3326 => x"7a",
          3327 => x"8d",
          3328 => x"82",
          3329 => x"d5",
          3330 => x"df",
          3331 => x"55",
          3332 => x"38",
          3333 => x"57",
          3334 => x"17",
          3335 => x"73",
          3336 => x"17",
          3337 => x"83",
          3338 => x"1b",
          3339 => x"77",
          3340 => x"81",
          3341 => x"51",
          3342 => x"57",
          3343 => x"ff",
          3344 => x"1a",
          3345 => x"82",
          3346 => x"08",
          3347 => x"08",
          3348 => x"3f",
          3349 => x"08",
          3350 => x"ab",
          3351 => x"8c",
          3352 => x"76",
          3353 => x"3d",
          3354 => x"08",
          3355 => x"59",
          3356 => x"72",
          3357 => x"d5",
          3358 => x"80",
          3359 => x"51",
          3360 => x"54",
          3361 => x"15",
          3362 => x"83",
          3363 => x"a2",
          3364 => x"51",
          3365 => x"54",
          3366 => x"38",
          3367 => x"38",
          3368 => x"88",
          3369 => x"60",
          3370 => x"96",
          3371 => x"83",
          3372 => x"81",
          3373 => x"05",
          3374 => x"57",
          3375 => x"10",
          3376 => x"53",
          3377 => x"70",
          3378 => x"8f",
          3379 => x"df",
          3380 => x"79",
          3381 => x"7a",
          3382 => x"84",
          3383 => x"ff",
          3384 => x"38",
          3385 => x"2a",
          3386 => x"34",
          3387 => x"30",
          3388 => x"25",
          3389 => x"85",
          3390 => x"34",
          3391 => x"8c",
          3392 => x"51",
          3393 => x"30",
          3394 => x"59",
          3395 => x"80",
          3396 => x"1a",
          3397 => x"70",
          3398 => x"a0",
          3399 => x"81",
          3400 => x"89",
          3401 => x"25",
          3402 => x"38",
          3403 => x"70",
          3404 => x"74",
          3405 => x"17",
          3406 => x"77",
          3407 => x"14",
          3408 => x"87",
          3409 => x"19",
          3410 => x"73",
          3411 => x"80",
          3412 => x"19",
          3413 => x"54",
          3414 => x"1c",
          3415 => x"79",
          3416 => x"85",
          3417 => x"06",
          3418 => x"15",
          3419 => x"74",
          3420 => x"19",
          3421 => x"59",
          3422 => x"17",
          3423 => x"34",
          3424 => x"53",
          3425 => x"9c",
          3426 => x"19",
          3427 => x"53",
          3428 => x"78",
          3429 => x"82",
          3430 => x"13",
          3431 => x"08",
          3432 => x"f0",
          3433 => x"80",
          3434 => x"af",
          3435 => x"dc",
          3436 => x"38",
          3437 => x"aa",
          3438 => x"33",
          3439 => x"81",
          3440 => x"dc",
          3441 => x"07",
          3442 => x"88",
          3443 => x"73",
          3444 => x"ab",
          3445 => x"ee",
          3446 => x"e1",
          3447 => x"08",
          3448 => x"05",
          3449 => x"08",
          3450 => x"ff",
          3451 => x"38",
          3452 => x"90",
          3453 => x"19",
          3454 => x"ff",
          3455 => x"73",
          3456 => x"55",
          3457 => x"2e",
          3458 => x"38",
          3459 => x"92",
          3460 => x"38",
          3461 => x"78",
          3462 => x"19",
          3463 => x"80",
          3464 => x"af",
          3465 => x"57",
          3466 => x"80",
          3467 => x"dc",
          3468 => x"2b",
          3469 => x"8c",
          3470 => x"a5",
          3471 => x"09",
          3472 => x"22",
          3473 => x"80",
          3474 => x"2e",
          3475 => x"1a",
          3476 => x"1f",
          3477 => x"83",
          3478 => x"05",
          3479 => x"27",
          3480 => x"ab",
          3481 => x"2e",
          3482 => x"55",
          3483 => x"32",
          3484 => x"53",
          3485 => x"38",
          3486 => x"e0",
          3487 => x"80",
          3488 => x"85",
          3489 => x"99",
          3490 => x"ff",
          3491 => x"09",
          3492 => x"10",
          3493 => x"a0",
          3494 => x"83",
          3495 => x"09",
          3496 => x"57",
          3497 => x"fe",
          3498 => x"2e",
          3499 => x"55",
          3500 => x"38",
          3501 => x"ae",
          3502 => x"53",
          3503 => x"3f",
          3504 => x"10",
          3505 => x"54",
          3506 => x"a0",
          3507 => x"30",
          3508 => x"79",
          3509 => x"38",
          3510 => x"54",
          3511 => x"81",
          3512 => x"72",
          3513 => x"51",
          3514 => x"7e",
          3515 => x"2e",
          3516 => x"79",
          3517 => x"58",
          3518 => x"5d",
          3519 => x"27",
          3520 => x"b5",
          3521 => x"82",
          3522 => x"70",
          3523 => x"56",
          3524 => x"ff",
          3525 => x"54",
          3526 => x"1f",
          3527 => x"83",
          3528 => x"7d",
          3529 => x"55",
          3530 => x"c3",
          3531 => x"52",
          3532 => x"82",
          3533 => x"80",
          3534 => x"39",
          3535 => x"85",
          3536 => x"16",
          3537 => x"81",
          3538 => x"06",
          3539 => x"54",
          3540 => x"de",
          3541 => x"e5",
          3542 => x"0b",
          3543 => x"81",
          3544 => x"fc",
          3545 => x"8c",
          3546 => x"73",
          3547 => x"76",
          3548 => x"81",
          3549 => x"81",
          3550 => x"76",
          3551 => x"81",
          3552 => x"38",
          3553 => x"34",
          3554 => x"e4",
          3555 => x"d5",
          3556 => x"d5",
          3557 => x"80",
          3558 => x"06",
          3559 => x"80",
          3560 => x"73",
          3561 => x"0b",
          3562 => x"39",
          3563 => x"85",
          3564 => x"81",
          3565 => x"1e",
          3566 => x"51",
          3567 => x"90",
          3568 => x"b8",
          3569 => x"82",
          3570 => x"a1",
          3571 => x"3d",
          3572 => x"ff",
          3573 => x"5c",
          3574 => x"38",
          3575 => x"9f",
          3576 => x"38",
          3577 => x"81",
          3578 => x"11",
          3579 => x"70",
          3580 => x"81",
          3581 => x"76",
          3582 => x"c7",
          3583 => x"57",
          3584 => x"70",
          3585 => x"53",
          3586 => x"e0",
          3587 => x"ff",
          3588 => x"38",
          3589 => x"51",
          3590 => x"72",
          3591 => x"70",
          3592 => x"32",
          3593 => x"73",
          3594 => x"70",
          3595 => x"19",
          3596 => x"38",
          3597 => x"74",
          3598 => x"39",
          3599 => x"d5",
          3600 => x"3d",
          3601 => x"34",
          3602 => x"75",
          3603 => x"d5",
          3604 => x"16",
          3605 => x"08",
          3606 => x"73",
          3607 => x"80",
          3608 => x"56",
          3609 => x"06",
          3610 => x"32",
          3611 => x"51",
          3612 => x"e8",
          3613 => x"53",
          3614 => x"51",
          3615 => x"55",
          3616 => x"38",
          3617 => x"8a",
          3618 => x"e4",
          3619 => x"2e",
          3620 => x"e4",
          3621 => x"0d",
          3622 => x"33",
          3623 => x"fc",
          3624 => x"8b",
          3625 => x"24",
          3626 => x"84",
          3627 => x"55",
          3628 => x"b1",
          3629 => x"06",
          3630 => x"ae",
          3631 => x"3f",
          3632 => x"70",
          3633 => x"76",
          3634 => x"2a",
          3635 => x"72",
          3636 => x"74",
          3637 => x"19",
          3638 => x"14",
          3639 => x"e4",
          3640 => x"54",
          3641 => x"76",
          3642 => x"70",
          3643 => x"86",
          3644 => x"5b",
          3645 => x"81",
          3646 => x"38",
          3647 => x"d5",
          3648 => x"81",
          3649 => x"83",
          3650 => x"53",
          3651 => x"15",
          3652 => x"08",
          3653 => x"0c",
          3654 => x"80",
          3655 => x"d9",
          3656 => x"72",
          3657 => x"05",
          3658 => x"59",
          3659 => x"2e",
          3660 => x"9e",
          3661 => x"06",
          3662 => x"33",
          3663 => x"06",
          3664 => x"91",
          3665 => x"16",
          3666 => x"c0",
          3667 => x"f9",
          3668 => x"f1",
          3669 => x"3f",
          3670 => x"06",
          3671 => x"06",
          3672 => x"c9",
          3673 => x"ff",
          3674 => x"dc",
          3675 => x"e4",
          3676 => x"c8",
          3677 => x"14",
          3678 => x"51",
          3679 => x"84",
          3680 => x"71",
          3681 => x"53",
          3682 => x"8b",
          3683 => x"80",
          3684 => x"39",
          3685 => x"82",
          3686 => x"08",
          3687 => x"8d",
          3688 => x"14",
          3689 => x"08",
          3690 => x"38",
          3691 => x"82",
          3692 => x"51",
          3693 => x"83",
          3694 => x"80",
          3695 => x"78",
          3696 => x"78",
          3697 => x"22",
          3698 => x"97",
          3699 => x"d5",
          3700 => x"82",
          3701 => x"f5",
          3702 => x"ff",
          3703 => x"9f",
          3704 => x"39",
          3705 => x"38",
          3706 => x"a4",
          3707 => x"0c",
          3708 => x"76",
          3709 => x"80",
          3710 => x"d5",
          3711 => x"8d",
          3712 => x"91",
          3713 => x"3f",
          3714 => x"74",
          3715 => x"79",
          3716 => x"ac",
          3717 => x"2e",
          3718 => x"2a",
          3719 => x"ff",
          3720 => x"a0",
          3721 => x"0b",
          3722 => x"0c",
          3723 => x"83",
          3724 => x"80",
          3725 => x"d5",
          3726 => x"72",
          3727 => x"38",
          3728 => x"3f",
          3729 => x"82",
          3730 => x"b6",
          3731 => x"e4",
          3732 => x"82",
          3733 => x"c8",
          3734 => x"82",
          3735 => x"d2",
          3736 => x"9c",
          3737 => x"e4",
          3738 => x"09",
          3739 => x"51",
          3740 => x"94",
          3741 => x"dc",
          3742 => x"0c",
          3743 => x"81",
          3744 => x"72",
          3745 => x"8c",
          3746 => x"80",
          3747 => x"3d",
          3748 => x"89",
          3749 => x"08",
          3750 => x"33",
          3751 => x"13",
          3752 => x"76",
          3753 => x"13",
          3754 => x"d5",
          3755 => x"38",
          3756 => x"80",
          3757 => x"82",
          3758 => x"fa",
          3759 => x"58",
          3760 => x"9a",
          3761 => x"e4",
          3762 => x"08",
          3763 => x"08",
          3764 => x"80",
          3765 => x"84",
          3766 => x"75",
          3767 => x"53",
          3768 => x"f6",
          3769 => x"73",
          3770 => x"04",
          3771 => x"80",
          3772 => x"78",
          3773 => x"06",
          3774 => x"9a",
          3775 => x"3f",
          3776 => x"e4",
          3777 => x"52",
          3778 => x"3f",
          3779 => x"e4",
          3780 => x"33",
          3781 => x"25",
          3782 => x"54",
          3783 => x"80",
          3784 => x"81",
          3785 => x"3f",
          3786 => x"02",
          3787 => x"81",
          3788 => x"06",
          3789 => x"88",
          3790 => x"58",
          3791 => x"70",
          3792 => x"81",
          3793 => x"ed",
          3794 => x"88",
          3795 => x"c2",
          3796 => x"15",
          3797 => x"d7",
          3798 => x"51",
          3799 => x"83",
          3800 => x"38",
          3801 => x"53",
          3802 => x"cc",
          3803 => x"82",
          3804 => x"39",
          3805 => x"33",
          3806 => x"55",
          3807 => x"55",
          3808 => x"81",
          3809 => x"38",
          3810 => x"a0",
          3811 => x"52",
          3812 => x"e4",
          3813 => x"55",
          3814 => x"38",
          3815 => x"54",
          3816 => x"c0",
          3817 => x"1b",
          3818 => x"70",
          3819 => x"e4",
          3820 => x"0c",
          3821 => x"3f",
          3822 => x"08",
          3823 => x"86",
          3824 => x"1a",
          3825 => x"0b",
          3826 => x"0c",
          3827 => x"54",
          3828 => x"d5",
          3829 => x"82",
          3830 => x"17",
          3831 => x"57",
          3832 => x"e7",
          3833 => x"d5",
          3834 => x"55",
          3835 => x"81",
          3836 => x"31",
          3837 => x"25",
          3838 => x"81",
          3839 => x"38",
          3840 => x"75",
          3841 => x"a2",
          3842 => x"3f",
          3843 => x"55",
          3844 => x"e4",
          3845 => x"80",
          3846 => x"e4",
          3847 => x"0d",
          3848 => x"59",
          3849 => x"52",
          3850 => x"e4",
          3851 => x"38",
          3852 => x"86",
          3853 => x"19",
          3854 => x"80",
          3855 => x"0b",
          3856 => x"39",
          3857 => x"82",
          3858 => x"08",
          3859 => x"74",
          3860 => x"94",
          3861 => x"56",
          3862 => x"22",
          3863 => x"55",
          3864 => x"19",
          3865 => x"52",
          3866 => x"e4",
          3867 => x"38",
          3868 => x"98",
          3869 => x"51",
          3870 => x"80",
          3871 => x"08",
          3872 => x"80",
          3873 => x"8a",
          3874 => x"27",
          3875 => x"54",
          3876 => x"51",
          3877 => x"08",
          3878 => x"56",
          3879 => x"16",
          3880 => x"95",
          3881 => x"b4",
          3882 => x"05",
          3883 => x"2b",
          3884 => x"94",
          3885 => x"71",
          3886 => x"38",
          3887 => x"51",
          3888 => x"fd",
          3889 => x"83",
          3890 => x"51",
          3891 => x"7e",
          3892 => x"1b",
          3893 => x"fd",
          3894 => x"e4",
          3895 => x"0d",
          3896 => x"58",
          3897 => x"52",
          3898 => x"e4",
          3899 => x"38",
          3900 => x"86",
          3901 => x"18",
          3902 => x"51",
          3903 => x"83",
          3904 => x"19",
          3905 => x"0b",
          3906 => x"39",
          3907 => x"74",
          3908 => x"7b",
          3909 => x"08",
          3910 => x"82",
          3911 => x"05",
          3912 => x"bf",
          3913 => x"55",
          3914 => x"98",
          3915 => x"3f",
          3916 => x"e4",
          3917 => x"81",
          3918 => x"ff",
          3919 => x"18",
          3920 => x"7e",
          3921 => x"2e",
          3922 => x"ff",
          3923 => x"fe",
          3924 => x"51",
          3925 => x"08",
          3926 => x"e4",
          3927 => x"78",
          3928 => x"7f",
          3929 => x"75",
          3930 => x"78",
          3931 => x"33",
          3932 => x"e4",
          3933 => x"08",
          3934 => x"9c",
          3935 => x"77",
          3936 => x"16",
          3937 => x"80",
          3938 => x"56",
          3939 => x"19",
          3940 => x"bb",
          3941 => x"de",
          3942 => x"76",
          3943 => x"ff",
          3944 => x"7b",
          3945 => x"18",
          3946 => x"3f",
          3947 => x"75",
          3948 => x"ff",
          3949 => x"d4",
          3950 => x"34",
          3951 => x"0c",
          3952 => x"94",
          3953 => x"5e",
          3954 => x"55",
          3955 => x"90",
          3956 => x"90",
          3957 => x"e4",
          3958 => x"0d",
          3959 => x"52",
          3960 => x"08",
          3961 => x"38",
          3962 => x"81",
          3963 => x"80",
          3964 => x"51",
          3965 => x"08",
          3966 => x"38",
          3967 => x"07",
          3968 => x"16",
          3969 => x"cc",
          3970 => x"15",
          3971 => x"b2",
          3972 => x"ed",
          3973 => x"b7",
          3974 => x"15",
          3975 => x"82",
          3976 => x"bf",
          3977 => x"76",
          3978 => x"04",
          3979 => x"fe",
          3980 => x"82",
          3981 => x"fc",
          3982 => x"82",
          3983 => x"08",
          3984 => x"0c",
          3985 => x"0d",
          3986 => x"e6",
          3987 => x"d5",
          3988 => x"e4",
          3989 => x"71",
          3990 => x"04",
          3991 => x"cc",
          3992 => x"3f",
          3993 => x"e4",
          3994 => x"52",
          3995 => x"3f",
          3996 => x"e4",
          3997 => x"33",
          3998 => x"25",
          3999 => x"54",
          4000 => x"84",
          4001 => x"73",
          4002 => x"70",
          4003 => x"e4",
          4004 => x"d5",
          4005 => x"83",
          4006 => x"0c",
          4007 => x"0d",
          4008 => x"08",
          4009 => x"80",
          4010 => x"e0",
          4011 => x"e4",
          4012 => x"a1",
          4013 => x"7c",
          4014 => x"55",
          4015 => x"80",
          4016 => x"d3",
          4017 => x"82",
          4018 => x"08",
          4019 => x"52",
          4020 => x"d5",
          4021 => x"82",
          4022 => x"7b",
          4023 => x"08",
          4024 => x"51",
          4025 => x"57",
          4026 => x"80",
          4027 => x"d5",
          4028 => x"a7",
          4029 => x"51",
          4030 => x"08",
          4031 => x"c4",
          4032 => x"82",
          4033 => x"76",
          4034 => x"82",
          4035 => x"38",
          4036 => x"74",
          4037 => x"78",
          4038 => x"56",
          4039 => x"c6",
          4040 => x"33",
          4041 => x"16",
          4042 => x"75",
          4043 => x"05",
          4044 => x"11",
          4045 => x"58",
          4046 => x"ff",
          4047 => x"58",
          4048 => x"7b",
          4049 => x"18",
          4050 => x"af",
          4051 => x"33",
          4052 => x"70",
          4053 => x"56",
          4054 => x"70",
          4055 => x"f5",
          4056 => x"a7",
          4057 => x"38",
          4058 => x"81",
          4059 => x"39",
          4060 => x"74",
          4061 => x"91",
          4062 => x"18",
          4063 => x"70",
          4064 => x"eb",
          4065 => x"e4",
          4066 => x"3d",
          4067 => x"54",
          4068 => x"82",
          4069 => x"08",
          4070 => x"72",
          4071 => x"73",
          4072 => x"70",
          4073 => x"57",
          4074 => x"08",
          4075 => x"75",
          4076 => x"11",
          4077 => x"73",
          4078 => x"16",
          4079 => x"e4",
          4080 => x"55",
          4081 => x"e4",
          4082 => x"70",
          4083 => x"71",
          4084 => x"53",
          4085 => x"a7",
          4086 => x"d3",
          4087 => x"d5",
          4088 => x"82",
          4089 => x"38",
          4090 => x"73",
          4091 => x"9f",
          4092 => x"75",
          4093 => x"17",
          4094 => x"70",
          4095 => x"80",
          4096 => x"ff",
          4097 => x"54",
          4098 => x"d5",
          4099 => x"74",
          4100 => x"e4",
          4101 => x"81",
          4102 => x"9c",
          4103 => x"16",
          4104 => x"16",
          4105 => x"53",
          4106 => x"79",
          4107 => x"e4",
          4108 => x"34",
          4109 => x"91",
          4110 => x"89",
          4111 => x"94",
          4112 => x"27",
          4113 => x"15",
          4114 => x"16",
          4115 => x"80",
          4116 => x"2e",
          4117 => x"53",
          4118 => x"0d",
          4119 => x"54",
          4120 => x"53",
          4121 => x"84",
          4122 => x"e4",
          4123 => x"eb",
          4124 => x"51",
          4125 => x"55",
          4126 => x"ab",
          4127 => x"80",
          4128 => x"70",
          4129 => x"57",
          4130 => x"08",
          4131 => x"d5",
          4132 => x"86",
          4133 => x"75",
          4134 => x"e4",
          4135 => x"06",
          4136 => x"80",
          4137 => x"54",
          4138 => x"0d",
          4139 => x"fc",
          4140 => x"3f",
          4141 => x"d5",
          4142 => x"04",
          4143 => x"fc",
          4144 => x"9a",
          4145 => x"d5",
          4146 => x"38",
          4147 => x"ff",
          4148 => x"53",
          4149 => x"52",
          4150 => x"e4",
          4151 => x"2e",
          4152 => x"87",
          4153 => x"74",
          4154 => x"52",
          4155 => x"d5",
          4156 => x"72",
          4157 => x"08",
          4158 => x"d5",
          4159 => x"3d",
          4160 => x"70",
          4161 => x"3f",
          4162 => x"e4",
          4163 => x"d2",
          4164 => x"82",
          4165 => x"cb",
          4166 => x"73",
          4167 => x"39",
          4168 => x"75",
          4169 => x"e4",
          4170 => x"0d",
          4171 => x"3d",
          4172 => x"c5",
          4173 => x"d5",
          4174 => x"0c",
          4175 => x"94",
          4176 => x"74",
          4177 => x"e6",
          4178 => x"5b",
          4179 => x"75",
          4180 => x"81",
          4181 => x"57",
          4182 => x"ff",
          4183 => x"ff",
          4184 => x"81",
          4185 => x"30",
          4186 => x"25",
          4187 => x"5a",
          4188 => x"38",
          4189 => x"d5",
          4190 => x"77",
          4191 => x"ad",
          4192 => x"82",
          4193 => x"70",
          4194 => x"56",
          4195 => x"9e",
          4196 => x"3f",
          4197 => x"06",
          4198 => x"19",
          4199 => x"14",
          4200 => x"e4",
          4201 => x"80",
          4202 => x"54",
          4203 => x"79",
          4204 => x"79",
          4205 => x"07",
          4206 => x"82",
          4207 => x"f9",
          4208 => x"53",
          4209 => x"d5",
          4210 => x"81",
          4211 => x"81",
          4212 => x"2a",
          4213 => x"55",
          4214 => x"17",
          4215 => x"81",
          4216 => x"e4",
          4217 => x"51",
          4218 => x"08",
          4219 => x"39",
          4220 => x"ad",
          4221 => x"2e",
          4222 => x"82",
          4223 => x"06",
          4224 => x"a1",
          4225 => x"9c",
          4226 => x"08",
          4227 => x"51",
          4228 => x"08",
          4229 => x"90",
          4230 => x"90",
          4231 => x"75",
          4232 => x"d5",
          4233 => x"3d",
          4234 => x"05",
          4235 => x"82",
          4236 => x"08",
          4237 => x"08",
          4238 => x"cf",
          4239 => x"d5",
          4240 => x"ff",
          4241 => x"06",
          4242 => x"cb",
          4243 => x"24",
          4244 => x"33",
          4245 => x"76",
          4246 => x"ff",
          4247 => x"74",
          4248 => x"56",
          4249 => x"54",
          4250 => x"2e",
          4251 => x"e4",
          4252 => x"52",
          4253 => x"e4",
          4254 => x"eb",
          4255 => x"51",
          4256 => x"08",
          4257 => x"87",
          4258 => x"08",
          4259 => x"08",
          4260 => x"3f",
          4261 => x"08",
          4262 => x"80",
          4263 => x"95",
          4264 => x"53",
          4265 => x"3f",
          4266 => x"38",
          4267 => x"d5",
          4268 => x"0c",
          4269 => x"82",
          4270 => x"9b",
          4271 => x"e4",
          4272 => x"b7",
          4273 => x"70",
          4274 => x"e4",
          4275 => x"38",
          4276 => x"e4",
          4277 => x"8f",
          4278 => x"85",
          4279 => x"74",
          4280 => x"8a",
          4281 => x"3f",
          4282 => x"82",
          4283 => x"82",
          4284 => x"06",
          4285 => x"08",
          4286 => x"81",
          4287 => x"38",
          4288 => x"ff",
          4289 => x"54",
          4290 => x"8b",
          4291 => x"a4",
          4292 => x"15",
          4293 => x"15",
          4294 => x"ce",
          4295 => x"53",
          4296 => x"ee",
          4297 => x"80",
          4298 => x"78",
          4299 => x"7f",
          4300 => x"ff",
          4301 => x"83",
          4302 => x"3f",
          4303 => x"e4",
          4304 => x"52",
          4305 => x"3f",
          4306 => x"b7",
          4307 => x"15",
          4308 => x"34",
          4309 => x"d5",
          4310 => x"75",
          4311 => x"73",
          4312 => x"04",
          4313 => x"51",
          4314 => x"fe",
          4315 => x"cd",
          4316 => x"d5",
          4317 => x"ab",
          4318 => x"58",
          4319 => x"55",
          4320 => x"02",
          4321 => x"54",
          4322 => x"53",
          4323 => x"80",
          4324 => x"53",
          4325 => x"ff",
          4326 => x"73",
          4327 => x"08",
          4328 => x"63",
          4329 => x"88",
          4330 => x"38",
          4331 => x"e4",
          4332 => x"bb",
          4333 => x"82",
          4334 => x"08",
          4335 => x"aa",
          4336 => x"51",
          4337 => x"33",
          4338 => x"84",
          4339 => x"73",
          4340 => x"8b",
          4341 => x"15",
          4342 => x"70",
          4343 => x"2e",
          4344 => x"e1",
          4345 => x"ad",
          4346 => x"51",
          4347 => x"d5",
          4348 => x"82",
          4349 => x"a3",
          4350 => x"80",
          4351 => x"e4",
          4352 => x"54",
          4353 => x"38",
          4354 => x"b4",
          4355 => x"15",
          4356 => x"9c",
          4357 => x"d5",
          4358 => x"8c",
          4359 => x"82",
          4360 => x"e4",
          4361 => x"0d",
          4362 => x"05",
          4363 => x"53",
          4364 => x"51",
          4365 => x"55",
          4366 => x"78",
          4367 => x"51",
          4368 => x"55",
          4369 => x"80",
          4370 => x"86",
          4371 => x"61",
          4372 => x"7a",
          4373 => x"74",
          4374 => x"83",
          4375 => x"3f",
          4376 => x"d5",
          4377 => x"3d",
          4378 => x"cc",
          4379 => x"3f",
          4380 => x"e4",
          4381 => x"52",
          4382 => x"3f",
          4383 => x"e4",
          4384 => x"33",
          4385 => x"a6",
          4386 => x"71",
          4387 => x"51",
          4388 => x"0b",
          4389 => x"a6",
          4390 => x"82",
          4391 => x"e9",
          4392 => x"53",
          4393 => x"51",
          4394 => x"82",
          4395 => x"e4",
          4396 => x"79",
          4397 => x"75",
          4398 => x"fa",
          4399 => x"8d",
          4400 => x"3f",
          4401 => x"e4",
          4402 => x"51",
          4403 => x"08",
          4404 => x"82",
          4405 => x"65",
          4406 => x"7b",
          4407 => x"34",
          4408 => x"38",
          4409 => x"34",
          4410 => x"70",
          4411 => x"a0",
          4412 => x"2e",
          4413 => x"34",
          4414 => x"80",
          4415 => x"c1",
          4416 => x"a4",
          4417 => x"3f",
          4418 => x"e4",
          4419 => x"55",
          4420 => x"38",
          4421 => x"38",
          4422 => x"ff",
          4423 => x"7b",
          4424 => x"3d",
          4425 => x"9c",
          4426 => x"51",
          4427 => x"82",
          4428 => x"e4",
          4429 => x"52",
          4430 => x"ef",
          4431 => x"56",
          4432 => x"57",
          4433 => x"82",
          4434 => x"80",
          4435 => x"96",
          4436 => x"e4",
          4437 => x"e4",
          4438 => x"80",
          4439 => x"f4",
          4440 => x"e4",
          4441 => x"88",
          4442 => x"39",
          4443 => x"81",
          4444 => x"38",
          4445 => x"81",
          4446 => x"77",
          4447 => x"6d",
          4448 => x"26",
          4449 => x"86",
          4450 => x"38",
          4451 => x"05",
          4452 => x"73",
          4453 => x"ff",
          4454 => x"80",
          4455 => x"55",
          4456 => x"08",
          4457 => x"38",
          4458 => x"3f",
          4459 => x"e4",
          4460 => x"66",
          4461 => x"82",
          4462 => x"06",
          4463 => x"2e",
          4464 => x"ff",
          4465 => x"54",
          4466 => x"53",
          4467 => x"ff",
          4468 => x"8b",
          4469 => x"51",
          4470 => x"0b",
          4471 => x"96",
          4472 => x"55",
          4473 => x"0d",
          4474 => x"88",
          4475 => x"fc",
          4476 => x"d2",
          4477 => x"82",
          4478 => x"1a",
          4479 => x"80",
          4480 => x"78",
          4481 => x"2a",
          4482 => x"90",
          4483 => x"58",
          4484 => x"39",
          4485 => x"70",
          4486 => x"af",
          4487 => x"30",
          4488 => x"e4",
          4489 => x"5a",
          4490 => x"38",
          4491 => x"82",
          4492 => x"74",
          4493 => x"81",
          4494 => x"75",
          4495 => x"e4",
          4496 => x"d5",
          4497 => x"82",
          4498 => x"56",
          4499 => x"38",
          4500 => x"77",
          4501 => x"87",
          4502 => x"ba",
          4503 => x"2e",
          4504 => x"2e",
          4505 => x"75",
          4506 => x"d0",
          4507 => x"d5",
          4508 => x"16",
          4509 => x"38",
          4510 => x"90",
          4511 => x"38",
          4512 => x"0c",
          4513 => x"73",
          4514 => x"05",
          4515 => x"26",
          4516 => x"0c",
          4517 => x"84",
          4518 => x"e4",
          4519 => x"0d",
          4520 => x"05",
          4521 => x"c4",
          4522 => x"d5",
          4523 => x"d5",
          4524 => x"05",
          4525 => x"84",
          4526 => x"08",
          4527 => x"d8",
          4528 => x"47",
          4529 => x"8e",
          4530 => x"ff",
          4531 => x"56",
          4532 => x"70",
          4533 => x"8c",
          4534 => x"83",
          4535 => x"82",
          4536 => x"74",
          4537 => x"80",
          4538 => x"55",
          4539 => x"78",
          4540 => x"26",
          4541 => x"8b",
          4542 => x"80",
          4543 => x"39",
          4544 => x"89",
          4545 => x"83",
          4546 => x"25",
          4547 => x"8b",
          4548 => x"38",
          4549 => x"51",
          4550 => x"d5",
          4551 => x"1b",
          4552 => x"e4",
          4553 => x"56",
          4554 => x"06",
          4555 => x"83",
          4556 => x"2e",
          4557 => x"ff",
          4558 => x"83",
          4559 => x"3f",
          4560 => x"9a",
          4561 => x"51",
          4562 => x"d5",
          4563 => x"2a",
          4564 => x"41",
          4565 => x"67",
          4566 => x"c5",
          4567 => x"80",
          4568 => x"56",
          4569 => x"62",
          4570 => x"74",
          4571 => x"55",
          4572 => x"81",
          4573 => x"38",
          4574 => x"5e",
          4575 => x"5a",
          4576 => x"e1",
          4577 => x"57",
          4578 => x"5a",
          4579 => x"26",
          4580 => x"10",
          4581 => x"74",
          4582 => x"ee",
          4583 => x"ef",
          4584 => x"84",
          4585 => x"a0",
          4586 => x"fc",
          4587 => x"f0",
          4588 => x"88",
          4589 => x"57",
          4590 => x"5a",
          4591 => x"26",
          4592 => x"10",
          4593 => x"74",
          4594 => x"ee",
          4595 => x"8f",
          4596 => x"05",
          4597 => x"26",
          4598 => x"08",
          4599 => x"11",
          4600 => x"83",
          4601 => x"a0",
          4602 => x"6a",
          4603 => x"72",
          4604 => x"59",
          4605 => x"89",
          4606 => x"84",
          4607 => x"18",
          4608 => x"74",
          4609 => x"31",
          4610 => x"52",
          4611 => x"e4",
          4612 => x"06",
          4613 => x"ff",
          4614 => x"b8",
          4615 => x"be",
          4616 => x"09",
          4617 => x"f5",
          4618 => x"38",
          4619 => x"80",
          4620 => x"96",
          4621 => x"2e",
          4622 => x"82",
          4623 => x"38",
          4624 => x"81",
          4625 => x"e0",
          4626 => x"81",
          4627 => x"78",
          4628 => x"8e",
          4629 => x"53",
          4630 => x"3f",
          4631 => x"51",
          4632 => x"8b",
          4633 => x"8d",
          4634 => x"52",
          4635 => x"81",
          4636 => x"70",
          4637 => x"54",
          4638 => x"ff",
          4639 => x"26",
          4640 => x"52",
          4641 => x"8a",
          4642 => x"8d",
          4643 => x"bf",
          4644 => x"3f",
          4645 => x"8d",
          4646 => x"ff",
          4647 => x"81",
          4648 => x"0a",
          4649 => x"c5",
          4650 => x"8d",
          4651 => x"ff",
          4652 => x"51",
          4653 => x"1b",
          4654 => x"0b",
          4655 => x"c2",
          4656 => x"52",
          4657 => x"88",
          4658 => x"8c",
          4659 => x"52",
          4660 => x"ff",
          4661 => x"a6",
          4662 => x"52",
          4663 => x"82",
          4664 => x"52",
          4665 => x"7e",
          4666 => x"ce",
          4667 => x"84",
          4668 => x"06",
          4669 => x"53",
          4670 => x"3f",
          4671 => x"ff",
          4672 => x"d2",
          4673 => x"86",
          4674 => x"1b",
          4675 => x"52",
          4676 => x"3f",
          4677 => x"8b",
          4678 => x"51",
          4679 => x"1f",
          4680 => x"de",
          4681 => x"52",
          4682 => x"53",
          4683 => x"3f",
          4684 => x"09",
          4685 => x"51",
          4686 => x"1b",
          4687 => x"52",
          4688 => x"ff",
          4689 => x"f8",
          4690 => x"fd",
          4691 => x"26",
          4692 => x"53",
          4693 => x"3f",
          4694 => x"84",
          4695 => x"7a",
          4696 => x"75",
          4697 => x"81",
          4698 => x"38",
          4699 => x"65",
          4700 => x"38",
          4701 => x"52",
          4702 => x"d5",
          4703 => x"75",
          4704 => x"8c",
          4705 => x"57",
          4706 => x"84",
          4707 => x"57",
          4708 => x"80",
          4709 => x"8c",
          4710 => x"81",
          4711 => x"76",
          4712 => x"d5",
          4713 => x"ff",
          4714 => x"83",
          4715 => x"38",
          4716 => x"ff",
          4717 => x"78",
          4718 => x"1b",
          4719 => x"16",
          4720 => x"83",
          4721 => x"1f",
          4722 => x"fe",
          4723 => x"34",
          4724 => x"07",
          4725 => x"e4",
          4726 => x"c6",
          4727 => x"52",
          4728 => x"3f",
          4729 => x"51",
          4730 => x"d5",
          4731 => x"52",
          4732 => x"56",
          4733 => x"39",
          4734 => x"39",
          4735 => x"d5",
          4736 => x"3d",
          4737 => x"60",
          4738 => x"25",
          4739 => x"55",
          4740 => x"c8",
          4741 => x"06",
          4742 => x"8d",
          4743 => x"05",
          4744 => x"2e",
          4745 => x"34",
          4746 => x"74",
          4747 => x"04",
          4748 => x"b3",
          4749 => x"09",
          4750 => x"51",
          4751 => x"76",
          4752 => x"17",
          4753 => x"81",
          4754 => x"8b",
          4755 => x"17",
          4756 => x"79",
          4757 => x"9f",
          4758 => x"75",
          4759 => x"0c",
          4760 => x"79",
          4761 => x"24",
          4762 => x"74",
          4763 => x"c9",
          4764 => x"38",
          4765 => x"06",
          4766 => x"39",
          4767 => x"89",
          4768 => x"54",
          4769 => x"ff",
          4770 => x"3d",
          4771 => x"e3",
          4772 => x"53",
          4773 => x"51",
          4774 => x"3f",
          4775 => x"75",
          4776 => x"53",
          4777 => x"38",
          4778 => x"c3",
          4779 => x"73",
          4780 => x"38",
          4781 => x"a8",
          4782 => x"81",
          4783 => x"51",
          4784 => x"10",
          4785 => x"51",
          4786 => x"ff",
          4787 => x"0c",
          4788 => x"02",
          4789 => x"05",
          4790 => x"ff",
          4791 => x"71",
          4792 => x"38",
          4793 => x"10",
          4794 => x"51",
          4795 => x"0d",
          4796 => x"83",
          4797 => x"83",
          4798 => x"52",
          4799 => x"cf",
          4800 => x"22",
          4801 => x"26",
          4802 => x"38",
          4803 => x"88",
          4804 => x"54",
          4805 => x"d7",
          4806 => x"73",
          4807 => x"70",
          4808 => x"11",
          4809 => x"39",
          4810 => x"31",
          4811 => x"9f",
          4812 => x"12",
          4813 => x"39",
          4814 => x"12",
          4815 => x"70",
          4816 => x"73",
          4817 => x"fe",
          4818 => x"e4",
          4819 => x"ff",
          4820 => x"00",
          4821 => x"2c",
          4822 => x"2b",
          4823 => x"2b",
          4824 => x"2b",
          4825 => x"2c",
          4826 => x"2c",
          4827 => x"2c",
          4828 => x"2c",
          4829 => x"2c",
          4830 => x"2c",
          4831 => x"42",
          4832 => x"42",
          4833 => x"42",
          4834 => x"49",
          4835 => x"4c",
          4836 => x"46",
          4837 => x"4c",
          4838 => x"4b",
          4839 => x"49",
          4840 => x"4a",
          4841 => x"4b",
          4842 => x"46",
          4843 => x"4b",
          4844 => x"4c",
          4845 => x"96",
          4846 => x"96",
          4847 => x"96",
          4848 => x"96",
          4849 => x"0e",
          4850 => x"17",
          4851 => x"17",
          4852 => x"17",
          4853 => x"17",
          4854 => x"17",
          4855 => x"17",
          4856 => x"0e",
          4857 => x"17",
          4858 => x"17",
          4859 => x"17",
          4860 => x"17",
          4861 => x"17",
          4862 => x"17",
          4863 => x"17",
          4864 => x"17",
          4865 => x"17",
          4866 => x"17",
          4867 => x"17",
          4868 => x"17",
          4869 => x"17",
          4870 => x"17",
          4871 => x"17",
          4872 => x"17",
          4873 => x"17",
          4874 => x"17",
          4875 => x"17",
          4876 => x"17",
          4877 => x"11",
          4878 => x"17",
          4879 => x"17",
          4880 => x"17",
          4881 => x"17",
          4882 => x"17",
          4883 => x"10",
          4884 => x"0e",
          4885 => x"17",
          4886 => x"17",
          4887 => x"0e",
          4888 => x"17",
          4889 => x"10",
          4890 => x"17",
          4891 => x"17",
          4892 => x"17",
          4893 => x"11",
          4894 => x"00",
          4895 => x"00",
          4896 => x"00",
          4897 => x"00",
          4898 => x"00",
          4899 => x"00",
          4900 => x"00",
          4901 => x"00",
          4902 => x"00",
          4903 => x"68",
          4904 => x"64",
          4905 => x"64",
          4906 => x"6c",
          4907 => x"70",
          4908 => x"74",
          4909 => x"00",
          4910 => x"00",
          4911 => x"00",
          4912 => x"00",
          4913 => x"00",
          4914 => x"00",
          4915 => x"73",
          4916 => x"00",
          4917 => x"61",
          4918 => x"2e",
          4919 => x"6f",
          4920 => x"2e",
          4921 => x"65",
          4922 => x"00",
          4923 => x"68",
          4924 => x"00",
          4925 => x"64",
          4926 => x"6d",
          4927 => x"63",
          4928 => x"69",
          4929 => x"6c",
          4930 => x"64",
          4931 => x"73",
          4932 => x"6c",
          4933 => x"65",
          4934 => x"64",
          4935 => x"20",
          4936 => x"65",
          4937 => x"74",
          4938 => x"69",
          4939 => x"65",
          4940 => x"76",
          4941 => x"00",
          4942 => x"6f",
          4943 => x"65",
          4944 => x"20",
          4945 => x"62",
          4946 => x"73",
          4947 => x"6f",
          4948 => x"64",
          4949 => x"72",
          4950 => x"72",
          4951 => x"6d",
          4952 => x"70",
          4953 => x"20",
          4954 => x"65",
          4955 => x"6c",
          4956 => x"63",
          4957 => x"73",
          4958 => x"6e",
          4959 => x"79",
          4960 => x"6f",
          4961 => x"70",
          4962 => x"73",
          4963 => x"72",
          4964 => x"20",
          4965 => x"63",
          4966 => x"63",
          4967 => x"00",
          4968 => x"6e",
          4969 => x"00",
          4970 => x"79",
          4971 => x"61",
          4972 => x"79",
          4973 => x"2e",
          4974 => x"61",
          4975 => x"38",
          4976 => x"20",
          4977 => x"00",
          4978 => x"20",
          4979 => x"32",
          4980 => x"00",
          4981 => x"00",
          4982 => x"2a",
          4983 => x"00",
          4984 => x"32",
          4985 => x"2e",
          4986 => x"50",
          4987 => x"25",
          4988 => x"20",
          4989 => x"00",
          4990 => x"74",
          4991 => x"48",
          4992 => x"00",
          4993 => x"69",
          4994 => x"74",
          4995 => x"74",
          4996 => x"00",
          4997 => x"52",
          4998 => x"72",
          4999 => x"43",
          5000 => x"6e",
          5001 => x"00",
          5002 => x"52",
          5003 => x"72",
          5004 => x"52",
          5005 => x"6e",
          5006 => x"00",
          5007 => x"52",
          5008 => x"72",
          5009 => x"52",
          5010 => x"6e",
          5011 => x"00",
          5012 => x"67",
          5013 => x"65",
          5014 => x"61",
          5015 => x"69",
          5016 => x"00",
          5017 => x"65",
          5018 => x"00",
          5019 => x"75",
          5020 => x"00",
          5021 => x"20",
          5022 => x"69",
          5023 => x"64",
          5024 => x"2c",
          5025 => x"20",
          5026 => x"6e",
          5027 => x"00",
          5028 => x"65",
          5029 => x"2e",
          5030 => x"70",
          5031 => x"00",
          5032 => x"69",
          5033 => x"00",
          5034 => x"25",
          5035 => x"30",
          5036 => x"78",
          5037 => x"6d",
          5038 => x"79",
          5039 => x"65",
          5040 => x"38",
          5041 => x"2d",
          5042 => x"38",
          5043 => x"2d",
          5044 => x"25",
          5045 => x"00",
          5046 => x"69",
          5047 => x"20",
          5048 => x"20",
          5049 => x"6c",
          5050 => x"64",
          5051 => x"6c",
          5052 => x"00",
          5053 => x"65",
          5054 => x"63",
          5055 => x"29",
          5056 => x"73",
          5057 => x"20",
          5058 => x"74",
          5059 => x"00",
          5060 => x"65",
          5061 => x"2e",
          5062 => x"55",
          5063 => x"3a",
          5064 => x"25",
          5065 => x"3a",
          5066 => x"00",
          5067 => x"00",
          5068 => x"6d",
          5069 => x"00",
          5070 => x"20",
          5071 => x"65",
          5072 => x"6f",
          5073 => x"73",
          5074 => x"6e",
          5075 => x"6e",
          5076 => x"00",
          5077 => x"6e",
          5078 => x"72",
          5079 => x"00",
          5080 => x"25",
          5081 => x"3a",
          5082 => x"0a",
          5083 => x"6e",
          5084 => x"69",
          5085 => x"66",
          5086 => x"20",
          5087 => x"00",
          5088 => x"63",
          5089 => x"65",
          5090 => x"00",
          5091 => x"20",
          5092 => x"28",
          5093 => x"38",
          5094 => x"20",
          5095 => x"20",
          5096 => x"58",
          5097 => x"0a",
          5098 => x"53",
          5099 => x"28",
          5100 => x"38",
          5101 => x"20",
          5102 => x"20",
          5103 => x"58",
          5104 => x"0a",
          5105 => x"4d",
          5106 => x"28",
          5107 => x"38",
          5108 => x"20",
          5109 => x"44",
          5110 => x"69",
          5111 => x"32",
          5112 => x"20",
          5113 => x"20",
          5114 => x"65",
          5115 => x"32",
          5116 => x"20",
          5117 => x"54",
          5118 => x"6e",
          5119 => x"32",
          5120 => x"20",
          5121 => x"4e",
          5122 => x"00",
          5123 => x"20",
          5124 => x"20",
          5125 => x"00",
          5126 => x"32",
          5127 => x"49",
          5128 => x"73",
          5129 => x"20",
          5130 => x"73",
          5131 => x"6f",
          5132 => x"73",
          5133 => x"58",
          5134 => x"20",
          5135 => x"6d",
          5136 => x"72",
          5137 => x"73",
          5138 => x"58",
          5139 => x"20",
          5140 => x"53",
          5141 => x"64",
          5142 => x"20",
          5143 => x"58",
          5144 => x"73",
          5145 => x"20",
          5146 => x"20",
          5147 => x"20",
          5148 => x"20",
          5149 => x"58",
          5150 => x"20",
          5151 => x"20",
          5152 => x"72",
          5153 => x"20",
          5154 => x"25",
          5155 => x"00",
          5156 => x"52",
          5157 => x"6b",
          5158 => x"20",
          5159 => x"20",
          5160 => x"4d",
          5161 => x"20",
          5162 => x"6e",
          5163 => x"20",
          5164 => x"72",
          5165 => x"25",
          5166 => x"00",
          5167 => x"00",
          5168 => x"00",
          5169 => x"00",
          5170 => x"4f",
          5171 => x"6b",
          5172 => x"a3",
          5173 => x"00",
          5174 => x"00",
          5175 => x"a2",
          5176 => x"00",
          5177 => x"00",
          5178 => x"a2",
          5179 => x"00",
          5180 => x"00",
          5181 => x"a2",
          5182 => x"00",
          5183 => x"00",
          5184 => x"a2",
          5185 => x"00",
          5186 => x"00",
          5187 => x"a2",
          5188 => x"00",
          5189 => x"00",
          5190 => x"a2",
          5191 => x"00",
          5192 => x"00",
          5193 => x"a2",
          5194 => x"00",
          5195 => x"00",
          5196 => x"a2",
          5197 => x"00",
          5198 => x"00",
          5199 => x"a2",
          5200 => x"00",
          5201 => x"00",
          5202 => x"a2",
          5203 => x"00",
          5204 => x"00",
          5205 => x"44",
          5206 => x"42",
          5207 => x"36",
          5208 => x"34",
          5209 => x"33",
          5210 => x"31",
          5211 => x"00",
          5212 => x"00",
          5213 => x"00",
          5214 => x"00",
          5215 => x"00",
          5216 => x"73",
          5217 => x"73",
          5218 => x"00",
          5219 => x"20",
          5220 => x"69",
          5221 => x"72",
          5222 => x"65",
          5223 => x"79",
          5224 => x"6f",
          5225 => x"00",
          5226 => x"20",
          5227 => x"65",
          5228 => x"74",
          5229 => x"65",
          5230 => x"6c",
          5231 => x"00",
          5232 => x"7c",
          5233 => x"3b",
          5234 => x"54",
          5235 => x"00",
          5236 => x"4f",
          5237 => x"20",
          5238 => x"20",
          5239 => x"20",
          5240 => x"45",
          5241 => x"20",
          5242 => x"a3",
          5243 => x"00",
          5244 => x"05",
          5245 => x"18",
          5246 => x"45",
          5247 => x"45",
          5248 => x"92",
          5249 => x"9a",
          5250 => x"4f",
          5251 => x"aa",
          5252 => x"b2",
          5253 => x"ba",
          5254 => x"c2",
          5255 => x"ca",
          5256 => x"d2",
          5257 => x"da",
          5258 => x"e2",
          5259 => x"ea",
          5260 => x"f2",
          5261 => x"fa",
          5262 => x"2c",
          5263 => x"2a",
          5264 => x"00",
          5265 => x"00",
          5266 => x"00",
          5267 => x"00",
          5268 => x"00",
          5269 => x"00",
          5270 => x"00",
          5271 => x"00",
          5272 => x"00",
          5273 => x"00",
          5274 => x"00",
          5275 => x"00",
          5276 => x"01",
          5277 => x"00",
          5278 => x"00",
          5279 => x"00",
          5280 => x"00",
          5281 => x"25",
          5282 => x"25",
          5283 => x"25",
          5284 => x"25",
          5285 => x"25",
          5286 => x"25",
          5287 => x"25",
          5288 => x"25",
          5289 => x"25",
          5290 => x"25",
          5291 => x"25",
          5292 => x"25",
          5293 => x"03",
          5294 => x"03",
          5295 => x"03",
          5296 => x"22",
          5297 => x"22",
          5298 => x"22",
          5299 => x"22",
          5300 => x"00",
          5301 => x"03",
          5302 => x"00",
          5303 => x"01",
          5304 => x"01",
          5305 => x"01",
          5306 => x"01",
          5307 => x"01",
          5308 => x"01",
          5309 => x"01",
          5310 => x"01",
          5311 => x"01",
          5312 => x"02",
          5313 => x"02",
          5314 => x"01",
          5315 => x"01",
          5316 => x"01",
          5317 => x"01",
          5318 => x"01",
          5319 => x"01",
          5320 => x"01",
          5321 => x"01",
          5322 => x"01",
          5323 => x"01",
          5324 => x"01",
          5325 => x"01",
          5326 => x"01",
          5327 => x"01",
          5328 => x"01",
          5329 => x"00",
          5330 => x"02",
          5331 => x"02",
          5332 => x"02",
          5333 => x"02",
          5334 => x"01",
          5335 => x"02",
          5336 => x"02",
          5337 => x"02",
          5338 => x"01",
          5339 => x"02",
          5340 => x"02",
          5341 => x"01",
          5342 => x"02",
          5343 => x"2c",
          5344 => x"02",
          5345 => x"02",
          5346 => x"02",
          5347 => x"02",
          5348 => x"02",
          5349 => x"03",
          5350 => x"00",
          5351 => x"03",
          5352 => x"00",
          5353 => x"03",
          5354 => x"03",
          5355 => x"03",
          5356 => x"03",
          5357 => x"03",
          5358 => x"04",
          5359 => x"04",
          5360 => x"04",
          5361 => x"04",
          5362 => x"04",
          5363 => x"00",
          5364 => x"1e",
          5365 => x"1f",
          5366 => x"1f",
          5367 => x"1f",
          5368 => x"1f",
          5369 => x"1f",
          5370 => x"00",
          5371 => x"1f",
          5372 => x"1f",
          5373 => x"1f",
          5374 => x"06",
          5375 => x"06",
          5376 => x"1f",
          5377 => x"00",
          5378 => x"1f",
          5379 => x"1f",
          5380 => x"21",
          5381 => x"02",
          5382 => x"24",
          5383 => x"2c",
          5384 => x"2c",
          5385 => x"2d",
          5386 => x"00",
          5387 => x"98",
          5388 => x"00",
          5389 => x"98",
          5390 => x"00",
          5391 => x"99",
          5392 => x"00",
          5393 => x"99",
          5394 => x"00",
          5395 => x"99",
          5396 => x"00",
          5397 => x"99",
          5398 => x"00",
          5399 => x"99",
          5400 => x"00",
          5401 => x"99",
          5402 => x"00",
          5403 => x"99",
          5404 => x"00",
          5405 => x"99",
          5406 => x"00",
          5407 => x"99",
          5408 => x"00",
          5409 => x"99",
          5410 => x"00",
          5411 => x"99",
          5412 => x"00",
          5413 => x"99",
          5414 => x"00",
          5415 => x"99",
          5416 => x"00",
          5417 => x"99",
          5418 => x"00",
          5419 => x"99",
          5420 => x"00",
          5421 => x"99",
          5422 => x"00",
          5423 => x"99",
          5424 => x"00",
          5425 => x"99",
          5426 => x"00",
          5427 => x"99",
          5428 => x"00",
          5429 => x"99",
          5430 => x"00",
          5431 => x"99",
          5432 => x"00",
          5433 => x"99",
          5434 => x"00",
          5435 => x"99",
          5436 => x"00",
          5437 => x"99",
          5438 => x"00",
          5439 => x"00",
          5440 => x"7f",
          5441 => x"7f",
          5442 => x"7f",
          5443 => x"00",
          5444 => x"ff",
          5445 => x"00",
          5446 => x"00",
          5447 => x"e1",
          5448 => x"00",
          5449 => x"01",
          5450 => x"00",
          5451 => x"00",
          5452 => x"00",
          5453 => x"00",
          5454 => x"00",
          5455 => x"00",
          5456 => x"00",
          5457 => x"00",
          5458 => x"00",
          5459 => x"00",
          5460 => x"00",
          5461 => x"00",
          5462 => x"00",
          5463 => x"00",
          5464 => x"00",
          5465 => x"00",
          5466 => x"00",
          5467 => x"00",
          5468 => x"00",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"85",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"90",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"91",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"82",
           193 => x"82",
           194 => x"82",
           195 => x"d5",
           196 => x"d5",
           197 => x"f0",
           198 => x"f0",
           199 => x"08",
           200 => x"0c",
           201 => x"84",
           202 => x"b1",
           203 => x"80",
           204 => x"d0",
           205 => x"80",
           206 => x"cb",
           207 => x"80",
           208 => x"d8",
           209 => x"90",
           210 => x"2d",
           211 => x"04",
           212 => x"82",
           213 => x"82",
           214 => x"82",
           215 => x"82",
           216 => x"82",
           217 => x"82",
           218 => x"82",
           219 => x"82",
           220 => x"82",
           221 => x"82",
           222 => x"82",
           223 => x"82",
           224 => x"82",
           225 => x"82",
           226 => x"82",
           227 => x"82",
           228 => x"82",
           229 => x"82",
           230 => x"82",
           231 => x"82",
           232 => x"82",
           233 => x"82",
           234 => x"82",
           235 => x"82",
           236 => x"82",
           237 => x"82",
           238 => x"82",
           239 => x"82",
           240 => x"82",
           241 => x"82",
           242 => x"82",
           243 => x"82",
           244 => x"82",
           245 => x"82",
           246 => x"82",
           247 => x"82",
           248 => x"82",
           249 => x"82",
           250 => x"82",
           251 => x"82",
           252 => x"82",
           253 => x"82",
           254 => x"82",
           255 => x"82",
           256 => x"82",
           257 => x"82",
           258 => x"82",
           259 => x"82",
           260 => x"82",
           261 => x"82",
           262 => x"82",
           263 => x"82",
           264 => x"82",
           265 => x"82",
           266 => x"82",
           267 => x"82",
           268 => x"82",
           269 => x"82",
           270 => x"82",
           271 => x"82",
           272 => x"82",
           273 => x"82",
           274 => x"82",
           275 => x"82",
           276 => x"82",
           277 => x"82",
           278 => x"82",
           279 => x"82",
           280 => x"82",
           281 => x"82",
           282 => x"82",
           283 => x"82",
           284 => x"82",
           285 => x"82",
           286 => x"82",
           287 => x"82",
           288 => x"82",
           289 => x"82",
           290 => x"82",
           291 => x"82",
           292 => x"82",
           293 => x"82",
           294 => x"82",
           295 => x"82",
           296 => x"82",
           297 => x"82",
           298 => x"82",
           299 => x"3c",
           300 => x"10",
           301 => x"10",
           302 => x"10",
           303 => x"10",
           304 => x"73",
           305 => x"81",
           306 => x"07",
           307 => x"72",
           308 => x"09",
           309 => x"0a",
           310 => x"51",
           311 => x"82",
           312 => x"70",
           313 => x"93",
           314 => x"c8",
           315 => x"82",
           316 => x"d5",
           317 => x"f0",
           318 => x"08",
           319 => x"08",
           320 => x"08",
           321 => x"e4",
           322 => x"05",
           323 => x"08",
           324 => x"87",
           325 => x"82",
           326 => x"0c",
           327 => x"90",
           328 => x"32",
           329 => x"71",
           330 => x"08",
           331 => x"39",
           332 => x"05",
           333 => x"08",
           334 => x"f0",
           335 => x"d5",
           336 => x"f0",
           337 => x"08",
           338 => x"f8",
           339 => x"80",
           340 => x"08",
           341 => x"08",
           342 => x"82",
           343 => x"08",
           344 => x"08",
           345 => x"06",
           346 => x"08",
           347 => x"d5",
           348 => x"f0",
           349 => x"73",
           350 => x"08",
           351 => x"05",
           352 => x"08",
           353 => x"05",
           354 => x"08",
           355 => x"82",
           356 => x"82",
           357 => x"82",
           358 => x"d5",
           359 => x"f0",
           360 => x"82",
           361 => x"0b",
           362 => x"82",
           363 => x"d5",
           364 => x"0b",
           365 => x"82",
           366 => x"d5",
           367 => x"f0",
           368 => x"f0",
           369 => x"f0",
           370 => x"81",
           371 => x"82",
           372 => x"d5",
           373 => x"f0",
           374 => x"80",
           375 => x"05",
           376 => x"8e",
           377 => x"82",
           378 => x"0c",
           379 => x"90",
           380 => x"05",
           381 => x"08",
           382 => x"08",
           383 => x"08",
           384 => x"08",
           385 => x"0c",
           386 => x"70",
           387 => x"3d",
           388 => x"d5",
           389 => x"ed",
           390 => x"08",
           391 => x"88",
           392 => x"0c",
           393 => x"85",
           394 => x"32",
           395 => x"53",
           396 => x"82",
           397 => x"ac",
           398 => x"08",
           399 => x"f0",
           400 => x"06",
           401 => x"82",
           402 => x"05",
           403 => x"82",
           404 => x"81",
           405 => x"8b",
           406 => x"33",
           407 => x"82",
           408 => x"72",
           409 => x"f0",
           410 => x"2e",
           411 => x"d5",
           412 => x"2b",
           413 => x"b2",
           414 => x"22",
           415 => x"81",
           416 => x"2e",
           417 => x"05",
           418 => x"72",
           419 => x"fe",
           420 => x"05",
           421 => x"70",
           422 => x"51",
           423 => x"82",
           424 => x"d5",
           425 => x"d5",
           426 => x"d0",
           427 => x"f0",
           428 => x"08",
           429 => x"98",
           430 => x"8b",
           431 => x"08",
           432 => x"e4",
           433 => x"06",
           434 => x"82",
           435 => x"88",
           436 => x"70",
           437 => x"72",
           438 => x"fd",
           439 => x"05",
           440 => x"51",
           441 => x"82",
           442 => x"98",
           443 => x"72",
           444 => x"08",
           445 => x"f8",
           446 => x"08",
           447 => x"08",
           448 => x"94",
           449 => x"08",
           450 => x"70",
           451 => x"82",
           452 => x"90",
           453 => x"08",
           454 => x"e4",
           455 => x"72",
           456 => x"fc",
           457 => x"05",
           458 => x"72",
           459 => x"fc",
           460 => x"05",
           461 => x"72",
           462 => x"fb",
           463 => x"05",
           464 => x"82",
           465 => x"0b",
           466 => x"fb",
           467 => x"05",
           468 => x"82",
           469 => x"c1",
           470 => x"fc",
           471 => x"05",
           472 => x"d5",
           473 => x"0b",
           474 => x"8d",
           475 => x"05",
           476 => x"08",
           477 => x"05",
           478 => x"d5",
           479 => x"f0",
           480 => x"53",
           481 => x"23",
           482 => x"90",
           483 => x"05",
           484 => x"90",
           485 => x"08",
           486 => x"e4",
           487 => x"06",
           488 => x"ab",
           489 => x"33",
           490 => x"53",
           491 => x"52",
           492 => x"08",
           493 => x"05",
           494 => x"fc",
           495 => x"d5",
           496 => x"08",
           497 => x"ec",
           498 => x"f4",
           499 => x"72",
           500 => x"8b",
           501 => x"05",
           502 => x"08",
           503 => x"05",
           504 => x"fc",
           505 => x"05",
           506 => x"51",
           507 => x"38",
           508 => x"70",
           509 => x"82",
           510 => x"53",
           511 => x"53",
           512 => x"23",
           513 => x"05",
           514 => x"e4",
           515 => x"f4",
           516 => x"05",
           517 => x"05",
           518 => x"82",
           519 => x"c1",
           520 => x"22",
           521 => x"51",
           522 => x"d5",
           523 => x"f0",
           524 => x"d5",
           525 => x"82",
           526 => x"a2",
           527 => x"08",
           528 => x"84",
           529 => x"0c",
           530 => x"05",
           531 => x"05",
           532 => x"0c",
           533 => x"80",
           534 => x"e4",
           535 => x"72",
           536 => x"82",
           537 => x"82",
           538 => x"d5",
           539 => x"bf",
           540 => x"08",
           541 => x"0b",
           542 => x"a9",
           543 => x"22",
           544 => x"82",
           545 => x"f8",
           546 => x"34",
           547 => x"05",
           548 => x"22",
           549 => x"51",
           550 => x"d5",
           551 => x"f0",
           552 => x"d5",
           553 => x"82",
           554 => x"a2",
           555 => x"08",
           556 => x"84",
           557 => x"0c",
           558 => x"05",
           559 => x"05",
           560 => x"0c",
           561 => x"70",
           562 => x"f0",
           563 => x"0b",
           564 => x"82",
           565 => x"d5",
           566 => x"f0",
           567 => x"54",
           568 => x"d5",
           569 => x"d5",
           570 => x"f0",
           571 => x"08",
           572 => x"89",
           573 => x"08",
           574 => x"82",
           575 => x"15",
           576 => x"d5",
           577 => x"82",
           578 => x"72",
           579 => x"d5",
           580 => x"f0",
           581 => x"f0",
           582 => x"d5",
           583 => x"82",
           584 => x"d5",
           585 => x"82",
           586 => x"53",
           587 => x"70",
           588 => x"53",
           589 => x"80",
           590 => x"d5",
           591 => x"f4",
           592 => x"31",
           593 => x"fc",
           594 => x"05",
           595 => x"80",
           596 => x"ec",
           597 => x"82",
           598 => x"d5",
           599 => x"2a",
           600 => x"80",
           601 => x"08",
           602 => x"d5",
           603 => x"f0",
           604 => x"d5",
           605 => x"f0",
           606 => x"90",
           607 => x"d5",
           608 => x"53",
           609 => x"23",
           610 => x"05",
           611 => x"f0",
           612 => x"08",
           613 => x"ec",
           614 => x"05",
           615 => x"51",
           616 => x"38",
           617 => x"70",
           618 => x"f0",
           619 => x"53",
           620 => x"f0",
           621 => x"51",
           622 => x"05",
           623 => x"e8",
           624 => x"fc",
           625 => x"72",
           626 => x"82",
           627 => x"83",
           628 => x"72",
           629 => x"08",
           630 => x"90",
           631 => x"51",
           632 => x"d5",
           633 => x"31",
           634 => x"ec",
           635 => x"08",
           636 => x"90",
           637 => x"51",
           638 => x"d5",
           639 => x"31",
           640 => x"ec",
           641 => x"05",
           642 => x"72",
           643 => x"05",
           644 => x"d5",
           645 => x"2b",
           646 => x"25",
           647 => x"05",
           648 => x"d2",
           649 => x"22",
           650 => x"51",
           651 => x"d5",
           652 => x"51",
           653 => x"d5",
           654 => x"2a",
           655 => x"80",
           656 => x"88",
           657 => x"3f",
           658 => x"05",
           659 => x"51",
           660 => x"82",
           661 => x"a0",
           662 => x"08",
           663 => x"81",
           664 => x"b1",
           665 => x"08",
           666 => x"d5",
           667 => x"90",
           668 => x"d5",
           669 => x"d5",
           670 => x"bc",
           671 => x"22",
           672 => x"51",
           673 => x"d5",
           674 => x"54",
           675 => x"05",
           676 => x"51",
           677 => x"d5",
           678 => x"51",
           679 => x"f0",
           680 => x"70",
           681 => x"2e",
           682 => x"05",
           683 => x"d5",
           684 => x"2b",
           685 => x"25",
           686 => x"05",
           687 => x"d2",
           688 => x"22",
           689 => x"51",
           690 => x"08",
           691 => x"72",
           692 => x"73",
           693 => x"80",
           694 => x"08",
           695 => x"f4",
           696 => x"f8",
           697 => x"09",
           698 => x"08",
           699 => x"08",
           700 => x"81",
           701 => x"05",
           702 => x"81",
           703 => x"08",
           704 => x"72",
           705 => x"72",
           706 => x"ff",
           707 => x"f0",
           708 => x"f0",
           709 => x"82",
           710 => x"05",
           711 => x"53",
           712 => x"d5",
           713 => x"80",
           714 => x"38",
           715 => x"ff",
           716 => x"08",
           717 => x"06",
           718 => x"df",
           719 => x"08",
           720 => x"08",
           721 => x"82",
           722 => x"05",
           723 => x"ff",
           724 => x"05",
           725 => x"82",
           726 => x"82",
           727 => x"05",
           728 => x"82",
           729 => x"33",
           730 => x"82",
           731 => x"87",
           732 => x"72",
           733 => x"f0",
           734 => x"54",
           735 => x"23",
           736 => x"53",
           737 => x"f0",
           738 => x"85",
           739 => x"08",
           740 => x"08",
           741 => x"80",
           742 => x"23",
           743 => x"f8",
           744 => x"81",
           745 => x"f0",
           746 => x"d5",
           747 => x"82",
           748 => x"0b",
           749 => x"ea",
           750 => x"05",
           751 => x"05",
           752 => x"39",
           753 => x"8c",
           754 => x"e0",
           755 => x"08",
           756 => x"95",
           757 => x"82",
           758 => x"0c",
           759 => x"53",
           760 => x"52",
           761 => x"51",
           762 => x"70",
           763 => x"0d",
           764 => x"f0",
           765 => x"3d",
           766 => x"f8",
           767 => x"11",
           768 => x"70",
           769 => x"72",
           770 => x"d5",
           771 => x"39",
           772 => x"53",
           773 => x"05",
           774 => x"88",
           775 => x"08",
           776 => x"53",
           777 => x"c8",
           778 => x"d5",
           779 => x"11",
           780 => x"e4",
           781 => x"38",
           782 => x"05",
           783 => x"08",
           784 => x"51",
           785 => x"d5",
           786 => x"38",
           787 => x"05",
           788 => x"08",
           789 => x"0c",
           790 => x"08",
           791 => x"82",
           792 => x"08",
           793 => x"0d",
           794 => x"05",
           795 => x"08",
           796 => x"81",
           797 => x"51",
           798 => x"0b",
           799 => x"80",
           800 => x"05",
           801 => x"08",
           802 => x"f0",
           803 => x"d5",
           804 => x"ff",
           805 => x"82",
           806 => x"d5",
           807 => x"d5",
           808 => x"11",
           809 => x"e4",
           810 => x"38",
           811 => x"05",
           812 => x"08",
           813 => x"08",
           814 => x"08",
           815 => x"87",
           816 => x"82",
           817 => x"0c",
           818 => x"52",
           819 => x"51",
           820 => x"82",
           821 => x"82",
           822 => x"08",
           823 => x"0d",
           824 => x"85",
           825 => x"32",
           826 => x"53",
           827 => x"82",
           828 => x"cb",
           829 => x"08",
           830 => x"81",
           831 => x"2e",
           832 => x"8c",
           833 => x"05",
           834 => x"14",
           835 => x"08",
           836 => x"d5",
           837 => x"54",
           838 => x"05",
           839 => x"05",
           840 => x"12",
           841 => x"08",
           842 => x"0c",
           843 => x"f0",
           844 => x"08",
           845 => x"08",
           846 => x"53",
           847 => x"2d",
           848 => x"38",
           849 => x"8c",
           850 => x"82",
           851 => x"82",
           852 => x"53",
           853 => x"08",
           854 => x"fc",
           855 => x"3d",
           856 => x"d5",
           857 => x"f9",
           858 => x"05",
           859 => x"70",
           860 => x"80",
           861 => x"f0",
           862 => x"82",
           863 => x"11",
           864 => x"51",
           865 => x"c5",
           866 => x"08",
           867 => x"53",
           868 => x"06",
           869 => x"d5",
           870 => x"08",
           871 => x"f0",
           872 => x"70",
           873 => x"51",
           874 => x"f0",
           875 => x"70",
           876 => x"51",
           877 => x"82",
           878 => x"08",
           879 => x"05",
           880 => x"fc",
           881 => x"08",
           882 => x"88",
           883 => x"70",
           884 => x"34",
           885 => x"05",
           886 => x"08",
           887 => x"71",
           888 => x"f0",
           889 => x"08",
           890 => x"51",
           891 => x"70",
           892 => x"52",
           893 => x"80",
           894 => x"08",
           895 => x"f4",
           896 => x"05",
           897 => x"08",
           898 => x"08",
           899 => x"06",
           900 => x"05",
           901 => x"f0",
           902 => x"d5",
           903 => x"52",
           904 => x"34",
           905 => x"52",
           906 => x"85",
           907 => x"08",
           908 => x"f0",
           909 => x"81",
           910 => x"08",
           911 => x"70",
           912 => x"51",
           913 => x"05",
           914 => x"0d",
           915 => x"f0",
           916 => x"3d",
           917 => x"08",
           918 => x"82",
           919 => x"d5",
           920 => x"f0",
           921 => x"a2",
           922 => x"08",
           923 => x"26",
           924 => x"f8",
           925 => x"05",
           926 => x"fc",
           927 => x"82",
           928 => x"d5",
           929 => x"d5",
           930 => x"f0",
           931 => x"08",
           932 => x"08",
           933 => x"90",
           934 => x"08",
           935 => x"90",
           936 => x"08",
           937 => x"90",
           938 => x"82",
           939 => x"05",
           940 => x"82",
           941 => x"05",
           942 => x"82",
           943 => x"d5",
           944 => x"71",
           945 => x"d5",
           946 => x"82",
           947 => x"d5",
           948 => x"82",
           949 => x"d5",
           950 => x"ba",
           951 => x"08",
           952 => x"f8",
           953 => x"08",
           954 => x"fc",
           955 => x"82",
           956 => x"05",
           957 => x"ff",
           958 => x"05",
           959 => x"85",
           960 => x"82",
           961 => x"0c",
           962 => x"88",
           963 => x"05",
           964 => x"08",
           965 => x"fc",
           966 => x"08",
           967 => x"51",
           968 => x"39",
           969 => x"ff",
           970 => x"0c",
           971 => x"82",
           972 => x"70",
           973 => x"0d",
           974 => x"f0",
           975 => x"3d",
           976 => x"08",
           977 => x"82",
           978 => x"71",
           979 => x"08",
           980 => x"05",
           981 => x"08",
           982 => x"f0",
           983 => x"d5",
           984 => x"ff",
           985 => x"ff",
           986 => x"05",
           987 => x"84",
           988 => x"82",
           989 => x"0c",
           990 => x"88",
           991 => x"05",
           992 => x"08",
           993 => x"82",
           994 => x"2e",
           995 => x"90",
           996 => x"08",
           997 => x"90",
           998 => x"08",
           999 => x"90",
          1000 => x"d5",
          1001 => x"33",
          1002 => x"81",
          1003 => x"0c",
          1004 => x"52",
          1005 => x"08",
          1006 => x"f0",
          1007 => x"82",
          1008 => x"82",
          1009 => x"82",
          1010 => x"08",
          1011 => x"0d",
          1012 => x"80",
          1013 => x"08",
          1014 => x"d5",
          1015 => x"82",
          1016 => x"d5",
          1017 => x"72",
          1018 => x"71",
          1019 => x"82",
          1020 => x"71",
          1021 => x"08",
          1022 => x"05",
          1023 => x"70",
          1024 => x"08",
          1025 => x"d5",
          1026 => x"82",
          1027 => x"d5",
          1028 => x"84",
          1029 => x"08",
          1030 => x"38",
          1031 => x"70",
          1032 => x"0b",
          1033 => x"80",
          1034 => x"05",
          1035 => x"8c",
          1036 => x"05",
          1037 => x"38",
          1038 => x"05",
          1039 => x"88",
          1040 => x"08",
          1041 => x"31",
          1042 => x"0c",
          1043 => x"80",
          1044 => x"0c",
          1045 => x"82",
          1046 => x"d5",
          1047 => x"02",
          1048 => x"82",
          1049 => x"82",
          1050 => x"81",
          1051 => x"82",
          1052 => x"d5",
          1053 => x"70",
          1054 => x"82",
          1055 => x"08",
          1056 => x"08",
          1057 => x"82",
          1058 => x"39",
          1059 => x"82",
          1060 => x"54",
          1061 => x"f8",
          1062 => x"88",
          1063 => x"fc",
          1064 => x"d5",
          1065 => x"f4",
          1066 => x"f4",
          1067 => x"3d",
          1068 => x"d5",
          1069 => x"fd",
          1070 => x"05",
          1071 => x"0c",
          1072 => x"8d",
          1073 => x"fc",
          1074 => x"f0",
          1075 => x"82",
          1076 => x"05",
          1077 => x"70",
          1078 => x"2e",
          1079 => x"05",
          1080 => x"8c",
          1081 => x"05",
          1082 => x"39",
          1083 => x"ff",
          1084 => x"0c",
          1085 => x"82",
          1086 => x"70",
          1087 => x"51",
          1088 => x"82",
          1089 => x"d5",
          1090 => x"02",
          1091 => x"82",
          1092 => x"d5",
          1093 => x"f0",
          1094 => x"d4",
          1095 => x"08",
          1096 => x"05",
          1097 => x"08",
          1098 => x"05",
          1099 => x"08",
          1100 => x"08",
          1101 => x"f0",
          1102 => x"71",
          1103 => x"08",
          1104 => x"05",
          1105 => x"08",
          1106 => x"0c",
          1107 => x"0c",
          1108 => x"d5",
          1109 => x"82",
          1110 => x"d5",
          1111 => x"b9",
          1112 => x"08",
          1113 => x"0c",
          1114 => x"05",
          1115 => x"08",
          1116 => x"08",
          1117 => x"f4",
          1118 => x"05",
          1119 => x"08",
          1120 => x"08",
          1121 => x"08",
          1122 => x"f0",
          1123 => x"08",
          1124 => x"82",
          1125 => x"d5",
          1126 => x"f0",
          1127 => x"d5",
          1128 => x"d5",
          1129 => x"c5",
          1130 => x"d5",
          1131 => x"d5",
          1132 => x"90",
          1133 => x"08",
          1134 => x"0c",
          1135 => x"70",
          1136 => x"0d",
          1137 => x"f0",
          1138 => x"3d",
          1139 => x"fc",
          1140 => x"05",
          1141 => x"f0",
          1142 => x"f0",
          1143 => x"d5",
          1144 => x"f0",
          1145 => x"38",
          1146 => x"30",
          1147 => x"81",
          1148 => x"08",
          1149 => x"08",
          1150 => x"08",
          1151 => x"0c",
          1152 => x"08",
          1153 => x"08",
          1154 => x"08",
          1155 => x"f8",
          1156 => x"54",
          1157 => x"04",
          1158 => x"f0",
          1159 => x"d5",
          1160 => x"d5",
          1161 => x"c5",
          1162 => x"d5",
          1163 => x"d5",
          1164 => x"02",
          1165 => x"81",
          1166 => x"08",
          1167 => x"08",
          1168 => x"70",
          1169 => x"0d",
          1170 => x"f0",
          1171 => x"3d",
          1172 => x"fc",
          1173 => x"08",
          1174 => x"8c",
          1175 => x"05",
          1176 => x"08",
          1177 => x"80",
          1178 => x"08",
          1179 => x"8c",
          1180 => x"8c",
          1181 => x"05",
          1182 => x"05",
          1183 => x"08",
          1184 => x"38",
          1185 => x"82",
          1186 => x"ad",
          1187 => x"08",
          1188 => x"31",
          1189 => x"82",
          1190 => x"d5",
          1191 => x"d5",
          1192 => x"f0",
          1193 => x"d5",
          1194 => x"f0",
          1195 => x"d5",
          1196 => x"39",
          1197 => x"80",
          1198 => x"88",
          1199 => x"f4",
          1200 => x"f0",
          1201 => x"f0",
          1202 => x"f0",
          1203 => x"0c",
          1204 => x"04",
          1205 => x"f0",
          1206 => x"d5",
          1207 => x"f0",
          1208 => x"0c",
          1209 => x"70",
          1210 => x"82",
          1211 => x"81",
          1212 => x"81",
          1213 => x"88",
          1214 => x"0c",
          1215 => x"f8",
          1216 => x"81",
          1217 => x"f0",
          1218 => x"08",
          1219 => x"71",
          1220 => x"82",
          1221 => x"d5",
          1222 => x"b0",
          1223 => x"82",
          1224 => x"08",
          1225 => x"53",
          1226 => x"05",
          1227 => x"33",
          1228 => x"82",
          1229 => x"e2",
          1230 => x"e8",
          1231 => x"80",
          1232 => x"08",
          1233 => x"88",
          1234 => x"0c",
          1235 => x"d5",
          1236 => x"39",
          1237 => x"05",
          1238 => x"08",
          1239 => x"08",
          1240 => x"08",
          1241 => x"d5",
          1242 => x"a0",
          1243 => x"f0",
          1244 => x"82",
          1245 => x"af",
          1246 => x"08",
          1247 => x"83",
          1248 => x"f0",
          1249 => x"88",
          1250 => x"34",
          1251 => x"05",
          1252 => x"82",
          1253 => x"72",
          1254 => x"0b",
          1255 => x"82",
          1256 => x"08",
          1257 => x"f0",
          1258 => x"08",
          1259 => x"81",
          1260 => x"05",
          1261 => x"38",
          1262 => x"e0",
          1263 => x"08",
          1264 => x"f8",
          1265 => x"82",
          1266 => x"d5",
          1267 => x"73",
          1268 => x"f8",
          1269 => x"82",
          1270 => x"d5",
          1271 => x"89",
          1272 => x"f0",
          1273 => x"82",
          1274 => x"d5",
          1275 => x"72",
          1276 => x"d5",
          1277 => x"39",
          1278 => x"70",
          1279 => x"29",
          1280 => x"70",
          1281 => x"0c",
          1282 => x"70",
          1283 => x"51",
          1284 => x"d5",
          1285 => x"39",
          1286 => x"53",
          1287 => x"f0",
          1288 => x"f0",
          1289 => x"08",
          1290 => x"fc",
          1291 => x"82",
          1292 => x"d5",
          1293 => x"e4",
          1294 => x"0c",
          1295 => x"d5",
          1296 => x"82",
          1297 => x"d5",
          1298 => x"73",
          1299 => x"08",
          1300 => x"72",
          1301 => x"72",
          1302 => x"09",
          1303 => x"08",
          1304 => x"71",
          1305 => x"08",
          1306 => x"09",
          1307 => x"d5",
          1308 => x"f0",
          1309 => x"05",
          1310 => x"33",
          1311 => x"82",
          1312 => x"72",
          1313 => x"38",
          1314 => x"70",
          1315 => x"51",
          1316 => x"f8",
          1317 => x"05",
          1318 => x"0c",
          1319 => x"80",
          1320 => x"08",
          1321 => x"38",
          1322 => x"f0",
          1323 => x"08",
          1324 => x"71",
          1325 => x"82",
          1326 => x"a4",
          1327 => x"f4",
          1328 => x"05",
          1329 => x"70",
          1330 => x"f0",
          1331 => x"82",
          1332 => x"72",
          1333 => x"d5",
          1334 => x"39",
          1335 => x"53",
          1336 => x"f0",
          1337 => x"26",
          1338 => x"d5",
          1339 => x"39",
          1340 => x"05",
          1341 => x"f8",
          1342 => x"38",
          1343 => x"53",
          1344 => x"80",
          1345 => x"0c",
          1346 => x"f0",
          1347 => x"d5",
          1348 => x"f0",
          1349 => x"27",
          1350 => x"f8",
          1351 => x"94",
          1352 => x"33",
          1353 => x"f0",
          1354 => x"08",
          1355 => x"72",
          1356 => x"82",
          1357 => x"90",
          1358 => x"08",
          1359 => x"72",
          1360 => x"82",
          1361 => x"72",
          1362 => x"d5",
          1363 => x"39",
          1364 => x"82",
          1365 => x"54",
          1366 => x"82",
          1367 => x"f7",
          1368 => x"33",
          1369 => x"08",
          1370 => x"33",
          1371 => x"05",
          1372 => x"08",
          1373 => x"08",
          1374 => x"82",
          1375 => x"a5",
          1376 => x"33",
          1377 => x"d5",
          1378 => x"d5",
          1379 => x"f0",
          1380 => x"08",
          1381 => x"0b",
          1382 => x"82",
          1383 => x"d5",
          1384 => x"f0",
          1385 => x"08",
          1386 => x"80",
          1387 => x"0c",
          1388 => x"74",
          1389 => x"06",
          1390 => x"80",
          1391 => x"05",
          1392 => x"82",
          1393 => x"54",
          1394 => x"fc",
          1395 => x"84",
          1396 => x"b4",
          1397 => x"58",
          1398 => x"54",
          1399 => x"0d",
          1400 => x"93",
          1401 => x"82",
          1402 => x"82",
          1403 => x"b3",
          1404 => x"b8",
          1405 => x"51",
          1406 => x"80",
          1407 => x"dd",
          1408 => x"39",
          1409 => x"82",
          1410 => x"b4",
          1411 => x"d4",
          1412 => x"b5",
          1413 => x"82",
          1414 => x"bc",
          1415 => x"9d",
          1416 => x"82",
          1417 => x"9c",
          1418 => x"85",
          1419 => x"3f",
          1420 => x"77",
          1421 => x"8a",
          1422 => x"51",
          1423 => x"ef",
          1424 => x"75",
          1425 => x"08",
          1426 => x"d0",
          1427 => x"0d",
          1428 => x"05",
          1429 => x"68",
          1430 => x"51",
          1431 => x"ff",
          1432 => x"07",
          1433 => x"56",
          1434 => x"52",
          1435 => x"f9",
          1436 => x"d5",
          1437 => x"08",
          1438 => x"e4",
          1439 => x"84",
          1440 => x"96",
          1441 => x"82",
          1442 => x"74",
          1443 => x"19",
          1444 => x"05",
          1445 => x"70",
          1446 => x"9f",
          1447 => x"74",
          1448 => x"53",
          1449 => x"51",
          1450 => x"d5",
          1451 => x"3d",
          1452 => x"33",
          1453 => x"52",
          1454 => x"e4",
          1455 => x"38",
          1456 => x"82",
          1457 => x"82",
          1458 => x"78",
          1459 => x"39",
          1460 => x"8a",
          1461 => x"61",
          1462 => x"33",
          1463 => x"5c",
          1464 => x"fc",
          1465 => x"84",
          1466 => x"74",
          1467 => x"2e",
          1468 => x"80",
          1469 => x"27",
          1470 => x"88",
          1471 => x"82",
          1472 => x"82",
          1473 => x"53",
          1474 => x"52",
          1475 => x"3f",
          1476 => x"b7",
          1477 => x"74",
          1478 => x"72",
          1479 => x"b7",
          1480 => x"51",
          1481 => x"82",
          1482 => x"dc",
          1483 => x"51",
          1484 => x"79",
          1485 => x"33",
          1486 => x"83",
          1487 => x"27",
          1488 => x"70",
          1489 => x"2e",
          1490 => x"38",
          1491 => x"88",
          1492 => x"51",
          1493 => x"b6",
          1494 => x"3f",
          1495 => x"8a",
          1496 => x"70",
          1497 => x"09",
          1498 => x"82",
          1499 => x"2c",
          1500 => x"32",
          1501 => x"07",
          1502 => x"57",
          1503 => x"2e",
          1504 => x"8c",
          1505 => x"fd",
          1506 => x"e4",
          1507 => x"0d",
          1508 => x"53",
          1509 => x"aa",
          1510 => x"e3",
          1511 => x"cc",
          1512 => x"b7",
          1513 => x"80",
          1514 => x"3d",
          1515 => x"96",
          1516 => x"51",
          1517 => x"99",
          1518 => x"72",
          1519 => x"71",
          1520 => x"af",
          1521 => x"3f",
          1522 => x"2a",
          1523 => x"2e",
          1524 => x"82",
          1525 => x"51",
          1526 => x"81",
          1527 => x"38",
          1528 => x"a8",
          1529 => x"e7",
          1530 => x"51",
          1531 => x"51",
          1532 => x"98",
          1533 => x"72",
          1534 => x"71",
          1535 => x"b7",
          1536 => x"3f",
          1537 => x"2a",
          1538 => x"2e",
          1539 => x"82",
          1540 => x"51",
          1541 => x"81",
          1542 => x"38",
          1543 => x"f8",
          1544 => x"ef",
          1545 => x"51",
          1546 => x"51",
          1547 => x"97",
          1548 => x"a4",
          1549 => x"3d",
          1550 => x"33",
          1551 => x"51",
          1552 => x"d8",
          1553 => x"82",
          1554 => x"81",
          1555 => x"30",
          1556 => x"25",
          1557 => x"0b",
          1558 => x"82",
          1559 => x"09",
          1560 => x"53",
          1561 => x"3f",
          1562 => x"38",
          1563 => x"3f",
          1564 => x"96",
          1565 => x"d0",
          1566 => x"33",
          1567 => x"8c",
          1568 => x"75",
          1569 => x"d5",
          1570 => x"3d",
          1571 => x"82",
          1572 => x"51",
          1573 => x"08",
          1574 => x"09",
          1575 => x"83",
          1576 => x"db",
          1577 => x"d7",
          1578 => x"d5",
          1579 => x"b9",
          1580 => x"41",
          1581 => x"ea",
          1582 => x"f8",
          1583 => x"3d",
          1584 => x"82",
          1585 => x"2c",
          1586 => x"a3",
          1587 => x"78",
          1588 => x"24",
          1589 => x"38",
          1590 => x"d6",
          1591 => x"38",
          1592 => x"78",
          1593 => x"39",
          1594 => x"78",
          1595 => x"c3",
          1596 => x"2e",
          1597 => x"81",
          1598 => x"83",
          1599 => x"89",
          1600 => x"85",
          1601 => x"b5",
          1602 => x"05",
          1603 => x"08",
          1604 => x"fe",
          1605 => x"ec",
          1606 => x"2e",
          1607 => x"11",
          1608 => x"3f",
          1609 => x"d5",
          1610 => x"ff",
          1611 => x"79",
          1612 => x"78",
          1613 => x"7a",
          1614 => x"3d",
          1615 => x"51",
          1616 => x"80",
          1617 => x"fc",
          1618 => x"e1",
          1619 => x"fd",
          1620 => x"53",
          1621 => x"82",
          1622 => x"38",
          1623 => x"3f",
          1624 => x"38",
          1625 => x"33",
          1626 => x"39",
          1627 => x"84",
          1628 => x"e4",
          1629 => x"3d",
          1630 => x"51",
          1631 => x"80",
          1632 => x"f8",
          1633 => x"e9",
          1634 => x"fc",
          1635 => x"ad",
          1636 => x"a8",
          1637 => x"5a",
          1638 => x"55",
          1639 => x"82",
          1640 => x"81",
          1641 => x"39",
          1642 => x"39",
          1643 => x"84",
          1644 => x"e4",
          1645 => x"33",
          1646 => x"d4",
          1647 => x"d4",
          1648 => x"38",
          1649 => x"82",
          1650 => x"88",
          1651 => x"39",
          1652 => x"2e",
          1653 => x"9a",
          1654 => x"80",
          1655 => x"45",
          1656 => x"80",
          1657 => x"53",
          1658 => x"82",
          1659 => x"d4",
          1660 => x"38",
          1661 => x"39",
          1662 => x"2e",
          1663 => x"bb",
          1664 => x"80",
          1665 => x"44",
          1666 => x"78",
          1667 => x"08",
          1668 => x"59",
          1669 => x"a4",
          1670 => x"08",
          1671 => x"11",
          1672 => x"3f",
          1673 => x"38",
          1674 => x"83",
          1675 => x"30",
          1676 => x"06",
          1677 => x"88",
          1678 => x"43",
          1679 => x"a0",
          1680 => x"64",
          1681 => x"51",
          1682 => x"11",
          1683 => x"3f",
          1684 => x"c1",
          1685 => x"ff",
          1686 => x"d5",
          1687 => x"59",
          1688 => x"64",
          1689 => x"11",
          1690 => x"3f",
          1691 => x"89",
          1692 => x"bb",
          1693 => x"f1",
          1694 => x"51",
          1695 => x"33",
          1696 => x"9f",
          1697 => x"fc",
          1698 => x"e1",
          1699 => x"91",
          1700 => x"33",
          1701 => x"b1",
          1702 => x"3f",
          1703 => x"11",
          1704 => x"3f",
          1705 => x"99",
          1706 => x"ff",
          1707 => x"d5",
          1708 => x"59",
          1709 => x"82",
          1710 => x"fe",
          1711 => x"e0",
          1712 => x"38",
          1713 => x"52",
          1714 => x"3f",
          1715 => x"52",
          1716 => x"46",
          1717 => x"b9",
          1718 => x"82",
          1719 => x"f0",
          1720 => x"e0",
          1721 => x"93",
          1722 => x"22",
          1723 => x"42",
          1724 => x"c3",
          1725 => x"fe",
          1726 => x"df",
          1727 => x"2e",
          1728 => x"11",
          1729 => x"3f",
          1730 => x"38",
          1731 => x"05",
          1732 => x"ff",
          1733 => x"d5",
          1734 => x"61",
          1735 => x"51",
          1736 => x"08",
          1737 => x"a7",
          1738 => x"78",
          1739 => x"27",
          1740 => x"53",
          1741 => x"82",
          1742 => x"61",
          1743 => x"42",
          1744 => x"c2",
          1745 => x"ff",
          1746 => x"e3",
          1747 => x"2e",
          1748 => x"b0",
          1749 => x"78",
          1750 => x"ff",
          1751 => x"d5",
          1752 => x"64",
          1753 => x"8a",
          1754 => x"e4",
          1755 => x"d5",
          1756 => x"ff",
          1757 => x"bc",
          1758 => x"c3",
          1759 => x"51",
          1760 => x"39",
          1761 => x"3d",
          1762 => x"38",
          1763 => x"3f",
          1764 => x"e4",
          1765 => x"d5",
          1766 => x"05",
          1767 => x"08",
          1768 => x"2e",
          1769 => x"51",
          1770 => x"8f",
          1771 => x"82",
          1772 => x"38",
          1773 => x"39",
          1774 => x"39",
          1775 => x"bc",
          1776 => x"52",
          1777 => x"a7",
          1778 => x"3d",
          1779 => x"ab",
          1780 => x"80",
          1781 => x"ff",
          1782 => x"93",
          1783 => x"d8",
          1784 => x"ff",
          1785 => x"82",
          1786 => x"80",
          1787 => x"80",
          1788 => x"ea",
          1789 => x"d5",
          1790 => x"07",
          1791 => x"5a",
          1792 => x"78",
          1793 => x"38",
          1794 => x"59",
          1795 => x"7e",
          1796 => x"7e",
          1797 => x"82",
          1798 => x"7c",
          1799 => x"82",
          1800 => x"f2",
          1801 => x"82",
          1802 => x"70",
          1803 => x"72",
          1804 => x"08",
          1805 => x"84",
          1806 => x"72",
          1807 => x"87",
          1808 => x"87",
          1809 => x"3f",
          1810 => x"08",
          1811 => x"51",
          1812 => x"08",
          1813 => x"87",
          1814 => x"0b",
          1815 => x"cd",
          1816 => x"84",
          1817 => x"f1",
          1818 => x"0c",
          1819 => x"54",
          1820 => x"bd",
          1821 => x"bd",
          1822 => x"de",
          1823 => x"ec",
          1824 => x"fe",
          1825 => x"88",
          1826 => x"e4",
          1827 => x"14",
          1828 => x"71",
          1829 => x"04",
          1830 => x"55",
          1831 => x"81",
          1832 => x"2e",
          1833 => x"53",
          1834 => x"2e",
          1835 => x"53",
          1836 => x"09",
          1837 => x"12",
          1838 => x"a2",
          1839 => x"2e",
          1840 => x"81",
          1841 => x"70",
          1842 => x"80",
          1843 => x"72",
          1844 => x"81",
          1845 => x"32",
          1846 => x"51",
          1847 => x"80",
          1848 => x"75",
          1849 => x"0c",
          1850 => x"76",
          1851 => x"86",
          1852 => x"c0",
          1853 => x"80",
          1854 => x"d5",
          1855 => x"3d",
          1856 => x"52",
          1857 => x"98",
          1858 => x"82",
          1859 => x"84",
          1860 => x"26",
          1861 => x"84",
          1862 => x"86",
          1863 => x"26",
          1864 => x"86",
          1865 => x"38",
          1866 => x"87",
          1867 => x"87",
          1868 => x"c0",
          1869 => x"c0",
          1870 => x"c0",
          1871 => x"c0",
          1872 => x"c0",
          1873 => x"c0",
          1874 => x"a4",
          1875 => x"80",
          1876 => x"52",
          1877 => x"0d",
          1878 => x"c0",
          1879 => x"c0",
          1880 => x"87",
          1881 => x"1c",
          1882 => x"79",
          1883 => x"08",
          1884 => x"98",
          1885 => x"87",
          1886 => x"1c",
          1887 => x"7b",
          1888 => x"08",
          1889 => x"0c",
          1890 => x"83",
          1891 => x"57",
          1892 => x"55",
          1893 => x"53",
          1894 => x"bd",
          1895 => x"3d",
          1896 => x"05",
          1897 => x"ff",
          1898 => x"84",
          1899 => x"c0",
          1900 => x"2a",
          1901 => x"80",
          1902 => x"81",
          1903 => x"81",
          1904 => x"80",
          1905 => x"81",
          1906 => x"73",
          1907 => x"80",
          1908 => x"c0",
          1909 => x"82",
          1910 => x"ff",
          1911 => x"30",
          1912 => x"82",
          1913 => x"f9",
          1914 => x"77",
          1915 => x"7a",
          1916 => x"fc",
          1917 => x"87",
          1918 => x"86",
          1919 => x"08",
          1920 => x"56",
          1921 => x"91",
          1922 => x"d7",
          1923 => x"51",
          1924 => x"93",
          1925 => x"ff",
          1926 => x"87",
          1927 => x"86",
          1928 => x"74",
          1929 => x"89",
          1930 => x"54",
          1931 => x"53",
          1932 => x"38",
          1933 => x"d3",
          1934 => x"57",
          1935 => x"75",
          1936 => x"94",
          1937 => x"81",
          1938 => x"8c",
          1939 => x"51",
          1940 => x"70",
          1941 => x"8d",
          1942 => x"51",
          1943 => x"ff",
          1944 => x"70",
          1945 => x"90",
          1946 => x"33",
          1947 => x"70",
          1948 => x"0c",
          1949 => x"82",
          1950 => x"54",
          1951 => x"80",
          1952 => x"51",
          1953 => x"06",
          1954 => x"38",
          1955 => x"94",
          1956 => x"87",
          1957 => x"81",
          1958 => x"84",
          1959 => x"d5",
          1960 => x"e4",
          1961 => x"fc",
          1962 => x"87",
          1963 => x"86",
          1964 => x"08",
          1965 => x"51",
          1966 => x"38",
          1967 => x"94",
          1968 => x"87",
          1969 => x"98",
          1970 => x"71",
          1971 => x"04",
          1972 => x"08",
          1973 => x"70",
          1974 => x"9e",
          1975 => x"c0",
          1976 => x"87",
          1977 => x"0c",
          1978 => x"8c",
          1979 => x"d4",
          1980 => x"82",
          1981 => x"08",
          1982 => x"b0",
          1983 => x"9e",
          1984 => x"c0",
          1985 => x"87",
          1986 => x"0c",
          1987 => x"ac",
          1988 => x"d4",
          1989 => x"51",
          1990 => x"9e",
          1991 => x"c0",
          1992 => x"87",
          1993 => x"0c",
          1994 => x"0b",
          1995 => x"80",
          1996 => x"2e",
          1997 => x"c5",
          1998 => x"08",
          1999 => x"52",
          2000 => x"71",
          2001 => x"c0",
          2002 => x"06",
          2003 => x"38",
          2004 => x"80",
          2005 => x"88",
          2006 => x"80",
          2007 => x"d4",
          2008 => x"90",
          2009 => x"52",
          2010 => x"52",
          2011 => x"87",
          2012 => x"80",
          2013 => x"83",
          2014 => x"34",
          2015 => x"70",
          2016 => x"70",
          2017 => x"82",
          2018 => x"9e",
          2019 => x"51",
          2020 => x"81",
          2021 => x"0b",
          2022 => x"80",
          2023 => x"2e",
          2024 => x"cd",
          2025 => x"08",
          2026 => x"52",
          2027 => x"71",
          2028 => x"c0",
          2029 => x"51",
          2030 => x"81",
          2031 => x"c0",
          2032 => x"70",
          2033 => x"d4",
          2034 => x"90",
          2035 => x"52",
          2036 => x"71",
          2037 => x"90",
          2038 => x"2a",
          2039 => x"34",
          2040 => x"70",
          2041 => x"2e",
          2042 => x"d3",
          2043 => x"87",
          2044 => x"34",
          2045 => x"82",
          2046 => x"82",
          2047 => x"89",
          2048 => x"d2",
          2049 => x"d5",
          2050 => x"80",
          2051 => x"82",
          2052 => x"be",
          2053 => x"d4",
          2054 => x"38",
          2055 => x"08",
          2056 => x"ff",
          2057 => x"54",
          2058 => x"80",
          2059 => x"52",
          2060 => x"3f",
          2061 => x"2e",
          2062 => x"d4",
          2063 => x"ec",
          2064 => x"ca",
          2065 => x"82",
          2066 => x"11",
          2067 => x"92",
          2068 => x"73",
          2069 => x"33",
          2070 => x"a2",
          2071 => x"80",
          2072 => x"52",
          2073 => x"3f",
          2074 => x"2e",
          2075 => x"82",
          2076 => x"82",
          2077 => x"89",
          2078 => x"ed",
          2079 => x"80",
          2080 => x"ff",
          2081 => x"54",
          2082 => x"a4",
          2083 => x"cd",
          2084 => x"82",
          2085 => x"82",
          2086 => x"89",
          2087 => x"a5",
          2088 => x"9d",
          2089 => x"c0",
          2090 => x"d4",
          2091 => x"ff",
          2092 => x"52",
          2093 => x"3f",
          2094 => x"3f",
          2095 => x"cc",
          2096 => x"b8",
          2097 => x"51",
          2098 => x"bd",
          2099 => x"54",
          2100 => x"f4",
          2101 => x"cb",
          2102 => x"82",
          2103 => x"52",
          2104 => x"e4",
          2105 => x"31",
          2106 => x"82",
          2107 => x"82",
          2108 => x"a9",
          2109 => x"84",
          2110 => x"82",
          2111 => x"76",
          2112 => x"08",
          2113 => x"ca",
          2114 => x"87",
          2115 => x"92",
          2116 => x"26",
          2117 => x"fc",
          2118 => x"f8",
          2119 => x"97",
          2120 => x"82",
          2121 => x"94",
          2122 => x"ff",
          2123 => x"71",
          2124 => x"c0",
          2125 => x"08",
          2126 => x"3d",
          2127 => x"79",
          2128 => x"13",
          2129 => x"51",
          2130 => x"33",
          2131 => x"82",
          2132 => x"05",
          2133 => x"52",
          2134 => x"38",
          2135 => x"85",
          2136 => x"02",
          2137 => x"55",
          2138 => x"82",
          2139 => x"ad",
          2140 => x"a0",
          2141 => x"c8",
          2142 => x"3f",
          2143 => x"34",
          2144 => x"77",
          2145 => x"34",
          2146 => x"7c",
          2147 => x"88",
          2148 => x"33",
          2149 => x"70",
          2150 => x"74",
          2151 => x"fb",
          2152 => x"29",
          2153 => x"54",
          2154 => x"d5",
          2155 => x"33",
          2156 => x"70",
          2157 => x"a7",
          2158 => x"ff",
          2159 => x"81",
          2160 => x"74",
          2161 => x"87",
          2162 => x"77",
          2163 => x"08",
          2164 => x"d5",
          2165 => x"3d",
          2166 => x"75",
          2167 => x"b0",
          2168 => x"3f",
          2169 => x"e6",
          2170 => x"0d",
          2171 => x"08",
          2172 => x"51",
          2173 => x"14",
          2174 => x"e6",
          2175 => x"82",
          2176 => x"95",
          2177 => x"82",
          2178 => x"80",
          2179 => x"0d",
          2180 => x"52",
          2181 => x"e7",
          2182 => x"38",
          2183 => x"52",
          2184 => x"bf",
          2185 => x"ba",
          2186 => x"82",
          2187 => x"d5",
          2188 => x"e4",
          2189 => x"80",
          2190 => x"17",
          2191 => x"da",
          2192 => x"ff",
          2193 => x"3d",
          2194 => x"5a",
          2195 => x"82",
          2196 => x"3f",
          2197 => x"ff",
          2198 => x"80",
          2199 => x"81",
          2200 => x"80",
          2201 => x"b7",
          2202 => x"58",
          2203 => x"25",
          2204 => x"05",
          2205 => x"74",
          2206 => x"2a",
          2207 => x"38",
          2208 => x"08",
          2209 => x"87",
          2210 => x"89",
          2211 => x"ba",
          2212 => x"9b",
          2213 => x"c5",
          2214 => x"ab",
          2215 => x"74",
          2216 => x"0c",
          2217 => x"7c",
          2218 => x"59",
          2219 => x"06",
          2220 => x"77",
          2221 => x"5b",
          2222 => x"a0",
          2223 => x"75",
          2224 => x"29",
          2225 => x"55",
          2226 => x"08",
          2227 => x"b3",
          2228 => x"c5",
          2229 => x"2e",
          2230 => x"b5",
          2231 => x"1a",
          2232 => x"05",
          2233 => x"08",
          2234 => x"78",
          2235 => x"d5",
          2236 => x"85",
          2237 => x"70",
          2238 => x"27",
          2239 => x"d5",
          2240 => x"3d",
          2241 => x"b4",
          2242 => x"af",
          2243 => x"d5",
          2244 => x"38",
          2245 => x"73",
          2246 => x"81",
          2247 => x"56",
          2248 => x"51",
          2249 => x"82",
          2250 => x"80",
          2251 => x"52",
          2252 => x"f1",
          2253 => x"8c",
          2254 => x"ed",
          2255 => x"08",
          2256 => x"f8",
          2257 => x"9a",
          2258 => x"82",
          2259 => x"06",
          2260 => x"51",
          2261 => x"08",
          2262 => x"25",
          2263 => x"05",
          2264 => x"80",
          2265 => x"51",
          2266 => x"ff",
          2267 => x"38",
          2268 => x"06",
          2269 => x"d5",
          2270 => x"b0",
          2271 => x"3f",
          2272 => x"d5",
          2273 => x"51",
          2274 => x"81",
          2275 => x"98",
          2276 => x"33",
          2277 => x"98",
          2278 => x"a4",
          2279 => x"51",
          2280 => x"58",
          2281 => x"38",
          2282 => x"80",
          2283 => x"98",
          2284 => x"ce",
          2285 => x"f6",
          2286 => x"ff",
          2287 => x"74",
          2288 => x"39",
          2289 => x"0a",
          2290 => x"06",
          2291 => x"38",
          2292 => x"ce",
          2293 => x"06",
          2294 => x"56",
          2295 => x"1c",
          2296 => x"98",
          2297 => x"33",
          2298 => x"10",
          2299 => x"11",
          2300 => x"51",
          2301 => x"fe",
          2302 => x"7d",
          2303 => x"80",
          2304 => x"75",
          2305 => x"9c",
          2306 => x"0c",
          2307 => x"38",
          2308 => x"54",
          2309 => x"54",
          2310 => x"ed",
          2311 => x"38",
          2312 => x"55",
          2313 => x"54",
          2314 => x"80",
          2315 => x"98",
          2316 => x"55",
          2317 => x"11",
          2318 => x"73",
          2319 => x"82",
          2320 => x"89",
          2321 => x"a4",
          2322 => x"80",
          2323 => x"98",
          2324 => x"56",
          2325 => x"f1",
          2326 => x"52",
          2327 => x"80",
          2328 => x"98",
          2329 => x"55",
          2330 => x"a8",
          2331 => x"82",
          2332 => x"74",
          2333 => x"c8",
          2334 => x"3f",
          2335 => x"0a",
          2336 => x"33",
          2337 => x"38",
          2338 => x"0b",
          2339 => x"80",
          2340 => x"3f",
          2341 => x"70",
          2342 => x"2e",
          2343 => x"ff",
          2344 => x"ff",
          2345 => x"82",
          2346 => x"a0",
          2347 => x"98",
          2348 => x"33",
          2349 => x"ad",
          2350 => x"74",
          2351 => x"33",
          2352 => x"80",
          2353 => x"98",
          2354 => x"55",
          2355 => x"c8",
          2356 => x"3f",
          2357 => x"70",
          2358 => x"51",
          2359 => x"38",
          2360 => x"ff",
          2361 => x"29",
          2362 => x"82",
          2363 => x"75",
          2364 => x"ed",
          2365 => x"34",
          2366 => x"ff",
          2367 => x"79",
          2368 => x"08",
          2369 => x"82",
          2370 => x"8f",
          2371 => x"f1",
          2372 => x"80",
          2373 => x"82",
          2374 => x"0c",
          2375 => x"33",
          2376 => x"82",
          2377 => x"9e",
          2378 => x"05",
          2379 => x"81",
          2380 => x"a8",
          2381 => x"73",
          2382 => x"54",
          2383 => x"2b",
          2384 => x"56",
          2385 => x"74",
          2386 => x"82",
          2387 => x"ff",
          2388 => x"29",
          2389 => x"82",
          2390 => x"75",
          2391 => x"52",
          2392 => x"ed",
          2393 => x"2c",
          2394 => x"57",
          2395 => x"f1",
          2396 => x"cc",
          2397 => x"80",
          2398 => x"a4",
          2399 => x"de",
          2400 => x"33",
          2401 => x"33",
          2402 => x"e8",
          2403 => x"14",
          2404 => x"1a",
          2405 => x"3f",
          2406 => x"06",
          2407 => x"75",
          2408 => x"82",
          2409 => x"f0",
          2410 => x"ed",
          2411 => x"34",
          2412 => x"d5",
          2413 => x"38",
          2414 => x"d5",
          2415 => x"d5",
          2416 => x"53",
          2417 => x"3f",
          2418 => x"29",
          2419 => x"56",
          2420 => x"51",
          2421 => x"08",
          2422 => x"08",
          2423 => x"52",
          2424 => x"1b",
          2425 => x"74",
          2426 => x"ff",
          2427 => x"2e",
          2428 => x"dc",
          2429 => x"74",
          2430 => x"e4",
          2431 => x"e4",
          2432 => x"74",
          2433 => x"80",
          2434 => x"e0",
          2435 => x"2e",
          2436 => x"3f",
          2437 => x"34",
          2438 => x"81",
          2439 => x"a5",
          2440 => x"ff",
          2441 => x"a4",
          2442 => x"53",
          2443 => x"ec",
          2444 => x"a8",
          2445 => x"a4",
          2446 => x"f5",
          2447 => x"81",
          2448 => x"74",
          2449 => x"a4",
          2450 => x"33",
          2451 => x"82",
          2452 => x"9a",
          2453 => x"05",
          2454 => x"c8",
          2455 => x"0b",
          2456 => x"82",
          2457 => x"80",
          2458 => x"bb",
          2459 => x"58",
          2460 => x"15",
          2461 => x"84",
          2462 => x"d5",
          2463 => x"76",
          2464 => x"82",
          2465 => x"80",
          2466 => x"88",
          2467 => x"17",
          2468 => x"d0",
          2469 => x"08",
          2470 => x"82",
          2471 => x"3d",
          2472 => x"81",
          2473 => x"12",
          2474 => x"ff",
          2475 => x"e4",
          2476 => x"0d",
          2477 => x"aa",
          2478 => x"08",
          2479 => x"2b",
          2480 => x"71",
          2481 => x"05",
          2482 => x"70",
          2483 => x"5b",
          2484 => x"34",
          2485 => x"08",
          2486 => x"82",
          2487 => x"d5",
          2488 => x"12",
          2489 => x"2b",
          2490 => x"52",
          2491 => x"70",
          2492 => x"12",
          2493 => x"83",
          2494 => x"56",
          2495 => x"89",
          2496 => x"d5",
          2497 => x"22",
          2498 => x"33",
          2499 => x"83",
          2500 => x"52",
          2501 => x"33",
          2502 => x"54",
          2503 => x"73",
          2504 => x"70",
          2505 => x"71",
          2506 => x"59",
          2507 => x"87",
          2508 => x"88",
          2509 => x"13",
          2510 => x"d4",
          2511 => x"71",
          2512 => x"06",
          2513 => x"53",
          2514 => x"87",
          2515 => x"a2",
          2516 => x"83",
          2517 => x"33",
          2518 => x"15",
          2519 => x"2b",
          2520 => x"55",
          2521 => x"80",
          2522 => x"ab",
          2523 => x"70",
          2524 => x"71",
          2525 => x"81",
          2526 => x"83",
          2527 => x"54",
          2528 => x"74",
          2529 => x"34",
          2530 => x"08",
          2531 => x"71",
          2532 => x"59",
          2533 => x"12",
          2534 => x"ff",
          2535 => x"52",
          2536 => x"15",
          2537 => x"0d",
          2538 => x"9e",
          2539 => x"82",
          2540 => x"2b",
          2541 => x"52",
          2542 => x"13",
          2543 => x"05",
          2544 => x"2a",
          2545 => x"34",
          2546 => x"08",
          2547 => x"71",
          2548 => x"59",
          2549 => x"83",
          2550 => x"88",
          2551 => x"13",
          2552 => x"d4",
          2553 => x"33",
          2554 => x"0c",
          2555 => x"3d",
          2556 => x"83",
          2557 => x"53",
          2558 => x"d4",
          2559 => x"11",
          2560 => x"71",
          2561 => x"81",
          2562 => x"2b",
          2563 => x"58",
          2564 => x"38",
          2565 => x"9d",
          2566 => x"85",
          2567 => x"2b",
          2568 => x"51",
          2569 => x"75",
          2570 => x"34",
          2571 => x"12",
          2572 => x"07",
          2573 => x"53",
          2574 => x"34",
          2575 => x"0b",
          2576 => x"34",
          2577 => x"14",
          2578 => x"d4",
          2579 => x"71",
          2580 => x"07",
          2581 => x"54",
          2582 => x"8b",
          2583 => x"52",
          2584 => x"f1",
          2585 => x"51",
          2586 => x"f5",
          2587 => x"e2",
          2588 => x"ff",
          2589 => x"33",
          2590 => x"70",
          2591 => x"ff",
          2592 => x"75",
          2593 => x"33",
          2594 => x"ff",
          2595 => x"06",
          2596 => x"59",
          2597 => x"80",
          2598 => x"84",
          2599 => x"2b",
          2600 => x"81",
          2601 => x"59",
          2602 => x"d4",
          2603 => x"71",
          2604 => x"06",
          2605 => x"75",
          2606 => x"79",
          2607 => x"74",
          2608 => x"2e",
          2609 => x"f8",
          2610 => x"80",
          2611 => x"3f",
          2612 => x"11",
          2613 => x"71",
          2614 => x"74",
          2615 => x"06",
          2616 => x"78",
          2617 => x"57",
          2618 => x"08",
          2619 => x"86",
          2620 => x"2b",
          2621 => x"53",
          2622 => x"75",
          2623 => x"70",
          2624 => x"71",
          2625 => x"5d",
          2626 => x"15",
          2627 => x"d4",
          2628 => x"33",
          2629 => x"70",
          2630 => x"54",
          2631 => x"34",
          2632 => x"54",
          2633 => x"0d",
          2634 => x"d5",
          2635 => x"71",
          2636 => x"51",
          2637 => x"53",
          2638 => x"0d",
          2639 => x"5c",
          2640 => x"08",
          2641 => x"f4",
          2642 => x"ff",
          2643 => x"83",
          2644 => x"fc",
          2645 => x"7e",
          2646 => x"08",
          2647 => x"08",
          2648 => x"ff",
          2649 => x"70",
          2650 => x"07",
          2651 => x"06",
          2652 => x"29",
          2653 => x"88",
          2654 => x"4e",
          2655 => x"41",
          2656 => x"8f",
          2657 => x"31",
          2658 => x"82",
          2659 => x"2b",
          2660 => x"81",
          2661 => x"2b",
          2662 => x"73",
          2663 => x"70",
          2664 => x"7b",
          2665 => x"73",
          2666 => x"78",
          2667 => x"ff",
          2668 => x"38",
          2669 => x"f6",
          2670 => x"55",
          2671 => x"1d",
          2672 => x"88",
          2673 => x"3f",
          2674 => x"82",
          2675 => x"7e",
          2676 => x"d5",
          2677 => x"59",
          2678 => x"08",
          2679 => x"06",
          2680 => x"54",
          2681 => x"51",
          2682 => x"1d",
          2683 => x"88",
          2684 => x"3f",
          2685 => x"82",
          2686 => x"7e",
          2687 => x"d5",
          2688 => x"59",
          2689 => x"08",
          2690 => x"55",
          2691 => x"a9",
          2692 => x"3f",
          2693 => x"e4",
          2694 => x"73",
          2695 => x"95",
          2696 => x"7a",
          2697 => x"53",
          2698 => x"7a",
          2699 => x"05",
          2700 => x"54",
          2701 => x"0d",
          2702 => x"70",
          2703 => x"e4",
          2704 => x"2e",
          2705 => x"d5",
          2706 => x"74",
          2707 => x"04",
          2708 => x"51",
          2709 => x"82",
          2710 => x"d5",
          2711 => x"3d",
          2712 => x"05",
          2713 => x"72",
          2714 => x"2b",
          2715 => x"88",
          2716 => x"88",
          2717 => x"8c",
          2718 => x"87",
          2719 => x"08",
          2720 => x"2e",
          2721 => x"51",
          2722 => x"80",
          2723 => x"98",
          2724 => x"38",
          2725 => x"d5",
          2726 => x"e4",
          2727 => x"0d",
          2728 => x"05",
          2729 => x"52",
          2730 => x"08",
          2731 => x"be",
          2732 => x"c0",
          2733 => x"12",
          2734 => x"40",
          2735 => x"98",
          2736 => x"0c",
          2737 => x"06",
          2738 => x"38",
          2739 => x"05",
          2740 => x"a2",
          2741 => x"38",
          2742 => x"38",
          2743 => x"98",
          2744 => x"c0",
          2745 => x"87",
          2746 => x"81",
          2747 => x"53",
          2748 => x"71",
          2749 => x"84",
          2750 => x"06",
          2751 => x"38",
          2752 => x"87",
          2753 => x"73",
          2754 => x"2e",
          2755 => x"82",
          2756 => x"f3",
          2757 => x"05",
          2758 => x"83",
          2759 => x"3f",
          2760 => x"54",
          2761 => x"81",
          2762 => x"c0",
          2763 => x"12",
          2764 => x"5f",
          2765 => x"8c",
          2766 => x"80",
          2767 => x"81",
          2768 => x"8c",
          2769 => x"7c",
          2770 => x"70",
          2771 => x"8a",
          2772 => x"71",
          2773 => x"52",
          2774 => x"80",
          2775 => x"c0",
          2776 => x"82",
          2777 => x"19",
          2778 => x"ff",
          2779 => x"78",
          2780 => x"80",
          2781 => x"26",
          2782 => x"06",
          2783 => x"52",
          2784 => x"8f",
          2785 => x"02",
          2786 => x"05",
          2787 => x"57",
          2788 => x"81",
          2789 => x"38",
          2790 => x"81",
          2791 => x"71",
          2792 => x"87",
          2793 => x"80",
          2794 => x"83",
          2795 => x"72",
          2796 => x"51",
          2797 => x"87",
          2798 => x"38",
          2799 => x"96",
          2800 => x"8c",
          2801 => x"51",
          2802 => x"56",
          2803 => x"85",
          2804 => x"83",
          2805 => x"d5",
          2806 => x"3d",
          2807 => x"71",
          2808 => x"53",
          2809 => x"0d",
          2810 => x"71",
          2811 => x"14",
          2812 => x"33",
          2813 => x"53",
          2814 => x"04",
          2815 => x"92",
          2816 => x"81",
          2817 => x"70",
          2818 => x"3d",
          2819 => x"70",
          2820 => x"51",
          2821 => x"70",
          2822 => x"05",
          2823 => x"72",
          2824 => x"0d",
          2825 => x"80",
          2826 => x"53",
          2827 => x"ff",
          2828 => x"04",
          2829 => x"52",
          2830 => x"34",
          2831 => x"3d",
          2832 => x"79",
          2833 => x"56",
          2834 => x"71",
          2835 => x"52",
          2836 => x"2e",
          2837 => x"86",
          2838 => x"76",
          2839 => x"8a",
          2840 => x"71",
          2841 => x"0c",
          2842 => x"d5",
          2843 => x"70",
          2844 => x"70",
          2845 => x"55",
          2846 => x"80",
          2847 => x"51",
          2848 => x"08",
          2849 => x"2e",
          2850 => x"74",
          2851 => x"04",
          2852 => x"83",
          2853 => x"80",
          2854 => x"53",
          2855 => x"52",
          2856 => x"08",
          2857 => x"82",
          2858 => x"16",
          2859 => x"18",
          2860 => x"9f",
          2861 => x"2e",
          2862 => x"76",
          2863 => x"51",
          2864 => x"79",
          2865 => x"04",
          2866 => x"80",
          2867 => x"38",
          2868 => x"e4",
          2869 => x"38",
          2870 => x"81",
          2871 => x"d5",
          2872 => x"55",
          2873 => x"82",
          2874 => x"f8",
          2875 => x"c0",
          2876 => x"d5",
          2877 => x"55",
          2878 => x"f0",
          2879 => x"2e",
          2880 => x"80",
          2881 => x"17",
          2882 => x"d4",
          2883 => x"d8",
          2884 => x"75",
          2885 => x"e4",
          2886 => x"de",
          2887 => x"17",
          2888 => x"52",
          2889 => x"a4",
          2890 => x"0c",
          2891 => x"33",
          2892 => x"34",
          2893 => x"51",
          2894 => x"80",
          2895 => x"d5",
          2896 => x"3d",
          2897 => x"fe",
          2898 => x"73",
          2899 => x"71",
          2900 => x"75",
          2901 => x"04",
          2902 => x"56",
          2903 => x"38",
          2904 => x"38",
          2905 => x"2e",
          2906 => x"38",
          2907 => x"39",
          2908 => x"b6",
          2909 => x"2a",
          2910 => x"55",
          2911 => x"81",
          2912 => x"b8",
          2913 => x"a8",
          2914 => x"57",
          2915 => x"08",
          2916 => x"14",
          2917 => x"07",
          2918 => x"52",
          2919 => x"75",
          2920 => x"76",
          2921 => x"73",
          2922 => x"08",
          2923 => x"06",
          2924 => x"3f",
          2925 => x"06",
          2926 => x"15",
          2927 => x"3f",
          2928 => x"82",
          2929 => x"05",
          2930 => x"08",
          2931 => x"58",
          2932 => x"0d",
          2933 => x"5a",
          2934 => x"82",
          2935 => x"82",
          2936 => x"2e",
          2937 => x"38",
          2938 => x"39",
          2939 => x"f7",
          2940 => x"2a",
          2941 => x"55",
          2942 => x"59",
          2943 => x"74",
          2944 => x"16",
          2945 => x"53",
          2946 => x"2b",
          2947 => x"71",
          2948 => x"0b",
          2949 => x"17",
          2950 => x"3f",
          2951 => x"e4",
          2952 => x"06",
          2953 => x"54",
          2954 => x"33",
          2955 => x"51",
          2956 => x"76",
          2957 => x"75",
          2958 => x"08",
          2959 => x"38",
          2960 => x"10",
          2961 => x"51",
          2962 => x"2a",
          2963 => x"f9",
          2964 => x"82",
          2965 => x"0a",
          2966 => x"70",
          2967 => x"54",
          2968 => x"8f",
          2969 => x"f6",
          2970 => x"78",
          2971 => x"04",
          2972 => x"08",
          2973 => x"a4",
          2974 => x"38",
          2975 => x"73",
          2976 => x"d5",
          2977 => x"80",
          2978 => x"eb",
          2979 => x"d5",
          2980 => x"52",
          2981 => x"e4",
          2982 => x"2e",
          2983 => x"81",
          2984 => x"ff",
          2985 => x"75",
          2986 => x"08",
          2987 => x"94",
          2988 => x"27",
          2989 => x"84",
          2990 => x"17",
          2991 => x"a6",
          2992 => x"0c",
          2993 => x"7c",
          2994 => x"95",
          2995 => x"2e",
          2996 => x"b2",
          2997 => x"7a",
          2998 => x"82",
          2999 => x"82",
          3000 => x"08",
          3001 => x"08",
          3002 => x"38",
          3003 => x"54",
          3004 => x"7a",
          3005 => x"81",
          3006 => x"83",
          3007 => x"f9",
          3008 => x"08",
          3009 => x"82",
          3010 => x"08",
          3011 => x"25",
          3012 => x"54",
          3013 => x"38",
          3014 => x"38",
          3015 => x"90",
          3016 => x"38",
          3017 => x"38",
          3018 => x"08",
          3019 => x"78",
          3020 => x"51",
          3021 => x"80",
          3022 => x"e4",
          3023 => x"38",
          3024 => x"e4",
          3025 => x"80",
          3026 => x"55",
          3027 => x"09",
          3028 => x"80",
          3029 => x"51",
          3030 => x"82",
          3031 => x"e4",
          3032 => x"79",
          3033 => x"8f",
          3034 => x"f9",
          3035 => x"74",
          3036 => x"17",
          3037 => x"54",
          3038 => x"94",
          3039 => x"54",
          3040 => x"56",
          3041 => x"80",
          3042 => x"55",
          3043 => x"82",
          3044 => x"f8",
          3045 => x"f0",
          3046 => x"56",
          3047 => x"7b",
          3048 => x"d5",
          3049 => x"17",
          3050 => x"b8",
          3051 => x"77",
          3052 => x"15",
          3053 => x"81",
          3054 => x"15",
          3055 => x"e4",
          3056 => x"22",
          3057 => x"70",
          3058 => x"82",
          3059 => x"f8",
          3060 => x"56",
          3061 => x"f1",
          3062 => x"e9",
          3063 => x"08",
          3064 => x"82",
          3065 => x"54",
          3066 => x"82",
          3067 => x"79",
          3068 => x"98",
          3069 => x"22",
          3070 => x"26",
          3071 => x"b0",
          3072 => x"d5",
          3073 => x"0b",
          3074 => x"9c",
          3075 => x"85",
          3076 => x"31",
          3077 => x"f4",
          3078 => x"18",
          3079 => x"08",
          3080 => x"38",
          3081 => x"89",
          3082 => x"ff",
          3083 => x"80",
          3084 => x"3d",
          3085 => x"08",
          3086 => x"54",
          3087 => x"80",
          3088 => x"53",
          3089 => x"38",
          3090 => x"b5",
          3091 => x"14",
          3092 => x"2a",
          3093 => x"26",
          3094 => x"16",
          3095 => x"53",
          3096 => x"51",
          3097 => x"53",
          3098 => x"08",
          3099 => x"d5",
          3100 => x"9c",
          3101 => x"80",
          3102 => x"15",
          3103 => x"14",
          3104 => x"82",
          3105 => x"d5",
          3106 => x"82",
          3107 => x"ba",
          3108 => x"ff",
          3109 => x"52",
          3110 => x"e4",
          3111 => x"72",
          3112 => x"d5",
          3113 => x"15",
          3114 => x"0c",
          3115 => x"8a",
          3116 => x"7d",
          3117 => x"76",
          3118 => x"08",
          3119 => x"38",
          3120 => x"08",
          3121 => x"d5",
          3122 => x"80",
          3123 => x"18",
          3124 => x"81",
          3125 => x"81",
          3126 => x"83",
          3127 => x"72",
          3128 => x"75",
          3129 => x"a5",
          3130 => x"52",
          3131 => x"e4",
          3132 => x"2e",
          3133 => x"81",
          3134 => x"d5",
          3135 => x"3d",
          3136 => x"ae",
          3137 => x"ff",
          3138 => x"71",
          3139 => x"94",
          3140 => x"e4",
          3141 => x"82",
          3142 => x"fc",
          3143 => x"ff",
          3144 => x"eb",
          3145 => x"72",
          3146 => x"73",
          3147 => x"98",
          3148 => x"0d",
          3149 => x"81",
          3150 => x"70",
          3151 => x"81",
          3152 => x"51",
          3153 => x"0c",
          3154 => x"60",
          3155 => x"5b",
          3156 => x"08",
          3157 => x"08",
          3158 => x"d5",
          3159 => x"82",
          3160 => x"55",
          3161 => x"dc",
          3162 => x"81",
          3163 => x"34",
          3164 => x"e5",
          3165 => x"56",
          3166 => x"2e",
          3167 => x"75",
          3168 => x"d5",
          3169 => x"72",
          3170 => x"81",
          3171 => x"ff",
          3172 => x"09",
          3173 => x"2a",
          3174 => x"2e",
          3175 => x"bf",
          3176 => x"0c",
          3177 => x"81",
          3178 => x"53",
          3179 => x"8f",
          3180 => x"5a",
          3181 => x"83",
          3182 => x"38",
          3183 => x"29",
          3184 => x"58",
          3185 => x"51",
          3186 => x"83",
          3187 => x"96",
          3188 => x"38",
          3189 => x"73",
          3190 => x"83",
          3191 => x"38",
          3192 => x"38",
          3193 => x"06",
          3194 => x"38",
          3195 => x"10",
          3196 => x"70",
          3197 => x"81",
          3198 => x"93",
          3199 => x"d5",
          3200 => x"7d",
          3201 => x"0c",
          3202 => x"d2",
          3203 => x"d5",
          3204 => x"fd",
          3205 => x"1a",
          3206 => x"3d",
          3207 => x"08",
          3208 => x"d7",
          3209 => x"d5",
          3210 => x"70",
          3211 => x"98",
          3212 => x"3f",
          3213 => x"e4",
          3214 => x"70",
          3215 => x"58",
          3216 => x"06",
          3217 => x"86",
          3218 => x"c3",
          3219 => x"51",
          3220 => x"82",
          3221 => x"06",
          3222 => x"86",
          3223 => x"73",
          3224 => x"81",
          3225 => x"38",
          3226 => x"70",
          3227 => x"5d",
          3228 => x"81",
          3229 => x"76",
          3230 => x"8c",
          3231 => x"b6",
          3232 => x"ff",
          3233 => x"33",
          3234 => x"59",
          3235 => x"e4",
          3236 => x"3f",
          3237 => x"06",
          3238 => x"81",
          3239 => x"80",
          3240 => x"78",
          3241 => x"19",
          3242 => x"82",
          3243 => x"80",
          3244 => x"83",
          3245 => x"38",
          3246 => x"a5",
          3247 => x"81",
          3248 => x"90",
          3249 => x"10",
          3250 => x"38",
          3251 => x"54",
          3252 => x"bb",
          3253 => x"b5",
          3254 => x"06",
          3255 => x"19",
          3256 => x"8b",
          3257 => x"51",
          3258 => x"80",
          3259 => x"0b",
          3260 => x"f5",
          3261 => x"82",
          3262 => x"38",
          3263 => x"0d",
          3264 => x"ab",
          3265 => x"5a",
          3266 => x"8c",
          3267 => x"73",
          3268 => x"10",
          3269 => x"39",
          3270 => x"3d",
          3271 => x"02",
          3272 => x"73",
          3273 => x"0b",
          3274 => x"08",
          3275 => x"78",
          3276 => x"80",
          3277 => x"83",
          3278 => x"2e",
          3279 => x"82",
          3280 => x"06",
          3281 => x"90",
          3282 => x"56",
          3283 => x"a0",
          3284 => x"80",
          3285 => x"87",
          3286 => x"74",
          3287 => x"27",
          3288 => x"34",
          3289 => x"57",
          3290 => x"ec",
          3291 => x"80",
          3292 => x"73",
          3293 => x"33",
          3294 => x"e4",
          3295 => x"54",
          3296 => x"55",
          3297 => x"38",
          3298 => x"39",
          3299 => x"78",
          3300 => x"76",
          3301 => x"15",
          3302 => x"34",
          3303 => x"f9",
          3304 => x"38",
          3305 => x"fe",
          3306 => x"2e",
          3307 => x"55",
          3308 => x"81",
          3309 => x"05",
          3310 => x"05",
          3311 => x"51",
          3312 => x"90",
          3313 => x"f9",
          3314 => x"59",
          3315 => x"82",
          3316 => x"08",
          3317 => x"80",
          3318 => x"90",
          3319 => x"51",
          3320 => x"57",
          3321 => x"a0",
          3322 => x"e4",
          3323 => x"08",
          3324 => x"d5",
          3325 => x"81",
          3326 => x"08",
          3327 => x"7c",
          3328 => x"34",
          3329 => x"82",
          3330 => x"df",
          3331 => x"77",
          3332 => x"8b",
          3333 => x"17",
          3334 => x"e4",
          3335 => x"3f",
          3336 => x"81",
          3337 => x"73",
          3338 => x"10",
          3339 => x"38",
          3340 => x"34",
          3341 => x"79",
          3342 => x"08",
          3343 => x"38",
          3344 => x"98",
          3345 => x"3f",
          3346 => x"e4",
          3347 => x"e4",
          3348 => x"c0",
          3349 => x"1a",
          3350 => x"08",
          3351 => x"73",
          3352 => x"34",
          3353 => x"94",
          3354 => x"70",
          3355 => x"56",
          3356 => x"38",
          3357 => x"82",
          3358 => x"08",
          3359 => x"75",
          3360 => x"08",
          3361 => x"9c",
          3362 => x"0b",
          3363 => x"27",
          3364 => x"74",
          3365 => x"08",
          3366 => x"c3",
          3367 => x"83",
          3368 => x"0c",
          3369 => x"7e",
          3370 => x"0b",
          3371 => x"2e",
          3372 => x"2e",
          3373 => x"8c",
          3374 => x"5c",
          3375 => x"78",
          3376 => x"56",
          3377 => x"15",
          3378 => x"72",
          3379 => x"80",
          3380 => x"ff",
          3381 => x"52",
          3382 => x"d7",
          3383 => x"ff",
          3384 => x"95",
          3385 => x"88",
          3386 => x"15",
          3387 => x"76",
          3388 => x"80",
          3389 => x"2e",
          3390 => x"7a",
          3391 => x"5b",
          3392 => x"22",
          3393 => x"7a",
          3394 => x"06",
          3395 => x"53",
          3396 => x"89",
          3397 => x"19",
          3398 => x"74",
          3399 => x"09",
          3400 => x"78",
          3401 => x"80",
          3402 => x"90",
          3403 => x"76",
          3404 => x"57",
          3405 => x"81",
          3406 => x"38",
          3407 => x"81",
          3408 => x"81",
          3409 => x"96",
          3410 => x"72",
          3411 => x"72",
          3412 => x"89",
          3413 => x"11",
          3414 => x"9c",
          3415 => x"88",
          3416 => x"53",
          3417 => x"81",
          3418 => x"a0",
          3419 => x"53",
          3420 => x"81",
          3421 => x"56",
          3422 => x"77",
          3423 => x"14",
          3424 => x"51",
          3425 => x"34",
          3426 => x"88",
          3427 => x"52",
          3428 => x"08",
          3429 => x"3f",
          3430 => x"98",
          3431 => x"e4",
          3432 => x"04",
          3433 => x"5e",
          3434 => x"73",
          3435 => x"80",
          3436 => x"8d",
          3437 => x"0c",
          3438 => x"70",
          3439 => x"09",
          3440 => x"80",
          3441 => x"78",
          3442 => x"73",
          3443 => x"54",
          3444 => x"0b",
          3445 => x"e7",
          3446 => x"87",
          3447 => x"11",
          3448 => x"fc",
          3449 => x"e4",
          3450 => x"ff",
          3451 => x"92",
          3452 => x"08",
          3453 => x"81",
          3454 => x"ff",
          3455 => x"9f",
          3456 => x"51",
          3457 => x"dc",
          3458 => x"91",
          3459 => x"d9",
          3460 => x"de",
          3461 => x"38",
          3462 => x"81",
          3463 => x"41",
          3464 => x"73",
          3465 => x"81",
          3466 => x"70",
          3467 => x"73",
          3468 => x"82",
          3469 => x"06",
          3470 => x"2e",
          3471 => x"2e",
          3472 => x"1a",
          3473 => x"06",
          3474 => x"ae",
          3475 => x"10",
          3476 => x"a0",
          3477 => x"26",
          3478 => x"81",
          3479 => x"78",
          3480 => x"73",
          3481 => x"80",
          3482 => x"05",
          3483 => x"a0",
          3484 => x"51",
          3485 => x"84",
          3486 => x"78",
          3487 => x"56",
          3488 => x"56",
          3489 => x"83",
          3490 => x"ff",
          3491 => x"2e",
          3492 => x"70",
          3493 => x"73",
          3494 => x"74",
          3495 => x"2e",
          3496 => x"07",
          3497 => x"16",
          3498 => x"ae",
          3499 => x"05",
          3500 => x"8f",
          3501 => x"73",
          3502 => x"8b",
          3503 => x"e8",
          3504 => x"7c",
          3505 => x"57",
          3506 => x"75",
          3507 => x"70",
          3508 => x"7c",
          3509 => x"89",
          3510 => x"80",
          3511 => x"38",
          3512 => x"70",
          3513 => x"51",
          3514 => x"38",
          3515 => x"79",
          3516 => x"7c",
          3517 => x"88",
          3518 => x"06",
          3519 => x"76",
          3520 => x"83",
          3521 => x"3f",
          3522 => x"06",
          3523 => x"55",
          3524 => x"80",
          3525 => x"57",
          3526 => x"ff",
          3527 => x"76",
          3528 => x"39",
          3529 => x"55",
          3530 => x"80",
          3531 => x"75",
          3532 => x"3f",
          3533 => x"38",
          3534 => x"a4",
          3535 => x"26",
          3536 => x"9f",
          3537 => x"7b",
          3538 => x"ff",
          3539 => x"05",
          3540 => x"fd",
          3541 => x"81",
          3542 => x"85",
          3543 => x"09",
          3544 => x"81",
          3545 => x"73",
          3546 => x"54",
          3547 => x"38",
          3548 => x"70",
          3549 => x"7b",
          3550 => x"38",
          3551 => x"70",
          3552 => x"85",
          3553 => x"1f",
          3554 => x"d5",
          3555 => x"82",
          3556 => x"82",
          3557 => x"06",
          3558 => x"81",
          3559 => x"73",
          3560 => x"54",
          3561 => x"80",
          3562 => x"c2",
          3563 => x"38",
          3564 => x"70",
          3565 => x"86",
          3566 => x"06",
          3567 => x"38",
          3568 => x"05",
          3569 => x"3f",
          3570 => x"f8",
          3571 => x"92",
          3572 => x"5b",
          3573 => x"59",
          3574 => x"c6",
          3575 => x"70",
          3576 => x"8d",
          3577 => x"09",
          3578 => x"d0",
          3579 => x"53",
          3580 => x"73",
          3581 => x"71",
          3582 => x"82",
          3583 => x"55",
          3584 => x"74",
          3585 => x"12",
          3586 => x"38",
          3587 => x"51",
          3588 => x"89",
          3589 => x"53",
          3590 => x"51",
          3591 => x"38",
          3592 => x"77",
          3593 => x"2a",
          3594 => x"51",
          3595 => x"84",
          3596 => x"94",
          3597 => x"38",
          3598 => x"86",
          3599 => x"82",
          3600 => x"fa",
          3601 => x"17",
          3602 => x"52",
          3603 => x"82",
          3604 => x"b6",
          3605 => x"e4",
          3606 => x"55",
          3607 => x"06",
          3608 => x"33",
          3609 => x"81",
          3610 => x"eb",
          3611 => x"07",
          3612 => x"81",
          3613 => x"83",
          3614 => x"16",
          3615 => x"08",
          3616 => x"9d",
          3617 => x"81",
          3618 => x"d5",
          3619 => x"80",
          3620 => x"d5",
          3621 => x"3d",
          3622 => x"05",
          3623 => x"51",
          3624 => x"58",
          3625 => x"08",
          3626 => x"08",
          3627 => x"08",
          3628 => x"87",
          3629 => x"fe",
          3630 => x"2e",
          3631 => x"a0",
          3632 => x"06",
          3633 => x"38",
          3634 => x"82",
          3635 => x"56",
          3636 => x"80",
          3637 => x"d8",
          3638 => x"81",
          3639 => x"d5",
          3640 => x"06",
          3641 => x"38",
          3642 => x"2a",
          3643 => x"72",
          3644 => x"52",
          3645 => x"08",
          3646 => x"93",
          3647 => x"82",
          3648 => x"2e",
          3649 => x"59",
          3650 => x"58",
          3651 => x"fe",
          3652 => x"e4",
          3653 => x"5b",
          3654 => x"75",
          3655 => x"d5",
          3656 => x"2a",
          3657 => x"29",
          3658 => x"57",
          3659 => x"80",
          3660 => x"fc",
          3661 => x"ff",
          3662 => x"1a",
          3663 => x"81",
          3664 => x"27",
          3665 => x"81",
          3666 => x"27",
          3667 => x"84",
          3668 => x"84",
          3669 => x"86",
          3670 => x"ff",
          3671 => x"81",
          3672 => x"51",
          3673 => x"83",
          3674 => x"80",
          3675 => x"d5",
          3676 => x"80",
          3677 => x"c8",
          3678 => x"06",
          3679 => x"26",
          3680 => x"78",
          3681 => x"59",
          3682 => x"2e",
          3683 => x"72",
          3684 => x"f2",
          3685 => x"3f",
          3686 => x"e4",
          3687 => x"57",
          3688 => x"cb",
          3689 => x"e4",
          3690 => x"8d",
          3691 => x"3f",
          3692 => x"14",
          3693 => x"08",
          3694 => x"72",
          3695 => x"22",
          3696 => x"5a",
          3697 => x"14",
          3698 => x"e1",
          3699 => x"82",
          3700 => x"38",
          3701 => x"ff",
          3702 => x"83",
          3703 => x"74",
          3704 => x"89",
          3705 => x"ca",
          3706 => x"7b",
          3707 => x"17",
          3708 => x"55",
          3709 => x"38",
          3710 => x"82",
          3711 => x"53",
          3712 => x"82",
          3713 => x"bd",
          3714 => x"0c",
          3715 => x"56",
          3716 => x"13",
          3717 => x"82",
          3718 => x"81",
          3719 => x"83",
          3720 => x"72",
          3721 => x"ff",
          3722 => x"15",
          3723 => x"76",
          3724 => x"38",
          3725 => x"82",
          3726 => x"53",
          3727 => x"f9",
          3728 => x"88",
          3729 => x"38",
          3730 => x"84",
          3731 => x"d5",
          3732 => x"72",
          3733 => x"80",
          3734 => x"3f",
          3735 => x"a4",
          3736 => x"84",
          3737 => x"d5",
          3738 => x"2e",
          3739 => x"14",
          3740 => x"08",
          3741 => x"c5",
          3742 => x"15",
          3743 => x"22",
          3744 => x"23",
          3745 => x"0b",
          3746 => x"0c",
          3747 => x"90",
          3748 => x"54",
          3749 => x"73",
          3750 => x"72",
          3751 => x"86",
          3752 => x"71",
          3753 => x"81",
          3754 => x"82",
          3755 => x"88",
          3756 => x"39",
          3757 => x"74",
          3758 => x"04",
          3759 => x"7a",
          3760 => x"f4",
          3761 => x"d5",
          3762 => x"e4",
          3763 => x"70",
          3764 => x"38",
          3765 => x"2e",
          3766 => x"0c",
          3767 => x"80",
          3768 => x"51",
          3769 => x"54",
          3770 => x"0d",
          3771 => x"05",
          3772 => x"54",
          3773 => x"bf",
          3774 => x"53",
          3775 => x"ae",
          3776 => x"d5",
          3777 => x"69",
          3778 => x"b0",
          3779 => x"d5",
          3780 => x"05",
          3781 => x"80",
          3782 => x"06",
          3783 => x"74",
          3784 => x"09",
          3785 => x"b1",
          3786 => x"39",
          3787 => x"73",
          3788 => x"81",
          3789 => x"38",
          3790 => x"07",
          3791 => x"2a",
          3792 => x"2e",
          3793 => x"d6",
          3794 => x"82",
          3795 => x"51",
          3796 => x"8b",
          3797 => x"51",
          3798 => x"05",
          3799 => x"0b",
          3800 => x"f1",
          3801 => x"80",
          3802 => x"51",
          3803 => x"55",
          3804 => x"b7",
          3805 => x"05",
          3806 => x"51",
          3807 => x"84",
          3808 => x"70",
          3809 => x"a9",
          3810 => x"2e",
          3811 => x"73",
          3812 => x"d5",
          3813 => x"0c",
          3814 => x"f8",
          3815 => x"51",
          3816 => x"80",
          3817 => x"a0",
          3818 => x"53",
          3819 => x"d5",
          3820 => x"1b",
          3821 => x"dd",
          3822 => x"e4",
          3823 => x"56",
          3824 => x"90",
          3825 => x"80",
          3826 => x"1a",
          3827 => x"51",
          3828 => x"82",
          3829 => x"38",
          3830 => x"8a",
          3831 => x"59",
          3832 => x"c5",
          3833 => x"82",
          3834 => x"82",
          3835 => x"09",
          3836 => x"78",
          3837 => x"80",
          3838 => x"38",
          3839 => x"c3",
          3840 => x"38",
          3841 => x"2e",
          3842 => x"ee",
          3843 => x"82",
          3844 => x"d5",
          3845 => x"39",
          3846 => x"d5",
          3847 => x"3d",
          3848 => x"5d",
          3849 => x"05",
          3850 => x"d5",
          3851 => x"8a",
          3852 => x"2e",
          3853 => x"90",
          3854 => x"74",
          3855 => x"82",
          3856 => x"ad",
          3857 => x"56",
          3858 => x"1a",
          3859 => x"38",
          3860 => x"38",
          3861 => x"56",
          3862 => x"11",
          3863 => x"5b",
          3864 => x"88",
          3865 => x"08",
          3866 => x"d5",
          3867 => x"9f",
          3868 => x"74",
          3869 => x"7e",
          3870 => x"08",
          3871 => x"e4",
          3872 => x"77",
          3873 => x"7f",
          3874 => x"75",
          3875 => x"77",
          3876 => x"33",
          3877 => x"e4",
          3878 => x"33",
          3879 => x"b4",
          3880 => x"27",
          3881 => x"52",
          3882 => x"7d",
          3883 => x"89",
          3884 => x"0c",
          3885 => x"80",
          3886 => x"83",
          3887 => x"7e",
          3888 => x"08",
          3889 => x"08",
          3890 => x"7c",
          3891 => x"31",
          3892 => x"94",
          3893 => x"5c",
          3894 => x"d5",
          3895 => x"3d",
          3896 => x"5d",
          3897 => x"05",
          3898 => x"d5",
          3899 => x"8a",
          3900 => x"2e",
          3901 => x"90",
          3902 => x"06",
          3903 => x"2e",
          3904 => x"91",
          3905 => x"81",
          3906 => x"95",
          3907 => x"56",
          3908 => x"5c",
          3909 => x"18",
          3910 => x"74",
          3911 => x"ff",
          3912 => x"7a",
          3913 => x"08",
          3914 => x"39",
          3915 => x"ac",
          3916 => x"d5",
          3917 => x"74",
          3918 => x"2e",
          3919 => x"88",
          3920 => x"0c",
          3921 => x"08",
          3922 => x"51",
          3923 => x"08",
          3924 => x"7e",
          3925 => x"e4",
          3926 => x"d5",
          3927 => x"57",
          3928 => x"1b",
          3929 => x"75",
          3930 => x"59",
          3931 => x"1a",
          3932 => x"d5",
          3933 => x"11",
          3934 => x"27",
          3935 => x"08",
          3936 => x"b8",
          3937 => x"55",
          3938 => x"2b",
          3939 => x"94",
          3940 => x"ff",
          3941 => x"fd",
          3942 => x"55",
          3943 => x"83",
          3944 => x"55",
          3945 => x"9c",
          3946 => x"b8",
          3947 => x"38",
          3948 => x"83",
          3949 => x"b9",
          3950 => x"16",
          3951 => x"7f",
          3952 => x"70",
          3953 => x"58",
          3954 => x"75",
          3955 => x"39",
          3956 => x"74",
          3957 => x"d5",
          3958 => x"3d",
          3959 => x"70",
          3960 => x"e4",
          3961 => x"80",
          3962 => x"70",
          3963 => x"2e",
          3964 => x"78",
          3965 => x"e4",
          3966 => x"d8",
          3967 => x"a0",
          3968 => x"88",
          3969 => x"51",
          3970 => x"9c",
          3971 => x"88",
          3972 => x"b7",
          3973 => x"ff",
          3974 => x"83",
          3975 => x"3f",
          3976 => x"81",
          3977 => x"34",
          3978 => x"0d",
          3979 => x"54",
          3980 => x"53",
          3981 => x"3d",
          3982 => x"3f",
          3983 => x"e4",
          3984 => x"74",
          3985 => x"3d",
          3986 => x"51",
          3987 => x"82",
          3988 => x"d5",
          3989 => x"52",
          3990 => x"0d",
          3991 => x"3d",
          3992 => x"e6",
          3993 => x"d5",
          3994 => x"64",
          3995 => x"e8",
          3996 => x"d5",
          3997 => x"05",
          3998 => x"80",
          3999 => x"0c",
          4000 => x"70",
          4001 => x"56",
          4002 => x"53",
          4003 => x"d5",
          4004 => x"82",
          4005 => x"06",
          4006 => x"e4",
          4007 => x"3d",
          4008 => x"3d",
          4009 => x"53",
          4010 => x"80",
          4011 => x"d5",
          4012 => x"83",
          4013 => x"7a",
          4014 => x"0c",
          4015 => x"73",
          4016 => x"80",
          4017 => x"3f",
          4018 => x"e4",
          4019 => x"08",
          4020 => x"82",
          4021 => x"08",
          4022 => x"52",
          4023 => x"e4",
          4024 => x"74",
          4025 => x"08",
          4026 => x"38",
          4027 => x"82",
          4028 => x"08",
          4029 => x"7b",
          4030 => x"e4",
          4031 => x"51",
          4032 => x"57",
          4033 => x"38",
          4034 => x"38",
          4035 => x"ea",
          4036 => x"52",
          4037 => x"3d",
          4038 => x"5a",
          4039 => x"80",
          4040 => x"70",
          4041 => x"81",
          4042 => x"38",
          4043 => x"82",
          4044 => x"08",
          4045 => x"55",
          4046 => x"38",
          4047 => x"55",
          4048 => x"77",
          4049 => x"ff",
          4050 => x"58",
          4051 => x"c0",
          4052 => x"05",
          4053 => x"56",
          4054 => x"16",
          4055 => x"73",
          4056 => x"26",
          4057 => x"91",
          4058 => x"70",
          4059 => x"ec",
          4060 => x"34",
          4061 => x"38",
          4062 => x"08",
          4063 => x"7a",
          4064 => x"26",
          4065 => x"d5",
          4066 => x"f7",
          4067 => x"05",
          4068 => x"3f",
          4069 => x"e4",
          4070 => x"53",
          4071 => x"54",
          4072 => x"33",
          4073 => x"54",
          4074 => x"15",
          4075 => x"58",
          4076 => x"8a",
          4077 => x"53",
          4078 => x"ff",
          4079 => x"d5",
          4080 => x"53",
          4081 => x"d5",
          4082 => x"30",
          4083 => x"77",
          4084 => x"51",
          4085 => x"73",
          4086 => x"bb",
          4087 => x"82",
          4088 => x"38",
          4089 => x"9e",
          4090 => x"0c",
          4091 => x"81",
          4092 => x"38",
          4093 => x"94",
          4094 => x"2a",
          4095 => x"72",
          4096 => x"51",
          4097 => x"08",
          4098 => x"82",
          4099 => x"52",
          4100 => x"d5",
          4101 => x"38",
          4102 => x"73",
          4103 => x"98",
          4104 => x"08",
          4105 => x"06",
          4106 => x"52",
          4107 => x"d5",
          4108 => x"16",
          4109 => x"0b",
          4110 => x"75",
          4111 => x"58",
          4112 => x"74",
          4113 => x"90",
          4114 => x"90",
          4115 => x"72",
          4116 => x"08",
          4117 => x"80",
          4118 => x"3d",
          4119 => x"89",
          4120 => x"80",
          4121 => x"3d",
          4122 => x"d5",
          4123 => x"80",
          4124 => x"75",
          4125 => x"08",
          4126 => x"38",
          4127 => x"57",
          4128 => x"33",
          4129 => x"55",
          4130 => x"16",
          4131 => x"82",
          4132 => x"54",
          4133 => x"52",
          4134 => x"d5",
          4135 => x"81",
          4136 => x"74",
          4137 => x"74",
          4138 => x"3d",
          4139 => x"3d",
          4140 => x"bb",
          4141 => x"82",
          4142 => x"0d",
          4143 => x"3d",
          4144 => x"e7",
          4145 => x"82",
          4146 => x"94",
          4147 => x"51",
          4148 => x"08",
          4149 => x"08",
          4150 => x"d5",
          4151 => x"84",
          4152 => x"53",
          4153 => x"38",
          4154 => x"72",
          4155 => x"82",
          4156 => x"70",
          4157 => x"e4",
          4158 => x"82",
          4159 => x"ed",
          4160 => x"3d",
          4161 => x"9e",
          4162 => x"d5",
          4163 => x"51",
          4164 => x"55",
          4165 => x"80",
          4166 => x"58",
          4167 => x"8d",
          4168 => x"52",
          4169 => x"d5",
          4170 => x"3d",
          4171 => x"92",
          4172 => x"dd",
          4173 => x"82",
          4174 => x"74",
          4175 => x"11",
          4176 => x"75",
          4177 => x"81",
          4178 => x"82",
          4179 => x"08",
          4180 => x"09",
          4181 => x"5f",
          4182 => x"51",
          4183 => x"08",
          4184 => x"08",
          4185 => x"08",
          4186 => x"80",
          4187 => x"59",
          4188 => x"c9",
          4189 => x"82",
          4190 => x"38",
          4191 => x"ff",
          4192 => x"5b",
          4193 => x"7c",
          4194 => x"52",
          4195 => x"06",
          4196 => x"8e",
          4197 => x"ff",
          4198 => x"82",
          4199 => x"b8",
          4200 => x"d5",
          4201 => x"70",
          4202 => x"51",
          4203 => x"56",
          4204 => x"7c",
          4205 => x"81",
          4206 => x"7a",
          4207 => x"04",
          4208 => x"05",
          4209 => x"82",
          4210 => x"08",
          4211 => x"75",
          4212 => x"81",
          4213 => x"87",
          4214 => x"94",
          4215 => x"27",
          4216 => x"d5",
          4217 => x"76",
          4218 => x"e4",
          4219 => x"ca",
          4220 => x"ff",
          4221 => x"ff",
          4222 => x"56",
          4223 => x"81",
          4224 => x"75",
          4225 => x"08",
          4226 => x"17",
          4227 => x"76",
          4228 => x"e4",
          4229 => x"0c",
          4230 => x"73",
          4231 => x"38",
          4232 => x"82",
          4233 => x"e0",
          4234 => x"9c",
          4235 => x"3f",
          4236 => x"e4",
          4237 => x"3d",
          4238 => x"cd",
          4239 => x"82",
          4240 => x"80",
          4241 => x"81",
          4242 => x"81",
          4243 => x"74",
          4244 => x"05",
          4245 => x"55",
          4246 => x"51",
          4247 => x"08",
          4248 => x"55",
          4249 => x"78",
          4250 => x"08",
          4251 => x"d5",
          4252 => x"70",
          4253 => x"d5",
          4254 => x"80",
          4255 => x"73",
          4256 => x"e4",
          4257 => x"38",
          4258 => x"e4",
          4259 => x"e4",
          4260 => x"ab",
          4261 => x"e4",
          4262 => x"07",
          4263 => x"2e",
          4264 => x"80",
          4265 => x"90",
          4266 => x"8c",
          4267 => x"82",
          4268 => x"e4",
          4269 => x"0d",
          4270 => x"52",
          4271 => x"d5",
          4272 => x"82",
          4273 => x"3d",
          4274 => x"d5",
          4275 => x"86",
          4276 => x"d5",
          4277 => x"82",
          4278 => x"70",
          4279 => x"54",
          4280 => x"52",
          4281 => x"bc",
          4282 => x"56",
          4283 => x"54",
          4284 => x"81",
          4285 => x"e4",
          4286 => x"38",
          4287 => x"b6",
          4288 => x"51",
          4289 => x"08",
          4290 => x"38",
          4291 => x"ff",
          4292 => x"b8",
          4293 => x"c3",
          4294 => x"80",
          4295 => x"75",
          4296 => x"b7",
          4297 => x"53",
          4298 => x"3f",
          4299 => x"34",
          4300 => x"51",
          4301 => x"0b",
          4302 => x"89",
          4303 => x"d5",
          4304 => x"0a",
          4305 => x"86",
          4306 => x"ff",
          4307 => x"8b",
          4308 => x"15",
          4309 => x"82",
          4310 => x"53",
          4311 => x"3f",
          4312 => x"0d",
          4313 => x"05",
          4314 => x"3d",
          4315 => x"d4",
          4316 => x"82",
          4317 => x"4e",
          4318 => x"52",
          4319 => x"08",
          4320 => x"38",
          4321 => x"06",
          4322 => x"a0",
          4323 => x"ff",
          4324 => x"b0",
          4325 => x"54",
          4326 => x"52",
          4327 => x"e4",
          4328 => x"38",
          4329 => x"06",
          4330 => x"92",
          4331 => x"d5",
          4332 => x"81",
          4333 => x"3f",
          4334 => x"e4",
          4335 => x"53",
          4336 => x"16",
          4337 => x"05",
          4338 => x"70",
          4339 => x"55",
          4340 => x"73",
          4341 => x"83",
          4342 => x"2a",
          4343 => x"80",
          4344 => x"80",
          4345 => x"b4",
          4346 => x"78",
          4347 => x"82",
          4348 => x"38",
          4349 => x"ff",
          4350 => x"79",
          4351 => x"d5",
          4352 => x"33",
          4353 => x"9a",
          4354 => x"ff",
          4355 => x"83",
          4356 => x"08",
          4357 => x"82",
          4358 => x"08",
          4359 => x"3f",
          4360 => x"d5",
          4361 => x"3d",
          4362 => x"84",
          4363 => x"82",
          4364 => x"3d",
          4365 => x"08",
          4366 => x"38",
          4367 => x"05",
          4368 => x"08",
          4369 => x"02",
          4370 => x"54",
          4371 => x"06",
          4372 => x"06",
          4373 => x"56",
          4374 => x"0b",
          4375 => x"97",
          4376 => x"82",
          4377 => x"ee",
          4378 => x"3d",
          4379 => x"ce",
          4380 => x"d5",
          4381 => x"64",
          4382 => x"d0",
          4383 => x"d5",
          4384 => x"05",
          4385 => x"73",
          4386 => x"22",
          4387 => x"1f",
          4388 => x"81",
          4389 => x"a1",
          4390 => x"74",
          4391 => x"04",
          4392 => x"80",
          4393 => x"3d",
          4394 => x"08",
          4395 => x"d5",
          4396 => x"57",
          4397 => x"70",
          4398 => x"80",
          4399 => x"52",
          4400 => x"97",
          4401 => x"d5",
          4402 => x"73",
          4403 => x"e4",
          4404 => x"38",
          4405 => x"08",
          4406 => x"19",
          4407 => x"74",
          4408 => x"ec",
          4409 => x"74",
          4410 => x"16",
          4411 => x"73",
          4412 => x"84",
          4413 => x"7a",
          4414 => x"07",
          4415 => x"80",
          4416 => x"7b",
          4417 => x"80",
          4418 => x"d5",
          4419 => x"55",
          4420 => x"8b",
          4421 => x"83",
          4422 => x"51",
          4423 => x"08",
          4424 => x"99",
          4425 => x"53",
          4426 => x"3d",
          4427 => x"08",
          4428 => x"d5",
          4429 => x"a0",
          4430 => x"9b",
          4431 => x"55",
          4432 => x"77",
          4433 => x"3f",
          4434 => x"26",
          4435 => x"51",
          4436 => x"d5",
          4437 => x"d5",
          4438 => x"74",
          4439 => x"c8",
          4440 => x"d5",
          4441 => x"27",
          4442 => x"8b",
          4443 => x"55",
          4444 => x"8f",
          4445 => x"70",
          4446 => x"74",
          4447 => x"16",
          4448 => x"9f",
          4449 => x"54",
          4450 => x"b1",
          4451 => x"a3",
          4452 => x"54",
          4453 => x"38",
          4454 => x"40",
          4455 => x"52",
          4456 => x"e4",
          4457 => x"f7",
          4458 => x"bc",
          4459 => x"d5",
          4460 => x"38",
          4461 => x"39",
          4462 => x"81",
          4463 => x"74",
          4464 => x"51",
          4465 => x"08",
          4466 => x"a0",
          4467 => x"51",
          4468 => x"0b",
          4469 => x"66",
          4470 => x"81",
          4471 => x"9c",
          4472 => x"73",
          4473 => x"3d",
          4474 => x"02",
          4475 => x"3d",
          4476 => x"5a",
          4477 => x"58",
          4478 => x"91",
          4479 => x"7c",
          4480 => x"59",
          4481 => x"81",
          4482 => x"73",
          4483 => x"82",
          4484 => x"8b",
          4485 => x"2b",
          4486 => x"fe",
          4487 => x"70",
          4488 => x"d5",
          4489 => x"40",
          4490 => x"88",
          4491 => x"38",
          4492 => x"56",
          4493 => x"3f",
          4494 => x"08",
          4495 => x"d5",
          4496 => x"82",
          4497 => x"38",
          4498 => x"16",
          4499 => x"87",
          4500 => x"74",
          4501 => x"38",
          4502 => x"2e",
          4503 => x"80",
          4504 => x"81",
          4505 => x"56",
          4506 => x"9d",
          4507 => x"82",
          4508 => x"81",
          4509 => x"d3",
          4510 => x"7c",
          4511 => x"b3",
          4512 => x"1b",
          4513 => x"54",
          4514 => x"fe",
          4515 => x"74",
          4516 => x"16",
          4517 => x"73",
          4518 => x"d5",
          4519 => x"3d",
          4520 => x"ef",
          4521 => x"59",
          4522 => x"82",
          4523 => x"82",
          4524 => x"ac",
          4525 => x"2e",
          4526 => x"e4",
          4527 => x"d5",
          4528 => x"33",
          4529 => x"ff",
          4530 => x"81",
          4531 => x"83",
          4532 => x"2a",
          4533 => x"74",
          4534 => x"53",
          4535 => x"3f",
          4536 => x"55",
          4537 => x"80",
          4538 => x"06",
          4539 => x"49",
          4540 => x"79",
          4541 => x"26",
          4542 => x"74",
          4543 => x"fe",
          4544 => x"70",
          4545 => x"7a",
          4546 => x"80",
          4547 => x"74",
          4548 => x"e0",
          4549 => x"7f",
          4550 => x"82",
          4551 => x"fe",
          4552 => x"d5",
          4553 => x"8e",
          4554 => x"81",
          4555 => x"1b",
          4556 => x"80",
          4557 => x"51",
          4558 => x"08",
          4559 => x"cd",
          4560 => x"39",
          4561 => x"7f",
          4562 => x"82",
          4563 => x"83",
          4564 => x"08",
          4565 => x"5f",
          4566 => x"8a",
          4567 => x"56",
          4568 => x"93",
          4569 => x"38",
          4570 => x"44",
          4571 => x"06",
          4572 => x"62",
          4573 => x"83",
          4574 => x"82",
          4575 => x"78",
          4576 => x"80",
          4577 => x"2a",
          4578 => x"56",
          4579 => x"77",
          4580 => x"79",
          4581 => x"5a",
          4582 => x"27",
          4583 => x"a9",
          4584 => x"29",
          4585 => x"55",
          4586 => x"08",
          4587 => x"ff",
          4588 => x"89",
          4589 => x"2a",
          4590 => x"56",
          4591 => x"77",
          4592 => x"79",
          4593 => x"5a",
          4594 => x"27",
          4595 => x"a9",
          4596 => x"84",
          4597 => x"f5",
          4598 => x"e4",
          4599 => x"71",
          4600 => x"5e",
          4601 => x"5c",
          4602 => x"05",
          4603 => x"70",
          4604 => x"57",
          4605 => x"06",
          4606 => x"5c",
          4607 => x"29",
          4608 => x"55",
          4609 => x"7c",
          4610 => x"31",
          4611 => x"d5",
          4612 => x"81",
          4613 => x"83",
          4614 => x"87",
          4615 => x"fd",
          4616 => x"2e",
          4617 => x"ff",
          4618 => x"a0",
          4619 => x"74",
          4620 => x"fd",
          4621 => x"80",
          4622 => x"39",
          4623 => x"92",
          4624 => x"59",
          4625 => x"86",
          4626 => x"09",
          4627 => x"f5",
          4628 => x"55",
          4629 => x"80",
          4630 => x"b0",
          4631 => x"7a",
          4632 => x"52",
          4633 => x"79",
          4634 => x"06",
          4635 => x"3f",
          4636 => x"32",
          4637 => x"06",
          4638 => x"8d",
          4639 => x"ff",
          4640 => x"06",
          4641 => x"3f",
          4642 => x"ff",
          4643 => x"34",
          4644 => x"d0",
          4645 => x"ff",
          4646 => x"51",
          4647 => x"09",
          4648 => x"b2",
          4649 => x"8d",
          4650 => x"ff",
          4651 => x"51",
          4652 => x"1b",
          4653 => x"b2",
          4654 => x"80",
          4655 => x"80",
          4656 => x"ac",
          4657 => x"82",
          4658 => x"ff",
          4659 => x"06",
          4660 => x"3f",
          4661 => x"0b",
          4662 => x"c0",
          4663 => x"3f",
          4664 => x"70",
          4665 => x"54",
          4666 => x"88",
          4667 => x"08",
          4668 => x"81",
          4669 => x"1f",
          4670 => x"af",
          4671 => x"51",
          4672 => x"a4",
          4673 => x"3f",
          4674 => x"e4",
          4675 => x"18",
          4676 => x"ee",
          4677 => x"ff",
          4678 => x"78",
          4679 => x"87",
          4680 => x"87",
          4681 => x"7a",
          4682 => x"66",
          4683 => x"88",
          4684 => x"2e",
          4685 => x"7a",
          4686 => x"84",
          4687 => x"0a",
          4688 => x"ff",
          4689 => x"38",
          4690 => x"8a",
          4691 => x"62",
          4692 => x"75",
          4693 => x"f7",
          4694 => x"38",
          4695 => x"52",
          4696 => x"16",
          4697 => x"38",
          4698 => x"8d",
          4699 => x"38",
          4700 => x"83",
          4701 => x"7a",
          4702 => x"82",
          4703 => x"16",
          4704 => x"38",
          4705 => x"86",
          4706 => x"38",
          4707 => x"81",
          4708 => x"54",
          4709 => x"84",
          4710 => x"08",
          4711 => x"55",
          4712 => x"82",
          4713 => x"51",
          4714 => x"62",
          4715 => x"fd",
          4716 => x"51",
          4717 => x"52",
          4718 => x"be",
          4719 => x"81",
          4720 => x"77",
          4721 => x"67",
          4722 => x"51",
          4723 => x"16",
          4724 => x"bf",
          4725 => x"d5",
          4726 => x"83",
          4727 => x"67",
          4728 => x"ce",
          4729 => x"7f",
          4730 => x"82",
          4731 => x"80",
          4732 => x"81",
          4733 => x"89",
          4734 => x"86",
          4735 => x"82",
          4736 => x"f5",
          4737 => x"79",
          4738 => x"78",
          4739 => x"55",
          4740 => x"51",
          4741 => x"81",
          4742 => x"74",
          4743 => x"81",
          4744 => x"8a",
          4745 => x"76",
          4746 => x"55",
          4747 => x"0d",
          4748 => x"05",
          4749 => x"2e",
          4750 => x"76",
          4751 => x"80",
          4752 => x"77",
          4753 => x"34",
          4754 => x"38",
          4755 => x"8c",
          4756 => x"3f",
          4757 => x"07",
          4758 => x"56",
          4759 => x"18",
          4760 => x"0d",
          4761 => x"75",
          4762 => x"54",
          4763 => x"51",
          4764 => x"91",
          4765 => x"81",
          4766 => x"83",
          4767 => x"0c",
          4768 => x"75",
          4769 => x"51",
          4770 => x"85",
          4771 => x"80",
          4772 => x"70",
          4773 => x"72",
          4774 => x"8d",
          4775 => x"0d",
          4776 => x"55",
          4777 => x"8a",
          4778 => x"80",
          4779 => x"51",
          4780 => x"b4",
          4781 => x"c9",
          4782 => x"38",
          4783 => x"53",
          4784 => x"71",
          4785 => x"51",
          4786 => x"81",
          4787 => x"e4",
          4788 => x"0d",
          4789 => x"96",
          4790 => x"80",
          4791 => x"39",
          4792 => x"91",
          4793 => x"70",
          4794 => x"54",
          4795 => x"3d",
          4796 => x"70",
          4797 => x"70",
          4798 => x"57",
          4799 => x"82",
          4800 => x"57",
          4801 => x"75",
          4802 => x"fb",
          4803 => x"70",
          4804 => x"18",
          4805 => x"80",
          4806 => x"38",
          4807 => x"51",
          4808 => x"76",
          4809 => x"c3",
          4810 => x"71",
          4811 => x"51",
          4812 => x"d0",
          4813 => x"90",
          4814 => x"b0",
          4815 => x"51",
          4816 => x"39",
          4817 => x"56",
          4818 => x"d5",
          4819 => x"ff",
          4820 => x"ff",
          4821 => x"00",
          4822 => x"00",
          4823 => x"00",
          4824 => x"00",
          4825 => x"00",
          4826 => x"00",
          4827 => x"00",
          4828 => x"00",
          4829 => x"00",
          4830 => x"00",
          4831 => x"00",
          4832 => x"00",
          4833 => x"00",
          4834 => x"00",
          4835 => x"00",
          4836 => x"00",
          4837 => x"00",
          4838 => x"00",
          4839 => x"00",
          4840 => x"00",
          4841 => x"00",
          4842 => x"00",
          4843 => x"00",
          4844 => x"00",
          4845 => x"00",
          4846 => x"00",
          4847 => x"00",
          4848 => x"00",
          4849 => x"00",
          4850 => x"00",
          4851 => x"00",
          4852 => x"00",
          4853 => x"00",
          4854 => x"00",
          4855 => x"00",
          4856 => x"00",
          4857 => x"00",
          4858 => x"00",
          4859 => x"00",
          4860 => x"00",
          4861 => x"00",
          4862 => x"00",
          4863 => x"00",
          4864 => x"00",
          4865 => x"00",
          4866 => x"00",
          4867 => x"00",
          4868 => x"00",
          4869 => x"00",
          4870 => x"00",
          4871 => x"00",
          4872 => x"00",
          4873 => x"00",
          4874 => x"00",
          4875 => x"00",
          4876 => x"00",
          4877 => x"00",
          4878 => x"00",
          4879 => x"00",
          4880 => x"00",
          4881 => x"00",
          4882 => x"00",
          4883 => x"00",
          4884 => x"00",
          4885 => x"00",
          4886 => x"00",
          4887 => x"00",
          4888 => x"00",
          4889 => x"00",
          4890 => x"00",
          4891 => x"00",
          4892 => x"00",
          4893 => x"00",
          4894 => x"00",
          4895 => x"6c",
          4896 => x"00",
          4897 => x"00",
          4898 => x"00",
          4899 => x"72",
          4900 => x"00",
          4901 => x"00",
          4902 => x"00",
          4903 => x"65",
          4904 => x"69",
          4905 => x"66",
          4906 => x"61",
          4907 => x"6d",
          4908 => x"72",
          4909 => x"00",
          4910 => x"00",
          4911 => x"00",
          4912 => x"63",
          4913 => x"63",
          4914 => x"00",
          4915 => x"69",
          4916 => x"72",
          4917 => x"6e",
          4918 => x"72",
          4919 => x"6e",
          4920 => x"79",
          4921 => x"6c",
          4922 => x"2e",
          4923 => x"74",
          4924 => x"2e",
          4925 => x"69",
          4926 => x"61",
          4927 => x"63",
          4928 => x"6e",
          4929 => x"69",
          4930 => x"61",
          4931 => x"74",
          4932 => x"69",
          4933 => x"6c",
          4934 => x"69",
          4935 => x"44",
          4936 => x"74",
          4937 => x"63",
          4938 => x"72",
          4939 => x"62",
          4940 => x"6e",
          4941 => x"00",
          4942 => x"6e",
          4943 => x"6c",
          4944 => x"6f",
          4945 => x"69",
          4946 => x"65",
          4947 => x"66",
          4948 => x"20",
          4949 => x"6f",
          4950 => x"6f",
          4951 => x"69",
          4952 => x"6f",
          4953 => x"6e",
          4954 => x"6c",
          4955 => x"69",
          4956 => x"6f",
          4957 => x"6e",
          4958 => x"65",
          4959 => x"72",
          4960 => x"6f",
          4961 => x"6f",
          4962 => x"65",
          4963 => x"61",
          4964 => x"73",
          4965 => x"65",
          4966 => x"75",
          4967 => x"00",
          4968 => x"77",
          4969 => x"2e",
          4970 => x"62",
          4971 => x"20",
          4972 => x"62",
          4973 => x"63",
          4974 => x"65",
          4975 => x"30",
          4976 => x"20",
          4977 => x"00",
          4978 => x"20",
          4979 => x"30",
          4980 => x"20",
          4981 => x"00",
          4982 => x"2a",
          4983 => x"00",
          4984 => x"2f",
          4985 => x"31",
          4986 => x"5a",
          4987 => x"20",
          4988 => x"73",
          4989 => x"0a",
          4990 => x"6e",
          4991 => x"20",
          4992 => x"00",
          4993 => x"20",
          4994 => x"70",
          4995 => x"6e",
          4996 => x"00",
          4997 => x"20",
          4998 => x"72",
          4999 => x"4f",
          5000 => x"69",
          5001 => x"74",
          5002 => x"20",
          5003 => x"72",
          5004 => x"41",
          5005 => x"69",
          5006 => x"74",
          5007 => x"20",
          5008 => x"72",
          5009 => x"41",
          5010 => x"69",
          5011 => x"74",
          5012 => x"6e",
          5013 => x"6d",
          5014 => x"6e",
          5015 => x"74",
          5016 => x"00",
          5017 => x"78",
          5018 => x"00",
          5019 => x"70",
          5020 => x"3a",
          5021 => x"64",
          5022 => x"74",
          5023 => x"73",
          5024 => x"30",
          5025 => x"65",
          5026 => x"61",
          5027 => x"00",
          5028 => x"6c",
          5029 => x"2e",
          5030 => x"6f",
          5031 => x"2e",
          5032 => x"72",
          5033 => x"00",
          5034 => x"28",
          5035 => x"25",
          5036 => x"38",
          5037 => x"75",
          5038 => x"72",
          5039 => x"6c",
          5040 => x"30",
          5041 => x"58",
          5042 => x"30",
          5043 => x"58",
          5044 => x"20",
          5045 => x"00",
          5046 => x"74",
          5047 => x"65",
          5048 => x"78",
          5049 => x"61",
          5050 => x"6f",
          5051 => x"38",
          5052 => x"00",
          5053 => x"72",
          5054 => x"20",
          5055 => x"64",
          5056 => x"65",
          5057 => x"67",
          5058 => x"61",
          5059 => x"00",
          5060 => x"72",
          5061 => x"67",
          5062 => x"50",
          5063 => x"64",
          5064 => x"2e",
          5065 => x"64",
          5066 => x"00",
          5067 => x"73",
          5068 => x"6f",
          5069 => x"00",
          5070 => x"79",
          5071 => x"74",
          5072 => x"6e",
          5073 => x"65",
          5074 => x"61",
          5075 => x"75",
          5076 => x"2e",
          5077 => x"69",
          5078 => x"72",
          5079 => x"2e",
          5080 => x"2f",
          5081 => x"64",
          5082 => x"64",
          5083 => x"6f",
          5084 => x"74",
          5085 => x"28",
          5086 => x"43",
          5087 => x"29",
          5088 => x"69",
          5089 => x"6c",
          5090 => x"3a",
          5091 => x"42",
          5092 => x"20",
          5093 => x"30",
          5094 => x"20",
          5095 => x"20",
          5096 => x"38",
          5097 => x"2e",
          5098 => x"4e",
          5099 => x"20",
          5100 => x"30",
          5101 => x"20",
          5102 => x"20",
          5103 => x"38",
          5104 => x"2e",
          5105 => x"41",
          5106 => x"20",
          5107 => x"30",
          5108 => x"20",
          5109 => x"52",
          5110 => x"76",
          5111 => x"30",
          5112 => x"20",
          5113 => x"31",
          5114 => x"6d",
          5115 => x"30",
          5116 => x"20",
          5117 => x"43",
          5118 => x"61",
          5119 => x"30",
          5120 => x"20",
          5121 => x"4f",
          5122 => x"00",
          5123 => x"42",
          5124 => x"20",
          5125 => x"00",
          5126 => x"53",
          5127 => x"50",
          5128 => x"73",
          5129 => x"20",
          5130 => x"65",
          5131 => x"74",
          5132 => x"65",
          5133 => x"38",
          5134 => x"20",
          5135 => x"65",
          5136 => x"61",
          5137 => x"65",
          5138 => x"38",
          5139 => x"20",
          5140 => x"20",
          5141 => x"64",
          5142 => x"20",
          5143 => x"38",
          5144 => x"69",
          5145 => x"20",
          5146 => x"64",
          5147 => x"20",
          5148 => x"20",
          5149 => x"34",
          5150 => x"20",
          5151 => x"6d",
          5152 => x"46",
          5153 => x"20",
          5154 => x"2e",
          5155 => x"0a",
          5156 => x"44",
          5157 => x"63",
          5158 => x"20",
          5159 => x"3d",
          5160 => x"64",
          5161 => x"20",
          5162 => x"6f",
          5163 => x"4d",
          5164 => x"46",
          5165 => x"2e",
          5166 => x"0a",
          5167 => x"00",
          5168 => x"6d",
          5169 => x"00",
          5170 => x"56",
          5171 => x"6e",
          5172 => x"00",
          5173 => x"00",
          5174 => x"00",
          5175 => x"00",
          5176 => x"00",
          5177 => x"00",
          5178 => x"00",
          5179 => x"00",
          5180 => x"00",
          5181 => x"00",
          5182 => x"00",
          5183 => x"00",
          5184 => x"00",
          5185 => x"00",
          5186 => x"00",
          5187 => x"00",
          5188 => x"00",
          5189 => x"00",
          5190 => x"00",
          5191 => x"00",
          5192 => x"00",
          5193 => x"00",
          5194 => x"00",
          5195 => x"00",
          5196 => x"00",
          5197 => x"00",
          5198 => x"00",
          5199 => x"00",
          5200 => x"00",
          5201 => x"00",
          5202 => x"00",
          5203 => x"00",
          5204 => x"00",
          5205 => x"5b",
          5206 => x"5b",
          5207 => x"5b",
          5208 => x"5b",
          5209 => x"5b",
          5210 => x"5b",
          5211 => x"00",
          5212 => x"00",
          5213 => x"00",
          5214 => x"00",
          5215 => x"00",
          5216 => x"69",
          5217 => x"69",
          5218 => x"00",
          5219 => x"20",
          5220 => x"61",
          5221 => x"20",
          5222 => x"68",
          5223 => x"72",
          5224 => x"74",
          5225 => x"00",
          5226 => x"74",
          5227 => x"72",
          5228 => x"73",
          5229 => x"6c",
          5230 => x"62",
          5231 => x"44",
          5232 => x"3f",
          5233 => x"2c",
          5234 => x"41",
          5235 => x"00",
          5236 => x"44",
          5237 => x"4f",
          5238 => x"20",
          5239 => x"20",
          5240 => x"4d",
          5241 => x"54",
          5242 => x"00",
          5243 => x"00",
          5244 => x"03",
          5245 => x"16",
          5246 => x"9a",
          5247 => x"45",
          5248 => x"92",
          5249 => x"99",
          5250 => x"49",
          5251 => x"a9",
          5252 => x"b1",
          5253 => x"b9",
          5254 => x"c1",
          5255 => x"c9",
          5256 => x"d1",
          5257 => x"d9",
          5258 => x"e1",
          5259 => x"e9",
          5260 => x"f1",
          5261 => x"f9",
          5262 => x"2e",
          5263 => x"22",
          5264 => x"00",
          5265 => x"10",
          5266 => x"00",
          5267 => x"04",
          5268 => x"00",
          5269 => x"e9",
          5270 => x"e5",
          5271 => x"e8",
          5272 => x"c4",
          5273 => x"c6",
          5274 => x"fb",
          5275 => x"dc",
          5276 => x"a7",
          5277 => x"f3",
          5278 => x"aa",
          5279 => x"ac",
          5280 => x"ab",
          5281 => x"93",
          5282 => x"62",
          5283 => x"51",
          5284 => x"5b",
          5285 => x"2c",
          5286 => x"5e",
          5287 => x"69",
          5288 => x"6c",
          5289 => x"65",
          5290 => x"53",
          5291 => x"0c",
          5292 => x"90",
          5293 => x"93",
          5294 => x"b5",
          5295 => x"a9",
          5296 => x"b5",
          5297 => x"65",
          5298 => x"f7",
          5299 => x"b7",
          5300 => x"a0",
          5301 => x"e0",
          5302 => x"ff",
          5303 => x"30",
          5304 => x"10",
          5305 => x"06",
          5306 => x"81",
          5307 => x"84",
          5308 => x"89",
          5309 => x"8d",
          5310 => x"91",
          5311 => x"f6",
          5312 => x"98",
          5313 => x"9d",
          5314 => x"a0",
          5315 => x"a4",
          5316 => x"a9",
          5317 => x"ac",
          5318 => x"b1",
          5319 => x"b5",
          5320 => x"b8",
          5321 => x"bc",
          5322 => x"c1",
          5323 => x"c5",
          5324 => x"c7",
          5325 => x"cd",
          5326 => x"8e",
          5327 => x"03",
          5328 => x"f8",
          5329 => x"3a",
          5330 => x"3b",
          5331 => x"40",
          5332 => x"0a",
          5333 => x"86",
          5334 => x"58",
          5335 => x"5c",
          5336 => x"93",
          5337 => x"64",
          5338 => x"97",
          5339 => x"6c",
          5340 => x"70",
          5341 => x"74",
          5342 => x"78",
          5343 => x"7c",
          5344 => x"a6",
          5345 => x"84",
          5346 => x"ae",
          5347 => x"45",
          5348 => x"90",
          5349 => x"03",
          5350 => x"ac",
          5351 => x"89",
          5352 => x"c2",
          5353 => x"c4",
          5354 => x"8c",
          5355 => x"18",
          5356 => x"f3",
          5357 => x"f7",
          5358 => x"fa",
          5359 => x"10",
          5360 => x"36",
          5361 => x"01",
          5362 => x"61",
          5363 => x"7d",
          5364 => x"96",
          5365 => x"08",
          5366 => x"08",
          5367 => x"06",
          5368 => x"52",
          5369 => x"56",
          5370 => x"70",
          5371 => x"c8",
          5372 => x"da",
          5373 => x"ea",
          5374 => x"80",
          5375 => x"a0",
          5376 => x"b8",
          5377 => x"cc",
          5378 => x"02",
          5379 => x"01",
          5380 => x"fc",
          5381 => x"70",
          5382 => x"83",
          5383 => x"2f",
          5384 => x"06",
          5385 => x"64",
          5386 => x"1a",
          5387 => x"00",
          5388 => x"00",
          5389 => x"00",
          5390 => x"00",
          5391 => x"00",
          5392 => x"00",
          5393 => x"00",
          5394 => x"00",
          5395 => x"00",
          5396 => x"00",
          5397 => x"00",
          5398 => x"00",
          5399 => x"00",
          5400 => x"00",
          5401 => x"00",
          5402 => x"00",
          5403 => x"00",
          5404 => x"00",
          5405 => x"00",
          5406 => x"00",
          5407 => x"00",
          5408 => x"00",
          5409 => x"00",
          5410 => x"00",
          5411 => x"00",
          5412 => x"00",
          5413 => x"00",
          5414 => x"00",
          5415 => x"00",
          5416 => x"00",
          5417 => x"00",
          5418 => x"00",
          5419 => x"00",
          5420 => x"00",
          5421 => x"00",
          5422 => x"00",
          5423 => x"00",
          5424 => x"00",
          5425 => x"00",
          5426 => x"00",
          5427 => x"00",
          5428 => x"00",
          5429 => x"00",
          5430 => x"00",
          5431 => x"00",
          5432 => x"00",
          5433 => x"00",
          5434 => x"00",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"81",
          5444 => x"7f",
          5445 => x"00",
          5446 => x"00",
          5447 => x"f5",
          5448 => x"00",
          5449 => x"01",
          5450 => x"00",
          5451 => x"00",
          5452 => x"00",
          5453 => x"00",
          5454 => x"00",
          5455 => x"00",
          5456 => x"00",
          5457 => x"00",
          5458 => x"00",
          5459 => x"00",
          5460 => x"00",
          5461 => x"00",
          5462 => x"00",
          5463 => x"00",
          5464 => x"00",
          5465 => x"00",
          5466 => x"00",
          5467 => x"03",
          5468 => x"03",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"9d",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"9f",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"8b",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b3",
           136 => x"0b",
           137 => x"0b",
           138 => x"f0",
           139 => x"0b",
           140 => x"0b",
           141 => x"ad",
           142 => x"0b",
           143 => x"0b",
           144 => x"ed",
           145 => x"0b",
           146 => x"0b",
           147 => x"ad",
           148 => x"0b",
           149 => x"0b",
           150 => x"ed",
           151 => x"0b",
           152 => x"0b",
           153 => x"ad",
           154 => x"0b",
           155 => x"0b",
           156 => x"ed",
           157 => x"0b",
           158 => x"0b",
           159 => x"ad",
           160 => x"0b",
           161 => x"0b",
           162 => x"ed",
           163 => x"0b",
           164 => x"0b",
           165 => x"ad",
           166 => x"0b",
           167 => x"0b",
           168 => x"ed",
           169 => x"0b",
           170 => x"0b",
           171 => x"ad",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"04",
           195 => x"82",
           196 => x"82",
           197 => x"d5",
           198 => x"d5",
           199 => x"f0",
           200 => x"f0",
           201 => x"08",
           202 => x"0c",
           203 => x"84",
           204 => x"80",
           205 => x"84",
           206 => x"80",
           207 => x"84",
           208 => x"93",
           209 => x"80",
           210 => x"c0",
           211 => x"90",
           212 => x"2d",
           213 => x"04",
           214 => x"2d",
           215 => x"04",
           216 => x"2d",
           217 => x"04",
           218 => x"2d",
           219 => x"04",
           220 => x"2d",
           221 => x"04",
           222 => x"2d",
           223 => x"04",
           224 => x"2d",
           225 => x"04",
           226 => x"2d",
           227 => x"04",
           228 => x"2d",
           229 => x"04",
           230 => x"2d",
           231 => x"04",
           232 => x"2d",
           233 => x"04",
           234 => x"2d",
           235 => x"04",
           236 => x"2d",
           237 => x"04",
           238 => x"2d",
           239 => x"04",
           240 => x"2d",
           241 => x"04",
           242 => x"2d",
           243 => x"04",
           244 => x"2d",
           245 => x"04",
           246 => x"2d",
           247 => x"04",
           248 => x"2d",
           249 => x"04",
           250 => x"2d",
           251 => x"04",
           252 => x"2d",
           253 => x"04",
           254 => x"2d",
           255 => x"04",
           256 => x"2d",
           257 => x"04",
           258 => x"2d",
           259 => x"04",
           260 => x"2d",
           261 => x"04",
           262 => x"2d",
           263 => x"04",
           264 => x"2d",
           265 => x"04",
           266 => x"2d",
           267 => x"04",
           268 => x"2d",
           269 => x"04",
           270 => x"2d",
           271 => x"04",
           272 => x"2d",
           273 => x"04",
           274 => x"2d",
           275 => x"04",
           276 => x"2d",
           277 => x"04",
           278 => x"2d",
           279 => x"04",
           280 => x"2d",
           281 => x"04",
           282 => x"2d",
           283 => x"04",
           284 => x"2d",
           285 => x"04",
           286 => x"2d",
           287 => x"04",
           288 => x"2d",
           289 => x"04",
           290 => x"2d",
           291 => x"04",
           292 => x"2d",
           293 => x"04",
           294 => x"2d",
           295 => x"04",
           296 => x"2d",
           297 => x"04",
           298 => x"2d",
           299 => x"04",
           300 => x"10",
           301 => x"10",
           302 => x"10",
           303 => x"10",
           304 => x"00",
           305 => x"09",
           306 => x"2b",
           307 => x"04",
           308 => x"05",
           309 => x"72",
           310 => x"51",
           311 => x"70",
           312 => x"71",
           313 => x"0b",
           314 => x"f0",
           315 => x"02",
           316 => x"82",
           317 => x"d5",
           318 => x"f0",
           319 => x"f0",
           320 => x"c8",
           321 => x"d5",
           322 => x"f8",
           323 => x"05",
           324 => x"54",
           325 => x"04",
           326 => x"f0",
           327 => x"08",
           328 => x"81",
           329 => x"52",
           330 => x"f0",
           331 => x"8d",
           332 => x"f4",
           333 => x"f0",
           334 => x"d5",
           335 => x"82",
           336 => x"d5",
           337 => x"f0",
           338 => x"08",
           339 => x"38",
           340 => x"05",
           341 => x"f0",
           342 => x"3f",
           343 => x"f0",
           344 => x"f0",
           345 => x"81",
           346 => x"f0",
           347 => x"82",
           348 => x"d5",
           349 => x"71",
           350 => x"05",
           351 => x"8c",
           352 => x"05",
           353 => x"fc",
           354 => x"f0",
           355 => x"34",
           356 => x"70",
           357 => x"52",
           358 => x"82",
           359 => x"d5",
           360 => x"02",
           361 => x"86",
           362 => x"34",
           363 => x"82",
           364 => x"0a",
           365 => x"0c",
           366 => x"82",
           367 => x"d5",
           368 => x"d5",
           369 => x"d5",
           370 => x"54",
           371 => x"70",
           372 => x"82",
           373 => x"d5",
           374 => x"54",
           375 => x"dc",
           376 => x"54",
           377 => x"04",
           378 => x"f0",
           379 => x"08",
           380 => x"fc",
           381 => x"05",
           382 => x"05",
           383 => x"05",
           384 => x"e4",
           385 => x"05",
           386 => x"08",
           387 => x"87",
           388 => x"82",
           389 => x"0c",
           390 => x"f0",
           391 => x"08",
           392 => x"14",
           393 => x"08",
           394 => x"81",
           395 => x"51",
           396 => x"0b",
           397 => x"96",
           398 => x"05",
           399 => x"d5",
           400 => x"ff",
           401 => x"38",
           402 => x"81",
           403 => x"0c",
           404 => x"70",
           405 => x"95",
           406 => x"05",
           407 => x"38",
           408 => x"53",
           409 => x"d5",
           410 => x"b0",
           411 => x"82",
           412 => x"98",
           413 => x"72",
           414 => x"05",
           415 => x"70",
           416 => x"80",
           417 => x"e4",
           418 => x"53",
           419 => x"23",
           420 => x"e8",
           421 => x"2c",
           422 => x"11",
           423 => x"72",
           424 => x"82",
           425 => x"82",
           426 => x"15",
           427 => x"d5",
           428 => x"f0",
           429 => x"70",
           430 => x"25",
           431 => x"f0",
           432 => x"08",
           433 => x"81",
           434 => x"38",
           435 => x"70",
           436 => x"2c",
           437 => x"53",
           438 => x"23",
           439 => x"e4",
           440 => x"06",
           441 => x"38",
           442 => x"70",
           443 => x"53",
           444 => x"f0",
           445 => x"08",
           446 => x"f0",
           447 => x"f0",
           448 => x"92",
           449 => x"05",
           450 => x"11",
           451 => x"04",
           452 => x"70",
           453 => x"f0",
           454 => x"08",
           455 => x"53",
           456 => x"23",
           457 => x"e4",
           458 => x"53",
           459 => x"23",
           460 => x"e4",
           461 => x"53",
           462 => x"23",
           463 => x"e4",
           464 => x"72",
           465 => x"80",
           466 => x"34",
           467 => x"e4",
           468 => x"72",
           469 => x"fb",
           470 => x"08",
           471 => x"ec",
           472 => x"82",
           473 => x"e3",
           474 => x"34",
           475 => x"90",
           476 => x"05",
           477 => x"90",
           478 => x"82",
           479 => x"d5",
           480 => x"51",
           481 => x"05",
           482 => x"08",
           483 => x"90",
           484 => x"08",
           485 => x"f0",
           486 => x"08",
           487 => x"81",
           488 => x"2e",
           489 => x"05",
           490 => x"2c",
           491 => x"08",
           492 => x"e4",
           493 => x"f4",
           494 => x"08",
           495 => x"82",
           496 => x"f0",
           497 => x"08",
           498 => x"08",
           499 => x"54",
           500 => x"23",
           501 => x"90",
           502 => x"05",
           503 => x"90",
           504 => x"08",
           505 => x"e4",
           506 => x"06",
           507 => x"ab",
           508 => x"33",
           509 => x"53",
           510 => x"52",
           511 => x"08",
           512 => x"05",
           513 => x"fc",
           514 => x"d5",
           515 => x"08",
           516 => x"ec",
           517 => x"f4",
           518 => x"72",
           519 => x"8a",
           520 => x"05",
           521 => x"51",
           522 => x"82",
           523 => x"d5",
           524 => x"82",
           525 => x"08",
           526 => x"53",
           527 => x"05",
           528 => x"08",
           529 => x"05",
           530 => x"dc",
           531 => x"dc",
           532 => x"05",
           533 => x"08",
           534 => x"08",
           535 => x"53",
           536 => x"23",
           537 => x"30",
           538 => x"82",
           539 => x"ff",
           540 => x"f0",
           541 => x"88",
           542 => x"23",
           543 => x"05",
           544 => x"72",
           545 => x"80",
           546 => x"05",
           547 => x"f4",
           548 => x"05",
           549 => x"51",
           550 => x"82",
           551 => x"d5",
           552 => x"82",
           553 => x"08",
           554 => x"53",
           555 => x"05",
           556 => x"08",
           557 => x"05",
           558 => x"d8",
           559 => x"d8",
           560 => x"05",
           561 => x"22",
           562 => x"d5",
           563 => x"f4",
           564 => x"0c",
           565 => x"82",
           566 => x"d5",
           567 => x"70",
           568 => x"82",
           569 => x"82",
           570 => x"d5",
           571 => x"f0",
           572 => x"53",
           573 => x"f0",
           574 => x"54",
           575 => x"70",
           576 => x"82",
           577 => x"39",
           578 => x"53",
           579 => x"82",
           580 => x"d5",
           581 => x"d5",
           582 => x"82",
           583 => x"05",
           584 => x"82",
           585 => x"53",
           586 => x"52",
           587 => x"08",
           588 => x"0c",
           589 => x"08",
           590 => x"82",
           591 => x"d5",
           592 => x"75",
           593 => x"08",
           594 => x"e4",
           595 => x"72",
           596 => x"08",
           597 => x"72",
           598 => x"82",
           599 => x"86",
           600 => x"72",
           601 => x"f0",
           602 => x"82",
           603 => x"d5",
           604 => x"82",
           605 => x"d5",
           606 => x"72",
           607 => x"82",
           608 => x"05",
           609 => x"05",
           610 => x"cc",
           611 => x"d5",
           612 => x"f0",
           613 => x"08",
           614 => x"e4",
           615 => x"06",
           616 => x"d0",
           617 => x"33",
           618 => x"d5",
           619 => x"51",
           620 => x"d5",
           621 => x"06",
           622 => x"e4",
           623 => x"08",
           624 => x"08",
           625 => x"54",
           626 => x"34",
           627 => x"70",
           628 => x"53",
           629 => x"f0",
           630 => x"70",
           631 => x"2c",
           632 => x"82",
           633 => x"75",
           634 => x"08",
           635 => x"f0",
           636 => x"70",
           637 => x"2c",
           638 => x"82",
           639 => x"75",
           640 => x"08",
           641 => x"e4",
           642 => x"53",
           643 => x"ec",
           644 => x"82",
           645 => x"90",
           646 => x"73",
           647 => x"88",
           648 => x"3f",
           649 => x"05",
           650 => x"51",
           651 => x"82",
           652 => x"ad",
           653 => x"82",
           654 => x"84",
           655 => x"72",
           656 => x"08",
           657 => x"a5",
           658 => x"e4",
           659 => x"06",
           660 => x"38",
           661 => x"52",
           662 => x"f0",
           663 => x"70",
           664 => x"2e",
           665 => x"05",
           666 => x"82",
           667 => x"72",
           668 => x"82",
           669 => x"82",
           670 => x"89",
           671 => x"05",
           672 => x"51",
           673 => x"82",
           674 => x"11",
           675 => x"ec",
           676 => x"2c",
           677 => x"82",
           678 => x"b0",
           679 => x"d5",
           680 => x"2a",
           681 => x"80",
           682 => x"e8",
           683 => x"82",
           684 => x"98",
           685 => x"73",
           686 => x"88",
           687 => x"3f",
           688 => x"05",
           689 => x"51",
           690 => x"f0",
           691 => x"54",
           692 => x"23",
           693 => x"53",
           694 => x"f0",
           695 => x"87",
           696 => x"08",
           697 => x"2e",
           698 => x"f0",
           699 => x"f0",
           700 => x"3f",
           701 => x"f8",
           702 => x"09",
           703 => x"f0",
           704 => x"53",
           705 => x"23",
           706 => x"83",
           707 => x"d5",
           708 => x"d5",
           709 => x"52",
           710 => x"81",
           711 => x"0c",
           712 => x"82",
           713 => x"72",
           714 => x"cb",
           715 => x"22",
           716 => x"f0",
           717 => x"ff",
           718 => x"80",
           719 => x"05",
           720 => x"05",
           721 => x"3f",
           722 => x"81",
           723 => x"0c",
           724 => x"f0",
           725 => x"38",
           726 => x"52",
           727 => x"ff",
           728 => x"0c",
           729 => x"70",
           730 => x"39",
           731 => x"70",
           732 => x"53",
           733 => x"d5",
           734 => x"54",
           735 => x"05",
           736 => x"51",
           737 => x"d5",
           738 => x"51",
           739 => x"f0",
           740 => x"f0",
           741 => x"3f",
           742 => x"05",
           743 => x"08",
           744 => x"09",
           745 => x"d5",
           746 => x"82",
           747 => x"0b",
           748 => x"8a",
           749 => x"23",
           750 => x"88",
           751 => x"f8",
           752 => x"ea",
           753 => x"08",
           754 => x"08",
           755 => x"f0",
           756 => x"0c",
           757 => x"04",
           758 => x"f0",
           759 => x"08",
           760 => x"08",
           761 => x"08",
           762 => x"08",
           763 => x"3d",
           764 => x"d5",
           765 => x"fb",
           766 => x"08",
           767 => x"85",
           768 => x"32",
           769 => x"53",
           770 => x"82",
           771 => x"92",
           772 => x"08",
           773 => x"88",
           774 => x"08",
           775 => x"f0",
           776 => x"06",
           777 => x"f1",
           778 => x"82",
           779 => x"90",
           780 => x"d5",
           781 => x"b1",
           782 => x"f8",
           783 => x"c8",
           784 => x"8a",
           785 => x"82",
           786 => x"8a",
           787 => x"f8",
           788 => x"05",
           789 => x"05",
           790 => x"05",
           791 => x"0d",
           792 => x"f0",
           793 => x"3d",
           794 => x"f8",
           795 => x"05",
           796 => x"70",
           797 => x"51",
           798 => x"ff",
           799 => x"0c",
           800 => x"88",
           801 => x"f0",
           802 => x"d5",
           803 => x"82",
           804 => x"81",
           805 => x"38",
           806 => x"82",
           807 => x"82",
           808 => x"90",
           809 => x"d5",
           810 => x"ab",
           811 => x"f8",
           812 => x"f0",
           813 => x"f0",
           814 => x"f0",
           815 => x"0c",
           816 => x"04",
           817 => x"f0",
           818 => x"08",
           819 => x"08",
           820 => x"70",
           821 => x"0d",
           822 => x"f0",
           823 => x"3d",
           824 => x"08",
           825 => x"81",
           826 => x"51",
           827 => x"0b",
           828 => x"81",
           829 => x"05",
           830 => x"70",
           831 => x"80",
           832 => x"08",
           833 => x"8c",
           834 => x"88",
           835 => x"f0",
           836 => x"82",
           837 => x"57",
           838 => x"81",
           839 => x"8c",
           840 => x"8c",
           841 => x"05",
           842 => x"05",
           843 => x"d5",
           844 => x"f0",
           845 => x"f0",
           846 => x"06",
           847 => x"72",
           848 => x"a3",
           849 => x"08",
           850 => x"0c",
           851 => x"70",
           852 => x"51",
           853 => x"f0",
           854 => x"08",
           855 => x"87",
           856 => x"82",
           857 => x"0c",
           858 => x"88",
           859 => x"32",
           860 => x"71",
           861 => x"d5",
           862 => x"39",
           863 => x"85",
           864 => x"06",
           865 => x"80",
           866 => x"05",
           867 => x"08",
           868 => x"bf",
           869 => x"82",
           870 => x"11",
           871 => x"d5",
           872 => x"33",
           873 => x"0c",
           874 => x"d5",
           875 => x"33",
           876 => x"51",
           877 => x"38",
           878 => x"70",
           879 => x"fc",
           880 => x"08",
           881 => x"f0",
           882 => x"08",
           883 => x"33",
           884 => x"14",
           885 => x"f8",
           886 => x"f0",
           887 => x"05",
           888 => x"d5",
           889 => x"f0",
           890 => x"08",
           891 => x"08",
           892 => x"0c",
           893 => x"08",
           894 => x"f0",
           895 => x"08",
           896 => x"88",
           897 => x"f0",
           898 => x"f0",
           899 => x"81",
           900 => x"f0",
           901 => x"d5",
           902 => x"82",
           903 => x"07",
           904 => x"05",
           905 => x"08",
           906 => x"33",
           907 => x"f0",
           908 => x"d5",
           909 => x"08",
           910 => x"f0",
           911 => x"06",
           912 => x"0c",
           913 => x"f8",
           914 => x"3d",
           915 => x"d5",
           916 => x"fd",
           917 => x"05",
           918 => x"0c",
           919 => x"82",
           920 => x"d5",
           921 => x"82",
           922 => x"05",
           923 => x"08",
           924 => x"08",
           925 => x"90",
           926 => x"08",
           927 => x"38",
           928 => x"82",
           929 => x"82",
           930 => x"d5",
           931 => x"f0",
           932 => x"f0",
           933 => x"08",
           934 => x"f0",
           935 => x"08",
           936 => x"f0",
           937 => x"08",
           938 => x"38",
           939 => x"ff",
           940 => x"0c",
           941 => x"ff",
           942 => x"0c",
           943 => x"82",
           944 => x"51",
           945 => x"82",
           946 => x"05",
           947 => x"82",
           948 => x"05",
           949 => x"82",
           950 => x"2e",
           951 => x"05",
           952 => x"08",
           953 => x"f0",
           954 => x"08",
           955 => x"34",
           956 => x"81",
           957 => x"0c",
           958 => x"88",
           959 => x"51",
           960 => x"04",
           961 => x"f0",
           962 => x"08",
           963 => x"fc",
           964 => x"05",
           965 => x"08",
           966 => x"f0",
           967 => x"06",
           968 => x"da",
           969 => x"08",
           970 => x"05",
           971 => x"08",
           972 => x"31",
           973 => x"3d",
           974 => x"d5",
           975 => x"fe",
           976 => x"05",
           977 => x"0c",
           978 => x"52",
           979 => x"05",
           980 => x"8c",
           981 => x"05",
           982 => x"d5",
           983 => x"82",
           984 => x"81",
           985 => x"38",
           986 => x"88",
           987 => x"51",
           988 => x"04",
           989 => x"f0",
           990 => x"08",
           991 => x"fc",
           992 => x"05",
           993 => x"0c",
           994 => x"80",
           995 => x"08",
           996 => x"f0",
           997 => x"08",
           998 => x"f0",
           999 => x"08",
          1000 => x"82",
          1001 => x"70",
          1002 => x"08",
          1003 => x"05",
          1004 => x"08",
          1005 => x"f0",
          1006 => x"d5",
          1007 => x"39",
          1008 => x"70",
          1009 => x"0d",
          1010 => x"f0",
          1011 => x"3d",
          1012 => x"08",
          1013 => x"f0",
          1014 => x"82",
          1015 => x"05",
          1016 => x"82",
          1017 => x"33",
          1018 => x"51",
          1019 => x"39",
          1020 => x"52",
          1021 => x"05",
          1022 => x"88",
          1023 => x"51",
          1024 => x"f0",
          1025 => x"82",
          1026 => x"05",
          1027 => x"82",
          1028 => x"2e",
          1029 => x"f0",
          1030 => x"e8",
          1031 => x"08",
          1032 => x"ff",
          1033 => x"0c",
          1034 => x"8c",
          1035 => x"08",
          1036 => x"8c",
          1037 => x"8c",
          1038 => x"fc",
          1039 => x"08",
          1040 => x"f0",
          1041 => x"71",
          1042 => x"05",
          1043 => x"39",
          1044 => x"05",
          1045 => x"08",
          1046 => x"82",
          1047 => x"08",
          1048 => x"0d",
          1049 => x"52",
          1050 => x"51",
          1051 => x"70",
          1052 => x"82",
          1053 => x"05",
          1054 => x"3f",
          1055 => x"f0",
          1056 => x"f0",
          1057 => x"0b",
          1058 => x"bc",
          1059 => x"08",
          1060 => x"05",
          1061 => x"08",
          1062 => x"08",
          1063 => x"08",
          1064 => x"82",
          1065 => x"08",
          1066 => x"08",
          1067 => x"88",
          1068 => x"82",
          1069 => x"0c",
          1070 => x"88",
          1071 => x"05",
          1072 => x"08",
          1073 => x"08",
          1074 => x"d5",
          1075 => x"33",
          1076 => x"81",
          1077 => x"0c",
          1078 => x"80",
          1079 => x"8c",
          1080 => x"08",
          1081 => x"8c",
          1082 => x"be",
          1083 => x"08",
          1084 => x"05",
          1085 => x"08",
          1086 => x"31",
          1087 => x"0c",
          1088 => x"08",
          1089 => x"82",
          1090 => x"08",
          1091 => x"0d",
          1092 => x"82",
          1093 => x"d5",
          1094 => x"80",
          1095 => x"05",
          1096 => x"90",
          1097 => x"05",
          1098 => x"90",
          1099 => x"05",
          1100 => x"f0",
          1101 => x"d5",
          1102 => x"71",
          1103 => x"05",
          1104 => x"fc",
          1105 => x"f0",
          1106 => x"e4",
          1107 => x"f0",
          1108 => x"82",
          1109 => x"0b",
          1110 => x"82",
          1111 => x"25",
          1112 => x"05",
          1113 => x"05",
          1114 => x"f4",
          1115 => x"05",
          1116 => x"f0",
          1117 => x"08",
          1118 => x"fc",
          1119 => x"05",
          1120 => x"f0",
          1121 => x"f0",
          1122 => x"d5",
          1123 => x"f0",
          1124 => x"0b",
          1125 => x"82",
          1126 => x"d5",
          1127 => x"82",
          1128 => x"82",
          1129 => x"82",
          1130 => x"82",
          1131 => x"82",
          1132 => x"2e",
          1133 => x"05",
          1134 => x"05",
          1135 => x"08",
          1136 => x"3d",
          1137 => x"d5",
          1138 => x"fb",
          1139 => x"08",
          1140 => x"88",
          1141 => x"d5",
          1142 => x"d5",
          1143 => x"82",
          1144 => x"d5",
          1145 => x"90",
          1146 => x"08",
          1147 => x"0c",
          1148 => x"05",
          1149 => x"05",
          1150 => x"e4",
          1151 => x"05",
          1152 => x"05",
          1153 => x"f0",
          1154 => x"f0",
          1155 => x"08",
          1156 => x"0c",
          1157 => x"0c",
          1158 => x"d5",
          1159 => x"82",
          1160 => x"82",
          1161 => x"80",
          1162 => x"82",
          1163 => x"82",
          1164 => x"08",
          1165 => x"0d",
          1166 => x"05",
          1167 => x"05",
          1168 => x"08",
          1169 => x"3d",
          1170 => x"d5",
          1171 => x"fd",
          1172 => x"08",
          1173 => x"f0",
          1174 => x"08",
          1175 => x"88",
          1176 => x"f0",
          1177 => x"38",
          1178 => x"05",
          1179 => x"08",
          1180 => x"08",
          1181 => x"fc",
          1182 => x"fc",
          1183 => x"f0",
          1184 => x"e1",
          1185 => x"08",
          1186 => x"26",
          1187 => x"05",
          1188 => x"08",
          1189 => x"0c",
          1190 => x"82",
          1191 => x"82",
          1192 => x"d5",
          1193 => x"82",
          1194 => x"d5",
          1195 => x"82",
          1196 => x"95",
          1197 => x"08",
          1198 => x"08",
          1199 => x"08",
          1200 => x"d5",
          1201 => x"d5",
          1202 => x"d5",
          1203 => x"e4",
          1204 => x"0c",
          1205 => x"d5",
          1206 => x"82",
          1207 => x"d5",
          1208 => x"73",
          1209 => x"08",
          1210 => x"72",
          1211 => x"72",
          1212 => x"09",
          1213 => x"08",
          1214 => x"71",
          1215 => x"08",
          1216 => x"09",
          1217 => x"d5",
          1218 => x"f0",
          1219 => x"05",
          1220 => x"33",
          1221 => x"82",
          1222 => x"72",
          1223 => x"38",
          1224 => x"70",
          1225 => x"51",
          1226 => x"f8",
          1227 => x"05",
          1228 => x"0c",
          1229 => x"80",
          1230 => x"08",
          1231 => x"38",
          1232 => x"f0",
          1233 => x"08",
          1234 => x"71",
          1235 => x"82",
          1236 => x"a4",
          1237 => x"f4",
          1238 => x"05",
          1239 => x"70",
          1240 => x"f0",
          1241 => x"82",
          1242 => x"72",
          1243 => x"d5",
          1244 => x"39",
          1245 => x"53",
          1246 => x"f0",
          1247 => x"26",
          1248 => x"d5",
          1249 => x"39",
          1250 => x"05",
          1251 => x"f8",
          1252 => x"38",
          1253 => x"53",
          1254 => x"80",
          1255 => x"0c",
          1256 => x"f0",
          1257 => x"d5",
          1258 => x"f0",
          1259 => x"27",
          1260 => x"f8",
          1261 => x"94",
          1262 => x"33",
          1263 => x"f0",
          1264 => x"08",
          1265 => x"72",
          1266 => x"82",
          1267 => x"90",
          1268 => x"08",
          1269 => x"72",
          1270 => x"82",
          1271 => x"72",
          1272 => x"d5",
          1273 => x"39",
          1274 => x"82",
          1275 => x"54",
          1276 => x"82",
          1277 => x"f7",
          1278 => x"33",
          1279 => x"08",
          1280 => x"33",
          1281 => x"05",
          1282 => x"08",
          1283 => x"08",
          1284 => x"82",
          1285 => x"a5",
          1286 => x"33",
          1287 => x"d5",
          1288 => x"d5",
          1289 => x"f0",
          1290 => x"08",
          1291 => x"0b",
          1292 => x"82",
          1293 => x"d5",
          1294 => x"f0",
          1295 => x"82",
          1296 => x"0b",
          1297 => x"82",
          1298 => x"80",
          1299 => x"05",
          1300 => x"53",
          1301 => x"34",
          1302 => x"2e",
          1303 => x"f0",
          1304 => x"05",
          1305 => x"f0",
          1306 => x"2e",
          1307 => x"82",
          1308 => x"d5",
          1309 => x"81",
          1310 => x"72",
          1311 => x"34",
          1312 => x"53",
          1313 => x"dc",
          1314 => x"08",
          1315 => x"08",
          1316 => x"08",
          1317 => x"f8",
          1318 => x"05",
          1319 => x"08",
          1320 => x"f0",
          1321 => x"84",
          1322 => x"d5",
          1323 => x"f0",
          1324 => x"05",
          1325 => x"33",
          1326 => x"81",
          1327 => x"08",
          1328 => x"88",
          1329 => x"0c",
          1330 => x"d5",
          1331 => x"39",
          1332 => x"53",
          1333 => x"82",
          1334 => x"80",
          1335 => x"33",
          1336 => x"d5",
          1337 => x"b9",
          1338 => x"82",
          1339 => x"d8",
          1340 => x"f4",
          1341 => x"08",
          1342 => x"90",
          1343 => x"33",
          1344 => x"39",
          1345 => x"05",
          1346 => x"d5",
          1347 => x"82",
          1348 => x"d5",
          1349 => x"73",
          1350 => x"08",
          1351 => x"27",
          1352 => x"05",
          1353 => x"d5",
          1354 => x"f0",
          1355 => x"53",
          1356 => x"34",
          1357 => x"53",
          1358 => x"f0",
          1359 => x"53",
          1360 => x"34",
          1361 => x"53",
          1362 => x"82",
          1363 => x"98",
          1364 => x"33",
          1365 => x"54",
          1366 => x"0b",
          1367 => x"80",
          1368 => x"05",
          1369 => x"05",
          1370 => x"05",
          1371 => x"fc",
          1372 => x"05",
          1373 => x"70",
          1374 => x"33",
          1375 => x"fe",
          1376 => x"05",
          1377 => x"82",
          1378 => x"82",
          1379 => x"d5",
          1380 => x"f0",
          1381 => x"81",
          1382 => x"0c",
          1383 => x"82",
          1384 => x"d5",
          1385 => x"70",
          1386 => x"2e",
          1387 => x"79",
          1388 => x"39",
          1389 => x"81",
          1390 => x"39",
          1391 => x"dc",
          1392 => x"3f",
          1393 => x"08",
          1394 => x"e7",
          1395 => x"38",
          1396 => x"ff",
          1397 => x"06",
          1398 => x"ff",
          1399 => x"3d",
          1400 => x"71",
          1401 => x"29",
          1402 => x"04",
          1403 => x"82",
          1404 => x"b3",
          1405 => x"c8",
          1406 => x"51",
          1407 => x"80",
          1408 => x"d6",
          1409 => x"39",
          1410 => x"82",
          1411 => x"b4",
          1412 => x"51",
          1413 => x"39",
          1414 => x"b5",
          1415 => x"51",
          1416 => x"39",
          1417 => x"b6",
          1418 => x"51",
          1419 => x"86",
          1420 => x"0d",
          1421 => x"26",
          1422 => x"29",
          1423 => x"51",
          1424 => x"52",
          1425 => x"e4",
          1426 => x"b6",
          1427 => x"3d",
          1428 => x"84",
          1429 => x"80",
          1430 => x"25",
          1431 => x"87",
          1432 => x"76",
          1433 => x"93",
          1434 => x"76",
          1435 => x"91",
          1436 => x"82",
          1437 => x"e4",
          1438 => x"d5",
          1439 => x"54",
          1440 => x"81",
          1441 => x"57",
          1442 => x"55",
          1443 => x"75",
          1444 => x"d8",
          1445 => x"30",
          1446 => x"70",
          1447 => x"56",
          1448 => x"f4",
          1449 => x"78",
          1450 => x"82",
          1451 => x"f8",
          1452 => x"05",
          1453 => x"7b",
          1454 => x"d5",
          1455 => x"88",
          1456 => x"39",
          1457 => x"54",
          1458 => x"51",
          1459 => x"83",
          1460 => x"0c",
          1461 => x"7f",
          1462 => x"05",
          1463 => x"5c",
          1464 => x"b6",
          1465 => x"b7",
          1466 => x"55",
          1467 => x"90",
          1468 => x"38",
          1469 => x"7a",
          1470 => x"b7",
          1471 => x"39",
          1472 => x"3f",
          1473 => x"18",
          1474 => x"08",
          1475 => x"bb",
          1476 => x"ff",
          1477 => x"39",
          1478 => x"38",
          1479 => x"ff",
          1480 => x"a4",
          1481 => x"55",
          1482 => x"d6",
          1483 => x"a8",
          1484 => x"74",
          1485 => x"70",
          1486 => x"27",
          1487 => x"74",
          1488 => x"06",
          1489 => x"80",
          1490 => x"8a",
          1491 => x"51",
          1492 => x"a0",
          1493 => x"ff",
          1494 => x"ae",
          1495 => x"9d",
          1496 => x"2b",
          1497 => x"2e",
          1498 => x"3f",
          1499 => x"98",
          1500 => x"9b",
          1501 => x"75",
          1502 => x"51",
          1503 => x"9b",
          1504 => x"53",
          1505 => x"26",
          1506 => x"d5",
          1507 => x"3d",
          1508 => x"b0",
          1509 => x"b5",
          1510 => x"a5",
          1511 => x"b7",
          1512 => x"82",
          1513 => x"74",
          1514 => x"86",
          1515 => x"c0",
          1516 => x"81",
          1517 => x"51",
          1518 => x"3f",
          1519 => x"52",
          1520 => x"98",
          1521 => x"c4",
          1522 => x"82",
          1523 => x"80",
          1524 => x"3f",
          1525 => x"80",
          1526 => x"70",
          1527 => x"92",
          1528 => x"b8",
          1529 => x"97",
          1530 => x"06",
          1531 => x"81",
          1532 => x"51",
          1533 => x"3f",
          1534 => x"52",
          1535 => x"97",
          1536 => x"cc",
          1537 => x"86",
          1538 => x"80",
          1539 => x"3f",
          1540 => x"80",
          1541 => x"70",
          1542 => x"92",
          1543 => x"b8",
          1544 => x"96",
          1545 => x"06",
          1546 => x"81",
          1547 => x"51",
          1548 => x"3f",
          1549 => x"fb",
          1550 => x"05",
          1551 => x"75",
          1552 => x"d0",
          1553 => x"53",
          1554 => x"51",
          1555 => x"08",
          1556 => x"80",
          1557 => x"73",
          1558 => x"0b",
          1559 => x"2e",
          1560 => x"f4",
          1561 => x"b8",
          1562 => x"8b",
          1563 => x"86",
          1564 => x"81",
          1565 => x"82",
          1566 => x"d8",
          1567 => x"06",
          1568 => x"52",
          1569 => x"82",
          1570 => x"cd",
          1571 => x"7e",
          1572 => x"7d",
          1573 => x"e4",
          1574 => x"2e",
          1575 => x"59",
          1576 => x"51",
          1577 => x"82",
          1578 => x"82",
          1579 => x"82",
          1580 => x"70",
          1581 => x"b0",
          1582 => x"80",
          1583 => x"b5",
          1584 => x"3f",
          1585 => x"90",
          1586 => x"87",
          1587 => x"38",
          1588 => x"bd",
          1589 => x"ba",
          1590 => x"8a",
          1591 => x"99",
          1592 => x"38",
          1593 => x"bf",
          1594 => x"38",
          1595 => x"80",
          1596 => x"f8",
          1597 => x"78",
          1598 => x"81",
          1599 => x"2e",
          1600 => x"81",
          1601 => x"39",
          1602 => x"84",
          1603 => x"e4",
          1604 => x"3d",
          1605 => x"51",
          1606 => x"80",
          1607 => x"f8",
          1608 => x"b2",
          1609 => x"82",
          1610 => x"51",
          1611 => x"5a",
          1612 => x"59",
          1613 => x"7a",
          1614 => x"b5",
          1615 => x"05",
          1616 => x"08",
          1617 => x"fe",
          1618 => x"eb",
          1619 => x"2e",
          1620 => x"11",
          1621 => x"3f",
          1622 => x"b2",
          1623 => x"9b",
          1624 => x"89",
          1625 => x"5b",
          1626 => x"eb",
          1627 => x"ff",
          1628 => x"d5",
          1629 => x"b5",
          1630 => x"05",
          1631 => x"08",
          1632 => x"fe",
          1633 => x"ea",
          1634 => x"2e",
          1635 => x"ff",
          1636 => x"27",
          1637 => x"5e",
          1638 => x"78",
          1639 => x"52",
          1640 => x"3f",
          1641 => x"d5",
          1642 => x"92",
          1643 => x"ff",
          1644 => x"d5",
          1645 => x"c8",
          1646 => x"82",
          1647 => x"82",
          1648 => x"88",
          1649 => x"39",
          1650 => x"2e",
          1651 => x"ab",
          1652 => x"80",
          1653 => x"45",
          1654 => x"78",
          1655 => x"08",
          1656 => x"fc",
          1657 => x"11",
          1658 => x"3f",
          1659 => x"82",
          1660 => x"89",
          1661 => x"cc",
          1662 => x"80",
          1663 => x"44",
          1664 => x"78",
          1665 => x"08",
          1666 => x"59",
          1667 => x"9c",
          1668 => x"33",
          1669 => x"d4",
          1670 => x"b0",
          1671 => x"f8",
          1672 => x"b2",
          1673 => x"a7",
          1674 => x"2e",
          1675 => x"70",
          1676 => x"7f",
          1677 => x"2e",
          1678 => x"88",
          1679 => x"3f",
          1680 => x"52",
          1681 => x"f8",
          1682 => x"80",
          1683 => x"da",
          1684 => x"f9",
          1685 => x"53",
          1686 => x"82",
          1687 => x"64",
          1688 => x"34",
          1689 => x"fc",
          1690 => x"a2",
          1691 => x"f9",
          1692 => x"82",
          1693 => x"82",
          1694 => x"79",
          1695 => x"79",
          1696 => x"38",
          1697 => x"fe",
          1698 => x"e6",
          1699 => x"2e",
          1700 => x"05",
          1701 => x"ff",
          1702 => x"ae",
          1703 => x"f4",
          1704 => x"e1",
          1705 => x"f8",
          1706 => x"53",
          1707 => x"82",
          1708 => x"61",
          1709 => x"70",
          1710 => x"3d",
          1711 => x"51",
          1712 => x"df",
          1713 => x"54",
          1714 => x"c3",
          1715 => x"f8",
          1716 => x"79",
          1717 => x"f7",
          1718 => x"61",
          1719 => x"fe",
          1720 => x"df",
          1721 => x"2e",
          1722 => x"05",
          1723 => x"78",
          1724 => x"51",
          1725 => x"3d",
          1726 => x"51",
          1727 => x"80",
          1728 => x"f0",
          1729 => x"99",
          1730 => x"a0",
          1731 => x"84",
          1732 => x"53",
          1733 => x"82",
          1734 => x"39",
          1735 => x"a0",
          1736 => x"c4",
          1737 => x"ff",
          1738 => x"59",
          1739 => x"79",
          1740 => x"11",
          1741 => x"3f",
          1742 => x"38",
          1743 => x"05",
          1744 => x"51",
          1745 => x"3d",
          1746 => x"51",
          1747 => x"80",
          1748 => x"bb",
          1749 => x"59",
          1750 => x"53",
          1751 => x"82",
          1752 => x"38",
          1753 => x"a6",
          1754 => x"d5",
          1755 => x"82",
          1756 => x"51",
          1757 => x"82",
          1758 => x"a5",
          1759 => x"a0",
          1760 => x"a8",
          1761 => x"97",
          1762 => x"d2",
          1763 => x"9c",
          1764 => x"d5",
          1765 => x"82",
          1766 => x"84",
          1767 => x"e4",
          1768 => x"80",
          1769 => x"08",
          1770 => x"08",
          1771 => x"7a",
          1772 => x"89",
          1773 => x"ca",
          1774 => x"c2",
          1775 => x"82",
          1776 => x"bc",
          1777 => x"ff",
          1778 => x"b5",
          1779 => x"3f",
          1780 => x"54",
          1781 => x"3d",
          1782 => x"3f",
          1783 => x"bc",
          1784 => x"51",
          1785 => x"58",
          1786 => x"55",
          1787 => x"80",
          1788 => x"51",
          1789 => x"82",
          1790 => x"72",
          1791 => x"80",
          1792 => x"5a",
          1793 => x"8d",
          1794 => x"5c",
          1795 => x"32",
          1796 => x"38",
          1797 => x"38",
          1798 => x"3f",
          1799 => x"39",
          1800 => x"3f",
          1801 => x"0b",
          1802 => x"8c",
          1803 => x"52",
          1804 => x"e4",
          1805 => x"87",
          1806 => x"3f",
          1807 => x"0c",
          1808 => x"55",
          1809 => x"a1",
          1810 => x"75",
          1811 => x"73",
          1812 => x"e4",
          1813 => x"0b",
          1814 => x"83",
          1815 => x"f7",
          1816 => x"02",
          1817 => x"82",
          1818 => x"13",
          1819 => x"0c",
          1820 => x"82",
          1821 => x"82",
          1822 => x"80",
          1823 => x"51",
          1824 => x"04",
          1825 => x"71",
          1826 => x"d5",
          1827 => x"ff",
          1828 => x"38",
          1829 => x"0d",
          1830 => x"54",
          1831 => x"2e",
          1832 => x"a0",
          1833 => x"13",
          1834 => x"a2",
          1835 => x"13",
          1836 => x"2e",
          1837 => x"81",
          1838 => x"70",
          1839 => x"80",
          1840 => x"39",
          1841 => x"54",
          1842 => x"70",
          1843 => x"80",
          1844 => x"09",
          1845 => x"a2",
          1846 => x"07",
          1847 => x"38",
          1848 => x"71",
          1849 => x"e4",
          1850 => x"0d",
          1851 => x"38",
          1852 => x"d7",
          1853 => x"38",
          1854 => x"82",
          1855 => x"fc",
          1856 => x"05",
          1857 => x"81",
          1858 => x"51",
          1859 => x"38",
          1860 => x"97",
          1861 => x"51",
          1862 => x"38",
          1863 => x"bb",
          1864 => x"55",
          1865 => x"d9",
          1866 => x"73",
          1867 => x"0b",
          1868 => x"87",
          1869 => x"87",
          1870 => x"87",
          1871 => x"87",
          1872 => x"87",
          1873 => x"87",
          1874 => x"98",
          1875 => x"0c",
          1876 => x"80",
          1877 => x"3d",
          1878 => x"87",
          1879 => x"87",
          1880 => x"23",
          1881 => x"82",
          1882 => x"5a",
          1883 => x"b0",
          1884 => x"c0",
          1885 => x"34",
          1886 => x"86",
          1887 => x"5c",
          1888 => x"a0",
          1889 => x"7d",
          1890 => x"7b",
          1891 => x"33",
          1892 => x"33",
          1893 => x"33",
          1894 => x"82",
          1895 => x"8f",
          1896 => x"9f",
          1897 => x"81",
          1898 => x"94",
          1899 => x"87",
          1900 => x"96",
          1901 => x"70",
          1902 => x"70",
          1903 => x"72",
          1904 => x"70",
          1905 => x"70",
          1906 => x"38",
          1907 => x"94",
          1908 => x"87",
          1909 => x"74",
          1910 => x"04",
          1911 => x"70",
          1912 => x"70",
          1913 => x"04",
          1914 => x"58",
          1915 => x"38",
          1916 => x"d3",
          1917 => x"56",
          1918 => x"2e",
          1919 => x"72",
          1920 => x"55",
          1921 => x"73",
          1922 => x"72",
          1923 => x"06",
          1924 => x"73",
          1925 => x"72",
          1926 => x"53",
          1927 => x"2e",
          1928 => x"77",
          1929 => x"0c",
          1930 => x"79",
          1931 => x"06",
          1932 => x"fc",
          1933 => x"82",
          1934 => x"59",
          1935 => x"51",
          1936 => x"94",
          1937 => x"70",
          1938 => x"2e",
          1939 => x"06",
          1940 => x"32",
          1941 => x"2e",
          1942 => x"06",
          1943 => x"81",
          1944 => x"52",
          1945 => x"94",
          1946 => x"74",
          1947 => x"57",
          1948 => x"e4",
          1949 => x"0d",
          1950 => x"06",
          1951 => x"72",
          1952 => x"94",
          1953 => x"81",
          1954 => x"e2",
          1955 => x"c0",
          1956 => x"38",
          1957 => x"70",
          1958 => x"51",
          1959 => x"82",
          1960 => x"d5",
          1961 => x"d3",
          1962 => x"53",
          1963 => x"2e",
          1964 => x"71",
          1965 => x"51",
          1966 => x"a0",
          1967 => x"c0",
          1968 => x"38",
          1969 => x"70",
          1970 => x"51",
          1971 => x"0d",
          1972 => x"80",
          1973 => x"51",
          1974 => x"c0",
          1975 => x"87",
          1976 => x"0c",
          1977 => x"88",
          1978 => x"d4",
          1979 => x"82",
          1980 => x"08",
          1981 => x"ac",
          1982 => x"9e",
          1983 => x"c0",
          1984 => x"87",
          1985 => x"0c",
          1986 => x"a8",
          1987 => x"d4",
          1988 => x"82",
          1989 => x"08",
          1990 => x"c0",
          1991 => x"87",
          1992 => x"0c",
          1993 => x"c0",
          1994 => x"80",
          1995 => x"84",
          1996 => x"80",
          1997 => x"d4",
          1998 => x"90",
          1999 => x"52",
          2000 => x"52",
          2001 => x"87",
          2002 => x"0a",
          2003 => x"83",
          2004 => x"34",
          2005 => x"70",
          2006 => x"70",
          2007 => x"82",
          2008 => x"9e",
          2009 => x"51",
          2010 => x"81",
          2011 => x"0b",
          2012 => x"80",
          2013 => x"2e",
          2014 => x"ca",
          2015 => x"08",
          2016 => x"52",
          2017 => x"71",
          2018 => x"c0",
          2019 => x"06",
          2020 => x"38",
          2021 => x"80",
          2022 => x"81",
          2023 => x"80",
          2024 => x"d4",
          2025 => x"90",
          2026 => x"52",
          2027 => x"52",
          2028 => x"87",
          2029 => x"06",
          2030 => x"38",
          2031 => x"87",
          2032 => x"06",
          2033 => x"82",
          2034 => x"9e",
          2035 => x"52",
          2036 => x"52",
          2037 => x"9e",
          2038 => x"84",
          2039 => x"d2",
          2040 => x"08",
          2041 => x"80",
          2042 => x"d4",
          2043 => x"70",
          2044 => x"d4",
          2045 => x"0d",
          2046 => x"3f",
          2047 => x"2e",
          2048 => x"93",
          2049 => x"af",
          2050 => x"73",
          2051 => x"08",
          2052 => x"82",
          2053 => x"82",
          2054 => x"94",
          2055 => x"9c",
          2056 => x"51",
          2057 => x"33",
          2058 => x"d4",
          2059 => x"54",
          2060 => x"f3",
          2061 => x"80",
          2062 => x"82",
          2063 => x"be",
          2064 => x"d4",
          2065 => x"38",
          2066 => x"08",
          2067 => x"ff",
          2068 => x"54",
          2069 => x"d0",
          2070 => x"92",
          2071 => x"73",
          2072 => x"33",
          2073 => x"8b",
          2074 => x"80",
          2075 => x"52",
          2076 => x"3f",
          2077 => x"2e",
          2078 => x"ad",
          2079 => x"73",
          2080 => x"51",
          2081 => x"33",
          2082 => x"c0",
          2083 => x"d4",
          2084 => x"38",
          2085 => x"3f",
          2086 => x"2e",
          2087 => x"ad",
          2088 => x"ad",
          2089 => x"82",
          2090 => x"82",
          2091 => x"51",
          2092 => x"08",
          2093 => x"eb",
          2094 => x"ee",
          2095 => x"c1",
          2096 => x"d4",
          2097 => x"75",
          2098 => x"08",
          2099 => x"54",
          2100 => x"c1",
          2101 => x"d4",
          2102 => x"38",
          2103 => x"c0",
          2104 => x"d5",
          2105 => x"71",
          2106 => x"52",
          2107 => x"3f",
          2108 => x"2e",
          2109 => x"bd",
          2110 => x"3f",
          2111 => x"29",
          2112 => x"e4",
          2113 => x"8f",
          2114 => x"3f",
          2115 => x"02",
          2116 => x"84",
          2117 => x"ad",
          2118 => x"c2",
          2119 => x"51",
          2120 => x"39",
          2121 => x"c3",
          2122 => x"51",
          2123 => x"04",
          2124 => x"87",
          2125 => x"d8",
          2126 => x"fd",
          2127 => x"2c",
          2128 => x"10",
          2129 => x"54",
          2130 => x"12",
          2131 => x"38",
          2132 => x"84",
          2133 => x"52",
          2134 => x"83",
          2135 => x"0c",
          2136 => x"79",
          2137 => x"33",
          2138 => x"38",
          2139 => x"ff",
          2140 => x"52",
          2141 => x"f1",
          2142 => x"bd",
          2143 => x"74",
          2144 => x"39",
          2145 => x"74",
          2146 => x"0d",
          2147 => x"02",
          2148 => x"b4",
          2149 => x"05",
          2150 => x"59",
          2151 => x"9a",
          2152 => x"84",
          2153 => x"70",
          2154 => x"82",
          2155 => x"b4",
          2156 => x"05",
          2157 => x"2e",
          2158 => x"51",
          2159 => x"33",
          2160 => x"34",
          2161 => x"27",
          2162 => x"34",
          2163 => x"b0",
          2164 => x"82",
          2165 => x"8c",
          2166 => x"52",
          2167 => x"d5",
          2168 => x"d4",
          2169 => x"ef",
          2170 => x"3d",
          2171 => x"72",
          2172 => x"71",
          2173 => x"ff",
          2174 => x"25",
          2175 => x"34",
          2176 => x"2e",
          2177 => x"3f",
          2178 => x"3f",
          2179 => x"3d",
          2180 => x"80",
          2181 => x"f5",
          2182 => x"d3",
          2183 => x"f8",
          2184 => x"9f",
          2185 => x"2e",
          2186 => x"3f",
          2187 => x"82",
          2188 => x"d5",
          2189 => x"55",
          2190 => x"81",
          2191 => x"8a",
          2192 => x"06",
          2193 => x"d9",
          2194 => x"08",
          2195 => x"52",
          2196 => x"f0",
          2197 => x"38",
          2198 => x"55",
          2199 => x"56",
          2200 => x"08",
          2201 => x"b2",
          2202 => x"18",
          2203 => x"08",
          2204 => x"ff",
          2205 => x"34",
          2206 => x"9f",
          2207 => x"85",
          2208 => x"b0",
          2209 => x"f4",
          2210 => x"2e",
          2211 => x"89",
          2212 => x"06",
          2213 => x"b2",
          2214 => x"3f",
          2215 => x"08",
          2216 => x"e4",
          2217 => x"0d",
          2218 => x"57",
          2219 => x"81",
          2220 => x"56",
          2221 => x"70",
          2222 => x"73",
          2223 => x"75",
          2224 => x"88",
          2225 => x"52",
          2226 => x"e4",
          2227 => x"ff",
          2228 => x"80",
          2229 => x"81",
          2230 => x"38",
          2231 => x"81",
          2232 => x"f8",
          2233 => x"e4",
          2234 => x"53",
          2235 => x"82",
          2236 => x"74",
          2237 => x"14",
          2238 => x"74",
          2239 => x"82",
          2240 => x"d3",
          2241 => x"08",
          2242 => x"0b",
          2243 => x"82",
          2244 => x"cb",
          2245 => x"55",
          2246 => x"2e",
          2247 => x"55",
          2248 => x"a8",
          2249 => x"08",
          2250 => x"08",
          2251 => x"76",
          2252 => x"de",
          2253 => x"2e",
          2254 => x"a2",
          2255 => x"e4",
          2256 => x"80",
          2257 => x"81",
          2258 => x"56",
          2259 => x"81",
          2260 => x"08",
          2261 => x"e4",
          2262 => x"08",
          2263 => x"ff",
          2264 => x"34",
          2265 => x"75",
          2266 => x"81",
          2267 => x"83",
          2268 => x"81",
          2269 => x"82",
          2270 => x"d5",
          2271 => x"d6",
          2272 => x"82",
          2273 => x"2c",
          2274 => x"78",
          2275 => x"70",
          2276 => x"9c",
          2277 => x"71",
          2278 => x"c3",
          2279 => x"51",
          2280 => x"5d",
          2281 => x"e9",
          2282 => x"81",
          2283 => x"70",
          2284 => x"80",
          2285 => x"51",
          2286 => x"81",
          2287 => x"38",
          2288 => x"b1",
          2289 => x"80",
          2290 => x"ff",
          2291 => x"97",
          2292 => x"f5",
          2293 => x"ff",
          2294 => x"80",
          2295 => x"81",
          2296 => x"74",
          2297 => x"9c",
          2298 => x"70",
          2299 => x"a8",
          2300 => x"58",
          2301 => x"06",
          2302 => x"08",
          2303 => x"34",
          2304 => x"39",
          2305 => x"ed",
          2306 => x"7d",
          2307 => x"e1",
          2308 => x"05",
          2309 => x"33",
          2310 => x"82",
          2311 => x"ab",
          2312 => x"51",
          2313 => x"1a",
          2314 => x"81",
          2315 => x"70",
          2316 => x"51",
          2317 => x"81",
          2318 => x"34",
          2319 => x"34",
          2320 => x"25",
          2321 => x"ed",
          2322 => x"81",
          2323 => x"70",
          2324 => x"51",
          2325 => x"82",
          2326 => x"33",
          2327 => x"81",
          2328 => x"70",
          2329 => x"51",
          2330 => x"ed",
          2331 => x"2c",
          2332 => x"56",
          2333 => x"f1",
          2334 => x"bd",
          2335 => x"80",
          2336 => x"a4",
          2337 => x"de",
          2338 => x"80",
          2339 => x"53",
          2340 => x"9c",
          2341 => x"33",
          2342 => x"80",
          2343 => x"33",
          2344 => x"34",
          2345 => x"34",
          2346 => x"ff",
          2347 => x"70",
          2348 => x"a4",
          2349 => x"25",
          2350 => x"33",
          2351 => x"73",
          2352 => x"81",
          2353 => x"70",
          2354 => x"51",
          2355 => x"f1",
          2356 => x"8d",
          2357 => x"2b",
          2358 => x"57",
          2359 => x"c1",
          2360 => x"51",
          2361 => x"0a",
          2362 => x"2c",
          2363 => x"75",
          2364 => x"82",
          2365 => x"74",
          2366 => x"51",
          2367 => x"52",
          2368 => x"e4",
          2369 => x"38",
          2370 => x"2e",
          2371 => x"51",
          2372 => x"34",
          2373 => x"0b",
          2374 => x"e4",
          2375 => x"a8",
          2376 => x"38",
          2377 => x"ff",
          2378 => x"ff",
          2379 => x"73",
          2380 => x"ed",
          2381 => x"55",
          2382 => x"14",
          2383 => x"98",
          2384 => x"06",
          2385 => x"38",
          2386 => x"34",
          2387 => x"51",
          2388 => x"0a",
          2389 => x"2c",
          2390 => x"75",
          2391 => x"08",
          2392 => x"82",
          2393 => x"98",
          2394 => x"56",
          2395 => x"82",
          2396 => x"9d",
          2397 => x"81",
          2398 => x"ed",
          2399 => x"25",
          2400 => x"a8",
          2401 => x"a4",
          2402 => x"f7",
          2403 => x"81",
          2404 => x"74",
          2405 => x"85",
          2406 => x"ff",
          2407 => x"54",
          2408 => x"39",
          2409 => x"b6",
          2410 => x"82",
          2411 => x"a4",
          2412 => x"82",
          2413 => x"a6",
          2414 => x"82",
          2415 => x"82",
          2416 => x"05",
          2417 => x"d8",
          2418 => x"84",
          2419 => x"08",
          2420 => x"74",
          2421 => x"e4",
          2422 => x"e4",
          2423 => x"74",
          2424 => x"ff",
          2425 => x"55",
          2426 => x"51",
          2427 => x"93",
          2428 => x"d4",
          2429 => x"38",
          2430 => x"d5",
          2431 => x"d5",
          2432 => x"53",
          2433 => x"3f",
          2434 => x"d4",
          2435 => x"80",
          2436 => x"e0",
          2437 => x"a4",
          2438 => x"06",
          2439 => x"ff",
          2440 => x"81",
          2441 => x"ed",
          2442 => x"a8",
          2443 => x"51",
          2444 => x"ed",
          2445 => x"ed",
          2446 => x"27",
          2447 => x"52",
          2448 => x"34",
          2449 => x"9a",
          2450 => x"a8",
          2451 => x"38",
          2452 => x"ff",
          2453 => x"ff",
          2454 => x"f4",
          2455 => x"f4",
          2456 => x"0b",
          2457 => x"53",
          2458 => x"aa",
          2459 => x"80",
          2460 => x"81",
          2461 => x"77",
          2462 => x"82",
          2463 => x"34",
          2464 => x"08",
          2465 => x"80",
          2466 => x"70",
          2467 => x"88",
          2468 => x"d5",
          2469 => x"d4",
          2470 => x"77",
          2471 => x"89",
          2472 => x"52",
          2473 => x"fb",
          2474 => x"ff",
          2475 => x"d5",
          2476 => x"3d",
          2477 => x"05",
          2478 => x"d4",
          2479 => x"83",
          2480 => x"33",
          2481 => x"ae",
          2482 => x"07",
          2483 => x"54",
          2484 => x"77",
          2485 => x"d4",
          2486 => x"70",
          2487 => x"82",
          2488 => x"81",
          2489 => x"83",
          2490 => x"56",
          2491 => x"06",
          2492 => x"82",
          2493 => x"72",
          2494 => x"16",
          2495 => x"34",
          2496 => x"82",
          2497 => x"05",
          2498 => x"11",
          2499 => x"71",
          2500 => x"55",
          2501 => x"13",
          2502 => x"2a",
          2503 => x"34",
          2504 => x"08",
          2505 => x"33",
          2506 => x"56",
          2507 => x"33",
          2508 => x"70",
          2509 => x"86",
          2510 => x"d5",
          2511 => x"33",
          2512 => x"ff",
          2513 => x"53",
          2514 => x"34",
          2515 => x"02",
          2516 => x"71",
          2517 => x"12",
          2518 => x"29",
          2519 => x"98",
          2520 => x"53",
          2521 => x"71",
          2522 => x"fe",
          2523 => x"16",
          2524 => x"2b",
          2525 => x"33",
          2526 => x"70",
          2527 => x"52",
          2528 => x"05",
          2529 => x"13",
          2530 => x"d4",
          2531 => x"33",
          2532 => x"56",
          2533 => x"81",
          2534 => x"81",
          2535 => x"51",
          2536 => x"81",
          2537 => x"3d",
          2538 => x"05",
          2539 => x"11",
          2540 => x"8b",
          2541 => x"59",
          2542 => x"81",
          2543 => x"8c",
          2544 => x"88",
          2545 => x"73",
          2546 => x"d4",
          2547 => x"33",
          2548 => x"56",
          2549 => x"33",
          2550 => x"70",
          2551 => x"82",
          2552 => x"d5",
          2553 => x"12",
          2554 => x"e4",
          2555 => x"f7",
          2556 => x"31",
          2557 => x"70",
          2558 => x"d5",
          2559 => x"82",
          2560 => x"2b",
          2561 => x"33",
          2562 => x"90",
          2563 => x"5b",
          2564 => x"8d",
          2565 => x"fe",
          2566 => x"33",
          2567 => x"83",
          2568 => x"53",
          2569 => x"34",
          2570 => x"14",
          2571 => x"84",
          2572 => x"2b",
          2573 => x"56",
          2574 => x"16",
          2575 => x"80",
          2576 => x"14",
          2577 => x"84",
          2578 => x"d5",
          2579 => x"33",
          2580 => x"80",
          2581 => x"56",
          2582 => x"34",
          2583 => x"73",
          2584 => x"f7",
          2585 => x"71",
          2586 => x"04",
          2587 => x"f8",
          2588 => x"ff",
          2589 => x"11",
          2590 => x"07",
          2591 => x"ff",
          2592 => x"38",
          2593 => x"12",
          2594 => x"ff",
          2595 => x"ff",
          2596 => x"56",
          2597 => x"73",
          2598 => x"5b",
          2599 => x"88",
          2600 => x"78",
          2601 => x"79",
          2602 => x"d5",
          2603 => x"33",
          2604 => x"ff",
          2605 => x"73",
          2606 => x"54",
          2607 => x"54",
          2608 => x"7a",
          2609 => x"51",
          2610 => x"80",
          2611 => x"c6",
          2612 => x"86",
          2613 => x"2b",
          2614 => x"55",
          2615 => x"ff",
          2616 => x"54",
          2617 => x"06",
          2618 => x"d4",
          2619 => x"1e",
          2620 => x"88",
          2621 => x"5e",
          2622 => x"34",
          2623 => x"08",
          2624 => x"33",
          2625 => x"53",
          2626 => x"86",
          2627 => x"d5",
          2628 => x"11",
          2629 => x"07",
          2630 => x"56",
          2631 => x"16",
          2632 => x"05",
          2633 => x"3d",
          2634 => x"82",
          2635 => x"3f",
          2636 => x"71",
          2637 => x"08",
          2638 => x"3d",
          2639 => x"40",
          2640 => x"d4",
          2641 => x"38",
          2642 => x"51",
          2643 => x"54",
          2644 => x"51",
          2645 => x"39",
          2646 => x"e4",
          2647 => x"d4",
          2648 => x"83",
          2649 => x"11",
          2650 => x"2b",
          2651 => x"ff",
          2652 => x"88",
          2653 => x"71",
          2654 => x"44",
          2655 => x"5b",
          2656 => x"25",
          2657 => x"75",
          2658 => x"54",
          2659 => x"88",
          2660 => x"33",
          2661 => x"90",
          2662 => x"54",
          2663 => x"31",
          2664 => x"77",
          2665 => x"54",
          2666 => x"38",
          2667 => x"ff",
          2668 => x"8e",
          2669 => x"51",
          2670 => x"18",
          2671 => x"79",
          2672 => x"71",
          2673 => x"f4",
          2674 => x"3f",
          2675 => x"06",
          2676 => x"82",
          2677 => x"55",
          2678 => x"d4",
          2679 => x"ff",
          2680 => x"15",
          2681 => x"78",
          2682 => x"08",
          2683 => x"71",
          2684 => x"9c",
          2685 => x"3f",
          2686 => x"06",
          2687 => x"82",
          2688 => x"55",
          2689 => x"d4",
          2690 => x"19",
          2691 => x"58",
          2692 => x"b0",
          2693 => x"d5",
          2694 => x"53",
          2695 => x"ff",
          2696 => x"3f",
          2697 => x"80",
          2698 => x"3f",
          2699 => x"08",
          2700 => x"7b",
          2701 => x"3d",
          2702 => x"29",
          2703 => x"d5",
          2704 => x"80",
          2705 => x"82",
          2706 => x"3f",
          2707 => x"0d",
          2708 => x"33",
          2709 => x"38",
          2710 => x"82",
          2711 => x"fc",
          2712 => x"84",
          2713 => x"51",
          2714 => x"84",
          2715 => x"51",
          2716 => x"81",
          2717 => x"92",
          2718 => x"0b",
          2719 => x"71",
          2720 => x"80",
          2721 => x"08",
          2722 => x"80",
          2723 => x"c0",
          2724 => x"87",
          2725 => x"82",
          2726 => x"d5",
          2727 => x"3d",
          2728 => x"bf",
          2729 => x"74",
          2730 => x"e4",
          2731 => x"81",
          2732 => x"87",
          2733 => x"8c",
          2734 => x"5a",
          2735 => x"c0",
          2736 => x"76",
          2737 => x"81",
          2738 => x"8e",
          2739 => x"81",
          2740 => x"74",
          2741 => x"83",
          2742 => x"8f",
          2743 => x"c0",
          2744 => x"87",
          2745 => x"2e",
          2746 => x"38",
          2747 => x"15",
          2748 => x"52",
          2749 => x"39",
          2750 => x"ff",
          2751 => x"90",
          2752 => x"71",
          2753 => x"38",
          2754 => x"80",
          2755 => x"72",
          2756 => x"04",
          2757 => x"8c",
          2758 => x"5b",
          2759 => x"e1",
          2760 => x"79",
          2761 => x"06",
          2762 => x"87",
          2763 => x"8c",
          2764 => x"59",
          2765 => x"98",
          2766 => x"0c",
          2767 => x"70",
          2768 => x"2e",
          2769 => x"33",
          2770 => x"2a",
          2771 => x"2e",
          2772 => x"52",
          2773 => x"08",
          2774 => x"84",
          2775 => x"87",
          2776 => x"70",
          2777 => x"ff",
          2778 => x"81",
          2779 => x"52",
          2780 => x"80",
          2781 => x"7a",
          2782 => x"80",
          2783 => x"81",
          2784 => x"0c",
          2785 => x"7a",
          2786 => x"88",
          2787 => x"56",
          2788 => x"08",
          2789 => x"fe",
          2790 => x"0c",
          2791 => x"38",
          2792 => x"2b",
          2793 => x"71",
          2794 => x"71",
          2795 => x"39",
          2796 => x"06",
          2797 => x"38",
          2798 => x"e8",
          2799 => x"71",
          2800 => x"92",
          2801 => x"06",
          2802 => x"80",
          2803 => x"0c",
          2804 => x"56",
          2805 => x"82",
          2806 => x"fe",
          2807 => x"33",
          2808 => x"0c",
          2809 => x"3d",
          2810 => x"33",
          2811 => x"81",
          2812 => x"75",
          2813 => x"52",
          2814 => x"0d",
          2815 => x"05",
          2816 => x"70",
          2817 => x"51",
          2818 => x"ff",
          2819 => x"72",
          2820 => x"2a",
          2821 => x"34",
          2822 => x"81",
          2823 => x"70",
          2824 => x"3d",
          2825 => x"70",
          2826 => x"05",
          2827 => x"34",
          2828 => x"0d",
          2829 => x"54",
          2830 => x"54",
          2831 => x"84",
          2832 => x"77",
          2833 => x"05",
          2834 => x"33",
          2835 => x"52",
          2836 => x"80",
          2837 => x"0c",
          2838 => x"74",
          2839 => x"2e",
          2840 => x"52",
          2841 => x"e4",
          2842 => x"82",
          2843 => x"77",
          2844 => x"33",
          2845 => x"ff",
          2846 => x"72",
          2847 => x"72",
          2848 => x"e4",
          2849 => x"80",
          2850 => x"55",
          2851 => x"0d",
          2852 => x"0b",
          2853 => x"2e",
          2854 => x"08",
          2855 => x"33",
          2856 => x"e4",
          2857 => x"38",
          2858 => x"b4",
          2859 => x"a0",
          2860 => x"27",
          2861 => x"82",
          2862 => x"54",
          2863 => x"33",
          2864 => x"5a",
          2865 => x"0d",
          2866 => x"56",
          2867 => x"af",
          2868 => x"d5",
          2869 => x"9f",
          2870 => x"52",
          2871 => x"82",
          2872 => x"ff",
          2873 => x"76",
          2874 => x"04",
          2875 => x"fe",
          2876 => x"82",
          2877 => x"33",
          2878 => x"80",
          2879 => x"81",
          2880 => x"84",
          2881 => x"b8",
          2882 => x"82",
          2883 => x"fb",
          2884 => x"52",
          2885 => x"85",
          2886 => x"fb",
          2887 => x"a0",
          2888 => x"08",
          2889 => x"3f",
          2890 => x"19",
          2891 => x"17",
          2892 => x"18",
          2893 => x"33",
          2894 => x"08",
          2895 => x"82",
          2896 => x"fb",
          2897 => x"08",
          2898 => x"74",
          2899 => x"75",
          2900 => x"53",
          2901 => x"0d",
          2902 => x"08",
          2903 => x"df",
          2904 => x"d7",
          2905 => x"82",
          2906 => x"89",
          2907 => x"bf",
          2908 => x"81",
          2909 => x"89",
          2910 => x"52",
          2911 => x"08",
          2912 => x"14",
          2913 => x"2a",
          2914 => x"57",
          2915 => x"e4",
          2916 => x"06",
          2917 => x"78",
          2918 => x"5c",
          2919 => x"38",
          2920 => x"39",
          2921 => x"52",
          2922 => x"e4",
          2923 => x"fe",
          2924 => x"cf",
          2925 => x"ff",
          2926 => x"a8",
          2927 => x"91",
          2928 => x"76",
          2929 => x"b8",
          2930 => x"e4",
          2931 => x"81",
          2932 => x"3d",
          2933 => x"7e",
          2934 => x"27",
          2935 => x"27",
          2936 => x"79",
          2937 => x"89",
          2938 => x"80",
          2939 => x"81",
          2940 => x"89",
          2941 => x"52",
          2942 => x"08",
          2943 => x"38",
          2944 => x"81",
          2945 => x"77",
          2946 => x"84",
          2947 => x"06",
          2948 => x"81",
          2949 => x"a8",
          2950 => x"d9",
          2951 => x"d5",
          2952 => x"ff",
          2953 => x"54",
          2954 => x"74",
          2955 => x"07",
          2956 => x"39",
          2957 => x"52",
          2958 => x"e4",
          2959 => x"d8",
          2960 => x"76",
          2961 => x"05",
          2962 => x"87",
          2963 => x"51",
          2964 => x"59",
          2965 => x"f0",
          2966 => x"06",
          2967 => x"54",
          2968 => x"08",
          2969 => x"51",
          2970 => x"34",
          2971 => x"0d",
          2972 => x"72",
          2973 => x"27",
          2974 => x"9d",
          2975 => x"53",
          2976 => x"82",
          2977 => x"08",
          2978 => x"80",
          2979 => x"82",
          2980 => x"74",
          2981 => x"d5",
          2982 => x"80",
          2983 => x"08",
          2984 => x"08",
          2985 => x"52",
          2986 => x"e4",
          2987 => x"11",
          2988 => x"74",
          2989 => x"0c",
          2990 => x"84",
          2991 => x"ff",
          2992 => x"e4",
          2993 => x"0d",
          2994 => x"79",
          2995 => x"80",
          2996 => x"26",
          2997 => x"52",
          2998 => x"74",
          2999 => x"38",
          3000 => x"e4",
          3001 => x"17",
          3002 => x"c7",
          3003 => x"56",
          3004 => x"77",
          3005 => x"38",
          3006 => x"26",
          3007 => x"51",
          3008 => x"e4",
          3009 => x"38",
          3010 => x"e4",
          3011 => x"80",
          3012 => x"08",
          3013 => x"ef",
          3014 => x"95",
          3015 => x"27",
          3016 => x"89",
          3017 => x"db",
          3018 => x"17",
          3019 => x"75",
          3020 => x"7a",
          3021 => x"08",
          3022 => x"d5",
          3023 => x"86",
          3024 => x"d5",
          3025 => x"07",
          3026 => x"55",
          3027 => x"2e",
          3028 => x"55",
          3029 => x"76",
          3030 => x"08",
          3031 => x"d5",
          3032 => x"55",
          3033 => x"2e",
          3034 => x"51",
          3035 => x"55",
          3036 => x"9c",
          3037 => x"56",
          3038 => x"15",
          3039 => x"07",
          3040 => x"ff",
          3041 => x"39",
          3042 => x"08",
          3043 => x"74",
          3044 => x"04",
          3045 => x"f3",
          3046 => x"81",
          3047 => x"38",
          3048 => x"82",
          3049 => x"b4",
          3050 => x"52",
          3051 => x"3f",
          3052 => x"8a",
          3053 => x"38",
          3054 => x"81",
          3055 => x"d5",
          3056 => x"15",
          3057 => x"07",
          3058 => x"75",
          3059 => x"04",
          3060 => x"58",
          3061 => x"80",
          3062 => x"80",
          3063 => x"17",
          3064 => x"53",
          3065 => x"08",
          3066 => x"53",
          3067 => x"72",
          3068 => x"08",
          3069 => x"16",
          3070 => x"75",
          3071 => x"f5",
          3072 => x"82",
          3073 => x"81",
          3074 => x"38",
          3075 => x"26",
          3076 => x"73",
          3077 => x"51",
          3078 => x"98",
          3079 => x"17",
          3080 => x"9a",
          3081 => x"74",
          3082 => x"83",
          3083 => x"0c",
          3084 => x"8a",
          3085 => x"70",
          3086 => x"57",
          3087 => x"38",
          3088 => x"08",
          3089 => x"cb",
          3090 => x"81",
          3091 => x"94",
          3092 => x"85",
          3093 => x"73",
          3094 => x"8a",
          3095 => x"06",
          3096 => x"73",
          3097 => x"08",
          3098 => x"e4",
          3099 => x"82",
          3100 => x"38",
          3101 => x"26",
          3102 => x"98",
          3103 => x"94",
          3104 => x"3f",
          3105 => x"82",
          3106 => x"38",
          3107 => x"2e",
          3108 => x"08",
          3109 => x"08",
          3110 => x"d5",
          3111 => x"0c",
          3112 => x"82",
          3113 => x"90",
          3114 => x"15",
          3115 => x"0c",
          3116 => x"7b",
          3117 => x"52",
          3118 => x"e4",
          3119 => x"ec",
          3120 => x"17",
          3121 => x"82",
          3122 => x"08",
          3123 => x"9c",
          3124 => x"72",
          3125 => x"38",
          3126 => x"72",
          3127 => x"53",
          3128 => x"56",
          3129 => x"38",
          3130 => x"81",
          3131 => x"d5",
          3132 => x"80",
          3133 => x"09",
          3134 => x"82",
          3135 => x"fd",
          3136 => x"eb",
          3137 => x"ff",
          3138 => x"53",
          3139 => x"38",
          3140 => x"d5",
          3141 => x"72",
          3142 => x"04",
          3143 => x"ff",
          3144 => x"55",
          3145 => x"53",
          3146 => x"38",
          3147 => x"eb",
          3148 => x"3d",
          3149 => x"70",
          3150 => x"74",
          3151 => x"70",
          3152 => x"51",
          3153 => x"e4",
          3154 => x"0d",
          3155 => x"5f",
          3156 => x"19",
          3157 => x"19",
          3158 => x"82",
          3159 => x"08",
          3160 => x"33",
          3161 => x"82",
          3162 => x"70",
          3163 => x"1a",
          3164 => x"81",
          3165 => x"81",
          3166 => x"ae",
          3167 => x"53",
          3168 => x"82",
          3169 => x"56",
          3170 => x"38",
          3171 => x"81",
          3172 => x"2e",
          3173 => x"86",
          3174 => x"80",
          3175 => x"81",
          3176 => x"1d",
          3177 => x"09",
          3178 => x"33",
          3179 => x"81",
          3180 => x"52",
          3181 => x"08",
          3182 => x"f8",
          3183 => x"8d",
          3184 => x"58",
          3185 => x"05",
          3186 => x"08",
          3187 => x"2e",
          3188 => x"c8",
          3189 => x"75",
          3190 => x"75",
          3191 => x"b0",
          3192 => x"c1",
          3193 => x"81",
          3194 => x"8e",
          3195 => x"73",
          3196 => x"1c",
          3197 => x"39",
          3198 => x"7b",
          3199 => x"82",
          3200 => x"72",
          3201 => x"1a",
          3202 => x"f8",
          3203 => x"82",
          3204 => x"08",
          3205 => x"98",
          3206 => x"90",
          3207 => x"70",
          3208 => x"f6",
          3209 => x"82",
          3210 => x"ff",
          3211 => x"0c",
          3212 => x"a9",
          3213 => x"d5",
          3214 => x"08",
          3215 => x"84",
          3216 => x"bf",
          3217 => x"73",
          3218 => x"82",
          3219 => x"06",
          3220 => x"73",
          3221 => x"81",
          3222 => x"70",
          3223 => x"55",
          3224 => x"70",
          3225 => x"92",
          3226 => x"06",
          3227 => x"58",
          3228 => x"06",
          3229 => x"7d",
          3230 => x"38",
          3231 => x"e5",
          3232 => x"ff",
          3233 => x"76",
          3234 => x"05",
          3235 => x"c7",
          3236 => x"8f",
          3237 => x"ff",
          3238 => x"77",
          3239 => x"51",
          3240 => x"08",
          3241 => x"81",
          3242 => x"74",
          3243 => x"06",
          3244 => x"75",
          3245 => x"b3",
          3246 => x"ff",
          3247 => x"70",
          3248 => x"2e",
          3249 => x"77",
          3250 => x"8b",
          3251 => x"51",
          3252 => x"5c",
          3253 => x"f9",
          3254 => x"ff",
          3255 => x"ab",
          3256 => x"38",
          3257 => x"08",
          3258 => x"08",
          3259 => x"ff",
          3260 => x"51",
          3261 => x"58",
          3262 => x"e8",
          3263 => x"3d",
          3264 => x"08",
          3265 => x"5d",
          3266 => x"73",
          3267 => x"5d",
          3268 => x"70",
          3269 => x"f0",
          3270 => x"92",
          3271 => x"3f",
          3272 => x"54",
          3273 => x"c0",
          3274 => x"1c",
          3275 => x"52",
          3276 => x"27",
          3277 => x"70",
          3278 => x"80",
          3279 => x"06",
          3280 => x"81",
          3281 => x"71",
          3282 => x"56",
          3283 => x"84",
          3284 => x"76",
          3285 => x"55",
          3286 => x"57",
          3287 => x"74",
          3288 => x"76",
          3289 => x"2a",
          3290 => x"3d",
          3291 => x"34",
          3292 => x"54",
          3293 => x"70",
          3294 => x"d5",
          3295 => x"17",
          3296 => x"15",
          3297 => x"89",
          3298 => x"d0",
          3299 => x"54",
          3300 => x"56",
          3301 => x"81",
          3302 => x"78",
          3303 => x"51",
          3304 => x"8b",
          3305 => x"27",
          3306 => x"e4",
          3307 => x"08",
          3308 => x"09",
          3309 => x"cb",
          3310 => x"cb",
          3311 => x"06",
          3312 => x"2e",
          3313 => x"fe",
          3314 => x"19",
          3315 => x"3f",
          3316 => x"e4",
          3317 => x"78",
          3318 => x"2b",
          3319 => x"79",
          3320 => x"08",
          3321 => x"38",
          3322 => x"d5",
          3323 => x"1a",
          3324 => x"82",
          3325 => x"08",
          3326 => x"1b",
          3327 => x"5b",
          3328 => x"17",
          3329 => x"34",
          3330 => x"51",
          3331 => x"05",
          3332 => x"2e",
          3333 => x"81",
          3334 => x"c7",
          3335 => x"b9",
          3336 => x"54",
          3337 => x"38",
          3338 => x"74",
          3339 => x"86",
          3340 => x"76",
          3341 => x"52",
          3342 => x"e4",
          3343 => x"c9",
          3344 => x"38",
          3345 => x"81",
          3346 => x"d5",
          3347 => x"d5",
          3348 => x"df",
          3349 => x"9c",
          3350 => x"1a",
          3351 => x"55",
          3352 => x"1d",
          3353 => x"0c",
          3354 => x"78",
          3355 => x"08",
          3356 => x"94",
          3357 => x"3f",
          3358 => x"e4",
          3359 => x"52",
          3360 => x"e4",
          3361 => x"38",
          3362 => x"81",
          3363 => x"77",
          3364 => x"52",
          3365 => x"e4",
          3366 => x"2e",
          3367 => x"06",
          3368 => x"e4",
          3369 => x"0d",
          3370 => x"80",
          3371 => x"80",
          3372 => x"ff",
          3373 => x"7f",
          3374 => x"5b",
          3375 => x"38",
          3376 => x"5b",
          3377 => x"80",
          3378 => x"53",
          3379 => x"5b",
          3380 => x"81",
          3381 => x"b5",
          3382 => x"80",
          3383 => x"83",
          3384 => x"27",
          3385 => x"74",
          3386 => x"97",
          3387 => x"30",
          3388 => x"72",
          3389 => x"80",
          3390 => x"74",
          3391 => x"80",
          3392 => x"70",
          3393 => x"38",
          3394 => x"79",
          3395 => x"05",
          3396 => x"70",
          3397 => x"08",
          3398 => x"53",
          3399 => x"2e",
          3400 => x"55",
          3401 => x"07",
          3402 => x"26",
          3403 => x"ae",
          3404 => x"17",
          3405 => x"34",
          3406 => x"b5",
          3407 => x"0b",
          3408 => x"72",
          3409 => x"0b",
          3410 => x"39",
          3411 => x"57",
          3412 => x"18",
          3413 => x"bf",
          3414 => x"38",
          3415 => x"53",
          3416 => x"2a",
          3417 => x"72",
          3418 => x"38",
          3419 => x"56",
          3420 => x"34",
          3421 => x"33",
          3422 => x"38",
          3423 => x"82",
          3424 => x"33",
          3425 => x"19",
          3426 => x"33",
          3427 => x"11",
          3428 => x"e4",
          3429 => x"87",
          3430 => x"23",
          3431 => x"d5",
          3432 => x"0d",
          3433 => x"41",
          3434 => x"55",
          3435 => x"73",
          3436 => x"2e",
          3437 => x"1f",
          3438 => x"64",
          3439 => x"2e",
          3440 => x"73",
          3441 => x"25",
          3442 => x"38",
          3443 => x"51",
          3444 => x"80",
          3445 => x"51",
          3446 => x"56",
          3447 => x"8c",
          3448 => x"3d",
          3449 => x"d5",
          3450 => x"83",
          3451 => x"27",
          3452 => x"e4",
          3453 => x"23",
          3454 => x"83",
          3455 => x"30",
          3456 => x"51",
          3457 => x"80",
          3458 => x"26",
          3459 => x"51",
          3460 => x"81",
          3461 => x"d7",
          3462 => x"23",
          3463 => x"15",
          3464 => x"57",
          3465 => x"38",
          3466 => x"30",
          3467 => x"54",
          3468 => x"27",
          3469 => x"81",
          3470 => x"ae",
          3471 => x"82",
          3472 => x"82",
          3473 => x"81",
          3474 => x"73",
          3475 => x"78",
          3476 => x"0b",
          3477 => x"78",
          3478 => x"70",
          3479 => x"8a",
          3480 => x"54",
          3481 => x"78",
          3482 => x"fe",
          3483 => x"72",
          3484 => x"51",
          3485 => x"2e",
          3486 => x"59",
          3487 => x"55",
          3488 => x"86",
          3489 => x"57",
          3490 => x"83",
          3491 => x"a0",
          3492 => x"1d",
          3493 => x"5d",
          3494 => x"38",
          3495 => x"ae",
          3496 => x"83",
          3497 => x"79",
          3498 => x"73",
          3499 => x"fe",
          3500 => x"2e",
          3501 => x"55",
          3502 => x"38",
          3503 => x"d5",
          3504 => x"5f",
          3505 => x"5f",
          3506 => x"38",
          3507 => x"32",
          3508 => x"54",
          3509 => x"2e",
          3510 => x"39",
          3511 => x"83",
          3512 => x"30",
          3513 => x"07",
          3514 => x"a6",
          3515 => x"7c",
          3516 => x"57",
          3517 => x"5d",
          3518 => x"fc",
          3519 => x"ff",
          3520 => x"57",
          3521 => x"ae",
          3522 => x"ff",
          3523 => x"51",
          3524 => x"75",
          3525 => x"33",
          3526 => x"38",
          3527 => x"38",
          3528 => x"c0",
          3529 => x"2a",
          3530 => x"58",
          3531 => x"38",
          3532 => x"cc",
          3533 => x"8a",
          3534 => x"56",
          3535 => x"99",
          3536 => x"ff",
          3537 => x"38",
          3538 => x"ff",
          3539 => x"a0",
          3540 => x"58",
          3541 => x"73",
          3542 => x"38",
          3543 => x"2e",
          3544 => x"2b",
          3545 => x"54",
          3546 => x"06",
          3547 => x"85",
          3548 => x"2a",
          3549 => x"38",
          3550 => x"85",
          3551 => x"2a",
          3552 => x"2e",
          3553 => x"ab",
          3554 => x"82",
          3555 => x"56",
          3556 => x"38",
          3557 => x"81",
          3558 => x"70",
          3559 => x"54",
          3560 => x"06",
          3561 => x"ff",
          3562 => x"80",
          3563 => x"bb",
          3564 => x"2a",
          3565 => x"38",
          3566 => x"81",
          3567 => x"e1",
          3568 => x"60",
          3569 => x"ef",
          3570 => x"0c",
          3571 => x"0c",
          3572 => x"7c",
          3573 => x"55",
          3574 => x"81",
          3575 => x"33",
          3576 => x"2e",
          3577 => x"2e",
          3578 => x"33",
          3579 => x"52",
          3580 => x"14",
          3581 => x"52",
          3582 => x"0b",
          3583 => x"7a",
          3584 => x"33",
          3585 => x"9f",
          3586 => x"89",
          3587 => x"54",
          3588 => x"26",
          3589 => x"06",
          3590 => x"51",
          3591 => x"85",
          3592 => x"74",
          3593 => x"9f",
          3594 => x"54",
          3595 => x"15",
          3596 => x"ff",
          3597 => x"86",
          3598 => x"51",
          3599 => x"70",
          3600 => x"04",
          3601 => x"83",
          3602 => x"79",
          3603 => x"55",
          3604 => x"84",
          3605 => x"d5",
          3606 => x"83",
          3607 => x"81",
          3608 => x"17",
          3609 => x"09",
          3610 => x"81",
          3611 => x"79",
          3612 => x"74",
          3613 => x"38",
          3614 => x"ee",
          3615 => x"e4",
          3616 => x"2e",
          3617 => x"52",
          3618 => x"82",
          3619 => x"08",
          3620 => x"82",
          3621 => x"f2",
          3622 => x"cb",
          3623 => x"60",
          3624 => x"08",
          3625 => x"e4",
          3626 => x"e4",
          3627 => x"70",
          3628 => x"2e",
          3629 => x"81",
          3630 => x"80",
          3631 => x"c6",
          3632 => x"ff",
          3633 => x"98",
          3634 => x"74",
          3635 => x"8a",
          3636 => x"39",
          3637 => x"d5",
          3638 => x"52",
          3639 => x"82",
          3640 => x"81",
          3641 => x"cb",
          3642 => x"82",
          3643 => x"56",
          3644 => x"74",
          3645 => x"e4",
          3646 => x"2e",
          3647 => x"38",
          3648 => x"7b",
          3649 => x"56",
          3650 => x"70",
          3651 => x"83",
          3652 => x"d5",
          3653 => x"05",
          3654 => x"56",
          3655 => x"82",
          3656 => x"9f",
          3657 => x"84",
          3658 => x"55",
          3659 => x"7a",
          3660 => x"51",
          3661 => x"81",
          3662 => x"d9",
          3663 => x"09",
          3664 => x"77",
          3665 => x"38",
          3666 => x"76",
          3667 => x"2e",
          3668 => x"26",
          3669 => x"ca",
          3670 => x"ff",
          3671 => x"09",
          3672 => x"14",
          3673 => x"08",
          3674 => x"38",
          3675 => x"82",
          3676 => x"0c",
          3677 => x"80",
          3678 => x"ff",
          3679 => x"81",
          3680 => x"06",
          3681 => x"52",
          3682 => x"80",
          3683 => x"53",
          3684 => x"83",
          3685 => x"87",
          3686 => x"d5",
          3687 => x"06",
          3688 => x"80",
          3689 => x"d5",
          3690 => x"74",
          3691 => x"ee",
          3692 => x"c6",
          3693 => x"e4",
          3694 => x"56",
          3695 => x"14",
          3696 => x"5a",
          3697 => x"8a",
          3698 => x"fe",
          3699 => x"55",
          3700 => x"f3",
          3701 => x"ff",
          3702 => x"74",
          3703 => x"57",
          3704 => x"57",
          3705 => x"82",
          3706 => x"0c",
          3707 => x"a8",
          3708 => x"54",
          3709 => x"af",
          3710 => x"3f",
          3711 => x"06",
          3712 => x"79",
          3713 => x"c7",
          3714 => x"15",
          3715 => x"8d",
          3716 => x"77",
          3717 => x"76",
          3718 => x"70",
          3719 => x"53",
          3720 => x"56",
          3721 => x"38",
          3722 => x"90",
          3723 => x"34",
          3724 => x"92",
          3725 => x"3f",
          3726 => x"06",
          3727 => x"80",
          3728 => x"ca",
          3729 => x"ea",
          3730 => x"34",
          3731 => x"82",
          3732 => x"53",
          3733 => x"06",
          3734 => x"96",
          3735 => x"85",
          3736 => x"38",
          3737 => x"82",
          3738 => x"f2",
          3739 => x"a0",
          3740 => x"e4",
          3741 => x"51",
          3742 => x"90",
          3743 => x"bc",
          3744 => x"bc",
          3745 => x"c4",
          3746 => x"15",
          3747 => x"0c",
          3748 => x"77",
          3749 => x"38",
          3750 => x"38",
          3751 => x"38",
          3752 => x"52",
          3753 => x"38",
          3754 => x"3f",
          3755 => x"71",
          3756 => x"83",
          3757 => x"52",
          3758 => x"0d",
          3759 => x"33",
          3760 => x"56",
          3761 => x"82",
          3762 => x"d5",
          3763 => x"05",
          3764 => x"84",
          3765 => x"80",
          3766 => x"75",
          3767 => x"38",
          3768 => x"05",
          3769 => x"08",
          3770 => x"3d",
          3771 => x"84",
          3772 => x"89",
          3773 => x"77",
          3774 => x"05",
          3775 => x"f6",
          3776 => x"82",
          3777 => x"5c",
          3778 => x"ea",
          3779 => x"82",
          3780 => x"d7",
          3781 => x"73",
          3782 => x"9c",
          3783 => x"38",
          3784 => x"2e",
          3785 => x"df",
          3786 => x"9e",
          3787 => x"54",
          3788 => x"70",
          3789 => x"8e",
          3790 => x"88",
          3791 => x"83",
          3792 => x"80",
          3793 => x"51",
          3794 => x"56",
          3795 => x"05",
          3796 => x"0b",
          3797 => x"7a",
          3798 => x"9c",
          3799 => x"81",
          3800 => x"80",
          3801 => x"54",
          3802 => x"05",
          3803 => x"08",
          3804 => x"38",
          3805 => x"b2",
          3806 => x"06",
          3807 => x"38",
          3808 => x"2a",
          3809 => x"2e",
          3810 => x"80",
          3811 => x"39",
          3812 => x"82",
          3813 => x"12",
          3814 => x"81",
          3815 => x"06",
          3816 => x"77",
          3817 => x"08",
          3818 => x"63",
          3819 => x"82",
          3820 => x"88",
          3821 => x"c0",
          3822 => x"d5",
          3823 => x"0c",
          3824 => x"77",
          3825 => x"34",
          3826 => x"94",
          3827 => x"06",
          3828 => x"38",
          3829 => x"84",
          3830 => x"0c",
          3831 => x"52",
          3832 => x"51",
          3833 => x"57",
          3834 => x"38",
          3835 => x"2e",
          3836 => x"75",
          3837 => x"07",
          3838 => x"8a",
          3839 => x"73",
          3840 => x"a9",
          3841 => x"80",
          3842 => x"c4",
          3843 => x"38",
          3844 => x"82",
          3845 => x"84",
          3846 => x"82",
          3847 => x"f2",
          3848 => x"40",
          3849 => x"fc",
          3850 => x"82",
          3851 => x"08",
          3852 => x"80",
          3853 => x"39",
          3854 => x"56",
          3855 => x"39",
          3856 => x"82",
          3857 => x"81",
          3858 => x"94",
          3859 => x"83",
          3860 => x"8c",
          3861 => x"06",
          3862 => x"8a",
          3863 => x"06",
          3864 => x"38",
          3865 => x"19",
          3866 => x"82",
          3867 => x"ff",
          3868 => x"38",
          3869 => x"52",
          3870 => x"e4",
          3871 => x"d5",
          3872 => x"57",
          3873 => x"1a",
          3874 => x"75",
          3875 => x"58",
          3876 => x"1b",
          3877 => x"d5",
          3878 => x"11",
          3879 => x"38",
          3880 => x"78",
          3881 => x"16",
          3882 => x"2b",
          3883 => x"77",
          3884 => x"1a",
          3885 => x"84",
          3886 => x"27",
          3887 => x"52",
          3888 => x"e4",
          3889 => x"19",
          3890 => x"52",
          3891 => x"76",
          3892 => x"1e",
          3893 => x"5e",
          3894 => x"82",
          3895 => x"f2",
          3896 => x"40",
          3897 => x"fc",
          3898 => x"82",
          3899 => x"08",
          3900 => x"80",
          3901 => x"39",
          3902 => x"81",
          3903 => x"80",
          3904 => x"0b",
          3905 => x"39",
          3906 => x"83",
          3907 => x"56",
          3908 => x"09",
          3909 => x"94",
          3910 => x"56",
          3911 => x"22",
          3912 => x"55",
          3913 => x"18",
          3914 => x"85",
          3915 => x"c6",
          3916 => x"82",
          3917 => x"38",
          3918 => x"ff",
          3919 => x"0c",
          3920 => x"19",
          3921 => x"19",
          3922 => x"74",
          3923 => x"e4",
          3924 => x"52",
          3925 => x"d5",
          3926 => x"82",
          3927 => x"5a",
          3928 => x"78",
          3929 => x"55",
          3930 => x"31",
          3931 => x"81",
          3932 => x"82",
          3933 => x"b4",
          3934 => x"79",
          3935 => x"16",
          3936 => x"52",
          3937 => x"7e",
          3938 => x"89",
          3939 => x"08",
          3940 => x"51",
          3941 => x"08",
          3942 => x"0c",
          3943 => x"08",
          3944 => x"57",
          3945 => x"56",
          3946 => x"bc",
          3947 => x"b0",
          3948 => x"08",
          3949 => x"ff",
          3950 => x"83",
          3951 => x"17",
          3952 => x"18",
          3953 => x"58",
          3954 => x"38",
          3955 => x"89",
          3956 => x"55",
          3957 => x"82",
          3958 => x"f8",
          3959 => x"53",
          3960 => x"d5",
          3961 => x"81",
          3962 => x"2a",
          3963 => x"80",
          3964 => x"52",
          3965 => x"d5",
          3966 => x"80",
          3967 => x"33",
          3968 => x"34",
          3969 => x"08",
          3970 => x"52",
          3971 => x"82",
          3972 => x"ff",
          3973 => x"51",
          3974 => x"0b",
          3975 => x"98",
          3976 => x"33",
          3977 => x"17",
          3978 => x"3d",
          3979 => x"52",
          3980 => x"08",
          3981 => x"86",
          3982 => x"ac",
          3983 => x"d5",
          3984 => x"08",
          3985 => x"86",
          3986 => x"3d",
          3987 => x"0b",
          3988 => x"82",
          3989 => x"80",
          3990 => x"3d",
          3991 => x"94",
          3992 => x"e8",
          3993 => x"82",
          3994 => x"58",
          3995 => x"dc",
          3996 => x"82",
          3997 => x"c7",
          3998 => x"73",
          3999 => x"12",
          4000 => x"33",
          4001 => x"55",
          4002 => x"7f",
          4003 => x"82",
          4004 => x"39",
          4005 => x"81",
          4006 => x"d5",
          4007 => x"a3",
          4008 => x"e1",
          4009 => x"80",
          4010 => x"52",
          4011 => x"82",
          4012 => x"08",
          4013 => x"0c",
          4014 => x"3d",
          4015 => x"54",
          4016 => x"52",
          4017 => x"90",
          4018 => x"d5",
          4019 => x"3d",
          4020 => x"3f",
          4021 => x"e4",
          4022 => x"08",
          4023 => x"d5",
          4024 => x"52",
          4025 => x"e4",
          4026 => x"b3",
          4027 => x"3f",
          4028 => x"e4",
          4029 => x"52",
          4030 => x"d5",
          4031 => x"74",
          4032 => x"08",
          4033 => x"c9",
          4034 => x"86",
          4035 => x"81",
          4036 => x"05",
          4037 => x"93",
          4038 => x"56",
          4039 => x"02",
          4040 => x"16",
          4041 => x"38",
          4042 => x"99",
          4043 => x"16",
          4044 => x"3d",
          4045 => x"58",
          4046 => x"eb",
          4047 => x"11",
          4048 => x"39",
          4049 => x"38",
          4050 => x"55",
          4051 => x"ed",
          4052 => x"d4",
          4053 => x"56",
          4054 => x"81",
          4055 => x"56",
          4056 => x"78",
          4057 => x"27",
          4058 => x"7a",
          4059 => x"55",
          4060 => x"5c",
          4061 => x"85",
          4062 => x"3d",
          4063 => x"33",
          4064 => x"78",
          4065 => x"82",
          4066 => x"04",
          4067 => x"fc",
          4068 => x"fc",
          4069 => x"d5",
          4070 => x"33",
          4071 => x"08",
          4072 => x"15",
          4073 => x"51",
          4074 => x"94",
          4075 => x"0c",
          4076 => x"79",
          4077 => x"51",
          4078 => x"52",
          4079 => x"82",
          4080 => x"70",
          4081 => x"82",
          4082 => x"76",
          4083 => x"0c",
          4084 => x"58",
          4085 => x"54",
          4086 => x"ff",
          4087 => x"54",
          4088 => x"9d",
          4089 => x"81",
          4090 => x"16",
          4091 => x"2e",
          4092 => x"de",
          4093 => x"18",
          4094 => x"81",
          4095 => x"56",
          4096 => x"74",
          4097 => x"e4",
          4098 => x"38",
          4099 => x"73",
          4100 => x"82",
          4101 => x"bf",
          4102 => x"53",
          4103 => x"73",
          4104 => x"15",
          4105 => x"ff",
          4106 => x"73",
          4107 => x"82",
          4108 => x"91",
          4109 => x"81",
          4110 => x"39",
          4111 => x"05",
          4112 => x"08",
          4113 => x"0c",
          4114 => x"72",
          4115 => x"53",
          4116 => x"16",
          4117 => x"0c",
          4118 => x"8b",
          4119 => x"56",
          4120 => x"38",
          4121 => x"8a",
          4122 => x"82",
          4123 => x"08",
          4124 => x"52",
          4125 => x"e4",
          4126 => x"c4",
          4127 => x"55",
          4128 => x"16",
          4129 => x"51",
          4130 => x"9c",
          4131 => x"3f",
          4132 => x"77",
          4133 => x"74",
          4134 => x"82",
          4135 => x"09",
          4136 => x"39",
          4137 => x"0c",
          4138 => x"89",
          4139 => x"87",
          4140 => x"e7",
          4141 => x"38",
          4142 => x"3d",
          4143 => x"89",
          4144 => x"54",
          4145 => x"53",
          4146 => x"74",
          4147 => x"73",
          4148 => x"e4",
          4149 => x"e4",
          4150 => x"82",
          4151 => x"08",
          4152 => x"80",
          4153 => x"a7",
          4154 => x"3f",
          4155 => x"3f",
          4156 => x"30",
          4157 => x"d5",
          4158 => x"72",
          4159 => x"04",
          4160 => x"89",
          4161 => x"de",
          4162 => x"82",
          4163 => x"75",
          4164 => x"08",
          4165 => x"02",
          4166 => x"55",
          4167 => x"55",
          4168 => x"76",
          4169 => x"82",
          4170 => x"f0",
          4171 => x"53",
          4172 => x"51",
          4173 => x"5b",
          4174 => x"7c",
          4175 => x"fe",
          4176 => x"55",
          4177 => x"0c",
          4178 => x"39",
          4179 => x"e4",
          4180 => x"2e",
          4181 => x"75",
          4182 => x"05",
          4183 => x"e4",
          4184 => x"e4",
          4185 => x"e4",
          4186 => x"07",
          4187 => x"53",
          4188 => x"26",
          4189 => x"08",
          4190 => x"98",
          4191 => x"58",
          4192 => x"08",
          4193 => x"38",
          4194 => x"5d",
          4195 => x"81",
          4196 => x"a9",
          4197 => x"ff",
          4198 => x"1b",
          4199 => x"39",
          4200 => x"82",
          4201 => x"30",
          4202 => x"5b",
          4203 => x"58",
          4204 => x"0c",
          4205 => x"33",
          4206 => x"34",
          4207 => x"0d",
          4208 => x"fc",
          4209 => x"3f",
          4210 => x"e4",
          4211 => x"56",
          4212 => x"70",
          4213 => x"55",
          4214 => x"38",
          4215 => x"08",
          4216 => x"82",
          4217 => x"52",
          4218 => x"d5",
          4219 => x"80",
          4220 => x"51",
          4221 => x"08",
          4222 => x"81",
          4223 => x"09",
          4224 => x"39",
          4225 => x"e4",
          4226 => x"98",
          4227 => x"52",
          4228 => x"d5",
          4229 => x"18",
          4230 => x"54",
          4231 => x"85",
          4232 => x"74",
          4233 => x"04",
          4234 => x"ff",
          4235 => x"cf",
          4236 => x"d5",
          4237 => x"a3",
          4238 => x"58",
          4239 => x"55",
          4240 => x"02",
          4241 => x"70",
          4242 => x"73",
          4243 => x"80",
          4244 => x"da",
          4245 => x"87",
          4246 => x"78",
          4247 => x"e4",
          4248 => x"51",
          4249 => x"38",
          4250 => x"15",
          4251 => x"82",
          4252 => x"3d",
          4253 => x"82",
          4254 => x"08",
          4255 => x"52",
          4256 => x"d5",
          4257 => x"86",
          4258 => x"d5",
          4259 => x"d5",
          4260 => x"c7",
          4261 => x"d5",
          4262 => x"08",
          4263 => x"80",
          4264 => x"38",
          4265 => x"af",
          4266 => x"74",
          4267 => x"3f",
          4268 => x"d5",
          4269 => x"3d",
          4270 => x"05",
          4271 => x"82",
          4272 => x"08",
          4273 => x"8e",
          4274 => x"82",
          4275 => x"08",
          4276 => x"82",
          4277 => x"06",
          4278 => x"33",
          4279 => x"86",
          4280 => x"74",
          4281 => x"af",
          4282 => x"55",
          4283 => x"87",
          4284 => x"09",
          4285 => x"d5",
          4286 => x"86",
          4287 => x"81",
          4288 => x"78",
          4289 => x"e4",
          4290 => x"9f",
          4291 => x"51",
          4292 => x"0b",
          4293 => x"80",
          4294 => x"52",
          4295 => x"3f",
          4296 => x"ff",
          4297 => x"11",
          4298 => x"ee",
          4299 => x"15",
          4300 => x"53",
          4301 => x"81",
          4302 => x"bf",
          4303 => x"82",
          4304 => x"b2",
          4305 => x"a3",
          4306 => x"51",
          4307 => x"0b",
          4308 => x"83",
          4309 => x"3f",
          4310 => x"80",
          4311 => x"a1",
          4312 => x"3d",
          4313 => x"84",
          4314 => x"aa",
          4315 => x"51",
          4316 => x"55",
          4317 => x"78",
          4318 => x"70",
          4319 => x"e4",
          4320 => x"be",
          4321 => x"a0",
          4322 => x"38",
          4323 => x"3d",
          4324 => x"3f",
          4325 => x"52",
          4326 => x"08",
          4327 => x"d5",
          4328 => x"97",
          4329 => x"81",
          4330 => x"2e",
          4331 => x"82",
          4332 => x"06",
          4333 => x"92",
          4334 => x"d5",
          4335 => x"93",
          4336 => x"8d",
          4337 => x"af",
          4338 => x"33",
          4339 => x"55",
          4340 => x"54",
          4341 => x"0b",
          4342 => x"84",
          4343 => x"73",
          4344 => x"2e",
          4345 => x"ff",
          4346 => x"52",
          4347 => x"55",
          4348 => x"de",
          4349 => x"51",
          4350 => x"08",
          4351 => x"82",
          4352 => x"16",
          4353 => x"06",
          4354 => x"51",
          4355 => x"0b",
          4356 => x"e4",
          4357 => x"3f",
          4358 => x"e4",
          4359 => x"98",
          4360 => x"82",
          4361 => x"ec",
          4362 => x"02",
          4363 => x"57",
          4364 => x"97",
          4365 => x"e4",
          4366 => x"cf",
          4367 => x"d0",
          4368 => x"e4",
          4369 => x"38",
          4370 => x"06",
          4371 => x"a7",
          4372 => x"71",
          4373 => x"55",
          4374 => x"81",
          4375 => x"a2",
          4376 => x"74",
          4377 => x"04",
          4378 => x"94",
          4379 => x"d0",
          4380 => x"82",
          4381 => x"58",
          4382 => x"c4",
          4383 => x"82",
          4384 => x"c7",
          4385 => x"55",
          4386 => x"17",
          4387 => x"96",
          4388 => x"54",
          4389 => x"ff",
          4390 => x"55",
          4391 => x"0d",
          4392 => x"5a",
          4393 => x"9a",
          4394 => x"e4",
          4395 => x"82",
          4396 => x"55",
          4397 => x"81",
          4398 => x"2e",
          4399 => x"80",
          4400 => x"ac",
          4401 => x"82",
          4402 => x"52",
          4403 => x"d5",
          4404 => x"bf",
          4405 => x"e4",
          4406 => x"81",
          4407 => x"33",
          4408 => x"27",
          4409 => x"80",
          4410 => x"ff",
          4411 => x"56",
          4412 => x"76",
          4413 => x"80",
          4414 => x"78",
          4415 => x"2e",
          4416 => x"38",
          4417 => x"9f",
          4418 => x"82",
          4419 => x"33",
          4420 => x"2e",
          4421 => x"2e",
          4422 => x"05",
          4423 => x"e4",
          4424 => x"0c",
          4425 => x"82",
          4426 => x"9d",
          4427 => x"e4",
          4428 => x"82",
          4429 => x"53",
          4430 => x"ff",
          4431 => x"51",
          4432 => x"38",
          4433 => x"cc",
          4434 => x"ff",
          4435 => x"08",
          4436 => x"82",
          4437 => x"82",
          4438 => x"55",
          4439 => x"82",
          4440 => x"82",
          4441 => x"75",
          4442 => x"38",
          4443 => x"86",
          4444 => x"27",
          4445 => x"77",
          4446 => x"56",
          4447 => x"81",
          4448 => x"73",
          4449 => x"33",
          4450 => x"81",
          4451 => x"02",
          4452 => x"51",
          4453 => x"87",
          4454 => x"78",
          4455 => x"70",
          4456 => x"d5",
          4457 => x"80",
          4458 => x"ae",
          4459 => x"82",
          4460 => x"c4",
          4461 => x"c6",
          4462 => x"09",
          4463 => x"75",
          4464 => x"74",
          4465 => x"e4",
          4466 => x"38",
          4467 => x"66",
          4468 => x"88",
          4469 => x"52",
          4470 => x"54",
          4471 => x"ff",
          4472 => x"54",
          4473 => x"9c",
          4474 => x"62",
          4475 => x"93",
          4476 => x"5e",
          4477 => x"08",
          4478 => x"38",
          4479 => x"38",
          4480 => x"08",
          4481 => x"70",
          4482 => x"55",
          4483 => x"39",
          4484 => x"82",
          4485 => x"89",
          4486 => x"56",
          4487 => x"06",
          4488 => x"82",
          4489 => x"7c",
          4490 => x"27",
          4491 => x"83",
          4492 => x"80",
          4493 => x"c1",
          4494 => x"14",
          4495 => x"82",
          4496 => x"38",
          4497 => x"95",
          4498 => x"81",
          4499 => x"06",
          4500 => x"56",
          4501 => x"b9",
          4502 => x"80",
          4503 => x"7a",
          4504 => x"73",
          4505 => x"ff",
          4506 => x"ff",
          4507 => x"58",
          4508 => x"74",
          4509 => x"73",
          4510 => x"7e",
          4511 => x"2e",
          4512 => x"8c",
          4513 => x"07",
          4514 => x"08",
          4515 => x"75",
          4516 => x"94",
          4517 => x"54",
          4518 => x"82",
          4519 => x"e8",
          4520 => x"80",
          4521 => x"5c",
          4522 => x"0b",
          4523 => x"38",
          4524 => x"ed",
          4525 => x"80",
          4526 => x"d5",
          4527 => x"82",
          4528 => x"12",
          4529 => x"51",
          4530 => x"08",
          4531 => x"57",
          4532 => x"82",
          4533 => x"56",
          4534 => x"05",
          4535 => x"cc",
          4536 => x"68",
          4537 => x"82",
          4538 => x"75",
          4539 => x"81",
          4540 => x"80",
          4541 => x"0a",
          4542 => x"55",
          4543 => x"8b",
          4544 => x"2a",
          4545 => x"59",
          4546 => x"70",
          4547 => x"56",
          4548 => x"80",
          4549 => x"52",
          4550 => x"56",
          4551 => x"83",
          4552 => x"82",
          4553 => x"55",
          4554 => x"09",
          4555 => x"29",
          4556 => x"74",
          4557 => x"17",
          4558 => x"e4",
          4559 => x"92",
          4560 => x"b7",
          4561 => x"52",
          4562 => x"56",
          4563 => x"62",
          4564 => x"e4",
          4565 => x"bf",
          4566 => x"26",
          4567 => x"8e",
          4568 => x"38",
          4569 => x"af",
          4570 => x"56",
          4571 => x"87",
          4572 => x"38",
          4573 => x"83",
          4574 => x"56",
          4575 => x"38",
          4576 => x"06",
          4577 => x"91",
          4578 => x"22",
          4579 => x"74",
          4580 => x"56",
          4581 => x"57",
          4582 => x"75",
          4583 => x"fe",
          4584 => x"84",
          4585 => x"5e",
          4586 => x"e4",
          4587 => x"fd",
          4588 => x"38",
          4589 => x"8c",
          4590 => x"22",
          4591 => x"74",
          4592 => x"56",
          4593 => x"57",
          4594 => x"75",
          4595 => x"fe",
          4596 => x"10",
          4597 => x"9f",
          4598 => x"d5",
          4599 => x"05",
          4600 => x"56",
          4601 => x"81",
          4602 => x"67",
          4603 => x"30",
          4604 => x"59",
          4605 => x"81",
          4606 => x"42",
          4607 => x"90",
          4608 => x"51",
          4609 => x"75",
          4610 => x"67",
          4611 => x"82",
          4612 => x"09",
          4613 => x"08",
          4614 => x"78",
          4615 => x"78",
          4616 => x"82",
          4617 => x"83",
          4618 => x"27",
          4619 => x"55",
          4620 => x"59",
          4621 => x"74",
          4622 => x"88",
          4623 => x"26",
          4624 => x"1a",
          4625 => x"38",
          4626 => x"2e",
          4627 => x"9f",
          4628 => x"06",
          4629 => x"84",
          4630 => x"8f",
          4631 => x"52",
          4632 => x"80",
          4633 => x"3f",
          4634 => x"ff",
          4635 => x"99",
          4636 => x"83",
          4637 => x"80",
          4638 => x"ff",
          4639 => x"ff",
          4640 => x"ff",
          4641 => x"e9",
          4642 => x"51",
          4643 => x"1c",
          4644 => x"8d",
          4645 => x"51",
          4646 => x"1b",
          4647 => x"2e",
          4648 => x"88",
          4649 => x"ff",
          4650 => x"51",
          4651 => x"1b",
          4652 => x"b0",
          4653 => x"52",
          4654 => x"ff",
          4655 => x"0b",
          4656 => x"c7",
          4657 => x"39",
          4658 => x"51",
          4659 => x"ff",
          4660 => x"d1",
          4661 => x"a9",
          4662 => x"c7",
          4663 => x"86",
          4664 => x"1b",
          4665 => x"81",
          4666 => x"ff",
          4667 => x"e4",
          4668 => x"09",
          4669 => x"86",
          4670 => x"88",
          4671 => x"7a",
          4672 => x"85",
          4673 => x"87",
          4674 => x"83",
          4675 => x"ff",
          4676 => x"8b",
          4677 => x"51",
          4678 => x"52",
          4679 => x"54",
          4680 => x"ff",
          4681 => x"53",
          4682 => x"3f",
          4683 => x"8c",
          4684 => x"83",
          4685 => x"52",
          4686 => x"52",
          4687 => x"f0",
          4688 => x"87",
          4689 => x"83",
          4690 => x"ff",
          4691 => x"74",
          4692 => x"54",
          4693 => x"86",
          4694 => x"be",
          4695 => x"08",
          4696 => x"76",
          4697 => x"cd",
          4698 => x"ff",
          4699 => x"83",
          4700 => x"26",
          4701 => x"53",
          4702 => x"3f",
          4703 => x"76",
          4704 => x"db",
          4705 => x"38",
          4706 => x"8a",
          4707 => x"38",
          4708 => x"81",
          4709 => x"ff",
          4710 => x"e4",
          4711 => x"1b",
          4712 => x"54",
          4713 => x"7f",
          4714 => x"39",
          4715 => x"80",
          4716 => x"7a",
          4717 => x"d5",
          4718 => x"83",
          4719 => x"0b",
          4720 => x"34",
          4721 => x"34",
          4722 => x"75",
          4723 => x"85",
          4724 => x"2a",
          4725 => x"82",
          4726 => x"52",
          4727 => x"3f",
          4728 => x"88",
          4729 => x"52",
          4730 => x"56",
          4731 => x"53",
          4732 => x"3f",
          4733 => x"38",
          4734 => x"56",
          4735 => x"75",
          4736 => x"04",
          4737 => x"80",
          4738 => x"76",
          4739 => x"11",
          4740 => x"79",
          4741 => x"09",
          4742 => x"55",
          4743 => x"70",
          4744 => x"74",
          4745 => x"80",
          4746 => x"76",
          4747 => x"3d",
          4748 => x"84",
          4749 => x"8a",
          4750 => x"52",
          4751 => x"56",
          4752 => x"08",
          4753 => x"75",
          4754 => x"a1",
          4755 => x"53",
          4756 => x"97",
          4757 => x"72",
          4758 => x"56",
          4759 => x"88",
          4760 => x"3d",
          4761 => x"80",
          4762 => x"05",
          4763 => x"08",
          4764 => x"08",
          4765 => x"09",
          4766 => x"55",
          4767 => x"e4",
          4768 => x"0d",
          4769 => x"73",
          4770 => x"0c",
          4771 => x"02",
          4772 => x"3d",
          4773 => x"52",
          4774 => x"ff",
          4775 => x"3d",
          4776 => x"22",
          4777 => x"26",
          4778 => x"52",
          4779 => x"27",
          4780 => x"06",
          4781 => x"82",
          4782 => x"9c",
          4783 => x"06",
          4784 => x"38",
          4785 => x"22",
          4786 => x"70",
          4787 => x"d5",
          4788 => x"3d",
          4789 => x"05",
          4790 => x"70",
          4791 => x"9a",
          4792 => x"06",
          4793 => x"38",
          4794 => x"22",
          4795 => x"84",
          4796 => x"51",
          4797 => x"38",
          4798 => x"a8",
          4799 => x"38",
          4800 => x"05",
          4801 => x"72",
          4802 => x"80",
          4803 => x"22",
          4804 => x"70",
          4805 => x"25",
          4806 => x"dc",
          4807 => x"05",
          4808 => x"10",
          4809 => x"80",
          4810 => x"72",
          4811 => x"12",
          4812 => x"39",
          4813 => x"51",
          4814 => x"ff",
          4815 => x"12",
          4816 => x"8c",
          4817 => x"16",
          4818 => x"82",
          4819 => x"00",
          4820 => x"ff",
          4821 => x"00",
          4822 => x"00",
          4823 => x"00",
          4824 => x"00",
          4825 => x"00",
          4826 => x"00",
          4827 => x"00",
          4828 => x"00",
          4829 => x"00",
          4830 => x"00",
          4831 => x"00",
          4832 => x"00",
          4833 => x"00",
          4834 => x"00",
          4835 => x"00",
          4836 => x"00",
          4837 => x"00",
          4838 => x"00",
          4839 => x"00",
          4840 => x"00",
          4841 => x"00",
          4842 => x"00",
          4843 => x"00",
          4844 => x"00",
          4845 => x"00",
          4846 => x"00",
          4847 => x"00",
          4848 => x"00",
          4849 => x"00",
          4850 => x"00",
          4851 => x"00",
          4852 => x"00",
          4853 => x"00",
          4854 => x"00",
          4855 => x"00",
          4856 => x"00",
          4857 => x"00",
          4858 => x"00",
          4859 => x"00",
          4860 => x"00",
          4861 => x"00",
          4862 => x"00",
          4863 => x"00",
          4864 => x"00",
          4865 => x"00",
          4866 => x"00",
          4867 => x"00",
          4868 => x"00",
          4869 => x"00",
          4870 => x"00",
          4871 => x"00",
          4872 => x"00",
          4873 => x"00",
          4874 => x"00",
          4875 => x"00",
          4876 => x"00",
          4877 => x"00",
          4878 => x"00",
          4879 => x"00",
          4880 => x"00",
          4881 => x"00",
          4882 => x"00",
          4883 => x"00",
          4884 => x"00",
          4885 => x"00",
          4886 => x"00",
          4887 => x"00",
          4888 => x"00",
          4889 => x"00",
          4890 => x"00",
          4891 => x"00",
          4892 => x"00",
          4893 => x"00",
          4894 => x"74",
          4895 => x"74",
          4896 => x"74",
          4897 => x"64",
          4898 => x"63",
          4899 => x"61",
          4900 => x"79",
          4901 => x"66",
          4902 => x"70",
          4903 => x"6d",
          4904 => x"68",
          4905 => x"68",
          4906 => x"63",
          4907 => x"6a",
          4908 => x"61",
          4909 => x"74",
          4910 => x"00",
          4911 => x"00",
          4912 => x"69",
          4913 => x"69",
          4914 => x"00",
          4915 => x"44",
          4916 => x"6f",
          4917 => x"72",
          4918 => x"6f",
          4919 => x"20",
          4920 => x"64",
          4921 => x"69",
          4922 => x"64",
          4923 => x"61",
          4924 => x"64",
          4925 => x"6c",
          4926 => x"6e",
          4927 => x"41",
          4928 => x"65",
          4929 => x"46",
          4930 => x"65",
          4931 => x"73",
          4932 => x"46",
          4933 => x"64",
          4934 => x"6c",
          4935 => x"53",
          4936 => x"69",
          4937 => x"65",
          4938 => x"44",
          4939 => x"6d",
          4940 => x"69",
          4941 => x"00",
          4942 => x"20",
          4943 => x"62",
          4944 => x"4e",
          4945 => x"74",
          4946 => x"6c",
          4947 => x"20",
          4948 => x"6e",
          4949 => x"46",
          4950 => x"62",
          4951 => x"54",
          4952 => x"20",
          4953 => x"6f",
          4954 => x"6c",
          4955 => x"46",
          4956 => x"6c",
          4957 => x"49",
          4958 => x"69",
          4959 => x"6f",
          4960 => x"54",
          4961 => x"20",
          4962 => x"6c",
          4963 => x"50",
          4964 => x"72",
          4965 => x"72",
          4966 => x"53",
          4967 => x"00",
          4968 => x"6f",
          4969 => x"72",
          4970 => x"20",
          4971 => x"73",
          4972 => x"20",
          4973 => x"65",
          4974 => x"72",
          4975 => x"25",
          4976 => x"3a",
          4977 => x"00",
          4978 => x"20",
          4979 => x"25",
          4980 => x"20",
          4981 => x"7c",
          4982 => x"0a",
          4983 => x"00",
          4984 => x"32",
          4985 => x"76",
          4986 => x"20",
          4987 => x"76",
          4988 => x"25",
          4989 => x"0a",
          4990 => x"49",
          4991 => x"74",
          4992 => x"72",
          4993 => x"72",
          4994 => x"75",
          4995 => x"69",
          4996 => x"74",
          4997 => x"4c",
          4998 => x"65",
          4999 => x"49",
          5000 => x"20",
          5001 => x"70",
          5002 => x"30",
          5003 => x"65",
          5004 => x"55",
          5005 => x"20",
          5006 => x"70",
          5007 => x"31",
          5008 => x"65",
          5009 => x"55",
          5010 => x"20",
          5011 => x"70",
          5012 => x"69",
          5013 => x"69",
          5014 => x"45",
          5015 => x"20",
          5016 => x"2e",
          5017 => x"65",
          5018 => x"00",
          5019 => x"7a",
          5020 => x"30",
          5021 => x"65",
          5022 => x"69",
          5023 => x"20",
          5024 => x"20",
          5025 => x"73",
          5026 => x"6d",
          5027 => x"2e",
          5028 => x"43",
          5029 => x"2e",
          5030 => x"43",
          5031 => x"2e",
          5032 => x"61",
          5033 => x"00",
          5034 => x"78",
          5035 => x"3e",
          5036 => x"30",
          5037 => x"44",
          5038 => x"6f",
          5039 => x"70",
          5040 => x"25",
          5041 => x"32",
          5042 => x"25",
          5043 => x"34",
          5044 => x"58",
          5045 => x"00",
          5046 => x"75",
          5047 => x"64",
          5048 => x"6c",
          5049 => x"43",
          5050 => x"63",
          5051 => x"30",
          5052 => x"0a",
          5053 => x"20",
          5054 => x"64",
          5055 => x"25",
          5056 => x"52",
          5057 => x"6e",
          5058 => x"63",
          5059 => x"2e",
          5060 => x"20",
          5061 => x"6e",
          5062 => x"5a",
          5063 => x"25",
          5064 => x"73",
          5065 => x"25",
          5066 => x"73",
          5067 => x"25",
          5068 => x"63",
          5069 => x"00",
          5070 => x"72",
          5071 => x"73",
          5072 => x"6e",
          5073 => x"63",
          5074 => x"6d",
          5075 => x"52",
          5076 => x"2e",
          5077 => x"6c",
          5078 => x"65",
          5079 => x"2e",
          5080 => x"64",
          5081 => x"25",
          5082 => x"25",
          5083 => x"43",
          5084 => x"61",
          5085 => x"20",
          5086 => x"6f",
          5087 => x"67",
          5088 => x"76",
          5089 => x"70",
          5090 => x"64",
          5091 => x"57",
          5092 => x"20",
          5093 => x"25",
          5094 => x"20",
          5095 => x"4d",
          5096 => x"30",
          5097 => x"29",
          5098 => x"49",
          5099 => x"4d",
          5100 => x"25",
          5101 => x"20",
          5102 => x"20",
          5103 => x"30",
          5104 => x"29",
          5105 => x"52",
          5106 => x"20",
          5107 => x"25",
          5108 => x"20",
          5109 => x"41",
          5110 => x"65",
          5111 => x"25",
          5112 => x"20",
          5113 => x"52",
          5114 => x"69",
          5115 => x"25",
          5116 => x"20",
          5117 => x"20",
          5118 => x"68",
          5119 => x"25",
          5120 => x"20",
          5121 => x"42",
          5122 => x"00",
          5123 => x"57",
          5124 => x"20",
          5125 => x"4c",
          5126 => x"50",
          5127 => x"53",
          5128 => x"65",
          5129 => x"20",
          5130 => x"52",
          5131 => x"63",
          5132 => x"72",
          5133 => x"30",
          5134 => x"20",
          5135 => x"4d",
          5136 => x"74",
          5137 => x"72",
          5138 => x"30",
          5139 => x"20",
          5140 => x"6b",
          5141 => x"41",
          5142 => x"20",
          5143 => x"30",
          5144 => x"4d",
          5145 => x"20",
          5146 => x"49",
          5147 => x"20",
          5148 => x"20",
          5149 => x"30",
          5150 => x"20",
          5151 => x"65",
          5152 => x"20",
          5153 => x"20",
          5154 => x"64",
          5155 => x"7a",
          5156 => x"53",
          5157 => x"6f",
          5158 => x"20",
          5159 => x"20",
          5160 => x"34",
          5161 => x"20",
          5162 => x"62",
          5163 => x"41",
          5164 => x"20",
          5165 => x"64",
          5166 => x"7a",
          5167 => x"6c",
          5168 => x"75",
          5169 => x"00",
          5170 => x"45",
          5171 => x"55",
          5172 => x"00",
          5173 => x"00",
          5174 => x"01",
          5175 => x"00",
          5176 => x"00",
          5177 => x"01",
          5178 => x"00",
          5179 => x"00",
          5180 => x"01",
          5181 => x"00",
          5182 => x"00",
          5183 => x"01",
          5184 => x"00",
          5185 => x"00",
          5186 => x"01",
          5187 => x"00",
          5188 => x"00",
          5189 => x"04",
          5190 => x"00",
          5191 => x"00",
          5192 => x"04",
          5193 => x"00",
          5194 => x"00",
          5195 => x"04",
          5196 => x"00",
          5197 => x"00",
          5198 => x"04",
          5199 => x"00",
          5200 => x"00",
          5201 => x"03",
          5202 => x"00",
          5203 => x"00",
          5204 => x"03",
          5205 => x"1b",
          5206 => x"1b",
          5207 => x"1b",
          5208 => x"1b",
          5209 => x"1b",
          5210 => x"1b",
          5211 => x"0e",
          5212 => x"0b",
          5213 => x"06",
          5214 => x"04",
          5215 => x"02",
          5216 => x"68",
          5217 => x"68",
          5218 => x"21",
          5219 => x"75",
          5220 => x"46",
          5221 => x"6f",
          5222 => x"74",
          5223 => x"6f",
          5224 => x"20",
          5225 => x"00",
          5226 => x"6f",
          5227 => x"63",
          5228 => x"69",
          5229 => x"69",
          5230 => x"61",
          5231 => x"53",
          5232 => x"3e",
          5233 => x"2b",
          5234 => x"46",
          5235 => x"32",
          5236 => x"53",
          5237 => x"4e",
          5238 => x"20",
          5239 => x"20",
          5240 => x"41",
          5241 => x"41",
          5242 => x"00",
          5243 => x"00",
          5244 => x"01",
          5245 => x"14",
          5246 => x"80",
          5247 => x"45",
          5248 => x"90",
          5249 => x"59",
          5250 => x"41",
          5251 => x"a8",
          5252 => x"b0",
          5253 => x"b8",
          5254 => x"c0",
          5255 => x"c8",
          5256 => x"d0",
          5257 => x"d8",
          5258 => x"e0",
          5259 => x"e8",
          5260 => x"f0",
          5261 => x"f8",
          5262 => x"2b",
          5263 => x"5c",
          5264 => x"7f",
          5265 => x"00",
          5266 => x"00",
          5267 => x"00",
          5268 => x"00",
          5269 => x"00",
          5270 => x"00",
          5271 => x"00",
          5272 => x"00",
          5273 => x"00",
          5274 => x"00",
          5275 => x"00",
          5276 => x"20",
          5277 => x"00",
          5278 => x"00",
          5279 => x"00",
          5280 => x"00",
          5281 => x"25",
          5282 => x"25",
          5283 => x"25",
          5284 => x"25",
          5285 => x"25",
          5286 => x"25",
          5287 => x"25",
          5288 => x"25",
          5289 => x"25",
          5290 => x"25",
          5291 => x"25",
          5292 => x"25",
          5293 => x"03",
          5294 => x"00",
          5295 => x"03",
          5296 => x"03",
          5297 => x"22",
          5298 => x"00",
          5299 => x"00",
          5300 => x"25",
          5301 => x"00",
          5302 => x"00",
          5303 => x"01",
          5304 => x"01",
          5305 => x"01",
          5306 => x"01",
          5307 => x"01",
          5308 => x"01",
          5309 => x"01",
          5310 => x"01",
          5311 => x"01",
          5312 => x"01",
          5313 => x"01",
          5314 => x"01",
          5315 => x"01",
          5316 => x"01",
          5317 => x"01",
          5318 => x"01",
          5319 => x"01",
          5320 => x"01",
          5321 => x"01",
          5322 => x"01",
          5323 => x"01",
          5324 => x"01",
          5325 => x"01",
          5326 => x"01",
          5327 => x"00",
          5328 => x"01",
          5329 => x"02",
          5330 => x"02",
          5331 => x"02",
          5332 => x"01",
          5333 => x"01",
          5334 => x"02",
          5335 => x"02",
          5336 => x"01",
          5337 => x"02",
          5338 => x"01",
          5339 => x"02",
          5340 => x"02",
          5341 => x"02",
          5342 => x"02",
          5343 => x"02",
          5344 => x"01",
          5345 => x"02",
          5346 => x"01",
          5347 => x"02",
          5348 => x"02",
          5349 => x"00",
          5350 => x"03",
          5351 => x"03",
          5352 => x"03",
          5353 => x"03",
          5354 => x"03",
          5355 => x"01",
          5356 => x"03",
          5357 => x"03",
          5358 => x"03",
          5359 => x"07",
          5360 => x"01",
          5361 => x"00",
          5362 => x"05",
          5363 => x"1d",
          5364 => x"01",
          5365 => x"06",
          5366 => x"06",
          5367 => x"06",
          5368 => x"1f",
          5369 => x"1f",
          5370 => x"1f",
          5371 => x"1f",
          5372 => x"1f",
          5373 => x"1f",
          5374 => x"1f",
          5375 => x"1f",
          5376 => x"1f",
          5377 => x"1f",
          5378 => x"06",
          5379 => x"00",
          5380 => x"1f",
          5381 => x"21",
          5382 => x"21",
          5383 => x"04",
          5384 => x"01",
          5385 => x"01",
          5386 => x"03",
          5387 => x"00",
          5388 => x"00",
          5389 => x"00",
          5390 => x"00",
          5391 => x"00",
          5392 => x"00",
          5393 => x"00",
          5394 => x"00",
          5395 => x"00",
          5396 => x"00",
          5397 => x"00",
          5398 => x"00",
          5399 => x"00",
          5400 => x"00",
          5401 => x"00",
          5402 => x"00",
          5403 => x"00",
          5404 => x"00",
          5405 => x"00",
          5406 => x"00",
          5407 => x"00",
          5408 => x"00",
          5409 => x"00",
          5410 => x"00",
          5411 => x"00",
          5412 => x"00",
          5413 => x"00",
          5414 => x"00",
          5415 => x"00",
          5416 => x"00",
          5417 => x"00",
          5418 => x"00",
          5419 => x"00",
          5420 => x"00",
          5421 => x"00",
          5422 => x"00",
          5423 => x"00",
          5424 => x"00",
          5425 => x"00",
          5426 => x"00",
          5427 => x"00",
          5428 => x"00",
          5429 => x"00",
          5430 => x"00",
          5431 => x"00",
          5432 => x"00",
          5433 => x"00",
          5434 => x"00",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"00",
          5444 => x"01",
          5445 => x"00",
          5446 => x"00",
          5447 => x"05",
          5448 => x"00",
          5449 => x"01",
          5450 => x"01",
          5451 => x"00",
          5452 => x"00",
          5453 => x"00",
          5454 => x"00",
          5455 => x"00",
          5456 => x"00",
          5457 => x"00",
          5458 => x"00",
          5459 => x"00",
          5460 => x"00",
          5461 => x"00",
          5462 => x"00",
          5463 => x"01",
          5464 => x"01",
          5465 => x"02",
          5466 => x"00",
          5467 => x"00",
          5468 => x"00",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assing the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0'.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
