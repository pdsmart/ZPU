-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87fa",
             1 => x"f80d0b0b",
             2 => x"0b93ed04",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"d1040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b93b4",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b82b7",
           162 => x"ec738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93b90400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80d2",
           171 => x"fe2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80cd",
           179 => x"fc2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"96040b0b",
           269 => x"0b8ca604",
           270 => x"0b0b0b8c",
           271 => x"b6040b0b",
           272 => x"0b8cc604",
           273 => x"0b0b0b8c",
           274 => x"d6040b0b",
           275 => x"0b8ce604",
           276 => x"0b0b0b8c",
           277 => x"f7040b0b",
           278 => x"0b8d8804",
           279 => x"0b0b0b8d",
           280 => x"98040b0b",
           281 => x"0b8da804",
           282 => x"0b0b0b8d",
           283 => x"b8040b0b",
           284 => x"0b8dc904",
           285 => x"0b0b0b8d",
           286 => x"da040b0b",
           287 => x"0b8deb04",
           288 => x"0b0b0b8d",
           289 => x"fc040b0b",
           290 => x"0b8e8d04",
           291 => x"0b0b0b8e",
           292 => x"9e040b0b",
           293 => x"0b8eaf04",
           294 => x"0b0b0b8e",
           295 => x"c0040b0b",
           296 => x"0b8ed104",
           297 => x"0b0b0b8e",
           298 => x"e2040b0b",
           299 => x"0b8ef304",
           300 => x"0b0b0b8f",
           301 => x"84040b0b",
           302 => x"0b8f9504",
           303 => x"0b0b0b8f",
           304 => x"a6040b0b",
           305 => x"0b8fb704",
           306 => x"0b0b0b8f",
           307 => x"c8040b0b",
           308 => x"0b8fd904",
           309 => x"0b0b0b8f",
           310 => x"ea040b0b",
           311 => x"0b8ffb04",
           312 => x"0b0b0b90",
           313 => x"8c040b0b",
           314 => x"0b909d04",
           315 => x"0b0b0b90",
           316 => x"ae040b0b",
           317 => x"0b90bf04",
           318 => x"0b0b0b90",
           319 => x"d0040b0b",
           320 => x"0b90e104",
           321 => x"0b0b0b90",
           322 => x"f2040b0b",
           323 => x"0b918304",
           324 => x"0b0b0b91",
           325 => x"94040b0b",
           326 => x"0b91a504",
           327 => x"0b0b0b91",
           328 => x"b6040b0b",
           329 => x"0b91c704",
           330 => x"0b0b0b91",
           331 => x"d8040b0b",
           332 => x"0b91e904",
           333 => x"0b0b0b91",
           334 => x"fa040b0b",
           335 => x"0b928b04",
           336 => x"0b0b0b92",
           337 => x"9c040b0b",
           338 => x"0b92ad04",
           339 => x"0b0b0b92",
           340 => x"be040b0b",
           341 => x"0b92cf04",
           342 => x"0b0b0b92",
           343 => x"e0040b0b",
           344 => x"0b92f104",
           345 => x"0b0b0b93",
           346 => x"8204ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482e0a4",
           386 => x"0c81818b",
           387 => x"2d82e0a4",
           388 => x"0880c080",
           389 => x"900482e0",
           390 => x"a40cb3e6",
           391 => x"2d82e0a4",
           392 => x"0880c080",
           393 => x"900482e0",
           394 => x"a40cb097",
           395 => x"2d82e0a4",
           396 => x"0880c080",
           397 => x"900482e0",
           398 => x"a40cafe1",
           399 => x"2d82e0a4",
           400 => x"0880c080",
           401 => x"900482e0",
           402 => x"a40c94e1",
           403 => x"2d82e0a4",
           404 => x"0880c080",
           405 => x"900482e0",
           406 => x"a40cb1f6",
           407 => x"2d82e0a4",
           408 => x"0880c080",
           409 => x"900482e0",
           410 => x"a40c80da",
           411 => x"9f2d82e0",
           412 => x"a40880c0",
           413 => x"80900482",
           414 => x"e0a40c80",
           415 => x"d4ce2d82",
           416 => x"e0a40880",
           417 => x"c0809004",
           418 => x"82e0a40c",
           419 => x"948c2d82",
           420 => x"e0a40880",
           421 => x"c0809004",
           422 => x"82e0a40c",
           423 => x"96f42d82",
           424 => x"e0a40880",
           425 => x"c0809004",
           426 => x"82e0a40c",
           427 => x"98812d82",
           428 => x"e0a40880",
           429 => x"c0809004",
           430 => x"82e0a40c",
           431 => x"80e0e72d",
           432 => x"82e0a408",
           433 => x"80c08090",
           434 => x"0482e0a4",
           435 => x"0c80fff6",
           436 => x"2d82e0a4",
           437 => x"0880c080",
           438 => x"900482e0",
           439 => x"a40c8180",
           440 => x"dd2d82e0",
           441 => x"a40880c0",
           442 => x"80900482",
           443 => x"e0a40c80",
           444 => x"fdb22d82",
           445 => x"e0a40880",
           446 => x"c0809004",
           447 => x"82e0a40c",
           448 => x"80fee52d",
           449 => x"82e0a408",
           450 => x"80c08090",
           451 => x"0482e0a4",
           452 => x"0c81f6a7",
           453 => x"2d82e0a4",
           454 => x"0880c080",
           455 => x"900482e0",
           456 => x"a40c8283",
           457 => x"a72d82e0",
           458 => x"a40880c0",
           459 => x"80900482",
           460 => x"e0a40c81",
           461 => x"fb8c2d82",
           462 => x"e0a40880",
           463 => x"c0809004",
           464 => x"82e0a40c",
           465 => x"81fe8c2d",
           466 => x"82e0a408",
           467 => x"80c08090",
           468 => x"0482e0a4",
           469 => x"0c8288e5",
           470 => x"2d82e0a4",
           471 => x"0880c080",
           472 => x"900482e0",
           473 => x"a40c8291",
           474 => x"ce2d82e0",
           475 => x"a40880c0",
           476 => x"80900482",
           477 => x"e0a40c82",
           478 => x"82842d82",
           479 => x"e0a40880",
           480 => x"c0809004",
           481 => x"82e0a40c",
           482 => x"828c882d",
           483 => x"82e0a408",
           484 => x"80c08090",
           485 => x"0482e0a4",
           486 => x"0c828da8",
           487 => x"2d82e0a4",
           488 => x"0880c080",
           489 => x"900482e0",
           490 => x"a40c828d",
           491 => x"c72d82e0",
           492 => x"a40880c0",
           493 => x"80900482",
           494 => x"e0a40c82",
           495 => x"95bb2d82",
           496 => x"e0a40880",
           497 => x"c0809004",
           498 => x"82e0a40c",
           499 => x"82939d2d",
           500 => x"82e0a408",
           501 => x"80c08090",
           502 => x"0482e0a4",
           503 => x"0c829897",
           504 => x"2d82e0a4",
           505 => x"0880c080",
           506 => x"900482e0",
           507 => x"a40c828e",
           508 => x"cd2d82e0",
           509 => x"a40880c0",
           510 => x"80900482",
           511 => x"e0a40c82",
           512 => x"9b9c2d82",
           513 => x"e0a40880",
           514 => x"c0809004",
           515 => x"82e0a40c",
           516 => x"829c9d2d",
           517 => x"82e0a408",
           518 => x"80c08090",
           519 => x"0482e0a4",
           520 => x"0c828487",
           521 => x"2d82e0a4",
           522 => x"0880c080",
           523 => x"900482e0",
           524 => x"a40c8283",
           525 => x"e02d82e0",
           526 => x"a40880c0",
           527 => x"80900482",
           528 => x"e0a40c82",
           529 => x"858b2d82",
           530 => x"e0a40880",
           531 => x"c0809004",
           532 => x"82e0a40c",
           533 => x"828fa42d",
           534 => x"82e0a408",
           535 => x"80c08090",
           536 => x"0482e0a4",
           537 => x"0c829d8e",
           538 => x"2d82e0a4",
           539 => x"0880c080",
           540 => x"900482e0",
           541 => x"a40c829f",
           542 => x"992d82e0",
           543 => x"a40880c0",
           544 => x"80900482",
           545 => x"e0a40c82",
           546 => x"a2a02d82",
           547 => x"e0a40880",
           548 => x"c0809004",
           549 => x"82e0a40c",
           550 => x"81f5c62d",
           551 => x"82e0a408",
           552 => x"80c08090",
           553 => x"0482e0a4",
           554 => x"0c82a58c",
           555 => x"2d82e0a4",
           556 => x"0880c080",
           557 => x"900482e0",
           558 => x"a40c82b4",
           559 => x"e92d82e0",
           560 => x"a40880c0",
           561 => x"80900482",
           562 => x"e0a40c82",
           563 => x"b2d52d82",
           564 => x"e0a40880",
           565 => x"c0809004",
           566 => x"82e0a40c",
           567 => x"81b58b2d",
           568 => x"82e0a408",
           569 => x"80c08090",
           570 => x"0482e0a4",
           571 => x"0c81b6f5",
           572 => x"2d82e0a4",
           573 => x"0880c080",
           574 => x"900482e0",
           575 => x"a40c81b8",
           576 => x"d92d82e0",
           577 => x"a40880c0",
           578 => x"80900482",
           579 => x"e0a40c80",
           580 => x"fbe42d82",
           581 => x"e0a40880",
           582 => x"c0809004",
           583 => x"82e0a40c",
           584 => x"80fd882d",
           585 => x"82e0a408",
           586 => x"80c08090",
           587 => x"0482e0a4",
           588 => x"0c818280",
           589 => x"2d82e0a4",
           590 => x"0880c080",
           591 => x"900482e0",
           592 => x"a40c80e0",
           593 => x"ef2d82e0",
           594 => x"a40880c0",
           595 => x"80900482",
           596 => x"e0a40c81",
           597 => x"af9f2d82",
           598 => x"e0a40880",
           599 => x"c0809004",
           600 => x"82e0a40c",
           601 => x"81afc72d",
           602 => x"82e0a408",
           603 => x"80c08090",
           604 => x"0482e0a4",
           605 => x"0c81b3bf",
           606 => x"2d82e0a4",
           607 => x"0880c080",
           608 => x"900482e0",
           609 => x"a40c81ac",
           610 => x"892d82e0",
           611 => x"a40880c0",
           612 => x"8090043c",
           613 => x"04101010",
           614 => x"10101010",
           615 => x"10101010",
           616 => x"10101010",
           617 => x"10101010",
           618 => x"10101010",
           619 => x"10101010",
           620 => x"10101010",
           621 => x"53510400",
           622 => x"007381ff",
           623 => x"06738306",
           624 => x"09810583",
           625 => x"05101010",
           626 => x"2b0772fc",
           627 => x"060c5151",
           628 => x"04727280",
           629 => x"728106ff",
           630 => x"05097206",
           631 => x"05711052",
           632 => x"720a100a",
           633 => x"5372ed38",
           634 => x"51515351",
           635 => x"0482e098",
           636 => x"7082fc84",
           637 => x"278e3880",
           638 => x"71708405",
           639 => x"530c0b0b",
           640 => x"0b93f004",
           641 => x"8c815180",
           642 => x"faa70400",
           643 => x"82e0a408",
           644 => x"0282e0a4",
           645 => x"0cfb3d0d",
           646 => x"82e0a408",
           647 => x"8c057082",
           648 => x"e0a408fc",
           649 => x"050c82e0",
           650 => x"a408fc05",
           651 => x"085482e0",
           652 => x"a4088805",
           653 => x"085382fb",
           654 => x"fc085254",
           655 => x"849a3f82",
           656 => x"e0980870",
           657 => x"82e0a408",
           658 => x"f8050c82",
           659 => x"e0a408f8",
           660 => x"05087082",
           661 => x"e0980c51",
           662 => x"54873d0d",
           663 => x"82e0a40c",
           664 => x"0482e0a4",
           665 => x"080282e0",
           666 => x"a40cfb3d",
           667 => x"0d82e0a4",
           668 => x"08900508",
           669 => x"85113370",
           670 => x"81327081",
           671 => x"06515151",
           672 => x"52718f38",
           673 => x"800b82e0",
           674 => x"a4088c05",
           675 => x"08258338",
           676 => x"8d39800b",
           677 => x"82e0a408",
           678 => x"f4050c81",
           679 => x"c43982e0",
           680 => x"a4088c05",
           681 => x"08ff0582",
           682 => x"e0a4088c",
           683 => x"050c800b",
           684 => x"82e0a408",
           685 => x"f8050c82",
           686 => x"e0a40888",
           687 => x"050882e0",
           688 => x"a408fc05",
           689 => x"0c82e0a4",
           690 => x"08f80508",
           691 => x"8a2e80f6",
           692 => x"38800b82",
           693 => x"e0a4088c",
           694 => x"05082580",
           695 => x"e93882e0",
           696 => x"a4089005",
           697 => x"0851a090",
           698 => x"3f82e098",
           699 => x"087082e0",
           700 => x"a408f805",
           701 => x"0c5282e0",
           702 => x"a408f805",
           703 => x"08ff2e09",
           704 => x"81068d38",
           705 => x"800b82e0",
           706 => x"a408f405",
           707 => x"0c80d239",
           708 => x"82e0a408",
           709 => x"fc050882",
           710 => x"e0a408f8",
           711 => x"05085353",
           712 => x"71733482",
           713 => x"e0a4088c",
           714 => x"0508ff05",
           715 => x"82e0a408",
           716 => x"8c050c82",
           717 => x"e0a408fc",
           718 => x"05088105",
           719 => x"82e0a408",
           720 => x"fc050cff",
           721 => x"803982e0",
           722 => x"a408fc05",
           723 => x"08528072",
           724 => x"3482e0a4",
           725 => x"08880508",
           726 => x"7082e0a4",
           727 => x"08f4050c",
           728 => x"5282e0a4",
           729 => x"08f40508",
           730 => x"82e0980c",
           731 => x"873d0d82",
           732 => x"e0a40c04",
           733 => x"82e0a408",
           734 => x"0282e0a4",
           735 => x"0cf43d0d",
           736 => x"860b82e0",
           737 => x"a408e505",
           738 => x"3482e0a4",
           739 => x"08880508",
           740 => x"82e0a408",
           741 => x"e0050cfe",
           742 => x"0a0b82e0",
           743 => x"a408e805",
           744 => x"0c82e0a4",
           745 => x"08900570",
           746 => x"82e0a408",
           747 => x"fc050c82",
           748 => x"e0a408fc",
           749 => x"05085482",
           750 => x"e0a4088c",
           751 => x"05085382",
           752 => x"e0a408e0",
           753 => x"05705351",
           754 => x"54818d3f",
           755 => x"82e09808",
           756 => x"7082e0a4",
           757 => x"08dc050c",
           758 => x"82e0a408",
           759 => x"ec050882",
           760 => x"e0a40888",
           761 => x"05080551",
           762 => x"54807434",
           763 => x"82e0a408",
           764 => x"dc050870",
           765 => x"82e0980c",
           766 => x"548e3d0d",
           767 => x"82e0a40c",
           768 => x"0482e0a4",
           769 => x"080282e0",
           770 => x"a40cfb3d",
           771 => x"0d82e0a4",
           772 => x"08900570",
           773 => x"82e0a408",
           774 => x"fc050c82",
           775 => x"e0a408fc",
           776 => x"05085482",
           777 => x"e0a4088c",
           778 => x"05085382",
           779 => x"e0a40888",
           780 => x"05085254",
           781 => x"a33f82e0",
           782 => x"98087082",
           783 => x"e0a408f8",
           784 => x"050c82e0",
           785 => x"a408f805",
           786 => x"087082e0",
           787 => x"980c5154",
           788 => x"873d0d82",
           789 => x"e0a40c04",
           790 => x"82e0a408",
           791 => x"0282e0a4",
           792 => x"0ced3d0d",
           793 => x"800b82e0",
           794 => x"a408e405",
           795 => x"2382e0a4",
           796 => x"08880508",
           797 => x"53800b8c",
           798 => x"140c82e0",
           799 => x"a4088805",
           800 => x"08851133",
           801 => x"70812a70",
           802 => x"81327081",
           803 => x"06515151",
           804 => x"51537280",
           805 => x"2e8d38ff",
           806 => x"0b82e0a4",
           807 => x"08e0050c",
           808 => x"96ac3982",
           809 => x"e0a4088c",
           810 => x"05085372",
           811 => x"33537282",
           812 => x"e0a408f8",
           813 => x"05347281",
           814 => x"ff065372",
           815 => x"802e95fa",
           816 => x"3882e0a4",
           817 => x"088c0508",
           818 => x"810582e0",
           819 => x"a4088c05",
           820 => x"0c82e0a4",
           821 => x"08e40522",
           822 => x"70810651",
           823 => x"5372802e",
           824 => x"958b3882",
           825 => x"e0a408f8",
           826 => x"053353af",
           827 => x"732781fc",
           828 => x"3882e0a4",
           829 => x"08f80533",
           830 => x"5372b926",
           831 => x"81ee3882",
           832 => x"e0a408f8",
           833 => x"05335372",
           834 => x"b02e0981",
           835 => x"0680c538",
           836 => x"82e0a408",
           837 => x"e8053370",
           838 => x"982b7098",
           839 => x"2c515153",
           840 => x"72b23882",
           841 => x"e0a408e4",
           842 => x"05227083",
           843 => x"2a708132",
           844 => x"70810651",
           845 => x"51515372",
           846 => x"802e9938",
           847 => x"82e0a408",
           848 => x"e4052270",
           849 => x"82800751",
           850 => x"537282e0",
           851 => x"a408e405",
           852 => x"23fed039",
           853 => x"82e0a408",
           854 => x"e8053370",
           855 => x"982b7098",
           856 => x"2c707083",
           857 => x"2b721173",
           858 => x"11515151",
           859 => x"53515553",
           860 => x"7282e0a4",
           861 => x"08e80534",
           862 => x"82e0a408",
           863 => x"e8053354",
           864 => x"82e0a408",
           865 => x"f8053370",
           866 => x"15d01151",
           867 => x"51537282",
           868 => x"e0a408e8",
           869 => x"053482e0",
           870 => x"a408e805",
           871 => x"3370982b",
           872 => x"70982c51",
           873 => x"51537280",
           874 => x"258b3880",
           875 => x"ff0b82e0",
           876 => x"a408e805",
           877 => x"3482e0a4",
           878 => x"08e40522",
           879 => x"70832a70",
           880 => x"81065151",
           881 => x"5372fddb",
           882 => x"3882e0a4",
           883 => x"08e80533",
           884 => x"70882b70",
           885 => x"902b7090",
           886 => x"2c70882c",
           887 => x"51515151",
           888 => x"537282e0",
           889 => x"a408ec05",
           890 => x"23fdb839",
           891 => x"82e0a408",
           892 => x"e4052270",
           893 => x"832a7081",
           894 => x"06515153",
           895 => x"72802e9d",
           896 => x"3882e0a4",
           897 => x"08e80533",
           898 => x"70982b70",
           899 => x"982c5151",
           900 => x"53728a38",
           901 => x"810b82e0",
           902 => x"a408e805",
           903 => x"3482e0a4",
           904 => x"08f80533",
           905 => x"e01182e0",
           906 => x"a408c405",
           907 => x"0c5382e0",
           908 => x"a408c405",
           909 => x"0880d826",
           910 => x"92943882",
           911 => x"e0a408c4",
           912 => x"05087082",
           913 => x"2b82b9dc",
           914 => x"11700851",
           915 => x"51515372",
           916 => x"0482e0a4",
           917 => x"08e40522",
           918 => x"70900751",
           919 => x"537282e0",
           920 => x"a408e405",
           921 => x"2382e0a4",
           922 => x"08e40522",
           923 => x"70a00751",
           924 => x"537282e0",
           925 => x"a408e405",
           926 => x"23fca839",
           927 => x"82e0a408",
           928 => x"e4052270",
           929 => x"81800751",
           930 => x"537282e0",
           931 => x"a408e405",
           932 => x"23fc9039",
           933 => x"82e0a408",
           934 => x"e4052270",
           935 => x"80c00751",
           936 => x"537282e0",
           937 => x"a408e405",
           938 => x"23fbf839",
           939 => x"82e0a408",
           940 => x"e4052270",
           941 => x"88075153",
           942 => x"7282e0a4",
           943 => x"08e40523",
           944 => x"800b82e0",
           945 => x"a408e805",
           946 => x"34fbd839",
           947 => x"82e0a408",
           948 => x"e4052270",
           949 => x"84075153",
           950 => x"7282e0a4",
           951 => x"08e40523",
           952 => x"fbc139bf",
           953 => x"0b82e0a4",
           954 => x"08fc0534",
           955 => x"82e0a408",
           956 => x"ec0522ff",
           957 => x"11515372",
           958 => x"82e0a408",
           959 => x"ec052380",
           960 => x"e30b82e0",
           961 => x"a408f805",
           962 => x"348da839",
           963 => x"82e0a408",
           964 => x"90050882",
           965 => x"e0a40890",
           966 => x"05088405",
           967 => x"82e0a408",
           968 => x"90050c70",
           969 => x"08515372",
           970 => x"82e0a408",
           971 => x"fc053482",
           972 => x"e0a408ec",
           973 => x"0522ff11",
           974 => x"51537282",
           975 => x"e0a408ec",
           976 => x"05238cef",
           977 => x"3982e0a4",
           978 => x"08900508",
           979 => x"82e0a408",
           980 => x"90050884",
           981 => x"0582e0a4",
           982 => x"0890050c",
           983 => x"700882e0",
           984 => x"a408fc05",
           985 => x"0c82e0a4",
           986 => x"08e40522",
           987 => x"70832a70",
           988 => x"81065151",
           989 => x"51537280",
           990 => x"2eab3882",
           991 => x"e0a408e8",
           992 => x"05337098",
           993 => x"2b537298",
           994 => x"2c5382e0",
           995 => x"a408fc05",
           996 => x"085253a4",
           997 => x"833f82e0",
           998 => x"98085372",
           999 => x"82e0a408",
          1000 => x"f4052399",
          1001 => x"3982e0a4",
          1002 => x"08fc0508",
          1003 => x"519d8a3f",
          1004 => x"82e09808",
          1005 => x"537282e0",
          1006 => x"a408f405",
          1007 => x"2382e0a4",
          1008 => x"08ec0522",
          1009 => x"5382e0a4",
          1010 => x"08f40522",
          1011 => x"73713154",
          1012 => x"547282e0",
          1013 => x"a408ec05",
          1014 => x"238bd839",
          1015 => x"82e0a408",
          1016 => x"90050882",
          1017 => x"e0a40890",
          1018 => x"05088405",
          1019 => x"82e0a408",
          1020 => x"90050c70",
          1021 => x"0882e0a4",
          1022 => x"08fc050c",
          1023 => x"82e0a408",
          1024 => x"e4052270",
          1025 => x"832a7081",
          1026 => x"06515151",
          1027 => x"5372802e",
          1028 => x"ab3882e0",
          1029 => x"a408e805",
          1030 => x"3370982b",
          1031 => x"5372982c",
          1032 => x"5382e0a4",
          1033 => x"08fc0508",
          1034 => x"5253a2ec",
          1035 => x"3f82e098",
          1036 => x"08537282",
          1037 => x"e0a408f4",
          1038 => x"05239939",
          1039 => x"82e0a408",
          1040 => x"fc050851",
          1041 => x"9bf33f82",
          1042 => x"e0980853",
          1043 => x"7282e0a4",
          1044 => x"08f40523",
          1045 => x"82e0a408",
          1046 => x"ec052253",
          1047 => x"82e0a408",
          1048 => x"f4052273",
          1049 => x"71315454",
          1050 => x"7282e0a4",
          1051 => x"08ec0523",
          1052 => x"8ac13982",
          1053 => x"e0a408e4",
          1054 => x"05227082",
          1055 => x"2a708106",
          1056 => x"51515372",
          1057 => x"802ea438",
          1058 => x"82e0a408",
          1059 => x"90050882",
          1060 => x"e0a40890",
          1061 => x"05088405",
          1062 => x"82e0a408",
          1063 => x"90050c70",
          1064 => x"0882e0a4",
          1065 => x"08dc050c",
          1066 => x"53a23982",
          1067 => x"e0a40890",
          1068 => x"050882e0",
          1069 => x"a4089005",
          1070 => x"08840582",
          1071 => x"e0a40890",
          1072 => x"050c7008",
          1073 => x"82e0a408",
          1074 => x"dc050c53",
          1075 => x"82e0a408",
          1076 => x"dc050882",
          1077 => x"e0a408fc",
          1078 => x"050c82e0",
          1079 => x"a408fc05",
          1080 => x"088025a4",
          1081 => x"3882e0a4",
          1082 => x"08e40522",
          1083 => x"70820751",
          1084 => x"537282e0",
          1085 => x"a408e405",
          1086 => x"2382e0a4",
          1087 => x"08fc0508",
          1088 => x"3082e0a4",
          1089 => x"08fc050c",
          1090 => x"82e0a408",
          1091 => x"e4052270",
          1092 => x"ffbf0651",
          1093 => x"537282e0",
          1094 => x"a408e405",
          1095 => x"2381af39",
          1096 => x"880b82e0",
          1097 => x"a408f405",
          1098 => x"23a93982",
          1099 => x"e0a408e4",
          1100 => x"05227080",
          1101 => x"c0075153",
          1102 => x"7282e0a4",
          1103 => x"08e40523",
          1104 => x"80f80b82",
          1105 => x"e0a408f8",
          1106 => x"0534900b",
          1107 => x"82e0a408",
          1108 => x"f4052382",
          1109 => x"e0a408e4",
          1110 => x"05227082",
          1111 => x"2a708106",
          1112 => x"51515372",
          1113 => x"802ea438",
          1114 => x"82e0a408",
          1115 => x"90050882",
          1116 => x"e0a40890",
          1117 => x"05088405",
          1118 => x"82e0a408",
          1119 => x"90050c70",
          1120 => x"0882e0a4",
          1121 => x"08d8050c",
          1122 => x"53a23982",
          1123 => x"e0a40890",
          1124 => x"050882e0",
          1125 => x"a4089005",
          1126 => x"08840582",
          1127 => x"e0a40890",
          1128 => x"050c7008",
          1129 => x"82e0a408",
          1130 => x"d8050c53",
          1131 => x"82e0a408",
          1132 => x"d8050882",
          1133 => x"e0a408fc",
          1134 => x"050c82e0",
          1135 => x"a408e405",
          1136 => x"2270cf06",
          1137 => x"51537282",
          1138 => x"e0a408e4",
          1139 => x"052382e0",
          1140 => x"a80b82e0",
          1141 => x"a408f005",
          1142 => x"0c82e0a4",
          1143 => x"08f00508",
          1144 => x"82e0a408",
          1145 => x"f4052282",
          1146 => x"e0a408fc",
          1147 => x"05087155",
          1148 => x"70545654",
          1149 => x"55aaca3f",
          1150 => x"82e09808",
          1151 => x"53727534",
          1152 => x"82e0a408",
          1153 => x"f0050882",
          1154 => x"e0a408d4",
          1155 => x"050c82e0",
          1156 => x"a408f005",
          1157 => x"08703351",
          1158 => x"53897327",
          1159 => x"a43882e0",
          1160 => x"a408f005",
          1161 => x"08537233",
          1162 => x"5482e0a4",
          1163 => x"08f80533",
          1164 => x"7015df11",
          1165 => x"51515372",
          1166 => x"82e0a408",
          1167 => x"d0053497",
          1168 => x"3982e0a4",
          1169 => x"08f00508",
          1170 => x"537233b0",
          1171 => x"11515372",
          1172 => x"82e0a408",
          1173 => x"d0053482",
          1174 => x"e0a408d4",
          1175 => x"05085382",
          1176 => x"e0a408d0",
          1177 => x"05337334",
          1178 => x"82e0a408",
          1179 => x"f0050881",
          1180 => x"0582e0a4",
          1181 => x"08f0050c",
          1182 => x"82e0a408",
          1183 => x"f4052270",
          1184 => x"5382e0a4",
          1185 => x"08fc0508",
          1186 => x"5253a0c7",
          1187 => x"3f82e098",
          1188 => x"087082e0",
          1189 => x"a408fc05",
          1190 => x"0c5382e0",
          1191 => x"a408fc05",
          1192 => x"08802e84",
          1193 => x"38feb239",
          1194 => x"82e0a408",
          1195 => x"f0050882",
          1196 => x"e0a85455",
          1197 => x"72547470",
          1198 => x"75315153",
          1199 => x"7282e0a4",
          1200 => x"08fc0534",
          1201 => x"82e0a408",
          1202 => x"e4052270",
          1203 => x"b2065153",
          1204 => x"72802e94",
          1205 => x"3882e0a4",
          1206 => x"08ec0522",
          1207 => x"ff115153",
          1208 => x"7282e0a4",
          1209 => x"08ec0523",
          1210 => x"82e0a408",
          1211 => x"e4052270",
          1212 => x"862a7081",
          1213 => x"06515153",
          1214 => x"72802e80",
          1215 => x"e73882e0",
          1216 => x"a408ec05",
          1217 => x"2270902b",
          1218 => x"82e0a408",
          1219 => x"cc050c82",
          1220 => x"e0a408cc",
          1221 => x"0508902c",
          1222 => x"82e0a408",
          1223 => x"cc050c82",
          1224 => x"e0a408f4",
          1225 => x"05225153",
          1226 => x"72902e09",
          1227 => x"81069538",
          1228 => x"82e0a408",
          1229 => x"cc0508fe",
          1230 => x"05537282",
          1231 => x"e0a408c8",
          1232 => x"05239339",
          1233 => x"82e0a408",
          1234 => x"cc0508ff",
          1235 => x"05537282",
          1236 => x"e0a408c8",
          1237 => x"052382e0",
          1238 => x"a408c805",
          1239 => x"2282e0a4",
          1240 => x"08ec0523",
          1241 => x"82e0a408",
          1242 => x"e4052270",
          1243 => x"832a7081",
          1244 => x"06515153",
          1245 => x"72802e80",
          1246 => x"d03882e0",
          1247 => x"a408e805",
          1248 => x"3370982b",
          1249 => x"70982c82",
          1250 => x"e0a408fc",
          1251 => x"05335751",
          1252 => x"51537274",
          1253 => x"24973882",
          1254 => x"e0a408e4",
          1255 => x"052270f7",
          1256 => x"06515372",
          1257 => x"82e0a408",
          1258 => x"e405239d",
          1259 => x"3982e0a4",
          1260 => x"08e80533",
          1261 => x"5382e0a4",
          1262 => x"08fc0533",
          1263 => x"73713154",
          1264 => x"547282e0",
          1265 => x"a408e805",
          1266 => x"3482e0a4",
          1267 => x"08e40522",
          1268 => x"70832a70",
          1269 => x"81065151",
          1270 => x"5372802e",
          1271 => x"b13882e0",
          1272 => x"a408e805",
          1273 => x"3370882b",
          1274 => x"70902b70",
          1275 => x"902c7088",
          1276 => x"2c515151",
          1277 => x"51537254",
          1278 => x"82e0a408",
          1279 => x"ec052270",
          1280 => x"75315153",
          1281 => x"7282e0a4",
          1282 => x"08ec0523",
          1283 => x"af3982e0",
          1284 => x"a408fc05",
          1285 => x"3370882b",
          1286 => x"70902b70",
          1287 => x"902c7088",
          1288 => x"2c515151",
          1289 => x"51537254",
          1290 => x"82e0a408",
          1291 => x"ec052270",
          1292 => x"75315153",
          1293 => x"7282e0a4",
          1294 => x"08ec0523",
          1295 => x"82e0a408",
          1296 => x"e4052270",
          1297 => x"83800651",
          1298 => x"5372b038",
          1299 => x"82e0a408",
          1300 => x"ec0522ff",
          1301 => x"11545472",
          1302 => x"82e0a408",
          1303 => x"ec052373",
          1304 => x"902b7090",
          1305 => x"2c515380",
          1306 => x"73259038",
          1307 => x"82e0a408",
          1308 => x"88050852",
          1309 => x"a0518aee",
          1310 => x"3fd23982",
          1311 => x"e0a408e4",
          1312 => x"05227081",
          1313 => x"2a708106",
          1314 => x"51515372",
          1315 => x"802e9138",
          1316 => x"82e0a408",
          1317 => x"88050852",
          1318 => x"ad518aca",
          1319 => x"3f80c739",
          1320 => x"82e0a408",
          1321 => x"e4052270",
          1322 => x"842a7081",
          1323 => x"06515153",
          1324 => x"72802e90",
          1325 => x"3882e0a4",
          1326 => x"08880508",
          1327 => x"52ab518a",
          1328 => x"a53fa339",
          1329 => x"82e0a408",
          1330 => x"e4052270",
          1331 => x"852a7081",
          1332 => x"06515153",
          1333 => x"72802e8e",
          1334 => x"3882e0a4",
          1335 => x"08880508",
          1336 => x"52a0518a",
          1337 => x"813f82e0",
          1338 => x"a408e405",
          1339 => x"2270862a",
          1340 => x"70810651",
          1341 => x"51537280",
          1342 => x"2eb13882",
          1343 => x"e0a40888",
          1344 => x"050852b0",
          1345 => x"5189df3f",
          1346 => x"82e0a408",
          1347 => x"f4052253",
          1348 => x"72902e09",
          1349 => x"81069438",
          1350 => x"82e0a408",
          1351 => x"88050852",
          1352 => x"82e0a408",
          1353 => x"f8053351",
          1354 => x"89bc3f82",
          1355 => x"e0a408e4",
          1356 => x"05227088",
          1357 => x"2a708106",
          1358 => x"51515372",
          1359 => x"802eb038",
          1360 => x"82e0a408",
          1361 => x"ec0522ff",
          1362 => x"11545472",
          1363 => x"82e0a408",
          1364 => x"ec052373",
          1365 => x"902b7090",
          1366 => x"2c515380",
          1367 => x"73259038",
          1368 => x"82e0a408",
          1369 => x"88050852",
          1370 => x"b05188fa",
          1371 => x"3fd23982",
          1372 => x"e0a408e4",
          1373 => x"05227083",
          1374 => x"2a708106",
          1375 => x"51515372",
          1376 => x"802eb038",
          1377 => x"82e0a408",
          1378 => x"e80533ff",
          1379 => x"11545472",
          1380 => x"82e0a408",
          1381 => x"e8053473",
          1382 => x"982b7098",
          1383 => x"2c515380",
          1384 => x"73259038",
          1385 => x"82e0a408",
          1386 => x"88050852",
          1387 => x"b05188b6",
          1388 => x"3fd23982",
          1389 => x"e0a408e4",
          1390 => x"05227087",
          1391 => x"2a708106",
          1392 => x"51515372",
          1393 => x"b03882e0",
          1394 => x"a408ec05",
          1395 => x"22ff1154",
          1396 => x"547282e0",
          1397 => x"a408ec05",
          1398 => x"2373902b",
          1399 => x"70902c51",
          1400 => x"53807325",
          1401 => x"903882e0",
          1402 => x"a4088805",
          1403 => x"0852a051",
          1404 => x"87f43fd2",
          1405 => x"3982e0a4",
          1406 => x"08f80533",
          1407 => x"537280e3",
          1408 => x"2e098106",
          1409 => x"973882e0",
          1410 => x"a4088805",
          1411 => x"085282e0",
          1412 => x"a408fc05",
          1413 => x"335187ce",
          1414 => x"3f81ee39",
          1415 => x"82e0a408",
          1416 => x"f8053353",
          1417 => x"7280f32e",
          1418 => x"09810680",
          1419 => x"cb3882e0",
          1420 => x"a408f405",
          1421 => x"22ff1151",
          1422 => x"537282e0",
          1423 => x"a408f405",
          1424 => x"237283ff",
          1425 => x"ff065372",
          1426 => x"83ffff2e",
          1427 => x"81bb3882",
          1428 => x"e0a40888",
          1429 => x"05085282",
          1430 => x"e0a408fc",
          1431 => x"05087033",
          1432 => x"5282e0a4",
          1433 => x"08fc0508",
          1434 => x"810582e0",
          1435 => x"a408fc05",
          1436 => x"0c5386f2",
          1437 => x"3fffb739",
          1438 => x"82e0a408",
          1439 => x"f8053353",
          1440 => x"7280d32e",
          1441 => x"09810680",
          1442 => x"cb3882e0",
          1443 => x"a408f405",
          1444 => x"22ff1151",
          1445 => x"537282e0",
          1446 => x"a408f405",
          1447 => x"237283ff",
          1448 => x"ff065372",
          1449 => x"83ffff2e",
          1450 => x"80df3882",
          1451 => x"e0a40888",
          1452 => x"05085282",
          1453 => x"e0a408fc",
          1454 => x"05087033",
          1455 => x"525386a6",
          1456 => x"3f82e0a4",
          1457 => x"08fc0508",
          1458 => x"810582e0",
          1459 => x"a408fc05",
          1460 => x"0cffb739",
          1461 => x"82e0a408",
          1462 => x"f0050882",
          1463 => x"e0a82ea9",
          1464 => x"3882e0a4",
          1465 => x"08880508",
          1466 => x"5282e0a4",
          1467 => x"08f00508",
          1468 => x"ff0582e0",
          1469 => x"a408f005",
          1470 => x"0c82e0a4",
          1471 => x"08f00508",
          1472 => x"70335253",
          1473 => x"85e03fcc",
          1474 => x"3982e0a4",
          1475 => x"08e40522",
          1476 => x"70872a70",
          1477 => x"81065151",
          1478 => x"5372802e",
          1479 => x"80c33882",
          1480 => x"e0a408ec",
          1481 => x"0522ff11",
          1482 => x"54547282",
          1483 => x"e0a408ec",
          1484 => x"05237390",
          1485 => x"2b70902c",
          1486 => x"51538073",
          1487 => x"25a33882",
          1488 => x"e0a40888",
          1489 => x"050852a0",
          1490 => x"51859b3f",
          1491 => x"d23982e0",
          1492 => x"a4088805",
          1493 => x"085282e0",
          1494 => x"a408f805",
          1495 => x"33518586",
          1496 => x"3f800b82",
          1497 => x"e0a408e4",
          1498 => x"0523eab7",
          1499 => x"3982e0a4",
          1500 => x"08f80533",
          1501 => x"5372a52e",
          1502 => x"098106a8",
          1503 => x"38810b82",
          1504 => x"e0a408e4",
          1505 => x"0523800b",
          1506 => x"82e0a408",
          1507 => x"ec052380",
          1508 => x"0b82e0a4",
          1509 => x"08e80534",
          1510 => x"8a0b82e0",
          1511 => x"a408f405",
          1512 => x"23ea8039",
          1513 => x"82e0a408",
          1514 => x"88050852",
          1515 => x"82e0a408",
          1516 => x"f8053351",
          1517 => x"84b03fe9",
          1518 => x"ea3982e0",
          1519 => x"a4088805",
          1520 => x"088c1108",
          1521 => x"7082e0a4",
          1522 => x"08e0050c",
          1523 => x"515382e0",
          1524 => x"a408e005",
          1525 => x"0882e098",
          1526 => x"0c953d0d",
          1527 => x"82e0a40c",
          1528 => x"0482e0a4",
          1529 => x"080282e0",
          1530 => x"a40cfd3d",
          1531 => x"0d82fbf8",
          1532 => x"085382e0",
          1533 => x"a4088c05",
          1534 => x"085282e0",
          1535 => x"a4088805",
          1536 => x"0851e4dd",
          1537 => x"3f82e098",
          1538 => x"087082e0",
          1539 => x"980c5485",
          1540 => x"3d0d82e0",
          1541 => x"a40c0482",
          1542 => x"e0a40802",
          1543 => x"82e0a40c",
          1544 => x"fb3d0d80",
          1545 => x"0b82e0a4",
          1546 => x"08f8050c",
          1547 => x"82fbfc08",
          1548 => x"85113370",
          1549 => x"812a7081",
          1550 => x"32708106",
          1551 => x"51515151",
          1552 => x"5372802e",
          1553 => x"8d38ff0b",
          1554 => x"82e0a408",
          1555 => x"f4050c81",
          1556 => x"923982e0",
          1557 => x"a4088805",
          1558 => x"08537233",
          1559 => x"82e0a408",
          1560 => x"88050881",
          1561 => x"0582e0a4",
          1562 => x"0888050c",
          1563 => x"537282e0",
          1564 => x"a408fc05",
          1565 => x"347281ff",
          1566 => x"06537280",
          1567 => x"2eb03882",
          1568 => x"fbfc0882",
          1569 => x"fbfc0853",
          1570 => x"82e0a408",
          1571 => x"fc053352",
          1572 => x"90110851",
          1573 => x"53722d82",
          1574 => x"e0980853",
          1575 => x"72802eff",
          1576 => x"b138ff0b",
          1577 => x"82e0a408",
          1578 => x"f8050cff",
          1579 => x"a53982fb",
          1580 => x"fc0882fb",
          1581 => x"fc085353",
          1582 => x"8a519013",
          1583 => x"0853722d",
          1584 => x"82e09808",
          1585 => x"5372802e",
          1586 => x"8a38ff0b",
          1587 => x"82e0a408",
          1588 => x"f8050c82",
          1589 => x"e0a408f8",
          1590 => x"05087082",
          1591 => x"e0a408f4",
          1592 => x"050c5382",
          1593 => x"e0a408f4",
          1594 => x"050882e0",
          1595 => x"980c873d",
          1596 => x"0d82e0a4",
          1597 => x"0c0482e0",
          1598 => x"a4080282",
          1599 => x"e0a40cfb",
          1600 => x"3d0d800b",
          1601 => x"82e0a408",
          1602 => x"f8050c82",
          1603 => x"e0a4088c",
          1604 => x"05088511",
          1605 => x"3370812a",
          1606 => x"70813270",
          1607 => x"81065151",
          1608 => x"51515372",
          1609 => x"802e8d38",
          1610 => x"ff0b82e0",
          1611 => x"a408f405",
          1612 => x"0c80f339",
          1613 => x"82e0a408",
          1614 => x"88050853",
          1615 => x"723382e0",
          1616 => x"a4088805",
          1617 => x"08810582",
          1618 => x"e0a40888",
          1619 => x"050c5372",
          1620 => x"82e0a408",
          1621 => x"fc053472",
          1622 => x"81ff0653",
          1623 => x"72802eb6",
          1624 => x"3882e0a4",
          1625 => x"088c0508",
          1626 => x"82e0a408",
          1627 => x"8c050853",
          1628 => x"82e0a408",
          1629 => x"fc053352",
          1630 => x"90110851",
          1631 => x"53722d82",
          1632 => x"e0980853",
          1633 => x"72802eff",
          1634 => x"ab38ff0b",
          1635 => x"82e0a408",
          1636 => x"f8050cff",
          1637 => x"9f3982e0",
          1638 => x"a408f805",
          1639 => x"087082e0",
          1640 => x"a408f405",
          1641 => x"0c5382e0",
          1642 => x"a408f405",
          1643 => x"0882e098",
          1644 => x"0c873d0d",
          1645 => x"82e0a40c",
          1646 => x"0482e0a4",
          1647 => x"080282e0",
          1648 => x"a40cfe3d",
          1649 => x"0d82fbfc",
          1650 => x"085282e0",
          1651 => x"a4088805",
          1652 => x"0851933f",
          1653 => x"82e09808",
          1654 => x"7082e098",
          1655 => x"0c53843d",
          1656 => x"0d82e0a4",
          1657 => x"0c0482e0",
          1658 => x"a4080282",
          1659 => x"e0a40cfb",
          1660 => x"3d0d82e0",
          1661 => x"a4088c05",
          1662 => x"08851133",
          1663 => x"70812a70",
          1664 => x"81327081",
          1665 => x"06515151",
          1666 => x"51537280",
          1667 => x"2e8d38ff",
          1668 => x"0b82e0a4",
          1669 => x"08fc050c",
          1670 => x"81cb3982",
          1671 => x"e0a4088c",
          1672 => x"05088511",
          1673 => x"3370822a",
          1674 => x"70810651",
          1675 => x"51515372",
          1676 => x"802e80db",
          1677 => x"3882e0a4",
          1678 => x"088c0508",
          1679 => x"82e0a408",
          1680 => x"8c050854",
          1681 => x"548c1408",
          1682 => x"88140825",
          1683 => x"9f3882e0",
          1684 => x"a4088c05",
          1685 => x"08700870",
          1686 => x"82e0a408",
          1687 => x"88050852",
          1688 => x"57545472",
          1689 => x"75347308",
          1690 => x"8105740c",
          1691 => x"82e0a408",
          1692 => x"8c05088c",
          1693 => x"11088105",
          1694 => x"8c120c82",
          1695 => x"e0a40888",
          1696 => x"05087082",
          1697 => x"e0a408fc",
          1698 => x"050c5153",
          1699 => x"80d73982",
          1700 => x"e0a4088c",
          1701 => x"050882e0",
          1702 => x"a4088c05",
          1703 => x"085382e0",
          1704 => x"a4088805",
          1705 => x"087081ff",
          1706 => x"06539012",
          1707 => x"08515454",
          1708 => x"722d82e0",
          1709 => x"98085372",
          1710 => x"a33882e0",
          1711 => x"a4088c05",
          1712 => x"088c1108",
          1713 => x"81058c12",
          1714 => x"0c82e0a4",
          1715 => x"08880508",
          1716 => x"7082e0a4",
          1717 => x"08fc050c",
          1718 => x"51538a39",
          1719 => x"ff0b82e0",
          1720 => x"a408fc05",
          1721 => x"0c82e0a4",
          1722 => x"08fc0508",
          1723 => x"82e0980c",
          1724 => x"873d0d82",
          1725 => x"e0a40c04",
          1726 => x"82e0a408",
          1727 => x"0282e0a4",
          1728 => x"0cf93d0d",
          1729 => x"82e0a408",
          1730 => x"88050885",
          1731 => x"11337081",
          1732 => x"32708106",
          1733 => x"51515152",
          1734 => x"71802e8d",
          1735 => x"38ff0b82",
          1736 => x"e0a408f8",
          1737 => x"050c8394",
          1738 => x"3982e0a4",
          1739 => x"08880508",
          1740 => x"85113370",
          1741 => x"862a7081",
          1742 => x"06515151",
          1743 => x"5271802e",
          1744 => x"80c53882",
          1745 => x"e0a40888",
          1746 => x"050882e0",
          1747 => x"a4088805",
          1748 => x"08535385",
          1749 => x"123370ff",
          1750 => x"bf065152",
          1751 => x"71851434",
          1752 => x"82e0a408",
          1753 => x"8805088c",
          1754 => x"11088105",
          1755 => x"8c120c82",
          1756 => x"e0a40888",
          1757 => x"05088411",
          1758 => x"337082e0",
          1759 => x"a408f805",
          1760 => x"0c515152",
          1761 => x"82b63982",
          1762 => x"e0a40888",
          1763 => x"05088511",
          1764 => x"3370822a",
          1765 => x"70810651",
          1766 => x"51515271",
          1767 => x"802e80d7",
          1768 => x"3882e0a4",
          1769 => x"08880508",
          1770 => x"70087033",
          1771 => x"82e0a408",
          1772 => x"fc050c51",
          1773 => x"5282e0a4",
          1774 => x"08fc0508",
          1775 => x"a93882e0",
          1776 => x"a4088805",
          1777 => x"0882e0a4",
          1778 => x"08880508",
          1779 => x"53538512",
          1780 => x"3370a007",
          1781 => x"51527185",
          1782 => x"1434ff0b",
          1783 => x"82e0a408",
          1784 => x"f8050c81",
          1785 => x"d73982e0",
          1786 => x"a4088805",
          1787 => x"08700881",
          1788 => x"05710c52",
          1789 => x"81a13982",
          1790 => x"e0a40888",
          1791 => x"050882e0",
          1792 => x"a4088805",
          1793 => x"08529411",
          1794 => x"08515271",
          1795 => x"2d82e098",
          1796 => x"087082e0",
          1797 => x"a408fc05",
          1798 => x"0c5282e0",
          1799 => x"a408fc05",
          1800 => x"08802580",
          1801 => x"f23882e0",
          1802 => x"a4088805",
          1803 => x"0882e0a4",
          1804 => x"08f4050c",
          1805 => x"82e0a408",
          1806 => x"88050885",
          1807 => x"113382e0",
          1808 => x"a408f005",
          1809 => x"0c5282e0",
          1810 => x"a408fc05",
          1811 => x"08ff2e09",
          1812 => x"81069538",
          1813 => x"82e0a408",
          1814 => x"f0050890",
          1815 => x"07527182",
          1816 => x"e0a408ec",
          1817 => x"05349339",
          1818 => x"82e0a408",
          1819 => x"f00508a0",
          1820 => x"07527182",
          1821 => x"e0a408ec",
          1822 => x"053482e0",
          1823 => x"a408f405",
          1824 => x"085282e0",
          1825 => x"a408ec05",
          1826 => x"33851334",
          1827 => x"ff0b82e0",
          1828 => x"a408f805",
          1829 => x"0ca63982",
          1830 => x"e0a40888",
          1831 => x"05088c11",
          1832 => x"0881058c",
          1833 => x"120c82e0",
          1834 => x"a408fc05",
          1835 => x"087081ff",
          1836 => x"067082e0",
          1837 => x"a408f805",
          1838 => x"0c515152",
          1839 => x"82e0a408",
          1840 => x"f8050882",
          1841 => x"e0980c89",
          1842 => x"3d0d82e0",
          1843 => x"a40c0482",
          1844 => x"e0a40802",
          1845 => x"82e0a40c",
          1846 => x"fd3d0d82",
          1847 => x"e0a40888",
          1848 => x"050882e0",
          1849 => x"a408fc05",
          1850 => x"0c82e0a4",
          1851 => x"088c0508",
          1852 => x"82e0a408",
          1853 => x"f8050c82",
          1854 => x"e0a40890",
          1855 => x"0508802e",
          1856 => x"82a23882",
          1857 => x"e0a408f8",
          1858 => x"050882e0",
          1859 => x"a408fc05",
          1860 => x"082681ac",
          1861 => x"3882e0a4",
          1862 => x"08f80508",
          1863 => x"82e0a408",
          1864 => x"90050805",
          1865 => x"5182e0a4",
          1866 => x"08fc0508",
          1867 => x"71278190",
          1868 => x"3882e0a4",
          1869 => x"08fc0508",
          1870 => x"82e0a408",
          1871 => x"90050805",
          1872 => x"82e0a408",
          1873 => x"fc050c82",
          1874 => x"e0a408f8",
          1875 => x"050882e0",
          1876 => x"a4089005",
          1877 => x"080582e0",
          1878 => x"a408f805",
          1879 => x"0c82e0a4",
          1880 => x"08900508",
          1881 => x"810582e0",
          1882 => x"a4089005",
          1883 => x"0c82e0a4",
          1884 => x"08900508",
          1885 => x"ff0582e0",
          1886 => x"a4089005",
          1887 => x"0c82e0a4",
          1888 => x"08900508",
          1889 => x"802e819c",
          1890 => x"3882e0a4",
          1891 => x"08fc0508",
          1892 => x"ff0582e0",
          1893 => x"a408fc05",
          1894 => x"0c82e0a4",
          1895 => x"08f80508",
          1896 => x"ff0582e0",
          1897 => x"a408f805",
          1898 => x"0c82e0a4",
          1899 => x"08fc0508",
          1900 => x"82e0a408",
          1901 => x"f8050853",
          1902 => x"51713371",
          1903 => x"34ffae39",
          1904 => x"82e0a408",
          1905 => x"90050881",
          1906 => x"0582e0a4",
          1907 => x"0890050c",
          1908 => x"82e0a408",
          1909 => x"900508ff",
          1910 => x"0582e0a4",
          1911 => x"0890050c",
          1912 => x"82e0a408",
          1913 => x"90050880",
          1914 => x"2eba3882",
          1915 => x"e0a408f8",
          1916 => x"05085170",
          1917 => x"3382e0a4",
          1918 => x"08f80508",
          1919 => x"810582e0",
          1920 => x"a408f805",
          1921 => x"0c82e0a4",
          1922 => x"08fc0508",
          1923 => x"52527171",
          1924 => x"3482e0a4",
          1925 => x"08fc0508",
          1926 => x"810582e0",
          1927 => x"a408fc05",
          1928 => x"0cffad39",
          1929 => x"82e0a408",
          1930 => x"88050870",
          1931 => x"82e0980c",
          1932 => x"51853d0d",
          1933 => x"82e0a40c",
          1934 => x"0482e0a4",
          1935 => x"080282e0",
          1936 => x"a40cfe3d",
          1937 => x"0d82e0a4",
          1938 => x"08880508",
          1939 => x"82e0a408",
          1940 => x"fc050c82",
          1941 => x"e0a408fc",
          1942 => x"05085271",
          1943 => x"3382e0a4",
          1944 => x"08fc0508",
          1945 => x"810582e0",
          1946 => x"a408fc05",
          1947 => x"0c7081ff",
          1948 => x"06515170",
          1949 => x"802e8338",
          1950 => x"da3982e0",
          1951 => x"a408fc05",
          1952 => x"08ff0582",
          1953 => x"e0a408fc",
          1954 => x"050c82e0",
          1955 => x"a408fc05",
          1956 => x"0882e0a4",
          1957 => x"08880508",
          1958 => x"317082e0",
          1959 => x"980c5184",
          1960 => x"3d0d82e0",
          1961 => x"a40c0482",
          1962 => x"e0a40802",
          1963 => x"82e0a40c",
          1964 => x"fe3d0d82",
          1965 => x"e0a40888",
          1966 => x"050882e0",
          1967 => x"a408fc05",
          1968 => x"0c82e0a4",
          1969 => x"088c0508",
          1970 => x"52713382",
          1971 => x"e0a4088c",
          1972 => x"05088105",
          1973 => x"82e0a408",
          1974 => x"8c050c82",
          1975 => x"e0a408fc",
          1976 => x"05085351",
          1977 => x"70723482",
          1978 => x"e0a408fc",
          1979 => x"05088105",
          1980 => x"82e0a408",
          1981 => x"fc050c70",
          1982 => x"81ff0651",
          1983 => x"70802e84",
          1984 => x"38ffbe39",
          1985 => x"82e0a408",
          1986 => x"88050870",
          1987 => x"82e0980c",
          1988 => x"51843d0d",
          1989 => x"82e0a40c",
          1990 => x"0482e0a4",
          1991 => x"080282e0",
          1992 => x"a40cfd3d",
          1993 => x"0d82e0a4",
          1994 => x"08880508",
          1995 => x"82e0a408",
          1996 => x"fc050c82",
          1997 => x"e0a4088c",
          1998 => x"050882e0",
          1999 => x"a408f805",
          2000 => x"0c82e0a4",
          2001 => x"08900508",
          2002 => x"802e80e5",
          2003 => x"3882e0a4",
          2004 => x"08900508",
          2005 => x"810582e0",
          2006 => x"a4089005",
          2007 => x"0c82e0a4",
          2008 => x"08900508",
          2009 => x"ff0582e0",
          2010 => x"a4089005",
          2011 => x"0c82e0a4",
          2012 => x"08900508",
          2013 => x"802eba38",
          2014 => x"82e0a408",
          2015 => x"f8050851",
          2016 => x"703382e0",
          2017 => x"a408f805",
          2018 => x"08810582",
          2019 => x"e0a408f8",
          2020 => x"050c82e0",
          2021 => x"a408fc05",
          2022 => x"08525271",
          2023 => x"713482e0",
          2024 => x"a408fc05",
          2025 => x"08810582",
          2026 => x"e0a408fc",
          2027 => x"050cffad",
          2028 => x"3982e0a4",
          2029 => x"08880508",
          2030 => x"7082e098",
          2031 => x"0c51853d",
          2032 => x"0d82e0a4",
          2033 => x"0c0482e0",
          2034 => x"a4080282",
          2035 => x"e0a40cfd",
          2036 => x"3d0d82e0",
          2037 => x"a4089005",
          2038 => x"08802e81",
          2039 => x"f43882e0",
          2040 => x"a4088c05",
          2041 => x"08527133",
          2042 => x"82e0a408",
          2043 => x"8c050881",
          2044 => x"0582e0a4",
          2045 => x"088c050c",
          2046 => x"82e0a408",
          2047 => x"88050870",
          2048 => x"337281ff",
          2049 => x"06535454",
          2050 => x"5171712e",
          2051 => x"843880ce",
          2052 => x"3982e0a4",
          2053 => x"08880508",
          2054 => x"52713382",
          2055 => x"e0a40888",
          2056 => x"05088105",
          2057 => x"82e0a408",
          2058 => x"88050c70",
          2059 => x"81ff0651",
          2060 => x"51708d38",
          2061 => x"800b82e0",
          2062 => x"a408fc05",
          2063 => x"0c819b39",
          2064 => x"82e0a408",
          2065 => x"900508ff",
          2066 => x"0582e0a4",
          2067 => x"0890050c",
          2068 => x"82e0a408",
          2069 => x"90050880",
          2070 => x"2e8438ff",
          2071 => x"813982e0",
          2072 => x"a4089005",
          2073 => x"08802e80",
          2074 => x"e83882e0",
          2075 => x"a4088805",
          2076 => x"08703352",
          2077 => x"53708d38",
          2078 => x"ff0b82e0",
          2079 => x"a408fc05",
          2080 => x"0c80d739",
          2081 => x"82e0a408",
          2082 => x"8c0508ff",
          2083 => x"0582e0a4",
          2084 => x"088c050c",
          2085 => x"82e0a408",
          2086 => x"8c050870",
          2087 => x"33525270",
          2088 => x"8c38810b",
          2089 => x"82e0a408",
          2090 => x"fc050cae",
          2091 => x"3982e0a4",
          2092 => x"08880508",
          2093 => x"703382e0",
          2094 => x"a4088c05",
          2095 => x"08703372",
          2096 => x"71317082",
          2097 => x"e0a408fc",
          2098 => x"050c5355",
          2099 => x"5252538a",
          2100 => x"39800b82",
          2101 => x"e0a408fc",
          2102 => x"050c82e0",
          2103 => x"a408fc05",
          2104 => x"0882e098",
          2105 => x"0c853d0d",
          2106 => x"82e0a40c",
          2107 => x"0482e0a4",
          2108 => x"080282e0",
          2109 => x"a40cfa3d",
          2110 => x"0d82e0a4",
          2111 => x"088c0508",
          2112 => x"5282e0a4",
          2113 => x"08880508",
          2114 => x"51818d3f",
          2115 => x"82e09808",
          2116 => x"7082e0a4",
          2117 => x"08f8050c",
          2118 => x"82e0a408",
          2119 => x"f8050881",
          2120 => x"05705351",
          2121 => x"5480ecf7",
          2122 => x"3f82e098",
          2123 => x"087082e0",
          2124 => x"a408fc05",
          2125 => x"0c5482e0",
          2126 => x"a408fc05",
          2127 => x"088c3880",
          2128 => x"0b82e0a4",
          2129 => x"08f4050c",
          2130 => x"bc3982e0",
          2131 => x"a408fc05",
          2132 => x"0882e0a4",
          2133 => x"08f80508",
          2134 => x"05548074",
          2135 => x"3482e0a4",
          2136 => x"08f80508",
          2137 => x"5382e0a4",
          2138 => x"08880508",
          2139 => x"5282e0a4",
          2140 => x"08fc0508",
          2141 => x"51fba23f",
          2142 => x"82e09808",
          2143 => x"7082e0a4",
          2144 => x"08f4050c",
          2145 => x"5482e0a4",
          2146 => x"08f40508",
          2147 => x"82e0980c",
          2148 => x"883d0d82",
          2149 => x"e0a40c04",
          2150 => x"82e0a408",
          2151 => x"0282e0a4",
          2152 => x"0cfd3d0d",
          2153 => x"82e0a408",
          2154 => x"88050882",
          2155 => x"e0a408f8",
          2156 => x"050c82e0",
          2157 => x"a4088c05",
          2158 => x"088d3880",
          2159 => x"0b82e0a4",
          2160 => x"08fc050c",
          2161 => x"80ec3982",
          2162 => x"e0a408f8",
          2163 => x"05085271",
          2164 => x"3382e0a4",
          2165 => x"08f80508",
          2166 => x"810582e0",
          2167 => x"a408f805",
          2168 => x"0c7081ff",
          2169 => x"06515170",
          2170 => x"802e9f38",
          2171 => x"82e0a408",
          2172 => x"8c0508ff",
          2173 => x"0582e0a4",
          2174 => x"088c050c",
          2175 => x"82e0a408",
          2176 => x"8c0508ff",
          2177 => x"2e8438ff",
          2178 => x"be3982e0",
          2179 => x"a408f805",
          2180 => x"08ff0582",
          2181 => x"e0a408f8",
          2182 => x"050c82e0",
          2183 => x"a408f805",
          2184 => x"0882e0a4",
          2185 => x"08880508",
          2186 => x"317082e0",
          2187 => x"a408fc05",
          2188 => x"0c5182e0",
          2189 => x"a408fc05",
          2190 => x"0882e098",
          2191 => x"0c853d0d",
          2192 => x"82e0a40c",
          2193 => x"0482e0a4",
          2194 => x"080282e0",
          2195 => x"a40cfe3d",
          2196 => x"0d82e0a4",
          2197 => x"08880508",
          2198 => x"82e0a408",
          2199 => x"fc050c82",
          2200 => x"e0a40890",
          2201 => x"0508802e",
          2202 => x"80d43882",
          2203 => x"e0a40890",
          2204 => x"05088105",
          2205 => x"82e0a408",
          2206 => x"90050c82",
          2207 => x"e0a40890",
          2208 => x"0508ff05",
          2209 => x"82e0a408",
          2210 => x"90050c82",
          2211 => x"e0a40890",
          2212 => x"0508802e",
          2213 => x"a93882e0",
          2214 => x"a4088c05",
          2215 => x"08517082",
          2216 => x"e0a408fc",
          2217 => x"05085252",
          2218 => x"71713482",
          2219 => x"e0a408fc",
          2220 => x"05088105",
          2221 => x"82e0a408",
          2222 => x"fc050cff",
          2223 => x"be3982e0",
          2224 => x"a4088805",
          2225 => x"087082e0",
          2226 => x"980c5184",
          2227 => x"3d0d82e0",
          2228 => x"a40c0482",
          2229 => x"e0a40802",
          2230 => x"82e0a40c",
          2231 => x"fe3d0d82",
          2232 => x"e0a4088c",
          2233 => x"05085282",
          2234 => x"e0a40888",
          2235 => x"05085193",
          2236 => x"3f82e098",
          2237 => x"087082e0",
          2238 => x"980c5384",
          2239 => x"3d0d82e0",
          2240 => x"a40c0482",
          2241 => x"e0a40802",
          2242 => x"82e0a40c",
          2243 => x"f63d0da0",
          2244 => x"0b82e0a4",
          2245 => x"08fc050c",
          2246 => x"82e0a408",
          2247 => x"8c050880",
          2248 => x"2e9b3882",
          2249 => x"e0a4088c",
          2250 => x"05085183",
          2251 => x"fc3f82e0",
          2252 => x"98087082",
          2253 => x"e0a408e4",
          2254 => x"050c528f",
          2255 => x"3982e0a4",
          2256 => x"08fc0508",
          2257 => x"82e0a408",
          2258 => x"e4050c82",
          2259 => x"e0a40888",
          2260 => x"0508802e",
          2261 => x"a33882e0",
          2262 => x"a4088805",
          2263 => x"085183c9",
          2264 => x"3f82e098",
          2265 => x"0882e0a4",
          2266 => x"08e40508",
          2267 => x"713182e0",
          2268 => x"a408e005",
          2269 => x"0c529739",
          2270 => x"82e0a408",
          2271 => x"e4050882",
          2272 => x"e0a408fc",
          2273 => x"05083182",
          2274 => x"e0a408e0",
          2275 => x"050c82e0",
          2276 => x"a408e005",
          2277 => x"0882e0a4",
          2278 => x"08f8050c",
          2279 => x"82e0a408",
          2280 => x"fc0508ff",
          2281 => x"05527182",
          2282 => x"e0a408f8",
          2283 => x"0508278d",
          2284 => x"38800b82",
          2285 => x"e0a408e8",
          2286 => x"050c82da",
          2287 => x"3982e0a4",
          2288 => x"08fc0508",
          2289 => x"ff055271",
          2290 => x"82e0a408",
          2291 => x"f805082e",
          2292 => x"09810694",
          2293 => x"3882e0a4",
          2294 => x"08880508",
          2295 => x"7082e0a4",
          2296 => x"08e8050c",
          2297 => x"5282af39",
          2298 => x"82e0a408",
          2299 => x"f8050881",
          2300 => x"0582e0a4",
          2301 => x"08f8050c",
          2302 => x"82e0a408",
          2303 => x"88050882",
          2304 => x"e0a408f8",
          2305 => x"05082a82",
          2306 => x"e0a408f4",
          2307 => x"050c82e0",
          2308 => x"a408fc05",
          2309 => x"0882e0a4",
          2310 => x"08f80508",
          2311 => x"3182e0a4",
          2312 => x"08880508",
          2313 => x"712b82e0",
          2314 => x"a4088805",
          2315 => x"0c52800b",
          2316 => x"82e0a408",
          2317 => x"f0050c82",
          2318 => x"e0a408f8",
          2319 => x"0508802e",
          2320 => x"81ab3882",
          2321 => x"e0a408f4",
          2322 => x"05081082",
          2323 => x"e0a408fc",
          2324 => x"0508ff05",
          2325 => x"82e0a408",
          2326 => x"88050871",
          2327 => x"2a707307",
          2328 => x"82e0a408",
          2329 => x"f4050c82",
          2330 => x"e0a40888",
          2331 => x"05081070",
          2332 => x"82e0a408",
          2333 => x"f0050807",
          2334 => x"82e0a408",
          2335 => x"88050c82",
          2336 => x"e0a4088c",
          2337 => x"050882e0",
          2338 => x"a408f405",
          2339 => x"0831ff11",
          2340 => x"82e0a408",
          2341 => x"fc0508ff",
          2342 => x"0571712c",
          2343 => x"82e0a408",
          2344 => x"ec050c82",
          2345 => x"e0a408ec",
          2346 => x"05088106",
          2347 => x"82e0a408",
          2348 => x"f0050c82",
          2349 => x"e0a4088c",
          2350 => x"050882e0",
          2351 => x"a408ec05",
          2352 => x"080682e0",
          2353 => x"a408f405",
          2354 => x"08713182",
          2355 => x"e0a408f4",
          2356 => x"050c82e0",
          2357 => x"a408f805",
          2358 => x"08ff0582",
          2359 => x"e0a408f8",
          2360 => x"050c5152",
          2361 => x"55515151",
          2362 => x"5353fecb",
          2363 => x"3982e0a4",
          2364 => x"08880508",
          2365 => x"107082e0",
          2366 => x"a408f005",
          2367 => x"080782e0",
          2368 => x"a4088805",
          2369 => x"0c82e0a4",
          2370 => x"08880508",
          2371 => x"7082e0a4",
          2372 => x"08e8050c",
          2373 => x"515282e0",
          2374 => x"a408e805",
          2375 => x"0882e098",
          2376 => x"0c8c3d0d",
          2377 => x"82e0a40c",
          2378 => x"0482e0a4",
          2379 => x"080282e0",
          2380 => x"a40cf83d",
          2381 => x"0d82e0a4",
          2382 => x"08880508",
          2383 => x"82e0a408",
          2384 => x"fc050c82",
          2385 => x"e0a408fc",
          2386 => x"0508fc80",
          2387 => x"80065170",
          2388 => x"8c38900b",
          2389 => x"82e0a408",
          2390 => x"f0050c8a",
          2391 => x"39800b82",
          2392 => x"e0a408f0",
          2393 => x"050c82e0",
          2394 => x"a408f005",
          2395 => x"0882e0a4",
          2396 => x"08f8050c",
          2397 => x"900b82e0",
          2398 => x"a408f805",
          2399 => x"083182e0",
          2400 => x"a408fc05",
          2401 => x"08712a82",
          2402 => x"e0a408fc",
          2403 => x"050c82e0",
          2404 => x"a408f805",
          2405 => x"0882e0a4",
          2406 => x"08f4050c",
          2407 => x"82e0a408",
          2408 => x"fc050883",
          2409 => x"fe800651",
          2410 => x"51708c38",
          2411 => x"880b82e0",
          2412 => x"a408ec05",
          2413 => x"0c8a3980",
          2414 => x"0b82e0a4",
          2415 => x"08ec050c",
          2416 => x"82e0a408",
          2417 => x"ec050882",
          2418 => x"e0a408f8",
          2419 => x"050c880b",
          2420 => x"82e0a408",
          2421 => x"f8050831",
          2422 => x"82e0a408",
          2423 => x"fc050871",
          2424 => x"2a82e0a4",
          2425 => x"08fc050c",
          2426 => x"82e0a408",
          2427 => x"f4050882",
          2428 => x"e0a408f8",
          2429 => x"05080582",
          2430 => x"e0a408f4",
          2431 => x"050c82e0",
          2432 => x"a408fc05",
          2433 => x"0881f006",
          2434 => x"5151708c",
          2435 => x"38840b82",
          2436 => x"e0a408e8",
          2437 => x"050c8a39",
          2438 => x"800b82e0",
          2439 => x"a408e805",
          2440 => x"0c82e0a4",
          2441 => x"08e80508",
          2442 => x"82e0a408",
          2443 => x"f8050c84",
          2444 => x"0b82e0a4",
          2445 => x"08f80508",
          2446 => x"3182e0a4",
          2447 => x"08fc0508",
          2448 => x"712a82e0",
          2449 => x"a408fc05",
          2450 => x"0c82e0a4",
          2451 => x"08f40508",
          2452 => x"82e0a408",
          2453 => x"f8050805",
          2454 => x"82e0a408",
          2455 => x"f4050c82",
          2456 => x"e0a408fc",
          2457 => x"05088c06",
          2458 => x"5151708c",
          2459 => x"38820b82",
          2460 => x"e0a408e4",
          2461 => x"050c8a39",
          2462 => x"800b82e0",
          2463 => x"a408e405",
          2464 => x"0c82e0a4",
          2465 => x"08e40508",
          2466 => x"82e0a408",
          2467 => x"f8050c82",
          2468 => x"0b82e0a4",
          2469 => x"08f80508",
          2470 => x"3182e0a4",
          2471 => x"08fc0508",
          2472 => x"712a82e0",
          2473 => x"a408fc05",
          2474 => x"0c82e0a4",
          2475 => x"08f40508",
          2476 => x"82e0a408",
          2477 => x"f8050805",
          2478 => x"82e0a408",
          2479 => x"f4050c82",
          2480 => x"0b82e0a4",
          2481 => x"08fc0508",
          2482 => x"3182e0a4",
          2483 => x"08fc0508",
          2484 => x"812a7081",
          2485 => x"32708106",
          2486 => x"70307075",
          2487 => x"0682e0a4",
          2488 => x"08f40508",
          2489 => x"11707082",
          2490 => x"e0980c53",
          2491 => x"51555151",
          2492 => x"51525351",
          2493 => x"8a3d0d82",
          2494 => x"e0a40c04",
          2495 => x"82e0a408",
          2496 => x"0282e0a4",
          2497 => x"0cfe3d0d",
          2498 => x"82e0a408",
          2499 => x"8c050852",
          2500 => x"82e0a408",
          2501 => x"88050851",
          2502 => x"84e43f82",
          2503 => x"e0980870",
          2504 => x"82e0a408",
          2505 => x"8c050829",
          2506 => x"82e0a408",
          2507 => x"88050871",
          2508 => x"317082e0",
          2509 => x"980c5151",
          2510 => x"53843d0d",
          2511 => x"82e0a40c",
          2512 => x"0482e0a4",
          2513 => x"080282e0",
          2514 => x"a40cfe3d",
          2515 => x"0d82e0a4",
          2516 => x"088c0508",
          2517 => x"5282e0a4",
          2518 => x"08880508",
          2519 => x"51933f82",
          2520 => x"e0980870",
          2521 => x"82e0980c",
          2522 => x"53843d0d",
          2523 => x"82e0a40c",
          2524 => x"0482e0a4",
          2525 => x"080282e0",
          2526 => x"a40cf63d",
          2527 => x"0da00b82",
          2528 => x"e0a408fc",
          2529 => x"050c82e0",
          2530 => x"a4088c05",
          2531 => x"08802e9b",
          2532 => x"3882e0a4",
          2533 => x"088c0508",
          2534 => x"51fb8e3f",
          2535 => x"82e09808",
          2536 => x"7082e0a4",
          2537 => x"08e4050c",
          2538 => x"528f3982",
          2539 => x"e0a408fc",
          2540 => x"050882e0",
          2541 => x"a408e405",
          2542 => x"0c82e0a4",
          2543 => x"08880508",
          2544 => x"802ea338",
          2545 => x"82e0a408",
          2546 => x"88050851",
          2547 => x"fadb3f82",
          2548 => x"e0980882",
          2549 => x"e0a408e4",
          2550 => x"05087131",
          2551 => x"82e0a408",
          2552 => x"e0050c52",
          2553 => x"973982e0",
          2554 => x"a408e405",
          2555 => x"0882e0a4",
          2556 => x"08fc0508",
          2557 => x"3182e0a4",
          2558 => x"08e0050c",
          2559 => x"82e0a408",
          2560 => x"e0050882",
          2561 => x"e0a408f8",
          2562 => x"050c82e0",
          2563 => x"a408fc05",
          2564 => x"08ff0552",
          2565 => x"7182e0a4",
          2566 => x"08f80508",
          2567 => x"27943882",
          2568 => x"e0a40888",
          2569 => x"05087082",
          2570 => x"e0a408e8",
          2571 => x"050c5282",
          2572 => x"ba3982e0",
          2573 => x"a408fc05",
          2574 => x"08ff0552",
          2575 => x"7182e0a4",
          2576 => x"08f80508",
          2577 => x"2e098106",
          2578 => x"8d38800b",
          2579 => x"82e0a408",
          2580 => x"e8050c82",
          2581 => x"963982e0",
          2582 => x"a408f805",
          2583 => x"08810582",
          2584 => x"e0a408f8",
          2585 => x"050c82e0",
          2586 => x"a4088805",
          2587 => x"0882e0a4",
          2588 => x"08f80508",
          2589 => x"2a82e0a4",
          2590 => x"08f4050c",
          2591 => x"82e0a408",
          2592 => x"fc050882",
          2593 => x"e0a408f8",
          2594 => x"05083182",
          2595 => x"e0a40888",
          2596 => x"0508712b",
          2597 => x"82e0a408",
          2598 => x"88050c52",
          2599 => x"800b82e0",
          2600 => x"a408f005",
          2601 => x"0c82e0a4",
          2602 => x"08f80508",
          2603 => x"802e81ab",
          2604 => x"3882e0a4",
          2605 => x"08f40508",
          2606 => x"1082e0a4",
          2607 => x"08fc0508",
          2608 => x"ff0582e0",
          2609 => x"a4088805",
          2610 => x"08712a70",
          2611 => x"730782e0",
          2612 => x"a408f405",
          2613 => x"0c82e0a4",
          2614 => x"08880508",
          2615 => x"107082e0",
          2616 => x"a408f005",
          2617 => x"080782e0",
          2618 => x"a4088805",
          2619 => x"0c82e0a4",
          2620 => x"088c0508",
          2621 => x"82e0a408",
          2622 => x"f4050831",
          2623 => x"ff1182e0",
          2624 => x"a408fc05",
          2625 => x"08ff0571",
          2626 => x"712c82e0",
          2627 => x"a408ec05",
          2628 => x"0c82e0a4",
          2629 => x"08ec0508",
          2630 => x"810682e0",
          2631 => x"a408f005",
          2632 => x"0c82e0a4",
          2633 => x"088c0508",
          2634 => x"82e0a408",
          2635 => x"ec050806",
          2636 => x"82e0a408",
          2637 => x"f4050871",
          2638 => x"3182e0a4",
          2639 => x"08f4050c",
          2640 => x"82e0a408",
          2641 => x"f80508ff",
          2642 => x"0582e0a4",
          2643 => x"08f8050c",
          2644 => x"51525551",
          2645 => x"51515353",
          2646 => x"fecb3982",
          2647 => x"e0a408f4",
          2648 => x"05087082",
          2649 => x"e0a408e8",
          2650 => x"050c5282",
          2651 => x"e0a408e8",
          2652 => x"050882e0",
          2653 => x"980c8c3d",
          2654 => x"0d82e0a4",
          2655 => x"0c0482e0",
          2656 => x"a4080282",
          2657 => x"e0a40cfb",
          2658 => x"3d0d9f0b",
          2659 => x"82e0a408",
          2660 => x"fc050c82",
          2661 => x"e0a40888",
          2662 => x"050882e0",
          2663 => x"a408fc05",
          2664 => x"082c82e0",
          2665 => x"a408f805",
          2666 => x"0c82e0a4",
          2667 => x"088c0508",
          2668 => x"82e0a408",
          2669 => x"fc05082c",
          2670 => x"82e0a408",
          2671 => x"f4050c82",
          2672 => x"e0a40888",
          2673 => x"050882e0",
          2674 => x"a408f805",
          2675 => x"08327082",
          2676 => x"e0a408f8",
          2677 => x"05083182",
          2678 => x"e0a40888",
          2679 => x"050c82e0",
          2680 => x"a4088c05",
          2681 => x"0882e0a4",
          2682 => x"08f40508",
          2683 => x"327082e0",
          2684 => x"a408f405",
          2685 => x"083182e0",
          2686 => x"a4088c05",
          2687 => x"0c82e0a4",
          2688 => x"08f80508",
          2689 => x"82e0a408",
          2690 => x"f4050832",
          2691 => x"82e0a408",
          2692 => x"f8050c82",
          2693 => x"e0a4088c",
          2694 => x"05085482",
          2695 => x"e0a40888",
          2696 => x"05085351",
          2697 => x"53f1ac3f",
          2698 => x"82e09808",
          2699 => x"7082e0a4",
          2700 => x"08f80508",
          2701 => x"327082e0",
          2702 => x"a408f805",
          2703 => x"08317082",
          2704 => x"e0980c51",
          2705 => x"5153873d",
          2706 => x"0d82e0a4",
          2707 => x"0c0482e0",
          2708 => x"a4080282",
          2709 => x"e0a40cf7",
          2710 => x"3d0d800b",
          2711 => x"82e0a408",
          2712 => x"f0053482",
          2713 => x"e0a4088c",
          2714 => x"05085380",
          2715 => x"730c82e0",
          2716 => x"a4088805",
          2717 => x"08700851",
          2718 => x"53723353",
          2719 => x"7282e0a4",
          2720 => x"08f80534",
          2721 => x"7281ff06",
          2722 => x"5372a02e",
          2723 => x"09810691",
          2724 => x"3882e0a4",
          2725 => x"08880508",
          2726 => x"70088105",
          2727 => x"710c53ce",
          2728 => x"3982e0a4",
          2729 => x"08f80533",
          2730 => x"5372ad2e",
          2731 => x"098106a4",
          2732 => x"38810b82",
          2733 => x"e0a408f0",
          2734 => x"053482e0",
          2735 => x"a4088805",
          2736 => x"08700881",
          2737 => x"05710c70",
          2738 => x"08515372",
          2739 => x"3382e0a4",
          2740 => x"08f80534",
          2741 => x"82e0a408",
          2742 => x"f8053353",
          2743 => x"72b02e09",
          2744 => x"810681dc",
          2745 => x"3882e0a4",
          2746 => x"08880508",
          2747 => x"70088105",
          2748 => x"710c7008",
          2749 => x"51537233",
          2750 => x"82e0a408",
          2751 => x"f8053482",
          2752 => x"e0a408f8",
          2753 => x"053382e0",
          2754 => x"a408e805",
          2755 => x"0c82e0a4",
          2756 => x"08e80508",
          2757 => x"80e22eb6",
          2758 => x"3882e0a4",
          2759 => x"08e80508",
          2760 => x"80f82e84",
          2761 => x"3880cd39",
          2762 => x"900b82e0",
          2763 => x"a408f405",
          2764 => x"3482e0a4",
          2765 => x"08880508",
          2766 => x"70088105",
          2767 => x"710c7008",
          2768 => x"51537233",
          2769 => x"82e0a408",
          2770 => x"f8053481",
          2771 => x"a439820b",
          2772 => x"82e0a408",
          2773 => x"f4053482",
          2774 => x"e0a40888",
          2775 => x"05087008",
          2776 => x"8105710c",
          2777 => x"70085153",
          2778 => x"723382e0",
          2779 => x"a408f805",
          2780 => x"3480fe39",
          2781 => x"82e0a408",
          2782 => x"f8053353",
          2783 => x"72a0268d",
          2784 => x"38810b82",
          2785 => x"e0a408ec",
          2786 => x"050c8380",
          2787 => x"3982e0a4",
          2788 => x"08f80533",
          2789 => x"53af7327",
          2790 => x"903882e0",
          2791 => x"a408f805",
          2792 => x"335372b9",
          2793 => x"2683388d",
          2794 => x"39800b82",
          2795 => x"e0a408ec",
          2796 => x"050c82d8",
          2797 => x"39880b82",
          2798 => x"e0a408f4",
          2799 => x"0534b239",
          2800 => x"82e0a408",
          2801 => x"f8053353",
          2802 => x"af732790",
          2803 => x"3882e0a4",
          2804 => x"08f80533",
          2805 => x"5372b926",
          2806 => x"83388d39",
          2807 => x"800b82e0",
          2808 => x"a408ec05",
          2809 => x"0c82a539",
          2810 => x"8a0b82e0",
          2811 => x"a408f405",
          2812 => x"34800b82",
          2813 => x"e0a408fc",
          2814 => x"050c82e0",
          2815 => x"a408f805",
          2816 => x"3353a073",
          2817 => x"2781cf38",
          2818 => x"82e0a408",
          2819 => x"f8053353",
          2820 => x"80e07327",
          2821 => x"943882e0",
          2822 => x"a408f805",
          2823 => x"33e01151",
          2824 => x"537282e0",
          2825 => x"a408f805",
          2826 => x"3482e0a4",
          2827 => x"08f80533",
          2828 => x"d0115153",
          2829 => x"7282e0a4",
          2830 => x"08f80534",
          2831 => x"82e0a408",
          2832 => x"f8053353",
          2833 => x"907327ad",
          2834 => x"3882e0a4",
          2835 => x"08f80533",
          2836 => x"f9115153",
          2837 => x"7282e0a4",
          2838 => x"08f80534",
          2839 => x"82e0a408",
          2840 => x"f8053353",
          2841 => x"7289268d",
          2842 => x"38800b82",
          2843 => x"e0a408ec",
          2844 => x"050c8198",
          2845 => x"3982e0a4",
          2846 => x"08f80533",
          2847 => x"82e0a408",
          2848 => x"f4053354",
          2849 => x"54727426",
          2850 => x"8d38800b",
          2851 => x"82e0a408",
          2852 => x"ec050c80",
          2853 => x"f73982e0",
          2854 => x"a408f405",
          2855 => x"337082e0",
          2856 => x"a408fc05",
          2857 => x"082982e0",
          2858 => x"a408f805",
          2859 => x"33701282",
          2860 => x"e0a408fc",
          2861 => x"050c82e0",
          2862 => x"a4088805",
          2863 => x"08700881",
          2864 => x"05710c70",
          2865 => x"08515152",
          2866 => x"55537233",
          2867 => x"82e0a408",
          2868 => x"f80534fe",
          2869 => x"a53982e0",
          2870 => x"a408f005",
          2871 => x"33537280",
          2872 => x"2e903882",
          2873 => x"e0a408fc",
          2874 => x"05083082",
          2875 => x"e0a408fc",
          2876 => x"050c82e0",
          2877 => x"a4088c05",
          2878 => x"0882e0a4",
          2879 => x"08fc0508",
          2880 => x"710c5381",
          2881 => x"0b82e0a4",
          2882 => x"08ec050c",
          2883 => x"82e0a408",
          2884 => x"ec050882",
          2885 => x"e0980c8b",
          2886 => x"3d0d82e0",
          2887 => x"a40c0482",
          2888 => x"e0a40802",
          2889 => x"82e0a40c",
          2890 => x"f73d0d80",
          2891 => x"0b82e0a4",
          2892 => x"08f00534",
          2893 => x"82e0a408",
          2894 => x"8c050853",
          2895 => x"80730c82",
          2896 => x"e0a40888",
          2897 => x"05087008",
          2898 => x"51537233",
          2899 => x"537282e0",
          2900 => x"a408f805",
          2901 => x"347281ff",
          2902 => x"065372a0",
          2903 => x"2e098106",
          2904 => x"913882e0",
          2905 => x"a4088805",
          2906 => x"08700881",
          2907 => x"05710c53",
          2908 => x"ce3982e0",
          2909 => x"a408f805",
          2910 => x"335372ad",
          2911 => x"2e098106",
          2912 => x"a438810b",
          2913 => x"82e0a408",
          2914 => x"f0053482",
          2915 => x"e0a40888",
          2916 => x"05087008",
          2917 => x"8105710c",
          2918 => x"70085153",
          2919 => x"723382e0",
          2920 => x"a408f805",
          2921 => x"3482e0a4",
          2922 => x"08f80533",
          2923 => x"5372b02e",
          2924 => x"09810681",
          2925 => x"dc3882e0",
          2926 => x"a4088805",
          2927 => x"08700881",
          2928 => x"05710c70",
          2929 => x"08515372",
          2930 => x"3382e0a4",
          2931 => x"08f80534",
          2932 => x"82e0a408",
          2933 => x"f8053382",
          2934 => x"e0a408e8",
          2935 => x"050c82e0",
          2936 => x"a408e805",
          2937 => x"0880e22e",
          2938 => x"b63882e0",
          2939 => x"a408e805",
          2940 => x"0880f82e",
          2941 => x"843880cd",
          2942 => x"39900b82",
          2943 => x"e0a408f4",
          2944 => x"053482e0",
          2945 => x"a4088805",
          2946 => x"08700881",
          2947 => x"05710c70",
          2948 => x"08515372",
          2949 => x"3382e0a4",
          2950 => x"08f80534",
          2951 => x"81a43982",
          2952 => x"0b82e0a4",
          2953 => x"08f40534",
          2954 => x"82e0a408",
          2955 => x"88050870",
          2956 => x"08810571",
          2957 => x"0c700851",
          2958 => x"53723382",
          2959 => x"e0a408f8",
          2960 => x"053480fe",
          2961 => x"3982e0a4",
          2962 => x"08f80533",
          2963 => x"5372a026",
          2964 => x"8d38810b",
          2965 => x"82e0a408",
          2966 => x"ec050c83",
          2967 => x"803982e0",
          2968 => x"a408f805",
          2969 => x"3353af73",
          2970 => x"27903882",
          2971 => x"e0a408f8",
          2972 => x"05335372",
          2973 => x"b9268338",
          2974 => x"8d39800b",
          2975 => x"82e0a408",
          2976 => x"ec050c82",
          2977 => x"d839880b",
          2978 => x"82e0a408",
          2979 => x"f40534b2",
          2980 => x"3982e0a4",
          2981 => x"08f80533",
          2982 => x"53af7327",
          2983 => x"903882e0",
          2984 => x"a408f805",
          2985 => x"335372b9",
          2986 => x"2683388d",
          2987 => x"39800b82",
          2988 => x"e0a408ec",
          2989 => x"050c82a5",
          2990 => x"398a0b82",
          2991 => x"e0a408f4",
          2992 => x"0534800b",
          2993 => x"82e0a408",
          2994 => x"fc050c82",
          2995 => x"e0a408f8",
          2996 => x"053353a0",
          2997 => x"732781cf",
          2998 => x"3882e0a4",
          2999 => x"08f80533",
          3000 => x"5380e073",
          3001 => x"27943882",
          3002 => x"e0a408f8",
          3003 => x"0533e011",
          3004 => x"51537282",
          3005 => x"e0a408f8",
          3006 => x"053482e0",
          3007 => x"a408f805",
          3008 => x"33d01151",
          3009 => x"537282e0",
          3010 => x"a408f805",
          3011 => x"3482e0a4",
          3012 => x"08f80533",
          3013 => x"53907327",
          3014 => x"ad3882e0",
          3015 => x"a408f805",
          3016 => x"33f91151",
          3017 => x"537282e0",
          3018 => x"a408f805",
          3019 => x"3482e0a4",
          3020 => x"08f80533",
          3021 => x"53728926",
          3022 => x"8d38800b",
          3023 => x"82e0a408",
          3024 => x"ec050c81",
          3025 => x"983982e0",
          3026 => x"a408f805",
          3027 => x"3382e0a4",
          3028 => x"08f40533",
          3029 => x"54547274",
          3030 => x"268d3880",
          3031 => x"0b82e0a4",
          3032 => x"08ec050c",
          3033 => x"80f73982",
          3034 => x"e0a408f4",
          3035 => x"05337082",
          3036 => x"e0a408fc",
          3037 => x"05082982",
          3038 => x"e0a408f8",
          3039 => x"05337012",
          3040 => x"82e0a408",
          3041 => x"fc050c82",
          3042 => x"e0a40888",
          3043 => x"05087008",
          3044 => x"8105710c",
          3045 => x"70085151",
          3046 => x"52555372",
          3047 => x"3382e0a4",
          3048 => x"08f80534",
          3049 => x"fea53982",
          3050 => x"e0a408f0",
          3051 => x"05335372",
          3052 => x"802e9038",
          3053 => x"82e0a408",
          3054 => x"fc050830",
          3055 => x"82e0a408",
          3056 => x"fc050c82",
          3057 => x"e0a4088c",
          3058 => x"050882e0",
          3059 => x"a408fc05",
          3060 => x"08710c53",
          3061 => x"810b82e0",
          3062 => x"a408ec05",
          3063 => x"0c82e0a4",
          3064 => x"08ec0508",
          3065 => x"82e0980c",
          3066 => x"8b3d0d82",
          3067 => x"e0a40c04",
          3068 => x"f83d0d7a",
          3069 => x"70087056",
          3070 => x"56597480",
          3071 => x"2e80df38",
          3072 => x"8c397715",
          3073 => x"790c8516",
          3074 => x"335480d2",
          3075 => x"39743354",
          3076 => x"73a02e09",
          3077 => x"81068638",
          3078 => x"811555f1",
          3079 => x"39805776",
          3080 => x"902982db",
          3081 => x"a0057008",
          3082 => x"5256dc8d",
          3083 => x"3f82e098",
          3084 => x"0882e098",
          3085 => x"08547553",
          3086 => x"76085258",
          3087 => x"df883f82",
          3088 => x"e098088b",
          3089 => x"38841633",
          3090 => x"5473812e",
          3091 => x"ffb43881",
          3092 => x"177081ff",
          3093 => x"06585498",
          3094 => x"7727c438",
          3095 => x"ff547382",
          3096 => x"e0980c8a",
          3097 => x"3d0d0481",
          3098 => x"a00b82e0",
          3099 => x"980c04ff",
          3100 => x"3d0d7352",
          3101 => x"71932681",
          3102 => x"8e387184",
          3103 => x"2982b7fc",
          3104 => x"05527108",
          3105 => x"0482bde4",
          3106 => x"51818039",
          3107 => x"82bdf051",
          3108 => x"80f93982",
          3109 => x"be805180",
          3110 => x"f23982be",
          3111 => x"905180eb",
          3112 => x"3982bea0",
          3113 => x"5180e439",
          3114 => x"82beb051",
          3115 => x"80dd3982",
          3116 => x"bec45180",
          3117 => x"d63982be",
          3118 => x"d45180cf",
          3119 => x"3982beec",
          3120 => x"5180c839",
          3121 => x"82bf8451",
          3122 => x"80c13982",
          3123 => x"bf9c51bb",
          3124 => x"3982bfb8",
          3125 => x"51b53982",
          3126 => x"bfcc51af",
          3127 => x"3982bff4",
          3128 => x"51a93982",
          3129 => x"c08451a3",
          3130 => x"3982c0a4",
          3131 => x"519d3982",
          3132 => x"c0b45197",
          3133 => x"3982c0cc",
          3134 => x"51913982",
          3135 => x"c0e4518b",
          3136 => x"3982c0fc",
          3137 => x"51853982",
          3138 => x"c18851ce",
          3139 => x"8a3f833d",
          3140 => x"0d04fb3d",
          3141 => x"0d777956",
          3142 => x"567487e7",
          3143 => x"268a3874",
          3144 => x"527587e8",
          3145 => x"29519039",
          3146 => x"87e85274",
          3147 => x"51e3a43f",
          3148 => x"82e09808",
          3149 => x"527551e3",
          3150 => x"9a3f82e0",
          3151 => x"98085479",
          3152 => x"53755282",
          3153 => x"c19851ff",
          3154 => x"b1c23f87",
          3155 => x"3d0d04ec",
          3156 => x"3d0d6602",
          3157 => x"840580e3",
          3158 => x"05335b57",
          3159 => x"80687830",
          3160 => x"707a0773",
          3161 => x"25515759",
          3162 => x"59785677",
          3163 => x"87ff2683",
          3164 => x"38815674",
          3165 => x"76077081",
          3166 => x"ff065155",
          3167 => x"93567481",
          3168 => x"82388153",
          3169 => x"76528c3d",
          3170 => x"70525681",
          3171 => x"93993f82",
          3172 => x"e0980857",
          3173 => x"82e09808",
          3174 => x"b93882e0",
          3175 => x"980887c0",
          3176 => x"98880c82",
          3177 => x"e0980859",
          3178 => x"963dd405",
          3179 => x"54848053",
          3180 => x"77527551",
          3181 => x"8197d53f",
          3182 => x"82e09808",
          3183 => x"5782e098",
          3184 => x"0890387a",
          3185 => x"5574802e",
          3186 => x"89387419",
          3187 => x"75195959",
          3188 => x"d739963d",
          3189 => x"d8055181",
          3190 => x"9fcd3f76",
          3191 => x"30707807",
          3192 => x"80257b30",
          3193 => x"709f2a72",
          3194 => x"06515751",
          3195 => x"5674802e",
          3196 => x"903882c1",
          3197 => x"bc5387c0",
          3198 => x"98880852",
          3199 => x"7851fe92",
          3200 => x"3f765675",
          3201 => x"82e0980c",
          3202 => x"963d0d04",
          3203 => x"f83d0d7c",
          3204 => x"028405b7",
          3205 => x"05335859",
          3206 => x"ff588053",
          3207 => x"7b527a51",
          3208 => x"fead3f82",
          3209 => x"e09808a8",
          3210 => x"3876802e",
          3211 => x"88387681",
          3212 => x"2e9c389c",
          3213 => x"3982fbf8",
          3214 => x"56615560",
          3215 => x"5482e098",
          3216 => x"537f527e",
          3217 => x"51782d82",
          3218 => x"e0980858",
          3219 => x"83397804",
          3220 => x"7782e098",
          3221 => x"0c8a3d0d",
          3222 => x"04f33d0d",
          3223 => x"7f616302",
          3224 => x"8c0580cf",
          3225 => x"05337373",
          3226 => x"1568415f",
          3227 => x"5d5b5e5e",
          3228 => x"5e77a438",
          3229 => x"fbf13f82",
          3230 => x"e0980881",
          3231 => x"ff065388",
          3232 => x"5872a82e",
          3233 => x"92389058",
          3234 => x"7280d02e",
          3235 => x"8a388639",
          3236 => x"805382d2",
          3237 => x"39a0587a",
          3238 => x"5282c1c4",
          3239 => x"51ffaeec",
          3240 => x"3f82c1cc",
          3241 => x"51ffaee4",
          3242 => x"3f805574",
          3243 => x"78278180",
          3244 => x"387b902e",
          3245 => x"89387ba0",
          3246 => x"2ea73880",
          3247 => x"c6397419",
          3248 => x"53727a27",
          3249 => x"8e387222",
          3250 => x"5282c1d0",
          3251 => x"51ffaebc",
          3252 => x"3f893982",
          3253 => x"c1dc51ff",
          3254 => x"aeb23f82",
          3255 => x"155580c3",
          3256 => x"39741953",
          3257 => x"727a278e",
          3258 => x"38720852",
          3259 => x"82c1c451",
          3260 => x"ffae993f",
          3261 => x"893982c1",
          3262 => x"d851ffae",
          3263 => x"8f3f8415",
          3264 => x"55a13974",
          3265 => x"1953727a",
          3266 => x"278e3872",
          3267 => x"335282c1",
          3268 => x"e451ffad",
          3269 => x"f73f8939",
          3270 => x"82c1ec51",
          3271 => x"ffaded3f",
          3272 => x"81155582",
          3273 => x"fbfc0852",
          3274 => x"a051cdba",
          3275 => x"3ffefc39",
          3276 => x"82c1f051",
          3277 => x"ffadd53f",
          3278 => x"80557478",
          3279 => x"2780c638",
          3280 => x"74197033",
          3281 => x"55538056",
          3282 => x"727a2783",
          3283 => x"38815680",
          3284 => x"539f7427",
          3285 => x"83388153",
          3286 => x"75730670",
          3287 => x"81ff0651",
          3288 => x"5372802e",
          3289 => x"90387380",
          3290 => x"fe268a38",
          3291 => x"82fbfc08",
          3292 => x"52735188",
          3293 => x"3982fbfc",
          3294 => x"0852a051",
          3295 => x"cce83f81",
          3296 => x"1555ffb6",
          3297 => x"3982c1f4",
          3298 => x"51c98c3f",
          3299 => x"7719781c",
          3300 => x"5c598051",
          3301 => x"98e03f82",
          3302 => x"e0980898",
          3303 => x"2b70982c",
          3304 => x"515776a0",
          3305 => x"2e098106",
          3306 => x"ac388051",
          3307 => x"98c83f82",
          3308 => x"e0980898",
          3309 => x"2b70982c",
          3310 => x"70a03270",
          3311 => x"30729b32",
          3312 => x"70307072",
          3313 => x"07737507",
          3314 => x"06515858",
          3315 => x"59575157",
          3316 => x"807324d6",
          3317 => x"38769b2e",
          3318 => x"fdb6387c",
          3319 => x"1e537279",
          3320 => x"26fdb438",
          3321 => x"ff537282",
          3322 => x"e0980c8f",
          3323 => x"3d0d04fc",
          3324 => x"3d0d029b",
          3325 => x"0533558a",
          3326 => x"51cbbe3f",
          3327 => x"82c1f852",
          3328 => x"82c1fc51",
          3329 => x"ffac853f",
          3330 => x"82dee822",
          3331 => x"51a6d83f",
          3332 => x"82c28454",
          3333 => x"82c29053",
          3334 => x"82dee933",
          3335 => x"5282c298",
          3336 => x"51ffabe8",
          3337 => x"3f74802e",
          3338 => x"8438a289",
          3339 => x"3f863d0d",
          3340 => x"04fe3d0d",
          3341 => x"87c09680",
          3342 => x"0853a6f4",
          3343 => x"3f815199",
          3344 => x"bf3f82c2",
          3345 => x"b4519ad4",
          3346 => x"3f805199",
          3347 => x"b33f7281",
          3348 => x"2a708106",
          3349 => x"51527180",
          3350 => x"2e923881",
          3351 => x"5199a13f",
          3352 => x"82c2cc51",
          3353 => x"9ab63f80",
          3354 => x"5199953f",
          3355 => x"72822a70",
          3356 => x"81065152",
          3357 => x"71802e92",
          3358 => x"38815199",
          3359 => x"833f82c2",
          3360 => x"dc519a98",
          3361 => x"3f805198",
          3362 => x"f73f7283",
          3363 => x"2a708106",
          3364 => x"51527180",
          3365 => x"2e923881",
          3366 => x"5198e53f",
          3367 => x"82c2ec51",
          3368 => x"99fa3f80",
          3369 => x"5198d93f",
          3370 => x"72842a70",
          3371 => x"81065152",
          3372 => x"71802e92",
          3373 => x"38815198",
          3374 => x"c73f82c3",
          3375 => x"805199dc",
          3376 => x"3f805198",
          3377 => x"bb3f7285",
          3378 => x"2a708106",
          3379 => x"51527180",
          3380 => x"2e923881",
          3381 => x"5198a93f",
          3382 => x"82c39451",
          3383 => x"99be3f80",
          3384 => x"51989d3f",
          3385 => x"72862a70",
          3386 => x"81065152",
          3387 => x"71802e92",
          3388 => x"38815198",
          3389 => x"8b3f82c3",
          3390 => x"a85199a0",
          3391 => x"3f805197",
          3392 => x"ff3f7287",
          3393 => x"2a708106",
          3394 => x"51527180",
          3395 => x"2e923881",
          3396 => x"5197ed3f",
          3397 => x"82c3bc51",
          3398 => x"99823f80",
          3399 => x"5197e13f",
          3400 => x"72882a70",
          3401 => x"81065152",
          3402 => x"71802e92",
          3403 => x"38815197",
          3404 => x"cf3f82c3",
          3405 => x"d05198e4",
          3406 => x"3f805197",
          3407 => x"c33fa4f8",
          3408 => x"3f843d0d",
          3409 => x"04fb3d0d",
          3410 => x"77028405",
          3411 => x"a3053370",
          3412 => x"55565680",
          3413 => x"527551d9",
          3414 => x"ec3f0b0b",
          3415 => x"82db9c33",
          3416 => x"5473a938",
          3417 => x"815382c4",
          3418 => x"8c5282f7",
          3419 => x"a851818b",
          3420 => x"b63f82e0",
          3421 => x"98083070",
          3422 => x"82e09808",
          3423 => x"07802582",
          3424 => x"71315151",
          3425 => x"54730b0b",
          3426 => x"82db9c34",
          3427 => x"0b0b82db",
          3428 => x"9c335473",
          3429 => x"812e0981",
          3430 => x"06af3882",
          3431 => x"f7a85374",
          3432 => x"52755181",
          3433 => x"c7af3f82",
          3434 => x"e0980880",
          3435 => x"2e8b3882",
          3436 => x"e0980851",
          3437 => x"c4e13f91",
          3438 => x"3982f7a8",
          3439 => x"518197e7",
          3440 => x"3f820b0b",
          3441 => x"0b82db9c",
          3442 => x"340b0b82",
          3443 => x"db9c3354",
          3444 => x"73822e09",
          3445 => x"81068c38",
          3446 => x"82c49c53",
          3447 => x"74527551",
          3448 => x"aaf03f80",
          3449 => x"0b82e098",
          3450 => x"0c873d0d",
          3451 => x"04cd3d0d",
          3452 => x"8070415e",
          3453 => x"ff7e82f7",
          3454 => x"a40c5f81",
          3455 => x"527d5180",
          3456 => x"c88a3f82",
          3457 => x"e0980881",
          3458 => x"ff065978",
          3459 => x"7e2e0981",
          3460 => x"06a33897",
          3461 => x"3d598353",
          3462 => x"82c4a852",
          3463 => x"7851d1f9",
          3464 => x"3f7d5378",
          3465 => x"5282e1c4",
          3466 => x"5181899a",
          3467 => x"3f82e098",
          3468 => x"087e2e88",
          3469 => x"3882c4ac",
          3470 => x"518de539",
          3471 => x"8170415e",
          3472 => x"82c4e451",
          3473 => x"ffa7c53f",
          3474 => x"973d7047",
          3475 => x"5a80f852",
          3476 => x"7951fdf1",
          3477 => x"3fb53dff",
          3478 => x"840551f3",
          3479 => x"933f82e0",
          3480 => x"9808902b",
          3481 => x"70902c51",
          3482 => x"597880c2",
          3483 => x"2e87a538",
          3484 => x"7880c224",
          3485 => x"b23878bd",
          3486 => x"2e81d238",
          3487 => x"78bd2490",
          3488 => x"3878802e",
          3489 => x"ffba3878",
          3490 => x"bc2e80da",
          3491 => x"388adc39",
          3492 => x"7880c02e",
          3493 => x"83993878",
          3494 => x"80c02485",
          3495 => x"ce3878bf",
          3496 => x"2e828c38",
          3497 => x"8ac53978",
          3498 => x"80f92e89",
          3499 => x"df387880",
          3500 => x"f9249238",
          3501 => x"7880c32e",
          3502 => x"888d3878",
          3503 => x"80f82e89",
          3504 => x"a7388aa7",
          3505 => x"39788183",
          3506 => x"2e8a8d38",
          3507 => x"78818324",
          3508 => x"8b387881",
          3509 => x"822e89f1",
          3510 => x"388a9039",
          3511 => x"7881852e",
          3512 => x"8a83388a",
          3513 => x"8639b53d",
          3514 => x"ff801153",
          3515 => x"ff840551",
          3516 => x"ecad3f82",
          3517 => x"e0980880",
          3518 => x"2efec538",
          3519 => x"b53dfefc",
          3520 => x"1153ff84",
          3521 => x"0551ec97",
          3522 => x"3f82e098",
          3523 => x"08802efe",
          3524 => x"af38b53d",
          3525 => x"fef81153",
          3526 => x"ff840551",
          3527 => x"ec813f82",
          3528 => x"e0980886",
          3529 => x"3882e098",
          3530 => x"084382c4",
          3531 => x"e851ffa5",
          3532 => x"db3f6464",
          3533 => x"5c5a797b",
          3534 => x"2781ec38",
          3535 => x"6259787a",
          3536 => x"7084055c",
          3537 => x"0c7a7a26",
          3538 => x"f53881db",
          3539 => x"39b53dff",
          3540 => x"801153ff",
          3541 => x"840551eb",
          3542 => x"c63f82e0",
          3543 => x"9808802e",
          3544 => x"fdde38b5",
          3545 => x"3dfefc11",
          3546 => x"53ff8405",
          3547 => x"51ebb03f",
          3548 => x"82e09808",
          3549 => x"802efdc8",
          3550 => x"38b53dfe",
          3551 => x"f81153ff",
          3552 => x"840551eb",
          3553 => x"9a3f82e0",
          3554 => x"9808802e",
          3555 => x"fdb23882",
          3556 => x"c4f851ff",
          3557 => x"a4f63f64",
          3558 => x"5a796427",
          3559 => x"81893862",
          3560 => x"59797081",
          3561 => x"055b3379",
          3562 => x"34628105",
          3563 => x"43eb39b5",
          3564 => x"3dff8011",
          3565 => x"53ff8405",
          3566 => x"51eae43f",
          3567 => x"82e09808",
          3568 => x"802efcfc",
          3569 => x"38b53dfe",
          3570 => x"fc1153ff",
          3571 => x"840551ea",
          3572 => x"ce3f82e0",
          3573 => x"9808802e",
          3574 => x"fce638b5",
          3575 => x"3dfef811",
          3576 => x"53ff8405",
          3577 => x"51eab83f",
          3578 => x"82e09808",
          3579 => x"802efcd0",
          3580 => x"3882c584",
          3581 => x"51ffa494",
          3582 => x"3f645a79",
          3583 => x"6427a838",
          3584 => x"6270337b",
          3585 => x"335e5a5b",
          3586 => x"787c2e92",
          3587 => x"3878557a",
          3588 => x"54793353",
          3589 => x"795282c5",
          3590 => x"9451ffa3",
          3591 => x"ef3f811a",
          3592 => x"63810544",
          3593 => x"5ad5398a",
          3594 => x"51c38e3f",
          3595 => x"fc9239b5",
          3596 => x"3dff8011",
          3597 => x"53ff8405",
          3598 => x"51e9e43f",
          3599 => x"82e09808",
          3600 => x"80df3882",
          3601 => x"defc3359",
          3602 => x"78802e89",
          3603 => x"3882deb4",
          3604 => x"084580cd",
          3605 => x"3982defd",
          3606 => x"33597880",
          3607 => x"2e883882",
          3608 => x"debc0845",
          3609 => x"bc3982de",
          3610 => x"fe335978",
          3611 => x"802e8838",
          3612 => x"82dec408",
          3613 => x"45ab3982",
          3614 => x"deff3359",
          3615 => x"78802e88",
          3616 => x"3882decc",
          3617 => x"08459a39",
          3618 => x"82defa33",
          3619 => x"5978802e",
          3620 => x"883882de",
          3621 => x"d4084589",
          3622 => x"3982dee4",
          3623 => x"08fc8005",
          3624 => x"45b53dfe",
          3625 => x"fc1153ff",
          3626 => x"840551e8",
          3627 => x"f23f82e0",
          3628 => x"980880de",
          3629 => x"3882defc",
          3630 => x"33597880",
          3631 => x"2e893882",
          3632 => x"deb80844",
          3633 => x"80cc3982",
          3634 => x"defd3359",
          3635 => x"78802e88",
          3636 => x"3882dec0",
          3637 => x"0844bb39",
          3638 => x"82defe33",
          3639 => x"5978802e",
          3640 => x"883882de",
          3641 => x"c80844aa",
          3642 => x"3982deff",
          3643 => x"33597880",
          3644 => x"2e883882",
          3645 => x"ded00844",
          3646 => x"993982de",
          3647 => x"fa335978",
          3648 => x"802e8838",
          3649 => x"82ded808",
          3650 => x"44883982",
          3651 => x"dee40888",
          3652 => x"0544b53d",
          3653 => x"fef81153",
          3654 => x"ff840551",
          3655 => x"e8813f82",
          3656 => x"e0980880",
          3657 => x"2ea73880",
          3658 => x"635c5c7a",
          3659 => x"882e8338",
          3660 => x"815c7a90",
          3661 => x"32703070",
          3662 => x"72079f2a",
          3663 => x"707f0651",
          3664 => x"515a5a78",
          3665 => x"802e8838",
          3666 => x"7aa02e83",
          3667 => x"38884382",
          3668 => x"c5b051ff",
          3669 => x"bdc13f80",
          3670 => x"55645462",
          3671 => x"53635264",
          3672 => x"51f1f63f",
          3673 => x"82c5bc51",
          3674 => x"87b639b5",
          3675 => x"3dff8011",
          3676 => x"53ff8405",
          3677 => x"51e7a83f",
          3678 => x"82e09808",
          3679 => x"802ef9c0",
          3680 => x"38b53dfe",
          3681 => x"fc1153ff",
          3682 => x"840551e7",
          3683 => x"923f82e0",
          3684 => x"9808802e",
          3685 => x"a4386459",
          3686 => x"0280cf05",
          3687 => x"33793464",
          3688 => x"810545b5",
          3689 => x"3dfefc11",
          3690 => x"53ff8405",
          3691 => x"51e6f03f",
          3692 => x"82e09808",
          3693 => x"e138f988",
          3694 => x"39647033",
          3695 => x"545282c5",
          3696 => x"c851ffa0",
          3697 => x"c73f82fb",
          3698 => x"f8085380",
          3699 => x"f8527951",
          3700 => x"ffa18e3f",
          3701 => x"79467933",
          3702 => x"5978ae2e",
          3703 => x"f8e2389f",
          3704 => x"79279f38",
          3705 => x"b53dfefc",
          3706 => x"1153ff84",
          3707 => x"0551e6af",
          3708 => x"3f82e098",
          3709 => x"08802e91",
          3710 => x"38645902",
          3711 => x"80cf0533",
          3712 => x"79346481",
          3713 => x"0545ffb1",
          3714 => x"3982c5d4",
          3715 => x"51ffbc87",
          3716 => x"3fffa639",
          3717 => x"b53dfef4",
          3718 => x"1153ff84",
          3719 => x"0551e0ae",
          3720 => x"3f82e098",
          3721 => x"08802ef8",
          3722 => x"9738b53d",
          3723 => x"fef01153",
          3724 => x"ff840551",
          3725 => x"e0983f82",
          3726 => x"e0980880",
          3727 => x"2ea63861",
          3728 => x"590280c2",
          3729 => x"05227970",
          3730 => x"82055b23",
          3731 => x"7842b53d",
          3732 => x"fef01153",
          3733 => x"ff840551",
          3734 => x"dff43f82",
          3735 => x"e09808df",
          3736 => x"38f7dd39",
          3737 => x"61702254",
          3738 => x"5282c5d8",
          3739 => x"51ff9f9c",
          3740 => x"3f82fbf8",
          3741 => x"085380f8",
          3742 => x"527951ff",
          3743 => x"9fe33f79",
          3744 => x"46793359",
          3745 => x"78ae2ef7",
          3746 => x"b738789f",
          3747 => x"26873861",
          3748 => x"820542d0",
          3749 => x"39b53dfe",
          3750 => x"f01153ff",
          3751 => x"840551df",
          3752 => x"ad3f82e0",
          3753 => x"9808802e",
          3754 => x"93386159",
          3755 => x"0280c205",
          3756 => x"22797082",
          3757 => x"055b2378",
          3758 => x"42ffa939",
          3759 => x"82c5d451",
          3760 => x"ffbad43f",
          3761 => x"ff9e39b5",
          3762 => x"3dfef411",
          3763 => x"53ff8405",
          3764 => x"51defb3f",
          3765 => x"82e09808",
          3766 => x"802ef6e4",
          3767 => x"38b53dfe",
          3768 => x"f01153ff",
          3769 => x"840551de",
          3770 => x"e53f82e0",
          3771 => x"9808802e",
          3772 => x"a0386161",
          3773 => x"710c5961",
          3774 => x"840542b5",
          3775 => x"3dfef011",
          3776 => x"53ff8405",
          3777 => x"51dec73f",
          3778 => x"82e09808",
          3779 => x"e538f6b0",
          3780 => x"39617008",
          3781 => x"545282c5",
          3782 => x"e451ff9d",
          3783 => x"ef3f82fb",
          3784 => x"f8085380",
          3785 => x"f8527951",
          3786 => x"ff9eb63f",
          3787 => x"79467933",
          3788 => x"5978ae2e",
          3789 => x"f68a389f",
          3790 => x"79279b38",
          3791 => x"b53dfef0",
          3792 => x"1153ff84",
          3793 => x"0551de86",
          3794 => x"3f82e098",
          3795 => x"08802e8d",
          3796 => x"38616171",
          3797 => x"0c596184",
          3798 => x"0542ffb5",
          3799 => x"3982c5d4",
          3800 => x"51ffb9b3",
          3801 => x"3fffaa39",
          3802 => x"b53dff80",
          3803 => x"1153ff84",
          3804 => x"0551e3ab",
          3805 => x"3f82e098",
          3806 => x"08802ef5",
          3807 => x"c3386452",
          3808 => x"82c5f451",
          3809 => x"ff9d853f",
          3810 => x"64597804",
          3811 => x"b53dff80",
          3812 => x"1153ff84",
          3813 => x"0551e387",
          3814 => x"3f82e098",
          3815 => x"08802ef5",
          3816 => x"9f386452",
          3817 => x"82c69051",
          3818 => x"ff9ce13f",
          3819 => x"6459782d",
          3820 => x"82e09808",
          3821 => x"802ef588",
          3822 => x"3882e098",
          3823 => x"085282c6",
          3824 => x"ac51ff9c",
          3825 => x"c73ff4f8",
          3826 => x"3982c6c8",
          3827 => x"51ffb8c7",
          3828 => x"3fff9c99",
          3829 => x"3ff4e939",
          3830 => x"82c6e451",
          3831 => x"ffb8b83f",
          3832 => x"8059ffa6",
          3833 => x"3992ce3f",
          3834 => x"f4d63997",
          3835 => x"3d335978",
          3836 => x"802ef4cc",
          3837 => x"3880f852",
          3838 => x"7951c9f1",
          3839 => x"3f82e098",
          3840 => x"085d82e0",
          3841 => x"9808802e",
          3842 => x"82923882",
          3843 => x"e0980846",
          3844 => x"b53dff84",
          3845 => x"055183cc",
          3846 => x"3f82e098",
          3847 => x"08607f06",
          3848 => x"5a5c7880",
          3849 => x"2e81d238",
          3850 => x"82e09808",
          3851 => x"51c48a3f",
          3852 => x"82e09808",
          3853 => x"8f2681c1",
          3854 => x"38815b7a",
          3855 => x"822eb238",
          3856 => x"7a822489",
          3857 => x"387a812e",
          3858 => x"8c3880ca",
          3859 => x"397a832e",
          3860 => x"ad3880c2",
          3861 => x"3982c6f8",
          3862 => x"567b5582",
          3863 => x"c6fc5480",
          3864 => x"5382c780",
          3865 => x"52b53dff",
          3866 => x"b00551ff",
          3867 => x"9e863fb8",
          3868 => x"397b52b5",
          3869 => x"3dffb005",
          3870 => x"51c4ac3f",
          3871 => x"ab397b55",
          3872 => x"82c6fc54",
          3873 => x"805382c7",
          3874 => x"9052b53d",
          3875 => x"ffb00551",
          3876 => x"ff9de13f",
          3877 => x"93397b54",
          3878 => x"805382c7",
          3879 => x"9c52b53d",
          3880 => x"ffb00551",
          3881 => x"ff9dcd3f",
          3882 => x"82deb458",
          3883 => x"82e0c857",
          3884 => x"7c566555",
          3885 => x"80549080",
          3886 => x"0a539080",
          3887 => x"0a52b53d",
          3888 => x"ffb00551",
          3889 => x"eac63f82",
          3890 => x"e0980882",
          3891 => x"e0980809",
          3892 => x"70307072",
          3893 => x"07802551",
          3894 => x"5b5b5f80",
          3895 => x"5a7a8326",
          3896 => x"8338815a",
          3897 => x"787a0659",
          3898 => x"78802e8d",
          3899 => x"38811b70",
          3900 => x"81ff065c",
          3901 => x"597afec3",
          3902 => x"387f8132",
          3903 => x"7e813207",
          3904 => x"59788938",
          3905 => x"7eff2e09",
          3906 => x"81068938",
          3907 => x"82c7a451",
          3908 => x"ffb6843f",
          3909 => x"7c51b1f1",
          3910 => x"3ff2a539",
          3911 => x"82c7b451",
          3912 => x"ffb5f43f",
          3913 => x"f29a39f5",
          3914 => x"3d0d800b",
          3915 => x"82e0c834",
          3916 => x"87c0948c",
          3917 => x"70085455",
          3918 => x"87848052",
          3919 => x"7251cb93",
          3920 => x"3f82e098",
          3921 => x"08902b75",
          3922 => x"08555387",
          3923 => x"84805273",
          3924 => x"51cb803f",
          3925 => x"7282e098",
          3926 => x"0807750c",
          3927 => x"87c0949c",
          3928 => x"70085455",
          3929 => x"87848052",
          3930 => x"7251cae7",
          3931 => x"3f82e098",
          3932 => x"08902b75",
          3933 => x"08555387",
          3934 => x"84805273",
          3935 => x"51cad43f",
          3936 => x"7282e098",
          3937 => x"0807750c",
          3938 => x"8c80830b",
          3939 => x"87c09484",
          3940 => x"0c8c8083",
          3941 => x"0b87c094",
          3942 => x"940c8182",
          3943 => x"985a8185",
          3944 => x"845b8302",
          3945 => x"84059905",
          3946 => x"34805c82",
          3947 => x"fbf80b87",
          3948 => x"3d708813",
          3949 => x"0c70720c",
          3950 => x"82fbfc0c",
          3951 => x"548aaa3f",
          3952 => x"93ee3f82",
          3953 => x"c7e051ff",
          3954 => x"b4cd3f82",
          3955 => x"c7ec51ff",
          3956 => x"b4c53f80",
          3957 => x"e8b15193",
          3958 => x"d23f8151",
          3959 => x"ec913ff0",
          3960 => x"8c3f8004",
          3961 => x"fc3d0d76",
          3962 => x"70085455",
          3963 => x"80735254",
          3964 => x"72742e81",
          3965 => x"8a387233",
          3966 => x"5170a02e",
          3967 => x"09810686",
          3968 => x"38811353",
          3969 => x"f1397233",
          3970 => x"5170a22e",
          3971 => x"09810686",
          3972 => x"38811353",
          3973 => x"81547252",
          3974 => x"73812e09",
          3975 => x"81069f38",
          3976 => x"84398112",
          3977 => x"52807233",
          3978 => x"525470a2",
          3979 => x"2e833881",
          3980 => x"5470802e",
          3981 => x"9d3873ea",
          3982 => x"38983981",
          3983 => x"12528072",
          3984 => x"33525470",
          3985 => x"a02e8338",
          3986 => x"81547080",
          3987 => x"2e843873",
          3988 => x"ea388072",
          3989 => x"33525470",
          3990 => x"a02e0981",
          3991 => x"06833881",
          3992 => x"5470a232",
          3993 => x"70307080",
          3994 => x"25760751",
          3995 => x"51517080",
          3996 => x"2e883880",
          3997 => x"72708105",
          3998 => x"54347175",
          3999 => x"0c725170",
          4000 => x"82e0980c",
          4001 => x"863d0d04",
          4002 => x"fc3d0d76",
          4003 => x"53720880",
          4004 => x"2e913886",
          4005 => x"3dfc0552",
          4006 => x"7251d7b2",
          4007 => x"3f82e098",
          4008 => x"08853880",
          4009 => x"53833974",
          4010 => x"537282e0",
          4011 => x"980c863d",
          4012 => x"0d04fc3d",
          4013 => x"0d768211",
          4014 => x"33ff0552",
          4015 => x"53815270",
          4016 => x"8b268198",
          4017 => x"38831333",
          4018 => x"ff055182",
          4019 => x"52709e26",
          4020 => x"818a3884",
          4021 => x"13335183",
          4022 => x"52709726",
          4023 => x"80fe3885",
          4024 => x"13335184",
          4025 => x"5270bb26",
          4026 => x"80f23886",
          4027 => x"13335185",
          4028 => x"5270bb26",
          4029 => x"80e63888",
          4030 => x"13225586",
          4031 => x"527487e7",
          4032 => x"2680d938",
          4033 => x"8a132254",
          4034 => x"87527387",
          4035 => x"e72680cc",
          4036 => x"38810b87",
          4037 => x"c0989c0c",
          4038 => x"722287c0",
          4039 => x"98bc0c82",
          4040 => x"133387c0",
          4041 => x"98b80c83",
          4042 => x"133387c0",
          4043 => x"98b40c84",
          4044 => x"133387c0",
          4045 => x"98b00c85",
          4046 => x"133387c0",
          4047 => x"98ac0c86",
          4048 => x"133387c0",
          4049 => x"98a80c74",
          4050 => x"87c098a4",
          4051 => x"0c7387c0",
          4052 => x"98a00c80",
          4053 => x"0b87c098",
          4054 => x"9c0c8052",
          4055 => x"7182e098",
          4056 => x"0c863d0d",
          4057 => x"04f33d0d",
          4058 => x"7f5b87c0",
          4059 => x"989c5d81",
          4060 => x"7d0c87c0",
          4061 => x"98bc085e",
          4062 => x"7d7b2387",
          4063 => x"c098b808",
          4064 => x"5a79821c",
          4065 => x"3487c098",
          4066 => x"b4085a79",
          4067 => x"831c3487",
          4068 => x"c098b008",
          4069 => x"5a79841c",
          4070 => x"3487c098",
          4071 => x"ac085a79",
          4072 => x"851c3487",
          4073 => x"c098a808",
          4074 => x"5a79861c",
          4075 => x"3487c098",
          4076 => x"a4085c7b",
          4077 => x"881c2387",
          4078 => x"c098a008",
          4079 => x"5a798a1c",
          4080 => x"23807d0c",
          4081 => x"7983ffff",
          4082 => x"06597b83",
          4083 => x"ffff0658",
          4084 => x"861b3357",
          4085 => x"851b3356",
          4086 => x"841b3355",
          4087 => x"831b3354",
          4088 => x"821b3353",
          4089 => x"7d83ffff",
          4090 => x"065282c8",
          4091 => x"8451ff94",
          4092 => x"9b3f8f3d",
          4093 => x"0d04fd3d",
          4094 => x"0d029705",
          4095 => x"33538052",
          4096 => x"72812e09",
          4097 => x"81068338",
          4098 => x"72527283",
          4099 => x"32703070",
          4100 => x"80257407",
          4101 => x"51515170",
          4102 => x"802e8638",
          4103 => x"84973f84",
          4104 => x"3984f03f",
          4105 => x"82e09808",
          4106 => x"982b7098",
          4107 => x"2c515271",
          4108 => x"ff2e0981",
          4109 => x"069e3880",
          4110 => x"5472812e",
          4111 => x"09810683",
          4112 => x"38725472",
          4113 => x"83327030",
          4114 => x"70802576",
          4115 => x"07515151",
          4116 => x"70ffab38",
          4117 => x"7182e098",
          4118 => x"0c853d0d",
          4119 => x"04fd3d0d",
          4120 => x"80538354",
          4121 => x"72882b53",
          4122 => x"8151ff8a",
          4123 => x"3f82e098",
          4124 => x"08982b70",
          4125 => x"982c7407",
          4126 => x"ff165654",
          4127 => x"52738025",
          4128 => x"e3387282",
          4129 => x"e0980c85",
          4130 => x"3d0d04fb",
          4131 => x"3d0d029f",
          4132 => x"053382de",
          4133 => x"b0337081",
          4134 => x"ff065855",
          4135 => x"5587c094",
          4136 => x"84517580",
          4137 => x"2e863887",
          4138 => x"c0949451",
          4139 => x"70087096",
          4140 => x"2a708106",
          4141 => x"53545270",
          4142 => x"802e8c38",
          4143 => x"71912a70",
          4144 => x"81065151",
          4145 => x"70d73872",
          4146 => x"81327081",
          4147 => x"06515170",
          4148 => x"802e8d38",
          4149 => x"71932a70",
          4150 => x"81065151",
          4151 => x"70ffbe38",
          4152 => x"7381ff06",
          4153 => x"5187c094",
          4154 => x"80527080",
          4155 => x"2e863887",
          4156 => x"c0949052",
          4157 => x"74720c74",
          4158 => x"82e0980c",
          4159 => x"873d0d04",
          4160 => x"ff3d0d02",
          4161 => x"8f053370",
          4162 => x"30709f2a",
          4163 => x"51525270",
          4164 => x"82deb034",
          4165 => x"833d0d04",
          4166 => x"f93d0d02",
          4167 => x"a7053358",
          4168 => x"778a2e09",
          4169 => x"81068738",
          4170 => x"7a528d51",
          4171 => x"eb3f82de",
          4172 => x"b0337081",
          4173 => x"ff065856",
          4174 => x"87c09484",
          4175 => x"5376802e",
          4176 => x"863887c0",
          4177 => x"94945372",
          4178 => x"0870962a",
          4179 => x"70810655",
          4180 => x"56547280",
          4181 => x"2e8c3873",
          4182 => x"912a7081",
          4183 => x"06515372",
          4184 => x"d7387481",
          4185 => x"32708106",
          4186 => x"51537280",
          4187 => x"2e8d3873",
          4188 => x"932a7081",
          4189 => x"06515372",
          4190 => x"ffbe3875",
          4191 => x"81ff0653",
          4192 => x"87c09480",
          4193 => x"5472802e",
          4194 => x"863887c0",
          4195 => x"94905477",
          4196 => x"740c800b",
          4197 => x"82e0980c",
          4198 => x"893d0d04",
          4199 => x"f93d0d79",
          4200 => x"54807433",
          4201 => x"7081ff06",
          4202 => x"53535770",
          4203 => x"772e80fc",
          4204 => x"387181ff",
          4205 => x"06811582",
          4206 => x"deb03370",
          4207 => x"81ff0659",
          4208 => x"57555887",
          4209 => x"c0948451",
          4210 => x"75802e86",
          4211 => x"3887c094",
          4212 => x"94517008",
          4213 => x"70962a70",
          4214 => x"81065354",
          4215 => x"5270802e",
          4216 => x"8c387191",
          4217 => x"2a708106",
          4218 => x"515170d7",
          4219 => x"38728132",
          4220 => x"70810651",
          4221 => x"5170802e",
          4222 => x"8d387193",
          4223 => x"2a708106",
          4224 => x"515170ff",
          4225 => x"be387481",
          4226 => x"ff065187",
          4227 => x"c0948052",
          4228 => x"70802e86",
          4229 => x"3887c094",
          4230 => x"90527772",
          4231 => x"0c811774",
          4232 => x"337081ff",
          4233 => x"06535357",
          4234 => x"70ff8638",
          4235 => x"7682e098",
          4236 => x"0c893d0d",
          4237 => x"04fe3d0d",
          4238 => x"82deb033",
          4239 => x"7081ff06",
          4240 => x"545287c0",
          4241 => x"94845172",
          4242 => x"802e8638",
          4243 => x"87c09494",
          4244 => x"51700870",
          4245 => x"822a7081",
          4246 => x"06515151",
          4247 => x"70802ee2",
          4248 => x"387181ff",
          4249 => x"065187c0",
          4250 => x"94805270",
          4251 => x"802e8638",
          4252 => x"87c09490",
          4253 => x"52710870",
          4254 => x"81ff0682",
          4255 => x"e0980c51",
          4256 => x"843d0d04",
          4257 => x"ffaf3f82",
          4258 => x"e0980881",
          4259 => x"ff0682e0",
          4260 => x"980c04fe",
          4261 => x"3d0d82de",
          4262 => x"b0337081",
          4263 => x"ff065253",
          4264 => x"87c09484",
          4265 => x"5270802e",
          4266 => x"863887c0",
          4267 => x"94945271",
          4268 => x"0870822a",
          4269 => x"70810651",
          4270 => x"5151ff52",
          4271 => x"70802ea0",
          4272 => x"387281ff",
          4273 => x"065187c0",
          4274 => x"94805270",
          4275 => x"802e8638",
          4276 => x"87c09490",
          4277 => x"52710870",
          4278 => x"982b7098",
          4279 => x"2c515351",
          4280 => x"7182e098",
          4281 => x"0c843d0d",
          4282 => x"04ff3d0d",
          4283 => x"87c09e80",
          4284 => x"08709c2a",
          4285 => x"8a065151",
          4286 => x"70802e84",
          4287 => x"b43887c0",
          4288 => x"9ea40882",
          4289 => x"deb40c87",
          4290 => x"c09ea808",
          4291 => x"82deb80c",
          4292 => x"87c09e94",
          4293 => x"0882debc",
          4294 => x"0c87c09e",
          4295 => x"980882de",
          4296 => x"c00c87c0",
          4297 => x"9e9c0882",
          4298 => x"dec40c87",
          4299 => x"c09ea008",
          4300 => x"82dec80c",
          4301 => x"87c09eac",
          4302 => x"0882decc",
          4303 => x"0c87c09e",
          4304 => x"b00882de",
          4305 => x"d00c87c0",
          4306 => x"9eb40882",
          4307 => x"ded40c87",
          4308 => x"c09eb808",
          4309 => x"82ded80c",
          4310 => x"87c09ebc",
          4311 => x"0882dedc",
          4312 => x"0c87c09e",
          4313 => x"c00882de",
          4314 => x"e00c87c0",
          4315 => x"9ec40882",
          4316 => x"dee40c87",
          4317 => x"c09e8008",
          4318 => x"517082de",
          4319 => x"e82387c0",
          4320 => x"9e840882",
          4321 => x"deec0c87",
          4322 => x"c09e8808",
          4323 => x"82def00c",
          4324 => x"87c09e8c",
          4325 => x"0882def4",
          4326 => x"0c810b82",
          4327 => x"def83480",
          4328 => x"0b87c09e",
          4329 => x"90087084",
          4330 => x"800a0651",
          4331 => x"52527080",
          4332 => x"2e833881",
          4333 => x"527182de",
          4334 => x"f934800b",
          4335 => x"87c09e90",
          4336 => x"08708880",
          4337 => x"0a065152",
          4338 => x"5270802e",
          4339 => x"83388152",
          4340 => x"7182defa",
          4341 => x"34800b87",
          4342 => x"c09e9008",
          4343 => x"7090800a",
          4344 => x"06515252",
          4345 => x"70802e83",
          4346 => x"38815271",
          4347 => x"82defb34",
          4348 => x"800b87c0",
          4349 => x"9e900870",
          4350 => x"88808006",
          4351 => x"51525270",
          4352 => x"802e8338",
          4353 => x"81527182",
          4354 => x"defc3480",
          4355 => x"0b87c09e",
          4356 => x"900870a0",
          4357 => x"80800651",
          4358 => x"52527080",
          4359 => x"2e833881",
          4360 => x"527182de",
          4361 => x"fd34800b",
          4362 => x"87c09e90",
          4363 => x"08709080",
          4364 => x"80065152",
          4365 => x"5270802e",
          4366 => x"83388152",
          4367 => x"7182defe",
          4368 => x"34800b87",
          4369 => x"c09e9008",
          4370 => x"70848080",
          4371 => x"06515252",
          4372 => x"70802e83",
          4373 => x"38815271",
          4374 => x"82deff34",
          4375 => x"800b87c0",
          4376 => x"9e900870",
          4377 => x"82808006",
          4378 => x"51525270",
          4379 => x"802e8338",
          4380 => x"81527182",
          4381 => x"df803480",
          4382 => x"0b87c09e",
          4383 => x"90087081",
          4384 => x"80800651",
          4385 => x"52527080",
          4386 => x"2e833881",
          4387 => x"527182df",
          4388 => x"8134800b",
          4389 => x"87c09e90",
          4390 => x"087080c0",
          4391 => x"80065152",
          4392 => x"5270802e",
          4393 => x"83388152",
          4394 => x"7182df82",
          4395 => x"34800b87",
          4396 => x"c09e9008",
          4397 => x"70a08006",
          4398 => x"51525270",
          4399 => x"802e8338",
          4400 => x"81527182",
          4401 => x"df833487",
          4402 => x"c09e9008",
          4403 => x"70988006",
          4404 => x"708a2a51",
          4405 => x"51517082",
          4406 => x"df843480",
          4407 => x"0b87c09e",
          4408 => x"90087084",
          4409 => x"80065152",
          4410 => x"5270802e",
          4411 => x"83388152",
          4412 => x"7182df85",
          4413 => x"3487c09e",
          4414 => x"90087083",
          4415 => x"f0067084",
          4416 => x"2a515151",
          4417 => x"7082df86",
          4418 => x"34800b87",
          4419 => x"c09e9008",
          4420 => x"70880651",
          4421 => x"52527080",
          4422 => x"2e833881",
          4423 => x"527182df",
          4424 => x"873487c0",
          4425 => x"9e900870",
          4426 => x"87065151",
          4427 => x"7082df88",
          4428 => x"34833d0d",
          4429 => x"04fb3d0d",
          4430 => x"82c89c51",
          4431 => x"ff89cd3f",
          4432 => x"82def833",
          4433 => x"5473802e",
          4434 => x"893882c8",
          4435 => x"b051ff89",
          4436 => x"bb3f82c8",
          4437 => x"c451ffa5",
          4438 => x"be3f82de",
          4439 => x"fa335473",
          4440 => x"802e9438",
          4441 => x"82ded408",
          4442 => x"82ded808",
          4443 => x"11545282",
          4444 => x"c8dc51ff",
          4445 => x"89963f82",
          4446 => x"deff3354",
          4447 => x"73802e94",
          4448 => x"3882decc",
          4449 => x"0882ded0",
          4450 => x"08115452",
          4451 => x"82c8f851",
          4452 => x"ff88f93f",
          4453 => x"82defc33",
          4454 => x"5473802e",
          4455 => x"943882de",
          4456 => x"b40882de",
          4457 => x"b8081154",
          4458 => x"5282c994",
          4459 => x"51ff88dc",
          4460 => x"3f82defd",
          4461 => x"33547380",
          4462 => x"2e943882",
          4463 => x"debc0882",
          4464 => x"dec00811",
          4465 => x"545282c9",
          4466 => x"b051ff88",
          4467 => x"bf3f82de",
          4468 => x"fe335473",
          4469 => x"802e9438",
          4470 => x"82dec408",
          4471 => x"82dec808",
          4472 => x"11545282",
          4473 => x"c9cc51ff",
          4474 => x"88a23f82",
          4475 => x"df833354",
          4476 => x"73802e8e",
          4477 => x"3882df84",
          4478 => x"335282c9",
          4479 => x"e851ff88",
          4480 => x"8b3f82df",
          4481 => x"87335473",
          4482 => x"802e8e38",
          4483 => x"82df8833",
          4484 => x"5282ca88",
          4485 => x"51ff87f4",
          4486 => x"3f82df85",
          4487 => x"33547380",
          4488 => x"2e8e3882",
          4489 => x"df863352",
          4490 => x"82caa851",
          4491 => x"ff87dd3f",
          4492 => x"82def933",
          4493 => x"5473802e",
          4494 => x"893882ca",
          4495 => x"c851ffa3",
          4496 => x"d63f82de",
          4497 => x"fb335473",
          4498 => x"802e8938",
          4499 => x"82cadc51",
          4500 => x"ffa3c43f",
          4501 => x"82df8033",
          4502 => x"5473802e",
          4503 => x"893882ca",
          4504 => x"e851ffa3",
          4505 => x"b23f82df",
          4506 => x"81335473",
          4507 => x"802e8938",
          4508 => x"82caf451",
          4509 => x"ffa3a03f",
          4510 => x"82df8233",
          4511 => x"5473802e",
          4512 => x"893882ca",
          4513 => x"fc51ffa3",
          4514 => x"8e3f82cb",
          4515 => x"8451ffa3",
          4516 => x"863f82de",
          4517 => x"dc085282",
          4518 => x"cb9051ff",
          4519 => x"86ee3f82",
          4520 => x"dee00852",
          4521 => x"82cbb851",
          4522 => x"ff86e13f",
          4523 => x"82dee408",
          4524 => x"5282cbe0",
          4525 => x"51ff86d4",
          4526 => x"3f82cc88",
          4527 => x"51ffa2d7",
          4528 => x"3f82dee8",
          4529 => x"225282cc",
          4530 => x"9051ff86",
          4531 => x"bf3f82de",
          4532 => x"ec0856bd",
          4533 => x"84c05275",
          4534 => x"51ffb7f7",
          4535 => x"3f82e098",
          4536 => x"08bd84c0",
          4537 => x"29767131",
          4538 => x"545482e0",
          4539 => x"98085282",
          4540 => x"ccb851ff",
          4541 => x"86963f82",
          4542 => x"deff3354",
          4543 => x"73802eaa",
          4544 => x"3882def0",
          4545 => x"0856bd84",
          4546 => x"c0527551",
          4547 => x"ffb7c43f",
          4548 => x"82e09808",
          4549 => x"bd84c029",
          4550 => x"76713154",
          4551 => x"5482e098",
          4552 => x"085282cc",
          4553 => x"e451ff85",
          4554 => x"e33f82de",
          4555 => x"fa335473",
          4556 => x"802eaa38",
          4557 => x"82def408",
          4558 => x"56bd84c0",
          4559 => x"527551ff",
          4560 => x"b7913f82",
          4561 => x"e09808bd",
          4562 => x"84c02976",
          4563 => x"71315454",
          4564 => x"82e09808",
          4565 => x"5282cd90",
          4566 => x"51ff85b0",
          4567 => x"3f8a51ff",
          4568 => x"a4d73f87",
          4569 => x"3d0d04fe",
          4570 => x"3d0d0292",
          4571 => x"0533ff05",
          4572 => x"52718426",
          4573 => x"aa387184",
          4574 => x"2982b8cc",
          4575 => x"05527108",
          4576 => x"0482cdbc",
          4577 => x"519d3982",
          4578 => x"cdc45197",
          4579 => x"3982cdcc",
          4580 => x"51913982",
          4581 => x"cdd4518b",
          4582 => x"3982cdd8",
          4583 => x"51853982",
          4584 => x"cde051ff",
          4585 => x"84e63f84",
          4586 => x"3d0d0471",
          4587 => x"88800c04",
          4588 => x"800b87c0",
          4589 => x"96840c04",
          4590 => x"82df8c08",
          4591 => x"87c09684",
          4592 => x"0c04fd3d",
          4593 => x"0d76982b",
          4594 => x"70982c79",
          4595 => x"982b7098",
          4596 => x"2c721013",
          4597 => x"70822b51",
          4598 => x"53515451",
          4599 => x"51800b82",
          4600 => x"cdec1233",
          4601 => x"55537174",
          4602 => x"259c3882",
          4603 => x"cde81108",
          4604 => x"12028405",
          4605 => x"97053371",
          4606 => x"33525252",
          4607 => x"70722e09",
          4608 => x"81068338",
          4609 => x"81537282",
          4610 => x"e0980c85",
          4611 => x"3d0d04fb",
          4612 => x"3d0d7902",
          4613 => x"8405a305",
          4614 => x"33713355",
          4615 => x"56547280",
          4616 => x"2eb13882",
          4617 => x"fbfc0852",
          4618 => x"8851ffa3",
          4619 => x"b93f82fb",
          4620 => x"fc0852a0",
          4621 => x"51ffa3ae",
          4622 => x"3f82fbfc",
          4623 => x"08528851",
          4624 => x"ffa3a33f",
          4625 => x"7333ff05",
          4626 => x"53727434",
          4627 => x"7281ff06",
          4628 => x"53cc3977",
          4629 => x"51ff83b4",
          4630 => x"3f747434",
          4631 => x"873d0d04",
          4632 => x"f63d0d7c",
          4633 => x"028405b7",
          4634 => x"05330288",
          4635 => x"05bb0533",
          4636 => x"82dfe833",
          4637 => x"70842982",
          4638 => x"df900570",
          4639 => x"08515959",
          4640 => x"5a585974",
          4641 => x"802e8638",
          4642 => x"74519afd",
          4643 => x"3f82dfe8",
          4644 => x"33708429",
          4645 => x"82df9005",
          4646 => x"81197054",
          4647 => x"58565a9d",
          4648 => x"fe3f82e0",
          4649 => x"9808750c",
          4650 => x"82dfe833",
          4651 => x"70842982",
          4652 => x"df900570",
          4653 => x"0851565a",
          4654 => x"74802ea7",
          4655 => x"38755378",
          4656 => x"527451ff",
          4657 => x"acd33f82",
          4658 => x"dfe83381",
          4659 => x"05557482",
          4660 => x"dfe83474",
          4661 => x"81ff0655",
          4662 => x"93752787",
          4663 => x"38800b82",
          4664 => x"dfe83477",
          4665 => x"802eb638",
          4666 => x"82dfe408",
          4667 => x"5675802e",
          4668 => x"ac3882df",
          4669 => x"e0335574",
          4670 => x"a4388c3d",
          4671 => x"fc055476",
          4672 => x"53785275",
          4673 => x"5180ec84",
          4674 => x"3f82dfe4",
          4675 => x"08528a51",
          4676 => x"81a2d63f",
          4677 => x"82dfe408",
          4678 => x"5180efe8",
          4679 => x"3f8c3d0d",
          4680 => x"04fd3d0d",
          4681 => x"82df9053",
          4682 => x"93547208",
          4683 => x"5271802e",
          4684 => x"89387151",
          4685 => x"99d33f80",
          4686 => x"730cff14",
          4687 => x"84145454",
          4688 => x"738025e6",
          4689 => x"38800b82",
          4690 => x"dfe83482",
          4691 => x"dfe40852",
          4692 => x"71802e95",
          4693 => x"38715180",
          4694 => x"f0cd3f82",
          4695 => x"dfe40851",
          4696 => x"99a73f80",
          4697 => x"0b82dfe4",
          4698 => x"0c853d0d",
          4699 => x"04dc3d0d",
          4700 => x"81578052",
          4701 => x"82dfe408",
          4702 => x"5180f5e9",
          4703 => x"3f82e098",
          4704 => x"0880d338",
          4705 => x"82dfe408",
          4706 => x"5380f852",
          4707 => x"883d7052",
          4708 => x"56819fc1",
          4709 => x"3f82e098",
          4710 => x"08802eba",
          4711 => x"387551ff",
          4712 => x"a9973f82",
          4713 => x"e0980855",
          4714 => x"800b82e0",
          4715 => x"9808259d",
          4716 => x"3882e098",
          4717 => x"08ff0570",
          4718 => x"17555580",
          4719 => x"74347553",
          4720 => x"76528117",
          4721 => x"82d0dc52",
          4722 => x"57ff80c0",
          4723 => x"3f74ff2e",
          4724 => x"098106ff",
          4725 => x"af38a63d",
          4726 => x"0d04d93d",
          4727 => x"0daa3d08",
          4728 => x"ad3d085a",
          4729 => x"5a817058",
          4730 => x"58805282",
          4731 => x"dfe40851",
          4732 => x"80f4f23f",
          4733 => x"82e09808",
          4734 => x"819538ff",
          4735 => x"0b82dfe4",
          4736 => x"08545580",
          4737 => x"f8528b3d",
          4738 => x"70525681",
          4739 => x"9ec73f82",
          4740 => x"e0980880",
          4741 => x"2ea53875",
          4742 => x"51ffa89d",
          4743 => x"3f82e098",
          4744 => x"08811858",
          4745 => x"55800b82",
          4746 => x"e0980825",
          4747 => x"8e3882e0",
          4748 => x"9808ff05",
          4749 => x"70175555",
          4750 => x"80743474",
          4751 => x"09703070",
          4752 => x"72079f2a",
          4753 => x"51555578",
          4754 => x"772e8538",
          4755 => x"73ffac38",
          4756 => x"82dfe408",
          4757 => x"8c110853",
          4758 => x"5180f489",
          4759 => x"3f82e098",
          4760 => x"08802e89",
          4761 => x"3882d0e8",
          4762 => x"51feffa0",
          4763 => x"3f78772e",
          4764 => x"0981069b",
          4765 => x"38755279",
          4766 => x"51ffa8ab",
          4767 => x"3f7951ff",
          4768 => x"a7b73fab",
          4769 => x"3d085482",
          4770 => x"e0980874",
          4771 => x"34805877",
          4772 => x"82e0980c",
          4773 => x"a93d0d04",
          4774 => x"f63d0d7c",
          4775 => x"7e715c71",
          4776 => x"72335759",
          4777 => x"5a5873a0",
          4778 => x"2e098106",
          4779 => x"a2387833",
          4780 => x"78055677",
          4781 => x"76279838",
          4782 => x"8117705b",
          4783 => x"70713356",
          4784 => x"585573a0",
          4785 => x"2e098106",
          4786 => x"86387575",
          4787 => x"26ea3880",
          4788 => x"54738829",
          4789 => x"82dfec05",
          4790 => x"70085255",
          4791 => x"ffa6da3f",
          4792 => x"82e09808",
          4793 => x"53795274",
          4794 => x"0851ffa9",
          4795 => x"d93f82e0",
          4796 => x"980880c5",
          4797 => x"38841533",
          4798 => x"5574812e",
          4799 => x"88387482",
          4800 => x"2e8838b5",
          4801 => x"39fce63f",
          4802 => x"ac39811a",
          4803 => x"5a8c3dfc",
          4804 => x"1153f805",
          4805 => x"51c4883f",
          4806 => x"82e09808",
          4807 => x"802e9a38",
          4808 => x"ff1b5378",
          4809 => x"527751fd",
          4810 => x"b13f82e0",
          4811 => x"980881ff",
          4812 => x"06557485",
          4813 => x"38745491",
          4814 => x"39811470",
          4815 => x"81ff0651",
          4816 => x"54827427",
          4817 => x"ff8b3880",
          4818 => x"547382e0",
          4819 => x"980c8c3d",
          4820 => x"0d04d33d",
          4821 => x"0db03d08",
          4822 => x"b23d08b4",
          4823 => x"3d08595f",
          4824 => x"5a800baf",
          4825 => x"3d3482df",
          4826 => x"e83382df",
          4827 => x"e408555b",
          4828 => x"7381cb38",
          4829 => x"7382dfe0",
          4830 => x"33555573",
          4831 => x"83388155",
          4832 => x"76802e81",
          4833 => x"bc388170",
          4834 => x"76065556",
          4835 => x"73802e81",
          4836 => x"ad38a851",
          4837 => x"98893f82",
          4838 => x"e0980882",
          4839 => x"dfe40c82",
          4840 => x"e0980880",
          4841 => x"2e819238",
          4842 => x"93537652",
          4843 => x"82e09808",
          4844 => x"5180def3",
          4845 => x"3f82e098",
          4846 => x"08802e8c",
          4847 => x"3882d194",
          4848 => x"51ff98d3",
          4849 => x"3f80f739",
          4850 => x"82e09808",
          4851 => x"5b82dfe4",
          4852 => x"085380f8",
          4853 => x"52903d70",
          4854 => x"5254819a",
          4855 => x"f83f82e0",
          4856 => x"98085682",
          4857 => x"e0980874",
          4858 => x"2e098106",
          4859 => x"80d03882",
          4860 => x"e0980851",
          4861 => x"ffa4c23f",
          4862 => x"82e09808",
          4863 => x"55800b82",
          4864 => x"e0980825",
          4865 => x"a93882e0",
          4866 => x"9808ff05",
          4867 => x"70175555",
          4868 => x"80743480",
          4869 => x"537481ff",
          4870 => x"06527551",
          4871 => x"f8c23f81",
          4872 => x"1b7081ff",
          4873 => x"065c5493",
          4874 => x"7b278338",
          4875 => x"805b74ff",
          4876 => x"2e098106",
          4877 => x"ff973886",
          4878 => x"397582df",
          4879 => x"e034768c",
          4880 => x"3882dfe4",
          4881 => x"08802e84",
          4882 => x"38f9d63f",
          4883 => x"8f3d5d80",
          4884 => x"51e7a33f",
          4885 => x"82e09808",
          4886 => x"982b7098",
          4887 => x"2c515978",
          4888 => x"ff2eec38",
          4889 => x"7881ff06",
          4890 => x"82f7d433",
          4891 => x"70982b70",
          4892 => x"982c82f7",
          4893 => x"d0337098",
          4894 => x"2b70972c",
          4895 => x"71982c05",
          4896 => x"70842982",
          4897 => x"cde80570",
          4898 => x"08157033",
          4899 => x"51515151",
          4900 => x"59595159",
          4901 => x"5d588156",
          4902 => x"73782e80",
          4903 => x"e9387774",
          4904 => x"27b43874",
          4905 => x"81800a29",
          4906 => x"81ff0a05",
          4907 => x"70982c51",
          4908 => x"55807524",
          4909 => x"80ce3876",
          4910 => x"53745277",
          4911 => x"51f6833f",
          4912 => x"82e09808",
          4913 => x"81ff0654",
          4914 => x"73802ed7",
          4915 => x"387482f7",
          4916 => x"d0348156",
          4917 => x"b1397481",
          4918 => x"800a2981",
          4919 => x"800a0570",
          4920 => x"982c7081",
          4921 => x"ff065651",
          4922 => x"55739526",
          4923 => x"97387653",
          4924 => x"74527751",
          4925 => x"f5cc3f82",
          4926 => x"e0980881",
          4927 => x"ff065473",
          4928 => x"cc38d339",
          4929 => x"80567580",
          4930 => x"2e80ca38",
          4931 => x"811c5574",
          4932 => x"82f7d434",
          4933 => x"74982b70",
          4934 => x"982c82f7",
          4935 => x"d0337098",
          4936 => x"2b70982c",
          4937 => x"70101170",
          4938 => x"822b82cd",
          4939 => x"ec11335e",
          4940 => x"51515157",
          4941 => x"58515574",
          4942 => x"772e0981",
          4943 => x"06fe9038",
          4944 => x"82cdf014",
          4945 => x"087d0c80",
          4946 => x"0b82f7d4",
          4947 => x"34800b82",
          4948 => x"f7d03492",
          4949 => x"397582f7",
          4950 => x"d4347582",
          4951 => x"f7d03478",
          4952 => x"af3d3475",
          4953 => x"7d0c7e54",
          4954 => x"739526fd",
          4955 => x"df387384",
          4956 => x"2982b8e0",
          4957 => x"05547308",
          4958 => x"0482f7dc",
          4959 => x"3354737e",
          4960 => x"2efdc938",
          4961 => x"82f7d833",
          4962 => x"55737527",
          4963 => x"ab387498",
          4964 => x"2b70982c",
          4965 => x"51557375",
          4966 => x"249e3874",
          4967 => x"1a547333",
          4968 => x"81153474",
          4969 => x"81800a29",
          4970 => x"81ff0a05",
          4971 => x"70982c82",
          4972 => x"f7dc3356",
          4973 => x"5155df39",
          4974 => x"82f7dc33",
          4975 => x"81115654",
          4976 => x"7482f7dc",
          4977 => x"34731a54",
          4978 => x"ae3d3374",
          4979 => x"3482f7d8",
          4980 => x"3354737e",
          4981 => x"25893881",
          4982 => x"14547382",
          4983 => x"f7d83482",
          4984 => x"f7dc3370",
          4985 => x"81800a29",
          4986 => x"81ff0a05",
          4987 => x"70982c82",
          4988 => x"f7d8335a",
          4989 => x"51565674",
          4990 => x"7725a838",
          4991 => x"82fbfc08",
          4992 => x"52741a70",
          4993 => x"335254ff",
          4994 => x"97dc3f74",
          4995 => x"81800a29",
          4996 => x"81800a05",
          4997 => x"70982c82",
          4998 => x"f7d83356",
          4999 => x"51557375",
          5000 => x"24da3882",
          5001 => x"f7dc3370",
          5002 => x"982b7098",
          5003 => x"2c82f7d8",
          5004 => x"335a5156",
          5005 => x"56747725",
          5006 => x"fc923882",
          5007 => x"fbfc0852",
          5008 => x"8851ff97",
          5009 => x"a13f7481",
          5010 => x"800a2981",
          5011 => x"800a0570",
          5012 => x"982c82f7",
          5013 => x"d8335651",
          5014 => x"55737524",
          5015 => x"de38fbec",
          5016 => x"39837a34",
          5017 => x"800b811b",
          5018 => x"3482f7dc",
          5019 => x"53805282",
          5020 => x"c1b851f3",
          5021 => x"9a3f81fd",
          5022 => x"3982f7dc",
          5023 => x"337081ff",
          5024 => x"06555573",
          5025 => x"802efbc4",
          5026 => x"3882f7d8",
          5027 => x"33ff0554",
          5028 => x"7382f7d8",
          5029 => x"34ff1554",
          5030 => x"7382f7dc",
          5031 => x"3482fbfc",
          5032 => x"08528851",
          5033 => x"ff96bf3f",
          5034 => x"82f7dc33",
          5035 => x"70982b70",
          5036 => x"982c82f7",
          5037 => x"d8335751",
          5038 => x"56577474",
          5039 => x"25ad3874",
          5040 => x"1a548114",
          5041 => x"33743482",
          5042 => x"fbfc0852",
          5043 => x"733351ff",
          5044 => x"96943f74",
          5045 => x"81800a29",
          5046 => x"81800a05",
          5047 => x"70982c82",
          5048 => x"f7d83358",
          5049 => x"51557575",
          5050 => x"24d53882",
          5051 => x"fbfc0852",
          5052 => x"a051ff95",
          5053 => x"f13f82f7",
          5054 => x"dc337098",
          5055 => x"2b70982c",
          5056 => x"82f7d833",
          5057 => x"57515657",
          5058 => x"747424fa",
          5059 => x"bf3882fb",
          5060 => x"fc085288",
          5061 => x"51ff95ce",
          5062 => x"3f748180",
          5063 => x"0a298180",
          5064 => x"0a057098",
          5065 => x"2c82f7d8",
          5066 => x"33585155",
          5067 => x"757525de",
          5068 => x"38fa9939",
          5069 => x"82f7d833",
          5070 => x"7a055480",
          5071 => x"743482fb",
          5072 => x"fc08528a",
          5073 => x"51ff959e",
          5074 => x"3f82f7d8",
          5075 => x"527951f6",
          5076 => x"c73f82e0",
          5077 => x"980881ff",
          5078 => x"06547396",
          5079 => x"3882f7d8",
          5080 => x"33547380",
          5081 => x"2e8f3881",
          5082 => x"53735279",
          5083 => x"51f1f13f",
          5084 => x"8439807a",
          5085 => x"34800b82",
          5086 => x"f7dc3480",
          5087 => x"0b82f7d8",
          5088 => x"347982e0",
          5089 => x"980caf3d",
          5090 => x"0d0482f7",
          5091 => x"dc335473",
          5092 => x"802ef9b8",
          5093 => x"3882fbfc",
          5094 => x"08528851",
          5095 => x"ff94c73f",
          5096 => x"82f7dc33",
          5097 => x"ff055473",
          5098 => x"82f7dc34",
          5099 => x"7381ff06",
          5100 => x"54dd3982",
          5101 => x"f7dc3382",
          5102 => x"f7d83355",
          5103 => x"5573752e",
          5104 => x"f98a38ff",
          5105 => x"14547382",
          5106 => x"f7d83474",
          5107 => x"982b7098",
          5108 => x"2c7581ff",
          5109 => x"06565155",
          5110 => x"747425ad",
          5111 => x"38741a54",
          5112 => x"81143374",
          5113 => x"3482fbfc",
          5114 => x"08527333",
          5115 => x"51ff93f6",
          5116 => x"3f748180",
          5117 => x"0a298180",
          5118 => x"0a057098",
          5119 => x"2c82f7d8",
          5120 => x"33585155",
          5121 => x"757524d5",
          5122 => x"3882fbfc",
          5123 => x"0852a051",
          5124 => x"ff93d33f",
          5125 => x"82f7dc33",
          5126 => x"70982b70",
          5127 => x"982c82f7",
          5128 => x"d8335751",
          5129 => x"56577474",
          5130 => x"24f8a138",
          5131 => x"82fbfc08",
          5132 => x"528851ff",
          5133 => x"93b03f74",
          5134 => x"81800a29",
          5135 => x"81800a05",
          5136 => x"70982c82",
          5137 => x"f7d83358",
          5138 => x"51557575",
          5139 => x"25de38f7",
          5140 => x"fb3982f7",
          5141 => x"dc337081",
          5142 => x"ff0682f7",
          5143 => x"d8335956",
          5144 => x"54747727",
          5145 => x"f7e63882",
          5146 => x"fbfc0852",
          5147 => x"81145473",
          5148 => x"82f7dc34",
          5149 => x"741a7033",
          5150 => x"5254ff92",
          5151 => x"e93f82f7",
          5152 => x"dc337081",
          5153 => x"ff0682f7",
          5154 => x"d8335856",
          5155 => x"54757526",
          5156 => x"d638f7b8",
          5157 => x"3982f7dc",
          5158 => x"53805282",
          5159 => x"c1b851ee",
          5160 => x"ee3f800b",
          5161 => x"82f7dc34",
          5162 => x"800b82f7",
          5163 => x"d834f79c",
          5164 => x"397ab038",
          5165 => x"82dfdc08",
          5166 => x"5574802e",
          5167 => x"a6387451",
          5168 => x"ff9af63f",
          5169 => x"82e09808",
          5170 => x"82f7d834",
          5171 => x"82e09808",
          5172 => x"81ff0681",
          5173 => x"05537452",
          5174 => x"7951ff9c",
          5175 => x"bc3f935b",
          5176 => x"81c0397a",
          5177 => x"842982df",
          5178 => x"9005fc11",
          5179 => x"08565474",
          5180 => x"802ea738",
          5181 => x"7451ff9a",
          5182 => x"c03f82e0",
          5183 => x"980882f7",
          5184 => x"d83482e0",
          5185 => x"980881ff",
          5186 => x"06810553",
          5187 => x"74527951",
          5188 => x"ff9c863f",
          5189 => x"ff1b5480",
          5190 => x"fa397308",
          5191 => x"5574802e",
          5192 => x"f6aa3874",
          5193 => x"51ff9a91",
          5194 => x"3f99397a",
          5195 => x"932e0981",
          5196 => x"06ae3882",
          5197 => x"df900855",
          5198 => x"74802ea4",
          5199 => x"387451ff",
          5200 => x"99f73f82",
          5201 => x"e0980882",
          5202 => x"f7d83482",
          5203 => x"e0980881",
          5204 => x"ff068105",
          5205 => x"53745279",
          5206 => x"51ff9bbd",
          5207 => x"3f80c339",
          5208 => x"7a842982",
          5209 => x"df940570",
          5210 => x"08565474",
          5211 => x"802eab38",
          5212 => x"7451ff99",
          5213 => x"c43f82e0",
          5214 => x"980882f7",
          5215 => x"d83482e0",
          5216 => x"980881ff",
          5217 => x"06810553",
          5218 => x"74527951",
          5219 => x"ff9b8a3f",
          5220 => x"811b5473",
          5221 => x"81ff065b",
          5222 => x"89397482",
          5223 => x"f7d83474",
          5224 => x"7a3482f7",
          5225 => x"dc5382f7",
          5226 => x"d8335279",
          5227 => x"51ece03f",
          5228 => x"f59a3982",
          5229 => x"f7dc3370",
          5230 => x"81ff0682",
          5231 => x"f7d83359",
          5232 => x"56547477",
          5233 => x"27f58538",
          5234 => x"82fbfc08",
          5235 => x"52811454",
          5236 => x"7382f7dc",
          5237 => x"34741a70",
          5238 => x"335254ff",
          5239 => x"90883ff4",
          5240 => x"eb3982f7",
          5241 => x"dc335473",
          5242 => x"802ef4e0",
          5243 => x"3882fbfc",
          5244 => x"08528851",
          5245 => x"ff8fef3f",
          5246 => x"82f7dc33",
          5247 => x"ff055473",
          5248 => x"82f7dc34",
          5249 => x"f4c639f9",
          5250 => x"3d0d84fa",
          5251 => x"f40b82e0",
          5252 => x"880ca080",
          5253 => x"0b82e084",
          5254 => x"23828080",
          5255 => x"53805284",
          5256 => x"faf451ff",
          5257 => x"a09f3f82",
          5258 => x"e0880854",
          5259 => x"80587774",
          5260 => x"34815776",
          5261 => x"81153482",
          5262 => x"e0880854",
          5263 => x"77841534",
          5264 => x"76851534",
          5265 => x"82e08808",
          5266 => x"54778615",
          5267 => x"34768715",
          5268 => x"3482e088",
          5269 => x"0882e084",
          5270 => x"22ff05fe",
          5271 => x"80800770",
          5272 => x"83ffff06",
          5273 => x"70882a58",
          5274 => x"51555674",
          5275 => x"88173473",
          5276 => x"89173482",
          5277 => x"e0842270",
          5278 => x"882982e0",
          5279 => x"880805f8",
          5280 => x"11515555",
          5281 => x"77821534",
          5282 => x"76831534",
          5283 => x"893d0d04",
          5284 => x"ff3d0d73",
          5285 => x"52815184",
          5286 => x"72278f38",
          5287 => x"fb12832a",
          5288 => x"82117083",
          5289 => x"ffff0651",
          5290 => x"51517082",
          5291 => x"e0980c83",
          5292 => x"3d0d04f9",
          5293 => x"3d0d02a6",
          5294 => x"05220284",
          5295 => x"05aa0522",
          5296 => x"710582e0",
          5297 => x"88087183",
          5298 => x"2b711174",
          5299 => x"832b7311",
          5300 => x"70338112",
          5301 => x"3371882b",
          5302 => x"0702a405",
          5303 => x"ae052271",
          5304 => x"81ffff06",
          5305 => x"0770882a",
          5306 => x"53515259",
          5307 => x"545b5b57",
          5308 => x"53545571",
          5309 => x"77347081",
          5310 => x"183482e0",
          5311 => x"88081475",
          5312 => x"882a5254",
          5313 => x"70821534",
          5314 => x"74831534",
          5315 => x"82e08808",
          5316 => x"70177033",
          5317 => x"81123371",
          5318 => x"882b0770",
          5319 => x"832b8fff",
          5320 => x"f8065152",
          5321 => x"56527105",
          5322 => x"7383ffff",
          5323 => x"0670882a",
          5324 => x"54545171",
          5325 => x"82123472",
          5326 => x"81ff0653",
          5327 => x"72831234",
          5328 => x"82e08808",
          5329 => x"16567176",
          5330 => x"34728117",
          5331 => x"34893d0d",
          5332 => x"04fb3d0d",
          5333 => x"82e08808",
          5334 => x"0284059e",
          5335 => x"05227083",
          5336 => x"2b721186",
          5337 => x"11338712",
          5338 => x"33718b2b",
          5339 => x"71832b07",
          5340 => x"585b5952",
          5341 => x"55527205",
          5342 => x"84123385",
          5343 => x"13337188",
          5344 => x"2b077088",
          5345 => x"2a545656",
          5346 => x"52708413",
          5347 => x"34738513",
          5348 => x"3482e088",
          5349 => x"08701484",
          5350 => x"11338512",
          5351 => x"33718b2b",
          5352 => x"71832b07",
          5353 => x"56595752",
          5354 => x"72058612",
          5355 => x"33871333",
          5356 => x"71882b07",
          5357 => x"70882a54",
          5358 => x"56565270",
          5359 => x"86133473",
          5360 => x"87133482",
          5361 => x"e0880813",
          5362 => x"70338112",
          5363 => x"3371882b",
          5364 => x"077081ff",
          5365 => x"ff067088",
          5366 => x"2a535153",
          5367 => x"53537173",
          5368 => x"34708114",
          5369 => x"34873d0d",
          5370 => x"04fa3d0d",
          5371 => x"02a20522",
          5372 => x"82e08808",
          5373 => x"71832b71",
          5374 => x"11703381",
          5375 => x"12337188",
          5376 => x"2b077088",
          5377 => x"29157033",
          5378 => x"81123371",
          5379 => x"982b7190",
          5380 => x"2b07535f",
          5381 => x"5355525a",
          5382 => x"56575354",
          5383 => x"71802580",
          5384 => x"f6387251",
          5385 => x"feab3f82",
          5386 => x"e0880870",
          5387 => x"16703381",
          5388 => x"1233718b",
          5389 => x"2b71832b",
          5390 => x"07741170",
          5391 => x"33811233",
          5392 => x"71882b07",
          5393 => x"70832b8f",
          5394 => x"fff80651",
          5395 => x"52545153",
          5396 => x"5a585372",
          5397 => x"0574882a",
          5398 => x"54527282",
          5399 => x"13347383",
          5400 => x"133482e0",
          5401 => x"88087016",
          5402 => x"70338112",
          5403 => x"33718b2b",
          5404 => x"71832b07",
          5405 => x"56595755",
          5406 => x"72057033",
          5407 => x"81123371",
          5408 => x"882b0770",
          5409 => x"81ffff06",
          5410 => x"70882a57",
          5411 => x"51525852",
          5412 => x"72743471",
          5413 => x"81153488",
          5414 => x"3d0d04fb",
          5415 => x"3d0d82e0",
          5416 => x"88080284",
          5417 => x"059e0522",
          5418 => x"70832b72",
          5419 => x"11821133",
          5420 => x"83123371",
          5421 => x"8b2b7183",
          5422 => x"2b07595b",
          5423 => x"59525652",
          5424 => x"73057133",
          5425 => x"81133371",
          5426 => x"882b0702",
          5427 => x"8c05a205",
          5428 => x"22710770",
          5429 => x"882a5351",
          5430 => x"53535371",
          5431 => x"73347081",
          5432 => x"143482e0",
          5433 => x"88087015",
          5434 => x"70338112",
          5435 => x"33718b2b",
          5436 => x"71832b07",
          5437 => x"56595752",
          5438 => x"72058212",
          5439 => x"33831333",
          5440 => x"71882b07",
          5441 => x"70882a54",
          5442 => x"55565270",
          5443 => x"82133472",
          5444 => x"83133482",
          5445 => x"e0880814",
          5446 => x"82113383",
          5447 => x"12337188",
          5448 => x"2b0782e0",
          5449 => x"980c5254",
          5450 => x"873d0d04",
          5451 => x"f73d0d7b",
          5452 => x"82e08808",
          5453 => x"31832a70",
          5454 => x"83ffff06",
          5455 => x"70535753",
          5456 => x"fda73f82",
          5457 => x"e0880876",
          5458 => x"832b7111",
          5459 => x"82113383",
          5460 => x"1233718b",
          5461 => x"2b71832b",
          5462 => x"07751170",
          5463 => x"33811233",
          5464 => x"71982b71",
          5465 => x"902b0753",
          5466 => x"42405153",
          5467 => x"5b585559",
          5468 => x"54728025",
          5469 => x"8d388280",
          5470 => x"80527551",
          5471 => x"fe9d3f81",
          5472 => x"84398414",
          5473 => x"33851533",
          5474 => x"718b2b71",
          5475 => x"832b0776",
          5476 => x"1179882a",
          5477 => x"53515558",
          5478 => x"55768614",
          5479 => x"347581ff",
          5480 => x"06567587",
          5481 => x"143482e0",
          5482 => x"88087019",
          5483 => x"84123385",
          5484 => x"13337188",
          5485 => x"2b077088",
          5486 => x"2a54575b",
          5487 => x"56537284",
          5488 => x"16347385",
          5489 => x"163482e0",
          5490 => x"88081853",
          5491 => x"800b8614",
          5492 => x"34800b87",
          5493 => x"143482e0",
          5494 => x"88085376",
          5495 => x"84143475",
          5496 => x"85143482",
          5497 => x"e0880818",
          5498 => x"70338112",
          5499 => x"3371882b",
          5500 => x"07708280",
          5501 => x"80077088",
          5502 => x"2a535155",
          5503 => x"56547474",
          5504 => x"34728115",
          5505 => x"348b3d0d",
          5506 => x"04ff3d0d",
          5507 => x"735282e0",
          5508 => x"88088438",
          5509 => x"f7f13f71",
          5510 => x"802e8638",
          5511 => x"7151fe8c",
          5512 => x"3f833d0d",
          5513 => x"04f53d0d",
          5514 => x"807e5258",
          5515 => x"f8e23f82",
          5516 => x"e0980883",
          5517 => x"ffff0682",
          5518 => x"e0880884",
          5519 => x"11338512",
          5520 => x"3371882b",
          5521 => x"07705f59",
          5522 => x"56585a81",
          5523 => x"ffff5975",
          5524 => x"782e80cb",
          5525 => x"38758829",
          5526 => x"17703381",
          5527 => x"12337188",
          5528 => x"2b077081",
          5529 => x"ffff0679",
          5530 => x"317083ff",
          5531 => x"ff06707f",
          5532 => x"27525351",
          5533 => x"56595577",
          5534 => x"79278a38",
          5535 => x"73802e85",
          5536 => x"3875785a",
          5537 => x"5b841533",
          5538 => x"85163371",
          5539 => x"882b0757",
          5540 => x"5475c238",
          5541 => x"7881ffff",
          5542 => x"2e85387a",
          5543 => x"79595680",
          5544 => x"76832b82",
          5545 => x"e0880811",
          5546 => x"70338112",
          5547 => x"3371882b",
          5548 => x"077081ff",
          5549 => x"ff065152",
          5550 => x"5a565c55",
          5551 => x"73752e83",
          5552 => x"38815580",
          5553 => x"54797826",
          5554 => x"81cc3874",
          5555 => x"5474802e",
          5556 => x"81c43877",
          5557 => x"7a2e0981",
          5558 => x"06893875",
          5559 => x"51f8f23f",
          5560 => x"81ac3982",
          5561 => x"80805379",
          5562 => x"527551f7",
          5563 => x"c63f82e0",
          5564 => x"8808701c",
          5565 => x"86113387",
          5566 => x"1233718b",
          5567 => x"2b71832b",
          5568 => x"07535a5e",
          5569 => x"5574057a",
          5570 => x"177083ff",
          5571 => x"ff067088",
          5572 => x"2a5c5956",
          5573 => x"54788415",
          5574 => x"347681ff",
          5575 => x"06577685",
          5576 => x"153482e0",
          5577 => x"88087583",
          5578 => x"2b711172",
          5579 => x"1e861133",
          5580 => x"87123371",
          5581 => x"882b0770",
          5582 => x"882a535b",
          5583 => x"5e535a56",
          5584 => x"54738619",
          5585 => x"34758719",
          5586 => x"3482e088",
          5587 => x"08701c84",
          5588 => x"11338512",
          5589 => x"33718b2b",
          5590 => x"71832b07",
          5591 => x"535d5a55",
          5592 => x"74055478",
          5593 => x"86153476",
          5594 => x"87153482",
          5595 => x"e0880870",
          5596 => x"16711d84",
          5597 => x"11338512",
          5598 => x"3371882b",
          5599 => x"0770882a",
          5600 => x"535a5f52",
          5601 => x"56547384",
          5602 => x"16347585",
          5603 => x"163482e0",
          5604 => x"88081b84",
          5605 => x"05547382",
          5606 => x"e0980c8d",
          5607 => x"3d0d04fe",
          5608 => x"3d0d7452",
          5609 => x"82e08808",
          5610 => x"8438f4db",
          5611 => x"3f715371",
          5612 => x"802e8b38",
          5613 => x"7151fced",
          5614 => x"3f82e098",
          5615 => x"08537282",
          5616 => x"e0980c84",
          5617 => x"3d0d04ee",
          5618 => x"3d0d6466",
          5619 => x"405c8070",
          5620 => x"424082e0",
          5621 => x"8808602e",
          5622 => x"09810684",
          5623 => x"38f4a83f",
          5624 => x"7b8e387e",
          5625 => x"51ffb83f",
          5626 => x"82e09808",
          5627 => x"5483c739",
          5628 => x"7e8b387b",
          5629 => x"51fc923f",
          5630 => x"7e5483ba",
          5631 => x"397e51f5",
          5632 => x"8f3f82e0",
          5633 => x"980883ff",
          5634 => x"ff0682e0",
          5635 => x"88087d71",
          5636 => x"31832a70",
          5637 => x"83ffff06",
          5638 => x"70832b73",
          5639 => x"11703381",
          5640 => x"12337188",
          5641 => x"2b077075",
          5642 => x"317083ff",
          5643 => x"ff067088",
          5644 => x"29fc0573",
          5645 => x"88291a70",
          5646 => x"33811233",
          5647 => x"71882b07",
          5648 => x"70902b53",
          5649 => x"444e5348",
          5650 => x"41525c54",
          5651 => x"5b415c56",
          5652 => x"5b5b7380",
          5653 => x"258f3876",
          5654 => x"81ffff06",
          5655 => x"75317083",
          5656 => x"ffff0642",
          5657 => x"54821633",
          5658 => x"83173371",
          5659 => x"882b0770",
          5660 => x"88291c70",
          5661 => x"33811233",
          5662 => x"71982b71",
          5663 => x"902b0753",
          5664 => x"47455256",
          5665 => x"54738025",
          5666 => x"8b387875",
          5667 => x"317083ff",
          5668 => x"ff064154",
          5669 => x"777b2781",
          5670 => x"fe386018",
          5671 => x"54737b2e",
          5672 => x"0981068f",
          5673 => x"387851f6",
          5674 => x"c03f7a83",
          5675 => x"ffff0658",
          5676 => x"81e5397f",
          5677 => x"8e387a74",
          5678 => x"24893878",
          5679 => x"51f6aa3f",
          5680 => x"81a5397f",
          5681 => x"18557a75",
          5682 => x"2480c838",
          5683 => x"791d8211",
          5684 => x"33831233",
          5685 => x"71882b07",
          5686 => x"535754f4",
          5687 => x"f43f8052",
          5688 => x"7851f7b7",
          5689 => x"3f82e098",
          5690 => x"0883ffff",
          5691 => x"067e547c",
          5692 => x"5370832b",
          5693 => x"82e08808",
          5694 => x"11840553",
          5695 => x"5559ff87",
          5696 => x"ce3f82e0",
          5697 => x"88081484",
          5698 => x"057583ff",
          5699 => x"ff06595c",
          5700 => x"81853960",
          5701 => x"15547a74",
          5702 => x"2480d438",
          5703 => x"7851f5c9",
          5704 => x"3f82e088",
          5705 => x"081d8211",
          5706 => x"33831233",
          5707 => x"71882b07",
          5708 => x"534354f4",
          5709 => x"9c3f8052",
          5710 => x"7851f6df",
          5711 => x"3f82e098",
          5712 => x"0883ffff",
          5713 => x"067e547c",
          5714 => x"5370832b",
          5715 => x"82e08808",
          5716 => x"11840553",
          5717 => x"5559ff86",
          5718 => x"f63f82e0",
          5719 => x"88081484",
          5720 => x"05606205",
          5721 => x"19555c73",
          5722 => x"83ffff06",
          5723 => x"58a9397b",
          5724 => x"7f5254f9",
          5725 => x"b03f82e0",
          5726 => x"98085c82",
          5727 => x"e0980880",
          5728 => x"2e93387d",
          5729 => x"53735282",
          5730 => x"e0980851",
          5731 => x"ff8b8a3f",
          5732 => x"7351f798",
          5733 => x"3f7a587a",
          5734 => x"78279938",
          5735 => x"80537a52",
          5736 => x"7851f28f",
          5737 => x"3f7a1983",
          5738 => x"2b82e088",
          5739 => x"08058405",
          5740 => x"51f6f93f",
          5741 => x"7b547382",
          5742 => x"e0980c94",
          5743 => x"3d0d04fc",
          5744 => x"3d0d7777",
          5745 => x"29705254",
          5746 => x"fbd53f82",
          5747 => x"e0980855",
          5748 => x"82e09808",
          5749 => x"802e8e38",
          5750 => x"73538052",
          5751 => x"82e09808",
          5752 => x"51ff90e1",
          5753 => x"3f7482e0",
          5754 => x"980c863d",
          5755 => x"0d04ff3d",
          5756 => x"0d028f05",
          5757 => x"33518152",
          5758 => x"70722687",
          5759 => x"3882e094",
          5760 => x"11335271",
          5761 => x"82e0980c",
          5762 => x"833d0d04",
          5763 => x"fc3d0d02",
          5764 => x"9b053302",
          5765 => x"84059f05",
          5766 => x"33565383",
          5767 => x"51728126",
          5768 => x"80e03872",
          5769 => x"842b87c0",
          5770 => x"928c1153",
          5771 => x"51885474",
          5772 => x"802e8438",
          5773 => x"81885473",
          5774 => x"720c87c0",
          5775 => x"928c1151",
          5776 => x"81710c85",
          5777 => x"0b87c098",
          5778 => x"8c0c7052",
          5779 => x"71087082",
          5780 => x"06515170",
          5781 => x"802e8a38",
          5782 => x"87c0988c",
          5783 => x"085170ec",
          5784 => x"387108fc",
          5785 => x"80800652",
          5786 => x"71923887",
          5787 => x"c0988c08",
          5788 => x"5170802e",
          5789 => x"87387182",
          5790 => x"e0941434",
          5791 => x"82e09413",
          5792 => x"33517082",
          5793 => x"e0980c86",
          5794 => x"3d0d04f3",
          5795 => x"3d0d6062",
          5796 => x"64028c05",
          5797 => x"bf053357",
          5798 => x"40585b83",
          5799 => x"74525afe",
          5800 => x"cd3f82e0",
          5801 => x"98088106",
          5802 => x"7a545271",
          5803 => x"81be3871",
          5804 => x"7275842b",
          5805 => x"87c09280",
          5806 => x"1187c092",
          5807 => x"8c1287c0",
          5808 => x"92841341",
          5809 => x"5a40575a",
          5810 => x"58850b87",
          5811 => x"c0988c0c",
          5812 => x"767d0c84",
          5813 => x"760c7508",
          5814 => x"70852a70",
          5815 => x"81065153",
          5816 => x"5471802e",
          5817 => x"8e387b08",
          5818 => x"52717b70",
          5819 => x"81055d34",
          5820 => x"81195980",
          5821 => x"74a20653",
          5822 => x"5371732e",
          5823 => x"83388153",
          5824 => x"7883ff26",
          5825 => x"8f387280",
          5826 => x"2e8a3887",
          5827 => x"c0988c08",
          5828 => x"5271c338",
          5829 => x"87c0988c",
          5830 => x"08527180",
          5831 => x"2e873878",
          5832 => x"84802e99",
          5833 => x"3881760c",
          5834 => x"87c0928c",
          5835 => x"15537208",
          5836 => x"70820651",
          5837 => x"5271f738",
          5838 => x"ff1a5a8d",
          5839 => x"39848017",
          5840 => x"81197081",
          5841 => x"ff065a53",
          5842 => x"5779802e",
          5843 => x"903873fc",
          5844 => x"80800652",
          5845 => x"7187387d",
          5846 => x"7826feed",
          5847 => x"3873fc80",
          5848 => x"80065271",
          5849 => x"802e8338",
          5850 => x"81527153",
          5851 => x"7282e098",
          5852 => x"0c8f3d0d",
          5853 => x"04f33d0d",
          5854 => x"60626402",
          5855 => x"8c05bf05",
          5856 => x"33574058",
          5857 => x"5b835980",
          5858 => x"745258fc",
          5859 => x"e13f82e0",
          5860 => x"98088106",
          5861 => x"79545271",
          5862 => x"782e0981",
          5863 => x"0681b138",
          5864 => x"7774842b",
          5865 => x"87c09280",
          5866 => x"1187c092",
          5867 => x"8c1287c0",
          5868 => x"92841340",
          5869 => x"595f565a",
          5870 => x"850b87c0",
          5871 => x"988c0c76",
          5872 => x"7d0c8276",
          5873 => x"0c805875",
          5874 => x"0870842a",
          5875 => x"70810651",
          5876 => x"53547180",
          5877 => x"2e8c387a",
          5878 => x"7081055c",
          5879 => x"337c0c81",
          5880 => x"18587381",
          5881 => x"2a708106",
          5882 => x"51527180",
          5883 => x"2e8a3887",
          5884 => x"c0988c08",
          5885 => x"5271d038",
          5886 => x"87c0988c",
          5887 => x"08527180",
          5888 => x"2e873877",
          5889 => x"84802e99",
          5890 => x"3881760c",
          5891 => x"87c0928c",
          5892 => x"15537208",
          5893 => x"70820651",
          5894 => x"5271f738",
          5895 => x"ff19598d",
          5896 => x"39811a70",
          5897 => x"81ff0684",
          5898 => x"8019595b",
          5899 => x"5278802e",
          5900 => x"903873fc",
          5901 => x"80800652",
          5902 => x"7187387d",
          5903 => x"7a26fef8",
          5904 => x"3873fc80",
          5905 => x"80065271",
          5906 => x"802e8338",
          5907 => x"81527153",
          5908 => x"7282e098",
          5909 => x"0c8f3d0d",
          5910 => x"04fa3d0d",
          5911 => x"7a028405",
          5912 => x"a3053302",
          5913 => x"8805a705",
          5914 => x"33715454",
          5915 => x"5657fafe",
          5916 => x"3f82e098",
          5917 => x"08810653",
          5918 => x"83547280",
          5919 => x"fe38850b",
          5920 => x"87c0988c",
          5921 => x"0c815671",
          5922 => x"762e80dc",
          5923 => x"38717624",
          5924 => x"93387484",
          5925 => x"2b87c092",
          5926 => x"8c115454",
          5927 => x"71802e8d",
          5928 => x"3880d439",
          5929 => x"71832e80",
          5930 => x"c63880cb",
          5931 => x"39720870",
          5932 => x"812a7081",
          5933 => x"06515152",
          5934 => x"71802e8a",
          5935 => x"3887c098",
          5936 => x"8c085271",
          5937 => x"e83887c0",
          5938 => x"988c0852",
          5939 => x"71963881",
          5940 => x"730c87c0",
          5941 => x"928c1453",
          5942 => x"72087082",
          5943 => x"06515271",
          5944 => x"f7389639",
          5945 => x"80569239",
          5946 => x"88800a77",
          5947 => x"0c853981",
          5948 => x"80770c72",
          5949 => x"56833984",
          5950 => x"56755473",
          5951 => x"82e0980c",
          5952 => x"883d0d04",
          5953 => x"fe3d0d74",
          5954 => x"81113371",
          5955 => x"3371882b",
          5956 => x"0782e098",
          5957 => x"0c535184",
          5958 => x"3d0d04fd",
          5959 => x"3d0d7583",
          5960 => x"11338212",
          5961 => x"3371902b",
          5962 => x"71882b07",
          5963 => x"81143370",
          5964 => x"7207882b",
          5965 => x"75337107",
          5966 => x"82e0980c",
          5967 => x"52535456",
          5968 => x"5452853d",
          5969 => x"0d04ff3d",
          5970 => x"0d730284",
          5971 => x"05920522",
          5972 => x"52527072",
          5973 => x"70810554",
          5974 => x"3470882a",
          5975 => x"51707234",
          5976 => x"833d0d04",
          5977 => x"ff3d0d73",
          5978 => x"75525270",
          5979 => x"72708105",
          5980 => x"54347088",
          5981 => x"2a517072",
          5982 => x"70810554",
          5983 => x"3470882a",
          5984 => x"51707270",
          5985 => x"81055434",
          5986 => x"70882a51",
          5987 => x"70723483",
          5988 => x"3d0d04fe",
          5989 => x"3d0d7675",
          5990 => x"77545451",
          5991 => x"70802e92",
          5992 => x"38717081",
          5993 => x"05533373",
          5994 => x"70810555",
          5995 => x"34ff1151",
          5996 => x"eb39843d",
          5997 => x"0d04fe3d",
          5998 => x"0d757776",
          5999 => x"54525372",
          6000 => x"72708105",
          6001 => x"5434ff11",
          6002 => x"5170f438",
          6003 => x"843d0d04",
          6004 => x"fc3d0d78",
          6005 => x"77795656",
          6006 => x"53747081",
          6007 => x"05563374",
          6008 => x"70810556",
          6009 => x"33717131",
          6010 => x"ff165652",
          6011 => x"52527280",
          6012 => x"2e863871",
          6013 => x"802ee238",
          6014 => x"7182e098",
          6015 => x"0c863d0d",
          6016 => x"04fe3d0d",
          6017 => x"74765451",
          6018 => x"89397173",
          6019 => x"2e8a3881",
          6020 => x"11517033",
          6021 => x"5271f338",
          6022 => x"703382e0",
          6023 => x"980c843d",
          6024 => x"0d04800b",
          6025 => x"82e0980c",
          6026 => x"04fb3d0d",
          6027 => x"77700870",
          6028 => x"70810552",
          6029 => x"33705455",
          6030 => x"5556e73f",
          6031 => x"ff5582e0",
          6032 => x"9808a238",
          6033 => x"72802e98",
          6034 => x"3883b552",
          6035 => x"725180f9",
          6036 => x"a23f82e0",
          6037 => x"980883ff",
          6038 => x"ff065372",
          6039 => x"802e8638",
          6040 => x"73760c72",
          6041 => x"557482e0",
          6042 => x"980c873d",
          6043 => x"0d04f73d",
          6044 => x"0d7b5680",
          6045 => x"0b831733",
          6046 => x"565a747a",
          6047 => x"2e80d638",
          6048 => x"8154b416",
          6049 => x"0853b816",
          6050 => x"70538117",
          6051 => x"335259f9",
          6052 => x"e43f82e0",
          6053 => x"98087a2e",
          6054 => x"098106b7",
          6055 => x"3882e098",
          6056 => x"08831734",
          6057 => x"b4160870",
          6058 => x"a8180831",
          6059 => x"a0180859",
          6060 => x"56587477",
          6061 => x"279f3882",
          6062 => x"16335574",
          6063 => x"822e0981",
          6064 => x"06933881",
          6065 => x"54761853",
          6066 => x"78528116",
          6067 => x"3351f9a5",
          6068 => x"3f833981",
          6069 => x"5a7982e0",
          6070 => x"980c8b3d",
          6071 => x"0d04fa3d",
          6072 => x"0d787a56",
          6073 => x"56805774",
          6074 => x"b417082e",
          6075 => x"af387551",
          6076 => x"fefc3f82",
          6077 => x"e0980857",
          6078 => x"82e09808",
          6079 => x"9f388154",
          6080 => x"7453b816",
          6081 => x"52811633",
          6082 => x"51f7803f",
          6083 => x"82e09808",
          6084 => x"802e8538",
          6085 => x"ff558157",
          6086 => x"74b4170c",
          6087 => x"7682e098",
          6088 => x"0c883d0d",
          6089 => x"04f83d0d",
          6090 => x"7a705257",
          6091 => x"fec03f82",
          6092 => x"e0980858",
          6093 => x"82e09808",
          6094 => x"81913876",
          6095 => x"33557483",
          6096 => x"2e098106",
          6097 => x"80f03884",
          6098 => x"17335978",
          6099 => x"812e0981",
          6100 => x"0680e338",
          6101 => x"84805382",
          6102 => x"e0980852",
          6103 => x"b8177052",
          6104 => x"56fcd33f",
          6105 => x"82d4d552",
          6106 => x"84b61751",
          6107 => x"fbd83f84",
          6108 => x"8b85a4d2",
          6109 => x"527551fb",
          6110 => x"eb3f868a",
          6111 => x"85e4f252",
          6112 => x"849c1751",
          6113 => x"fbde3f94",
          6114 => x"17085284",
          6115 => x"a01751fb",
          6116 => x"d33f9017",
          6117 => x"085284a4",
          6118 => x"1751fbc8",
          6119 => x"3fa41708",
          6120 => x"810570b4",
          6121 => x"190c7955",
          6122 => x"53755281",
          6123 => x"173351f7",
          6124 => x"c43f7784",
          6125 => x"18348053",
          6126 => x"80528117",
          6127 => x"3351f999",
          6128 => x"3f82e098",
          6129 => x"08802e83",
          6130 => x"38815877",
          6131 => x"82e0980c",
          6132 => x"8a3d0d04",
          6133 => x"fb3d0d77",
          6134 => x"fe1a9c12",
          6135 => x"08fe0555",
          6136 => x"56548056",
          6137 => x"7473278d",
          6138 => x"388a1422",
          6139 => x"757129b0",
          6140 => x"16080557",
          6141 => x"537582e0",
          6142 => x"980c873d",
          6143 => x"0d04f93d",
          6144 => x"0d7a7a70",
          6145 => x"08565457",
          6146 => x"81772781",
          6147 => x"df38769c",
          6148 => x"15082781",
          6149 => x"d738ff74",
          6150 => x"33545872",
          6151 => x"822e80f5",
          6152 => x"38728224",
          6153 => x"89387281",
          6154 => x"2e8d3881",
          6155 => x"bf397283",
          6156 => x"2e818e38",
          6157 => x"81b63976",
          6158 => x"812a1770",
          6159 => x"892aa816",
          6160 => x"08055374",
          6161 => x"5255fd96",
          6162 => x"3f82e098",
          6163 => x"08819f38",
          6164 => x"7483ff06",
          6165 => x"14b81133",
          6166 => x"81177089",
          6167 => x"2aa81808",
          6168 => x"05557654",
          6169 => x"575753fc",
          6170 => x"f53f82e0",
          6171 => x"980880fe",
          6172 => x"387483ff",
          6173 => x"0614b811",
          6174 => x"3370882b",
          6175 => x"78077981",
          6176 => x"0671842a",
          6177 => x"5c525851",
          6178 => x"537280e2",
          6179 => x"38759fff",
          6180 => x"065880da",
          6181 => x"3976882a",
          6182 => x"a8150805",
          6183 => x"527351fc",
          6184 => x"bd3f82e0",
          6185 => x"980880c6",
          6186 => x"38761083",
          6187 => x"fe067405",
          6188 => x"b80551f8",
          6189 => x"cf3f82e0",
          6190 => x"980883ff",
          6191 => x"ff0658ae",
          6192 => x"3976872a",
          6193 => x"a8150805",
          6194 => x"527351fc",
          6195 => x"913f82e0",
          6196 => x"98089b38",
          6197 => x"76822b83",
          6198 => x"fc067405",
          6199 => x"b80551f8",
          6200 => x"ba3f82e0",
          6201 => x"9808f00a",
          6202 => x"06588339",
          6203 => x"81587782",
          6204 => x"e0980c89",
          6205 => x"3d0d04f8",
          6206 => x"3d0d7a7c",
          6207 => x"7e5a5856",
          6208 => x"82598177",
          6209 => x"27829e38",
          6210 => x"769c1708",
          6211 => x"27829638",
          6212 => x"75335372",
          6213 => x"792e819d",
          6214 => x"38727924",
          6215 => x"89387281",
          6216 => x"2e8d3882",
          6217 => x"80397283",
          6218 => x"2e81b838",
          6219 => x"81f73976",
          6220 => x"812a1770",
          6221 => x"892aa818",
          6222 => x"08055376",
          6223 => x"5255fb9e",
          6224 => x"3f82e098",
          6225 => x"085982e0",
          6226 => x"980881d9",
          6227 => x"387483ff",
          6228 => x"0616b805",
          6229 => x"81167881",
          6230 => x"06595654",
          6231 => x"77537680",
          6232 => x"2e8f3877",
          6233 => x"842b9ff0",
          6234 => x"0674338f",
          6235 => x"06710751",
          6236 => x"53727434",
          6237 => x"810b8317",
          6238 => x"3474892a",
          6239 => x"a8170805",
          6240 => x"527551fa",
          6241 => x"d93f82e0",
          6242 => x"98085982",
          6243 => x"e0980881",
          6244 => x"94387483",
          6245 => x"ff0616b8",
          6246 => x"0578842a",
          6247 => x"5454768f",
          6248 => x"3877882a",
          6249 => x"743381f0",
          6250 => x"06718f06",
          6251 => x"07515372",
          6252 => x"743480ec",
          6253 => x"3976882a",
          6254 => x"a8170805",
          6255 => x"527551fa",
          6256 => x"9d3f82e0",
          6257 => x"98085982",
          6258 => x"e0980880",
          6259 => x"d8387783",
          6260 => x"ffff0652",
          6261 => x"761083fe",
          6262 => x"067605b8",
          6263 => x"0551f6e6",
          6264 => x"3fbe3976",
          6265 => x"872aa817",
          6266 => x"08055275",
          6267 => x"51f9ef3f",
          6268 => x"82e09808",
          6269 => x"5982e098",
          6270 => x"08ab3877",
          6271 => x"f00a0677",
          6272 => x"822b83fc",
          6273 => x"067018b8",
          6274 => x"05705451",
          6275 => x"5454f68b",
          6276 => x"3f82e098",
          6277 => x"088f0a06",
          6278 => x"74075272",
          6279 => x"51f6c53f",
          6280 => x"810b8317",
          6281 => x"347882e0",
          6282 => x"980c8a3d",
          6283 => x"0d04f83d",
          6284 => x"0d7a7c7e",
          6285 => x"72085956",
          6286 => x"56598175",
          6287 => x"27a43874",
          6288 => x"9c170827",
          6289 => x"9d387380",
          6290 => x"2eaa38ff",
          6291 => x"53735275",
          6292 => x"51fda43f",
          6293 => x"82e09808",
          6294 => x"5482e098",
          6295 => x"0880f238",
          6296 => x"93398254",
          6297 => x"80eb3981",
          6298 => x"5480e639",
          6299 => x"82e09808",
          6300 => x"5480de39",
          6301 => x"74527851",
          6302 => x"fb843f82",
          6303 => x"e0980858",
          6304 => x"82e09808",
          6305 => x"802e80c7",
          6306 => x"3882e098",
          6307 => x"08812ed2",
          6308 => x"3882e098",
          6309 => x"08ff2ecf",
          6310 => x"38805374",
          6311 => x"527551fc",
          6312 => x"d63f82e0",
          6313 => x"9808c538",
          6314 => x"9c1608fe",
          6315 => x"11941808",
          6316 => x"57555774",
          6317 => x"74279038",
          6318 => x"81159417",
          6319 => x"0c841633",
          6320 => x"81075473",
          6321 => x"84173477",
          6322 => x"55767826",
          6323 => x"ffa63880",
          6324 => x"547382e0",
          6325 => x"980c8a3d",
          6326 => x"0d04f63d",
          6327 => x"0d7c7e71",
          6328 => x"08595b5b",
          6329 => x"79953890",
          6330 => x"17085877",
          6331 => x"802e8838",
          6332 => x"9c170878",
          6333 => x"26b23881",
          6334 => x"58ae3979",
          6335 => x"527a51f9",
          6336 => x"fd3f8155",
          6337 => x"7482e098",
          6338 => x"082782e0",
          6339 => x"3882e098",
          6340 => x"085582e0",
          6341 => x"9808ff2e",
          6342 => x"82d2389c",
          6343 => x"170882e0",
          6344 => x"98082682",
          6345 => x"c7387958",
          6346 => x"94170870",
          6347 => x"56547380",
          6348 => x"2e82b938",
          6349 => x"777a2e09",
          6350 => x"810680e2",
          6351 => x"38811a56",
          6352 => x"9c170876",
          6353 => x"26833882",
          6354 => x"5675527a",
          6355 => x"51f9af3f",
          6356 => x"805982e0",
          6357 => x"9808812e",
          6358 => x"09810686",
          6359 => x"3882e098",
          6360 => x"085982e0",
          6361 => x"98080970",
          6362 => x"30707207",
          6363 => x"8025707c",
          6364 => x"0782e098",
          6365 => x"08545151",
          6366 => x"55557381",
          6367 => x"ef3882e0",
          6368 => x"9808802e",
          6369 => x"95389017",
          6370 => x"08548174",
          6371 => x"27903873",
          6372 => x"9c180827",
          6373 => x"89387358",
          6374 => x"85397580",
          6375 => x"db387756",
          6376 => x"8116569c",
          6377 => x"17087626",
          6378 => x"89388256",
          6379 => x"75782681",
          6380 => x"ac387552",
          6381 => x"7a51f8c6",
          6382 => x"3f82e098",
          6383 => x"08802eb8",
          6384 => x"38805982",
          6385 => x"e0980881",
          6386 => x"2e098106",
          6387 => x"863882e0",
          6388 => x"98085982",
          6389 => x"e0980809",
          6390 => x"70307072",
          6391 => x"07802570",
          6392 => x"7c075151",
          6393 => x"55557380",
          6394 => x"f8387578",
          6395 => x"2e098106",
          6396 => x"ffae3873",
          6397 => x"5580f539",
          6398 => x"ff537552",
          6399 => x"7651f9f7",
          6400 => x"3f82e098",
          6401 => x"0882e098",
          6402 => x"08307082",
          6403 => x"e0980807",
          6404 => x"80255155",
          6405 => x"5579802e",
          6406 => x"94387380",
          6407 => x"2e8f3875",
          6408 => x"53795276",
          6409 => x"51f9d03f",
          6410 => x"82e09808",
          6411 => x"5574a538",
          6412 => x"7590180c",
          6413 => x"9c1708fe",
          6414 => x"05941808",
          6415 => x"56547474",
          6416 => x"268638ff",
          6417 => x"1594180c",
          6418 => x"84173381",
          6419 => x"07547384",
          6420 => x"18349739",
          6421 => x"ff567481",
          6422 => x"2e90388c",
          6423 => x"3980558c",
          6424 => x"3982e098",
          6425 => x"08558539",
          6426 => x"81567555",
          6427 => x"7482e098",
          6428 => x"0c8c3d0d",
          6429 => x"04f83d0d",
          6430 => x"7a705255",
          6431 => x"f3f03f82",
          6432 => x"e0980858",
          6433 => x"815682e0",
          6434 => x"980880d8",
          6435 => x"387b5274",
          6436 => x"51f6c13f",
          6437 => x"82e09808",
          6438 => x"82e09808",
          6439 => x"b4170c59",
          6440 => x"84805377",
          6441 => x"52b81570",
          6442 => x"5257f28a",
          6443 => x"3f775684",
          6444 => x"39811656",
          6445 => x"8a152258",
          6446 => x"75782797",
          6447 => x"38815475",
          6448 => x"19537652",
          6449 => x"81153351",
          6450 => x"edab3f82",
          6451 => x"e0980880",
          6452 => x"2edf388a",
          6453 => x"15227632",
          6454 => x"70307072",
          6455 => x"07709f2a",
          6456 => x"53515656",
          6457 => x"7582e098",
          6458 => x"0c8a3d0d",
          6459 => x"04f83d0d",
          6460 => x"7a7c7108",
          6461 => x"58565774",
          6462 => x"f0800a26",
          6463 => x"80f13874",
          6464 => x"9f065372",
          6465 => x"80e93874",
          6466 => x"90180c88",
          6467 => x"17085473",
          6468 => x"aa387533",
          6469 => x"53827327",
          6470 => x"8838ac16",
          6471 => x"0854739b",
          6472 => x"3874852a",
          6473 => x"53820b88",
          6474 => x"17225a58",
          6475 => x"72792780",
          6476 => x"fe38ac16",
          6477 => x"0898180c",
          6478 => x"80cd398a",
          6479 => x"16227089",
          6480 => x"2b545872",
          6481 => x"7526b238",
          6482 => x"73527651",
          6483 => x"f5b03f82",
          6484 => x"e0980854",
          6485 => x"82e09808",
          6486 => x"ff2ebd38",
          6487 => x"810b82e0",
          6488 => x"9808278b",
          6489 => x"389c1608",
          6490 => x"82e09808",
          6491 => x"26853882",
          6492 => x"58bd3974",
          6493 => x"733155cb",
          6494 => x"39735275",
          6495 => x"51f4d53f",
          6496 => x"82e09808",
          6497 => x"98180c73",
          6498 => x"94180c98",
          6499 => x"17085382",
          6500 => x"5872802e",
          6501 => x"9a388539",
          6502 => x"81589439",
          6503 => x"74892a13",
          6504 => x"98180c74",
          6505 => x"83ff0616",
          6506 => x"b8059c18",
          6507 => x"0c805877",
          6508 => x"82e0980c",
          6509 => x"8a3d0d04",
          6510 => x"f83d0d7a",
          6511 => x"70089012",
          6512 => x"08a00559",
          6513 => x"5754f080",
          6514 => x"0a772786",
          6515 => x"38800b98",
          6516 => x"150c9814",
          6517 => x"08538455",
          6518 => x"72802e81",
          6519 => x"cb387683",
          6520 => x"ff065877",
          6521 => x"81b53881",
          6522 => x"1398150c",
          6523 => x"94140855",
          6524 => x"74923876",
          6525 => x"852a8817",
          6526 => x"22565374",
          6527 => x"7326819b",
          6528 => x"3880c039",
          6529 => x"8a1622ff",
          6530 => x"0577892a",
          6531 => x"06537281",
          6532 => x"8a387452",
          6533 => x"7351f3e6",
          6534 => x"3f82e098",
          6535 => x"08538255",
          6536 => x"810b82e0",
          6537 => x"98082780",
          6538 => x"ff388155",
          6539 => x"82e09808",
          6540 => x"ff2e80f4",
          6541 => x"389c1608",
          6542 => x"82e09808",
          6543 => x"2680ca38",
          6544 => x"7b8a3877",
          6545 => x"98150c84",
          6546 => x"5580dd39",
          6547 => x"94140852",
          6548 => x"7351f986",
          6549 => x"3f82e098",
          6550 => x"08538755",
          6551 => x"82e09808",
          6552 => x"802e80c4",
          6553 => x"38825582",
          6554 => x"e0980881",
          6555 => x"2eba3881",
          6556 => x"5582e098",
          6557 => x"08ff2eb0",
          6558 => x"3882e098",
          6559 => x"08527551",
          6560 => x"fbf33f82",
          6561 => x"e09808a0",
          6562 => x"38729415",
          6563 => x"0c725275",
          6564 => x"51f2c13f",
          6565 => x"82e09808",
          6566 => x"98150c76",
          6567 => x"90150c77",
          6568 => x"16b8059c",
          6569 => x"150c8055",
          6570 => x"7482e098",
          6571 => x"0c8a3d0d",
          6572 => x"04f73d0d",
          6573 => x"7b7d7108",
          6574 => x"5b5b5780",
          6575 => x"527651fc",
          6576 => x"ac3f82e0",
          6577 => x"98085482",
          6578 => x"e0980880",
          6579 => x"ec3882e0",
          6580 => x"98085698",
          6581 => x"17085278",
          6582 => x"51f0833f",
          6583 => x"82e09808",
          6584 => x"5482e098",
          6585 => x"0880d238",
          6586 => x"82e09808",
          6587 => x"9c180870",
          6588 => x"33515458",
          6589 => x"7281e52e",
          6590 => x"09810683",
          6591 => x"38815882",
          6592 => x"e0980855",
          6593 => x"72833881",
          6594 => x"55777507",
          6595 => x"5372802e",
          6596 => x"8e388116",
          6597 => x"56757a2e",
          6598 => x"09810688",
          6599 => x"38a53982",
          6600 => x"e0980856",
          6601 => x"81527651",
          6602 => x"fd8e3f82",
          6603 => x"e0980854",
          6604 => x"82e09808",
          6605 => x"802eff9b",
          6606 => x"3873842e",
          6607 => x"09810683",
          6608 => x"38875473",
          6609 => x"82e0980c",
          6610 => x"8b3d0d04",
          6611 => x"fd3d0d76",
          6612 => x"9a115254",
          6613 => x"ebae3f82",
          6614 => x"e0980883",
          6615 => x"ffff0676",
          6616 => x"70335153",
          6617 => x"5371832e",
          6618 => x"09810690",
          6619 => x"38941451",
          6620 => x"eb923f82",
          6621 => x"e0980890",
          6622 => x"2b730753",
          6623 => x"7282e098",
          6624 => x"0c853d0d",
          6625 => x"04fc3d0d",
          6626 => x"77797083",
          6627 => x"ffff0654",
          6628 => x"9a125355",
          6629 => x"55ebaf3f",
          6630 => x"76703351",
          6631 => x"5372832e",
          6632 => x"0981068b",
          6633 => x"3873902a",
          6634 => x"52941551",
          6635 => x"eb983f86",
          6636 => x"3d0d04fd",
          6637 => x"3d0d7554",
          6638 => x"80518b53",
          6639 => x"70812a71",
          6640 => x"81802905",
          6641 => x"74708105",
          6642 => x"56337105",
          6643 => x"7081ff06",
          6644 => x"ff165651",
          6645 => x"515172e4",
          6646 => x"387082e0",
          6647 => x"980c853d",
          6648 => x"0d04f23d",
          6649 => x"0d606240",
          6650 => x"59847908",
          6651 => x"5f5b81ff",
          6652 => x"705d5d98",
          6653 => x"1908802e",
          6654 => x"83803898",
          6655 => x"1908527d",
          6656 => x"51eddb3f",
          6657 => x"82e09808",
          6658 => x"5b82e098",
          6659 => x"0882eb38",
          6660 => x"9c190870",
          6661 => x"33555573",
          6662 => x"8638845b",
          6663 => x"82dc398b",
          6664 => x"1533bf06",
          6665 => x"7081ff06",
          6666 => x"58537286",
          6667 => x"1a3482e0",
          6668 => x"98085673",
          6669 => x"81e52e09",
          6670 => x"81068338",
          6671 => x"815682e0",
          6672 => x"98085373",
          6673 => x"ae2e0981",
          6674 => x"06833881",
          6675 => x"53757307",
          6676 => x"53729938",
          6677 => x"82e09808",
          6678 => x"77df0654",
          6679 => x"5672882e",
          6680 => x"09810683",
          6681 => x"38815675",
          6682 => x"7f2e8738",
          6683 => x"81ff5c81",
          6684 => x"ef39768f",
          6685 => x"2e098106",
          6686 => x"81ca3873",
          6687 => x"862a7081",
          6688 => x"06515372",
          6689 => x"802e9238",
          6690 => x"8d153374",
          6691 => x"81bf0670",
          6692 => x"901c08ac",
          6693 => x"1d0c565d",
          6694 => x"5d737c2e",
          6695 => x"09810681",
          6696 => x"9c388d15",
          6697 => x"33537c73",
          6698 => x"2e098106",
          6699 => x"818f388c",
          6700 => x"1e089a16",
          6701 => x"525ae8cc",
          6702 => x"3f82e098",
          6703 => x"0883ffff",
          6704 => x"06537280",
          6705 => x"f8387433",
          6706 => x"7081bf06",
          6707 => x"8d29f305",
          6708 => x"5154817b",
          6709 => x"585882d2",
          6710 => x"a8173375",
          6711 => x"0551e8a4",
          6712 => x"3f82e098",
          6713 => x"0883ffff",
          6714 => x"06567780",
          6715 => x"2e963873",
          6716 => x"81fe2680",
          6717 => x"c8387310",
          6718 => x"1a765953",
          6719 => x"75732381",
          6720 => x"14548b39",
          6721 => x"7583ffff",
          6722 => x"2e098106",
          6723 => x"b0388117",
          6724 => x"578c7727",
          6725 => x"c1387433",
          6726 => x"70862a70",
          6727 => x"81065154",
          6728 => x"5572802e",
          6729 => x"8e387381",
          6730 => x"fe269238",
          6731 => x"73101a53",
          6732 => x"807323ff",
          6733 => x"1c7081ff",
          6734 => x"06515384",
          6735 => x"3981ff53",
          6736 => x"725c9d39",
          6737 => x"7b933874",
          6738 => x"51fce83f",
          6739 => x"82e09808",
          6740 => x"81ff0653",
          6741 => x"727d2ea7",
          6742 => x"38ff0bac",
          6743 => x"1a0ca039",
          6744 => x"80527851",
          6745 => x"f8d23f82",
          6746 => x"e098085b",
          6747 => x"82e09808",
          6748 => x"89389819",
          6749 => x"08fd8438",
          6750 => x"8639800b",
          6751 => x"981a0c7a",
          6752 => x"82e0980c",
          6753 => x"903d0d04",
          6754 => x"f23d0d60",
          6755 => x"70084059",
          6756 => x"80527851",
          6757 => x"f6d73f82",
          6758 => x"e0980858",
          6759 => x"82e09808",
          6760 => x"83a43881",
          6761 => x"ff705f5c",
          6762 => x"ff0bac1a",
          6763 => x"0c981908",
          6764 => x"527e51ea",
          6765 => x"a93f82e0",
          6766 => x"98085882",
          6767 => x"e0980883",
          6768 => x"85389c19",
          6769 => x"08703357",
          6770 => x"57758638",
          6771 => x"845882f6",
          6772 => x"398b1733",
          6773 => x"bf067081",
          6774 => x"ff065654",
          6775 => x"73861a34",
          6776 => x"7581e52e",
          6777 => x"82c33874",
          6778 => x"832a7081",
          6779 => x"06515474",
          6780 => x"8f2e8e38",
          6781 => x"7382b238",
          6782 => x"748f2e09",
          6783 => x"810681f7",
          6784 => x"38ab1933",
          6785 => x"70862a70",
          6786 => x"81065155",
          6787 => x"557382a1",
          6788 => x"3875862a",
          6789 => x"70810651",
          6790 => x"5473802e",
          6791 => x"92388d17",
          6792 => x"337681bf",
          6793 => x"0670901c",
          6794 => x"08ac1d0c",
          6795 => x"585d5e75",
          6796 => x"7c2e0981",
          6797 => x"0681b938",
          6798 => x"8d173356",
          6799 => x"7d762e09",
          6800 => x"810681ac",
          6801 => x"388c1f08",
          6802 => x"9a18525d",
          6803 => x"e5b63f82",
          6804 => x"e0980883",
          6805 => x"ffff0655",
          6806 => x"74819538",
          6807 => x"763370bf",
          6808 => x"068d29f3",
          6809 => x"05595681",
          6810 => x"755c5a82",
          6811 => x"d2a81b33",
          6812 => x"770551e5",
          6813 => x"8f3f82e0",
          6814 => x"980883ff",
          6815 => x"ff065679",
          6816 => x"802eb138",
          6817 => x"7781fe26",
          6818 => x"80e63875",
          6819 => x"5180e1a0",
          6820 => x"3f82e098",
          6821 => x"0878101e",
          6822 => x"70225355",
          6823 => x"81195955",
          6824 => x"80e18d3f",
          6825 => x"7482e098",
          6826 => x"082e0981",
          6827 => x"0680c138",
          6828 => x"755a8b39",
          6829 => x"7583ffff",
          6830 => x"2e098106",
          6831 => x"b338811b",
          6832 => x"5b8c7b27",
          6833 => x"ffa53876",
          6834 => x"3370862a",
          6835 => x"70810651",
          6836 => x"55577980",
          6837 => x"2e903873",
          6838 => x"802e8b38",
          6839 => x"77101d70",
          6840 => x"22515473",
          6841 => x"8b38ff1c",
          6842 => x"7081ff06",
          6843 => x"51548439",
          6844 => x"81ff5473",
          6845 => x"5cbb397b",
          6846 => x"93387651",
          6847 => x"f9b53f82",
          6848 => x"e0980881",
          6849 => x"ff065473",
          6850 => x"7e2ebb38",
          6851 => x"ab193381",
          6852 => x"06547395",
          6853 => x"388b53a0",
          6854 => x"19529c19",
          6855 => x"0851e5b0",
          6856 => x"3f82e098",
          6857 => x"08802e9e",
          6858 => x"3881ff5c",
          6859 => x"ff0bac1a",
          6860 => x"0c805278",
          6861 => x"51f5813f",
          6862 => x"82e09808",
          6863 => x"5882e098",
          6864 => x"08802efc",
          6865 => x"e8387782",
          6866 => x"e0980c90",
          6867 => x"3d0d04ee",
          6868 => x"3d0d6470",
          6869 => x"08ab1233",
          6870 => x"81a00656",
          6871 => x"5d5a8655",
          6872 => x"7385b538",
          6873 => x"738c1d08",
          6874 => x"70225656",
          6875 => x"5d73802e",
          6876 => x"8d38811d",
          6877 => x"70101670",
          6878 => x"2251555d",
          6879 => x"f0398c53",
          6880 => x"a01a7053",
          6881 => x"923d7053",
          6882 => x"5f59e487",
          6883 => x"3f0280cb",
          6884 => x"05338106",
          6885 => x"5473802e",
          6886 => x"82a83880",
          6887 => x"c00bab1b",
          6888 => x"34815b8c",
          6889 => x"1c087b56",
          6890 => x"588b537d",
          6891 => x"527851e3",
          6892 => x"e23f857b",
          6893 => x"2780c638",
          6894 => x"7a567722",
          6895 => x"7083ffff",
          6896 => x"06555573",
          6897 => x"802eb438",
          6898 => x"7483ffff",
          6899 => x"06821959",
          6900 => x"558f5774",
          6901 => x"81067610",
          6902 => x"0775812a",
          6903 => x"71902a70",
          6904 => x"81065156",
          6905 => x"56567380",
          6906 => x"2e873875",
          6907 => x"84a0a132",
          6908 => x"56ff1757",
          6909 => x"768025db",
          6910 => x"38c03975",
          6911 => x"55870284",
          6912 => x"05bf0557",
          6913 => x"5774b007",
          6914 => x"bf0654b9",
          6915 => x"74278438",
          6916 => x"87145473",
          6917 => x"7634ff16",
          6918 => x"ff187684",
          6919 => x"2a575856",
          6920 => x"74e33894",
          6921 => x"3dec0517",
          6922 => x"5480fe74",
          6923 => x"34807727",
          6924 => x"b5387833",
          6925 => x"5473a02e",
          6926 => x"ad387419",
          6927 => x"70335254",
          6928 => x"e3e03f82",
          6929 => x"e0980880",
          6930 => x"2e8c38ff",
          6931 => x"17547474",
          6932 => x"2e943881",
          6933 => x"15558115",
          6934 => x"55747727",
          6935 => x"89387419",
          6936 => x"70335154",
          6937 => x"d039943d",
          6938 => x"7705eb05",
          6939 => x"54781581",
          6940 => x"165658a0",
          6941 => x"56768726",
          6942 => x"8a388117",
          6943 => x"81157033",
          6944 => x"58555775",
          6945 => x"78348775",
          6946 => x"27e33879",
          6947 => x"51f9f93f",
          6948 => x"82e09808",
          6949 => x"8b38811b",
          6950 => x"5b80e37b",
          6951 => x"27fe8438",
          6952 => x"87557a80",
          6953 => x"e42e82f0",
          6954 => x"3882e098",
          6955 => x"085582e0",
          6956 => x"9808842e",
          6957 => x"09810682",
          6958 => x"df380280",
          6959 => x"cb0533ab",
          6960 => x"1b340280",
          6961 => x"cb053370",
          6962 => x"812a7081",
          6963 => x"0651555e",
          6964 => x"81597380",
          6965 => x"2e90388d",
          6966 => x"528c1d51",
          6967 => x"feebf43f",
          6968 => x"82e09808",
          6969 => x"19597852",
          6970 => x"7951f3c5",
          6971 => x"3f82e098",
          6972 => x"085782e0",
          6973 => x"9808829e",
          6974 => x"38ff1959",
          6975 => x"78802e81",
          6976 => x"d4387885",
          6977 => x"2b901b08",
          6978 => x"71315354",
          6979 => x"7951efdd",
          6980 => x"3f82e098",
          6981 => x"085782e0",
          6982 => x"980881fa",
          6983 => x"38a01a51",
          6984 => x"f5913f82",
          6985 => x"e0980881",
          6986 => x"ff065d98",
          6987 => x"1a08527b",
          6988 => x"51e3ab3f",
          6989 => x"82e09808",
          6990 => x"5782e098",
          6991 => x"0881d738",
          6992 => x"8c1c089c",
          6993 => x"1b087a81",
          6994 => x"ff065a57",
          6995 => x"5b7c8d17",
          6996 => x"348f0b8b",
          6997 => x"173482e0",
          6998 => x"98088c17",
          6999 => x"3482e098",
          7000 => x"08529a16",
          7001 => x"51dfdf3f",
          7002 => x"778d29f3",
          7003 => x"05775555",
          7004 => x"7383ffff",
          7005 => x"2e8b3874",
          7006 => x"101b7022",
          7007 => x"81175751",
          7008 => x"54735282",
          7009 => x"d2a81733",
          7010 => x"760551df",
          7011 => x"b93f7385",
          7012 => x"3883ffff",
          7013 => x"54811757",
          7014 => x"8c7727d4",
          7015 => x"387383ff",
          7016 => x"ff2e8b38",
          7017 => x"74101b70",
          7018 => x"22515473",
          7019 => x"86387780",
          7020 => x"c0075877",
          7021 => x"7634810b",
          7022 => x"831d3480",
          7023 => x"527951ef",
          7024 => x"f73f82e0",
          7025 => x"98085782",
          7026 => x"e0980880",
          7027 => x"c938ff19",
          7028 => x"5978fed7",
          7029 => x"38981a08",
          7030 => x"527b51e2",
          7031 => x"813f82e0",
          7032 => x"98085782",
          7033 => x"e09808ae",
          7034 => x"38a05382",
          7035 => x"e0980852",
          7036 => x"9c1a0851",
          7037 => x"dfc03f8b",
          7038 => x"53a01a52",
          7039 => x"9c1a0851",
          7040 => x"df913f9c",
          7041 => x"1a08ab1b",
          7042 => x"33980655",
          7043 => x"55738c16",
          7044 => x"34810b83",
          7045 => x"1d347655",
          7046 => x"7482e098",
          7047 => x"0c943d0d",
          7048 => x"04fa3d0d",
          7049 => x"78700890",
          7050 => x"1208ac13",
          7051 => x"08565957",
          7052 => x"5572ff2e",
          7053 => x"94387252",
          7054 => x"7451edb1",
          7055 => x"3f82e098",
          7056 => x"085482e0",
          7057 => x"980880c9",
          7058 => x"38981508",
          7059 => x"527551e1",
          7060 => x"8d3f82e0",
          7061 => x"98085482",
          7062 => x"e09808ab",
          7063 => x"389c1508",
          7064 => x"53e57334",
          7065 => x"810b8317",
          7066 => x"34901508",
          7067 => x"7727a238",
          7068 => x"82e09808",
          7069 => x"527451ee",
          7070 => x"bf3f82e0",
          7071 => x"98085482",
          7072 => x"e0980880",
          7073 => x"2ec33873",
          7074 => x"842e0981",
          7075 => x"06833882",
          7076 => x"547382e0",
          7077 => x"980c883d",
          7078 => x"0d04f43d",
          7079 => x"0d7e6071",
          7080 => x"085f595c",
          7081 => x"800b9619",
          7082 => x"34981c08",
          7083 => x"802e83e2",
          7084 => x"38ac1c08",
          7085 => x"ff2e81bb",
          7086 => x"38807071",
          7087 => x"7f8c0508",
          7088 => x"70225757",
          7089 => x"5b5c5772",
          7090 => x"772e819d",
          7091 => x"38781014",
          7092 => x"7022811b",
          7093 => x"5b56537a",
          7094 => x"973880d0",
          7095 => x"80157083",
          7096 => x"ffff0651",
          7097 => x"53728fff",
          7098 => x"26863874",
          7099 => x"5b80df39",
          7100 => x"76189611",
          7101 => x"81ff7931",
          7102 => x"585b5483",
          7103 => x"b5527a90",
          7104 => x"2b750751",
          7105 => x"80d7843f",
          7106 => x"82e09808",
          7107 => x"83ffff06",
          7108 => x"5581ff75",
          7109 => x"27953881",
          7110 => x"7627a538",
          7111 => x"74882a53",
          7112 => x"727a3474",
          7113 => x"97153482",
          7114 => x"559f3974",
          7115 => x"30763070",
          7116 => x"78078025",
          7117 => x"72802507",
          7118 => x"52545473",
          7119 => x"802e8538",
          7120 => x"80579a39",
          7121 => x"747a3481",
          7122 => x"55741757",
          7123 => x"805b8c1d",
          7124 => x"08791011",
          7125 => x"70225154",
          7126 => x"5472fef1",
          7127 => x"387a3070",
          7128 => x"80257030",
          7129 => x"79065951",
          7130 => x"53771794",
          7131 => x"0553800b",
          7132 => x"82143480",
          7133 => x"70891a58",
          7134 => x"5a579c1c",
          7135 => x"08197033",
          7136 => x"811b5b56",
          7137 => x"5374a02e",
          7138 => x"b7387485",
          7139 => x"2e098106",
          7140 => x"843881e5",
          7141 => x"55788932",
          7142 => x"70307072",
          7143 => x"07802551",
          7144 => x"5454768b",
          7145 => x"26903872",
          7146 => x"802e8b38",
          7147 => x"ae767081",
          7148 => x"05583481",
          7149 => x"17577476",
          7150 => x"70810558",
          7151 => x"34811757",
          7152 => x"8a7927ff",
          7153 => x"b5387717",
          7154 => x"88055380",
          7155 => x"0b811434",
          7156 => x"96183353",
          7157 => x"72818738",
          7158 => x"768b38bf",
          7159 => x"0b961934",
          7160 => x"815780e1",
          7161 => x"39727389",
          7162 => x"1a33555a",
          7163 => x"5772802e",
          7164 => x"80d33896",
          7165 => x"18891955",
          7166 => x"567333ff",
          7167 => x"bf115455",
          7168 => x"729926aa",
          7169 => x"389c1c08",
          7170 => x"8c113351",
          7171 => x"53887927",
          7172 => x"87387284",
          7173 => x"2a538539",
          7174 => x"72832a53",
          7175 => x"72810653",
          7176 => x"72802e8a",
          7177 => x"38a01570",
          7178 => x"83ffff06",
          7179 => x"56537476",
          7180 => x"70810558",
          7181 => x"34811981",
          7182 => x"15811971",
          7183 => x"33565955",
          7184 => x"5972ffb5",
          7185 => x"38771794",
          7186 => x"0553800b",
          7187 => x"8214349c",
          7188 => x"1c088c11",
          7189 => x"33515372",
          7190 => x"85387289",
          7191 => x"19349c1c",
          7192 => x"08538b13",
          7193 => x"33881934",
          7194 => x"9c1c089c",
          7195 => x"115253d9",
          7196 => x"aa3f82e0",
          7197 => x"9808780c",
          7198 => x"961351d9",
          7199 => x"873f82e0",
          7200 => x"98088619",
          7201 => x"23981351",
          7202 => x"d8fa3f82",
          7203 => x"e0980884",
          7204 => x"19238e3d",
          7205 => x"0d04f03d",
          7206 => x"0d627008",
          7207 => x"415e8064",
          7208 => x"70335155",
          7209 => x"5573af2e",
          7210 => x"83388155",
          7211 => x"7380dc2e",
          7212 => x"92387480",
          7213 => x"2e8d387f",
          7214 => x"98050888",
          7215 => x"1f0caa39",
          7216 => x"81154480",
          7217 => x"64703356",
          7218 => x"565673af",
          7219 => x"2e098106",
          7220 => x"83388156",
          7221 => x"7380dc32",
          7222 => x"70307080",
          7223 => x"25780751",
          7224 => x"515473dc",
          7225 => x"3873881f",
          7226 => x"0c637033",
          7227 => x"5154739f",
          7228 => x"269638ff",
          7229 => x"800bab1f",
          7230 => x"3480527d",
          7231 => x"51e7ee3f",
          7232 => x"82e09808",
          7233 => x"5687e139",
          7234 => x"63417d08",
          7235 => x"8c11085b",
          7236 => x"54805992",
          7237 => x"3dfc0551",
          7238 => x"da8f3f82",
          7239 => x"e09808ff",
          7240 => x"2e82b138",
          7241 => x"83ffff0b",
          7242 => x"82e09808",
          7243 => x"27923878",
          7244 => x"101a82e0",
          7245 => x"9808902a",
          7246 => x"55557375",
          7247 => x"23811959",
          7248 => x"82e09808",
          7249 => x"83ffff06",
          7250 => x"70af3270",
          7251 => x"309f7327",
          7252 => x"71802507",
          7253 => x"51515556",
          7254 => x"73b43875",
          7255 => x"80dc2eae",
          7256 => x"387580ff",
          7257 => x"26913875",
          7258 => x"5282d1c4",
          7259 => x"51d9923f",
          7260 => x"82e09808",
          7261 => x"81de3878",
          7262 => x"81fe2681",
          7263 => x"d7387810",
          7264 => x"1a547574",
          7265 => x"23811959",
          7266 => x"ff893981",
          7267 => x"15418061",
          7268 => x"70335656",
          7269 => x"5773af2e",
          7270 => x"09810683",
          7271 => x"38815773",
          7272 => x"80dc3270",
          7273 => x"30708025",
          7274 => x"79075151",
          7275 => x"5473dc38",
          7276 => x"74449f76",
          7277 => x"27822b57",
          7278 => x"78812e09",
          7279 => x"81068c38",
          7280 => x"79225473",
          7281 => x"ae2ea538",
          7282 => x"80d23978",
          7283 => x"822e0981",
          7284 => x"0680c938",
          7285 => x"821a2254",
          7286 => x"73ae2e09",
          7287 => x"810680c1",
          7288 => x"38792254",
          7289 => x"73ae2e09",
          7290 => x"8106b638",
          7291 => x"78101a54",
          7292 => x"80742380",
          7293 => x"0ba01f56",
          7294 => x"58ae5478",
          7295 => x"78268338",
          7296 => x"a0547375",
          7297 => x"70810557",
          7298 => x"34811858",
          7299 => x"8a7827e9",
          7300 => x"3876a007",
          7301 => x"5473ab1f",
          7302 => x"3484c439",
          7303 => x"78802ea8",
          7304 => x"3878101a",
          7305 => x"fe055574",
          7306 => x"22fe1671",
          7307 => x"72a03270",
          7308 => x"30709f2a",
          7309 => x"51515358",
          7310 => x"565475ae",
          7311 => x"2e843873",
          7312 => x"8738ff19",
          7313 => x"5978e038",
          7314 => x"78197a11",
          7315 => x"55568074",
          7316 => x"23788d38",
          7317 => x"86568590",
          7318 => x"39768307",
          7319 => x"57839939",
          7320 => x"807a2270",
          7321 => x"83ffff06",
          7322 => x"56565d73",
          7323 => x"a02e0981",
          7324 => x"06933881",
          7325 => x"1d70101b",
          7326 => x"70225155",
          7327 => x"5d73a02e",
          7328 => x"f2387c8f",
          7329 => x"387483ff",
          7330 => x"ff065473",
          7331 => x"ae2e0981",
          7332 => x"06853876",
          7333 => x"83075778",
          7334 => x"802eaa38",
          7335 => x"7916fe05",
          7336 => x"70225154",
          7337 => x"73ae2e9d",
          7338 => x"3878101a",
          7339 => x"fe0555ff",
          7340 => x"19597880",
          7341 => x"2e8f38fe",
          7342 => x"15702255",
          7343 => x"5573ae2e",
          7344 => x"098106eb",
          7345 => x"388b53a0",
          7346 => x"52a01e51",
          7347 => x"d5e83f80",
          7348 => x"70595c88",
          7349 => x"5f7c101a",
          7350 => x"7022811f",
          7351 => x"5f575475",
          7352 => x"802e8294",
          7353 => x"3875a02e",
          7354 => x"963875ae",
          7355 => x"32703070",
          7356 => x"80255151",
          7357 => x"547c792e",
          7358 => x"8c387380",
          7359 => x"2e893876",
          7360 => x"830757d1",
          7361 => x"39805473",
          7362 => x"5b7e7826",
          7363 => x"8338815b",
          7364 => x"7c793270",
          7365 => x"30707207",
          7366 => x"8025707e",
          7367 => x"07515155",
          7368 => x"5573802e",
          7369 => x"a6387e8b",
          7370 => x"2efeae38",
          7371 => x"7c792e8b",
          7372 => x"38768307",
          7373 => x"577c7926",
          7374 => x"81be3878",
          7375 => x"5d88588b",
          7376 => x"7c822b81",
          7377 => x"fc065d5f",
          7378 => x"ff8b3980",
          7379 => x"ff7627af",
          7380 => x"38768207",
          7381 => x"5783b552",
          7382 => x"755180ce",
          7383 => x"ae3f82e0",
          7384 => x"980883ff",
          7385 => x"ff067087",
          7386 => x"2a708106",
          7387 => x"51555673",
          7388 => x"802e8c38",
          7389 => x"7580ff06",
          7390 => x"82d2b811",
          7391 => x"33575481",
          7392 => x"ff7627a4",
          7393 => x"38ff1f54",
          7394 => x"7378268a",
          7395 => x"38768307",
          7396 => x"7f5957fe",
          7397 => x"c0397d18",
          7398 => x"a0057688",
          7399 => x"2a555573",
          7400 => x"75348118",
          7401 => x"5880c339",
          7402 => x"75802e92",
          7403 => x"38755282",
          7404 => x"d1d051d4",
          7405 => x"cc3f82e0",
          7406 => x"9808802e",
          7407 => x"8a3880df",
          7408 => x"77830758",
          7409 => x"56a439ff",
          7410 => x"bf165473",
          7411 => x"99268538",
          7412 => x"7b82075c",
          7413 => x"ff9f1654",
          7414 => x"7399268e",
          7415 => x"387b8107",
          7416 => x"e0177083",
          7417 => x"ffff0658",
          7418 => x"555c7d18",
          7419 => x"a0055475",
          7420 => x"74348118",
          7421 => x"58fdde39",
          7422 => x"a01e3354",
          7423 => x"7381e52e",
          7424 => x"09810686",
          7425 => x"38850ba0",
          7426 => x"1f347e88",
          7427 => x"2e098106",
          7428 => x"88387b82",
          7429 => x"2b81fc06",
          7430 => x"5c7b8c06",
          7431 => x"54738c2e",
          7432 => x"8d387b83",
          7433 => x"06547383",
          7434 => x"2e098106",
          7435 => x"85387682",
          7436 => x"07577681",
          7437 => x"2a708106",
          7438 => x"5154739f",
          7439 => x"387b8106",
          7440 => x"5473802e",
          7441 => x"85387690",
          7442 => x"07577b82",
          7443 => x"2a708106",
          7444 => x"51547380",
          7445 => x"2e853876",
          7446 => x"88075776",
          7447 => x"ab1f347d",
          7448 => x"51eaa53f",
          7449 => x"82e09808",
          7450 => x"ab1f3356",
          7451 => x"5682e098",
          7452 => x"08802ebe",
          7453 => x"3882e098",
          7454 => x"08842e09",
          7455 => x"810680e8",
          7456 => x"3874852a",
          7457 => x"70810676",
          7458 => x"822a5751",
          7459 => x"5473802e",
          7460 => x"96387481",
          7461 => x"06547380",
          7462 => x"2ef8ed38",
          7463 => x"ff800bab",
          7464 => x"1f348056",
          7465 => x"80c23974",
          7466 => x"81065473",
          7467 => x"bb388556",
          7468 => x"b7397482",
          7469 => x"2a708106",
          7470 => x"515473ac",
          7471 => x"38861e33",
          7472 => x"70842a70",
          7473 => x"81065155",
          7474 => x"5573802e",
          7475 => x"e138901e",
          7476 => x"0883ff06",
          7477 => x"6005b805",
          7478 => x"527f51e4",
          7479 => x"ef3f82e0",
          7480 => x"9808881f",
          7481 => x"0cf8a139",
          7482 => x"7582e098",
          7483 => x"0c923d0d",
          7484 => x"04f63d0d",
          7485 => x"7c5bff7b",
          7486 => x"08707173",
          7487 => x"55595c55",
          7488 => x"5973802e",
          7489 => x"81c63875",
          7490 => x"70810557",
          7491 => x"33709f26",
          7492 => x"525271ba",
          7493 => x"2e8d3870",
          7494 => x"ee3871ba",
          7495 => x"2e098106",
          7496 => x"81a53873",
          7497 => x"33d01170",
          7498 => x"81ff0651",
          7499 => x"52537089",
          7500 => x"26913882",
          7501 => x"147381ff",
          7502 => x"06d00556",
          7503 => x"5271762e",
          7504 => x"80f73880",
          7505 => x"0b82d298",
          7506 => x"59557708",
          7507 => x"7a555776",
          7508 => x"70810558",
          7509 => x"33747081",
          7510 => x"055633ff",
          7511 => x"9f125353",
          7512 => x"53709926",
          7513 => x"8938e013",
          7514 => x"7081ff06",
          7515 => x"5451ff9f",
          7516 => x"12517099",
          7517 => x"268938e0",
          7518 => x"127081ff",
          7519 => x"06535172",
          7520 => x"30709f2a",
          7521 => x"51517272",
          7522 => x"2e098106",
          7523 => x"853870ff",
          7524 => x"be387230",
          7525 => x"74773270",
          7526 => x"30707207",
          7527 => x"9f2a739f",
          7528 => x"2a075354",
          7529 => x"54517080",
          7530 => x"2e8f3881",
          7531 => x"15841959",
          7532 => x"55837525",
          7533 => x"ff94388b",
          7534 => x"39748324",
          7535 => x"86387476",
          7536 => x"7c0c5978",
          7537 => x"51863982",
          7538 => x"f7f43351",
          7539 => x"7082e098",
          7540 => x"0c8c3d0d",
          7541 => x"04fa3d0d",
          7542 => x"7856800b",
          7543 => x"831734ff",
          7544 => x"0bb4170c",
          7545 => x"79527551",
          7546 => x"d1f43f84",
          7547 => x"5582e098",
          7548 => x"08818038",
          7549 => x"84b61651",
          7550 => x"ce8a3f82",
          7551 => x"e0980883",
          7552 => x"ffff0654",
          7553 => x"83557382",
          7554 => x"d4d52e09",
          7555 => x"810680e3",
          7556 => x"38800bb8",
          7557 => x"17335657",
          7558 => x"7481e92e",
          7559 => x"09810683",
          7560 => x"38815774",
          7561 => x"81eb3270",
          7562 => x"30708025",
          7563 => x"79075151",
          7564 => x"54738a38",
          7565 => x"7481e82e",
          7566 => x"098106b5",
          7567 => x"38835382",
          7568 => x"d1d85280",
          7569 => x"ee1651cf",
          7570 => x"873f82e0",
          7571 => x"98085582",
          7572 => x"e0980880",
          7573 => x"2e9d3885",
          7574 => x"5382d1dc",
          7575 => x"52818a16",
          7576 => x"51ceed3f",
          7577 => x"82e09808",
          7578 => x"5582e098",
          7579 => x"08802e83",
          7580 => x"38825574",
          7581 => x"82e0980c",
          7582 => x"883d0d04",
          7583 => x"f23d0d61",
          7584 => x"02840580",
          7585 => x"cb053358",
          7586 => x"5580750c",
          7587 => x"6051fce1",
          7588 => x"3f82e098",
          7589 => x"08588b56",
          7590 => x"800b82e0",
          7591 => x"98082487",
          7592 => x"c73882e0",
          7593 => x"98088429",
          7594 => x"82f7e005",
          7595 => x"70085553",
          7596 => x"8c567380",
          7597 => x"2e87b138",
          7598 => x"73750c76",
          7599 => x"81fe0674",
          7600 => x"33545772",
          7601 => x"802eae38",
          7602 => x"81143351",
          7603 => x"c6a03f82",
          7604 => x"e0980881",
          7605 => x"ff067081",
          7606 => x"06545572",
          7607 => x"98387680",
          7608 => x"2e878338",
          7609 => x"74822a70",
          7610 => x"81065153",
          7611 => x"8a567286",
          7612 => x"f73886f2",
          7613 => x"39807434",
          7614 => x"77185982",
          7615 => x"e08c1933",
          7616 => x"81153481",
          7617 => x"52811433",
          7618 => x"51c6813f",
          7619 => x"82e09808",
          7620 => x"81ff0670",
          7621 => x"81065455",
          7622 => x"83567286",
          7623 => x"cb387680",
          7624 => x"2e8f3874",
          7625 => x"822a7081",
          7626 => x"0651538a",
          7627 => x"567286b8",
          7628 => x"38807053",
          7629 => x"74525bfd",
          7630 => x"9c3f82e0",
          7631 => x"980881ff",
          7632 => x"06577682",
          7633 => x"2e933876",
          7634 => x"8126819c",
          7635 => x"3882e08d",
          7636 => x"19335372",
          7637 => x"7b2e8190",
          7638 => x"388c3d74",
          7639 => x"56598356",
          7640 => x"83fa1533",
          7641 => x"70585372",
          7642 => x"802e8d38",
          7643 => x"83fe1551",
          7644 => x"cba93f82",
          7645 => x"e0980857",
          7646 => x"76797084",
          7647 => x"055b0cff",
          7648 => x"16901656",
          7649 => x"56758025",
          7650 => x"d7387718",
          7651 => x"82e08d11",
          7652 => x"33703070",
          7653 => x"9f2a7271",
          7654 => x"31953d71",
          7655 => x"842905f0",
          7656 => x"055a5351",
          7657 => x"55575974",
          7658 => x"085b8357",
          7659 => x"7a802e90",
          7660 => x"387a5273",
          7661 => x"51fc9e3f",
          7662 => x"82e09808",
          7663 => x"81ff0657",
          7664 => x"800b82e0",
          7665 => x"8d1a3354",
          7666 => x"5872782e",
          7667 => x"09810683",
          7668 => x"38815881",
          7669 => x"77279138",
          7670 => x"77802e8c",
          7671 => x"38811684",
          7672 => x"16565683",
          7673 => x"7627c038",
          7674 => x"81567684",
          7675 => x"2e84f938",
          7676 => x"8d567681",
          7677 => x"2684f138",
          7678 => x"80c31451",
          7679 => x"ca863f82",
          7680 => x"e0980883",
          7681 => x"ffff0653",
          7682 => x"7284802e",
          7683 => x"09810684",
          7684 => x"d73880ce",
          7685 => x"1451c9ec",
          7686 => x"3f82e098",
          7687 => x"0883ffff",
          7688 => x"0658778d",
          7689 => x"3880dc14",
          7690 => x"51c9f03f",
          7691 => x"82e09808",
          7692 => x"5877a015",
          7693 => x"0c80c814",
          7694 => x"33821534",
          7695 => x"80c81433",
          7696 => x"ff117081",
          7697 => x"ff065154",
          7698 => x"558d5672",
          7699 => x"81268498",
          7700 => x"387481ff",
          7701 => x"06787129",
          7702 => x"80c51633",
          7703 => x"52595372",
          7704 => x"8a152372",
          7705 => x"802e8b38",
          7706 => x"ff137306",
          7707 => x"5372802e",
          7708 => x"86388d56",
          7709 => x"83f23980",
          7710 => x"c91451c9",
          7711 => x"873f82e0",
          7712 => x"98085382",
          7713 => x"e0980888",
          7714 => x"1523728f",
          7715 => x"06578d56",
          7716 => x"7683d538",
          7717 => x"80cb1451",
          7718 => x"c8ea3f82",
          7719 => x"e0980883",
          7720 => x"ffff0655",
          7721 => x"748d3880",
          7722 => x"d81451c8",
          7723 => x"ee3f82e0",
          7724 => x"98085580",
          7725 => x"c61451c8",
          7726 => x"cb3f82e0",
          7727 => x"980883ff",
          7728 => x"ff06538d",
          7729 => x"5672802e",
          7730 => x"839e3888",
          7731 => x"14227814",
          7732 => x"71842a05",
          7733 => x"5a5a7875",
          7734 => x"26838d38",
          7735 => x"8a142252",
          7736 => x"74793151",
          7737 => x"fed3ec3f",
          7738 => x"82e09808",
          7739 => x"5582e098",
          7740 => x"08802e82",
          7741 => x"f33882e0",
          7742 => x"980880ff",
          7743 => x"fffff526",
          7744 => x"83388357",
          7745 => x"7483fff5",
          7746 => x"26833882",
          7747 => x"57749ff5",
          7748 => x"26853881",
          7749 => x"5789398d",
          7750 => x"5676802e",
          7751 => x"82ca3882",
          7752 => x"15709c16",
          7753 => x"0c7ba416",
          7754 => x"0c731c70",
          7755 => x"a8170c7a",
          7756 => x"1db0170c",
          7757 => x"54557683",
          7758 => x"2e098106",
          7759 => x"af3880e2",
          7760 => x"1451c7c0",
          7761 => x"3f82e098",
          7762 => x"0883ffff",
          7763 => x"06538d56",
          7764 => x"72829538",
          7765 => x"79829138",
          7766 => x"80e41451",
          7767 => x"c7bd3f82",
          7768 => x"e09808ac",
          7769 => x"150c7482",
          7770 => x"2b53a239",
          7771 => x"8d567980",
          7772 => x"2e81f538",
          7773 => x"7713ac15",
          7774 => x"0c741553",
          7775 => x"76822e8d",
          7776 => x"38741015",
          7777 => x"70812a76",
          7778 => x"81060551",
          7779 => x"5383ff13",
          7780 => x"892a538d",
          7781 => x"5672a015",
          7782 => x"082681cc",
          7783 => x"38ff0b94",
          7784 => x"150cff0b",
          7785 => x"90150cff",
          7786 => x"800b8415",
          7787 => x"3476832e",
          7788 => x"09810681",
          7789 => x"923880e8",
          7790 => x"1451c6c8",
          7791 => x"3f82e098",
          7792 => x"0883ffff",
          7793 => x"06537281",
          7794 => x"2e098106",
          7795 => x"80f93881",
          7796 => x"1b527351",
          7797 => x"ca883f82",
          7798 => x"e0980880",
          7799 => x"ea3882e0",
          7800 => x"98088415",
          7801 => x"3484b614",
          7802 => x"51c6993f",
          7803 => x"82e09808",
          7804 => x"83ffff06",
          7805 => x"537282d4",
          7806 => x"d52e0981",
          7807 => x"0680c838",
          7808 => x"b81451c6",
          7809 => x"963f82e0",
          7810 => x"9808848b",
          7811 => x"85a4d22e",
          7812 => x"098106b3",
          7813 => x"38849c14",
          7814 => x"51c6803f",
          7815 => x"82e09808",
          7816 => x"868a85e4",
          7817 => x"f22e0981",
          7818 => x"069d3884",
          7819 => x"a01451c5",
          7820 => x"ea3f82e0",
          7821 => x"98089415",
          7822 => x"0c84a414",
          7823 => x"51c5dc3f",
          7824 => x"82e09808",
          7825 => x"90150c76",
          7826 => x"743482f7",
          7827 => x"f0228105",
          7828 => x"537282f7",
          7829 => x"f0237286",
          7830 => x"152382f7",
          7831 => x"f80b8c15",
          7832 => x"0c800b98",
          7833 => x"150c8056",
          7834 => x"7582e098",
          7835 => x"0c903d0d",
          7836 => x"04fb3d0d",
          7837 => x"77548955",
          7838 => x"73802eba",
          7839 => x"38730853",
          7840 => x"72802eb2",
          7841 => x"38723352",
          7842 => x"71802eaa",
          7843 => x"38861322",
          7844 => x"84152257",
          7845 => x"5271762e",
          7846 => x"0981069a",
          7847 => x"38811333",
          7848 => x"51ffbeca",
          7849 => x"3f82e098",
          7850 => x"08810652",
          7851 => x"71883871",
          7852 => x"74085455",
          7853 => x"83398053",
          7854 => x"7873710c",
          7855 => x"527482e0",
          7856 => x"980c873d",
          7857 => x"0d04fa3d",
          7858 => x"0d02ab05",
          7859 => x"337a5889",
          7860 => x"3dfc0552",
          7861 => x"56f49a3f",
          7862 => x"8b54800b",
          7863 => x"82e09808",
          7864 => x"24bc3882",
          7865 => x"e0980884",
          7866 => x"2982f7e0",
          7867 => x"05700855",
          7868 => x"5573802e",
          7869 => x"84388074",
          7870 => x"34785473",
          7871 => x"802e8438",
          7872 => x"80743478",
          7873 => x"750c7554",
          7874 => x"75802e92",
          7875 => x"38805389",
          7876 => x"3d705384",
          7877 => x"0551f6e4",
          7878 => x"3f82e098",
          7879 => x"08547382",
          7880 => x"e0980c88",
          7881 => x"3d0d04ea",
          7882 => x"3d0d6802",
          7883 => x"840580eb",
          7884 => x"05335959",
          7885 => x"89547880",
          7886 => x"2e84c838",
          7887 => x"77bf0670",
          7888 => x"54993dcc",
          7889 => x"05539a3d",
          7890 => x"84055258",
          7891 => x"f6ae3f82",
          7892 => x"e0980855",
          7893 => x"82e09808",
          7894 => x"84a4387a",
          7895 => x"5c69528c",
          7896 => x"3d705256",
          7897 => x"eab03f82",
          7898 => x"e0980855",
          7899 => x"82e09808",
          7900 => x"92380280",
          7901 => x"d7053370",
          7902 => x"982b5557",
          7903 => x"73802583",
          7904 => x"38865577",
          7905 => x"9c065473",
          7906 => x"802e81ab",
          7907 => x"3874802e",
          7908 => x"95387484",
          7909 => x"2e098106",
          7910 => x"aa387551",
          7911 => x"dfb13f82",
          7912 => x"e0980855",
          7913 => x"9e3902b2",
          7914 => x"05339106",
          7915 => x"547381b8",
          7916 => x"3877822a",
          7917 => x"70810651",
          7918 => x"5473802e",
          7919 => x"8e388855",
          7920 => x"83bc3977",
          7921 => x"88075874",
          7922 => x"83b43877",
          7923 => x"832a7081",
          7924 => x"06515473",
          7925 => x"802e81af",
          7926 => x"3862527a",
          7927 => x"51d6ed3f",
          7928 => x"82e09808",
          7929 => x"568288b2",
          7930 => x"0a52628e",
          7931 => x"0551c2f4",
          7932 => x"3f6254a0",
          7933 => x"0b8b1534",
          7934 => x"80536252",
          7935 => x"7a51d785",
          7936 => x"3f805262",
          7937 => x"9c0551c2",
          7938 => x"db3f7a54",
          7939 => x"810b8315",
          7940 => x"3475802e",
          7941 => x"80f1387a",
          7942 => x"b4110851",
          7943 => x"54805375",
          7944 => x"52983dd0",
          7945 => x"0551cc86",
          7946 => x"3f82e098",
          7947 => x"085582e0",
          7948 => x"980882ca",
          7949 => x"38b73974",
          7950 => x"82c43802",
          7951 => x"b2053370",
          7952 => x"842a7081",
          7953 => x"06515556",
          7954 => x"73802e86",
          7955 => x"38845582",
          7956 => x"ad397781",
          7957 => x"2a708106",
          7958 => x"51547380",
          7959 => x"2ea93875",
          7960 => x"81065473",
          7961 => x"802ea038",
          7962 => x"87558292",
          7963 => x"3973527a",
          7964 => x"51c4eb3f",
          7965 => x"82e09808",
          7966 => x"7bff1890",
          7967 => x"120c5555",
          7968 => x"82e09808",
          7969 => x"81f83877",
          7970 => x"832a7081",
          7971 => x"06515473",
          7972 => x"802e8638",
          7973 => x"7780c007",
          7974 => x"587ab411",
          7975 => x"08a01b0c",
          7976 => x"63a41b0c",
          7977 => x"63537052",
          7978 => x"57d5a13f",
          7979 => x"82e09808",
          7980 => x"82e09808",
          7981 => x"881b0c63",
          7982 => x"9c05525a",
          7983 => x"c0dd3f82",
          7984 => x"e0980882",
          7985 => x"e098088c",
          7986 => x"1b0c777a",
          7987 => x"0c568617",
          7988 => x"22841a23",
          7989 => x"77901a34",
          7990 => x"800b911a",
          7991 => x"34800b9c",
          7992 => x"1a0c800b",
          7993 => x"941a0c77",
          7994 => x"852a7081",
          7995 => x"06515473",
          7996 => x"802e818d",
          7997 => x"3882e098",
          7998 => x"08802e81",
          7999 => x"843882e0",
          8000 => x"9808941a",
          8001 => x"0c8a1722",
          8002 => x"70892b7b",
          8003 => x"525957a8",
          8004 => x"39765278",
          8005 => x"51c5e73f",
          8006 => x"82e09808",
          8007 => x"5782e098",
          8008 => x"08812683",
          8009 => x"38825582",
          8010 => x"e09808ff",
          8011 => x"2e098106",
          8012 => x"83387955",
          8013 => x"75783156",
          8014 => x"74307076",
          8015 => x"07802551",
          8016 => x"54777627",
          8017 => x"8a388170",
          8018 => x"7506555a",
          8019 => x"73c33876",
          8020 => x"981a0c74",
          8021 => x"a9387583",
          8022 => x"ff065473",
          8023 => x"802ea238",
          8024 => x"76527a51",
          8025 => x"c4ee3f82",
          8026 => x"e0980885",
          8027 => x"3882558e",
          8028 => x"3975892a",
          8029 => x"82e09808",
          8030 => x"059c1a0c",
          8031 => x"84398079",
          8032 => x"0c745473",
          8033 => x"82e0980c",
          8034 => x"983d0d04",
          8035 => x"f23d0d60",
          8036 => x"63656440",
          8037 => x"405d5980",
          8038 => x"7e0c903d",
          8039 => x"fc055278",
          8040 => x"51f9ce3f",
          8041 => x"82e09808",
          8042 => x"5582e098",
          8043 => x"088a3891",
          8044 => x"19335574",
          8045 => x"802e8638",
          8046 => x"745682c7",
          8047 => x"39901933",
          8048 => x"81065587",
          8049 => x"5674802e",
          8050 => x"82b93895",
          8051 => x"39820b91",
          8052 => x"1a348256",
          8053 => x"82ad3981",
          8054 => x"0b911a34",
          8055 => x"815682a3",
          8056 => x"398c1908",
          8057 => x"941a0831",
          8058 => x"55747c27",
          8059 => x"8338745c",
          8060 => x"7b802e82",
          8061 => x"8c389419",
          8062 => x"087083ff",
          8063 => x"06565674",
          8064 => x"81b4387e",
          8065 => x"8a1122ff",
          8066 => x"0577892a",
          8067 => x"065b5579",
          8068 => x"a8387587",
          8069 => x"38881908",
          8070 => x"558f3998",
          8071 => x"19085278",
          8072 => x"51c3db3f",
          8073 => x"82e09808",
          8074 => x"55817527",
          8075 => x"ff9f3874",
          8076 => x"ff2effa3",
          8077 => x"3874981a",
          8078 => x"0c981908",
          8079 => x"527e51c3",
          8080 => x"933f82e0",
          8081 => x"9808802e",
          8082 => x"ff833882",
          8083 => x"e098081a",
          8084 => x"7c892a59",
          8085 => x"5777802e",
          8086 => x"80d83877",
          8087 => x"1a7f8a11",
          8088 => x"22585c55",
          8089 => x"75752785",
          8090 => x"38757a31",
          8091 => x"58775476",
          8092 => x"537c5281",
          8093 => x"1b3351ff",
          8094 => x"b8913f82",
          8095 => x"e09808fe",
          8096 => x"d6387e83",
          8097 => x"11335656",
          8098 => x"74802ea0",
          8099 => x"38b41608",
          8100 => x"77315574",
          8101 => x"78279538",
          8102 => x"848053b8",
          8103 => x"1652b416",
          8104 => x"08773189",
          8105 => x"2b7d0551",
          8106 => x"ffbde83f",
          8107 => x"77892b56",
          8108 => x"ba39769c",
          8109 => x"1a0c9419",
          8110 => x"0883ff06",
          8111 => x"84807131",
          8112 => x"57557b76",
          8113 => x"2783387b",
          8114 => x"569c1908",
          8115 => x"527e51c0",
          8116 => x"8d3f82e0",
          8117 => x"9808fdff",
          8118 => x"38755394",
          8119 => x"190883ff",
          8120 => x"061fb805",
          8121 => x"527c51ff",
          8122 => x"bda93f7b",
          8123 => x"76317e08",
          8124 => x"177f0c76",
          8125 => x"1e941b08",
          8126 => x"18941c0c",
          8127 => x"5e5cfdf0",
          8128 => x"39805675",
          8129 => x"82e0980c",
          8130 => x"903d0d04",
          8131 => x"f23d0d60",
          8132 => x"63656440",
          8133 => x"405d5880",
          8134 => x"7e0c903d",
          8135 => x"fc055277",
          8136 => x"51f6ce3f",
          8137 => x"82e09808",
          8138 => x"5582e098",
          8139 => x"088a3891",
          8140 => x"18335574",
          8141 => x"802e8638",
          8142 => x"745683bf",
          8143 => x"39901833",
          8144 => x"70812a70",
          8145 => x"81065156",
          8146 => x"56875674",
          8147 => x"802e83ab",
          8148 => x"38953982",
          8149 => x"0b911934",
          8150 => x"8256839f",
          8151 => x"39810b91",
          8152 => x"19348156",
          8153 => x"83953994",
          8154 => x"18087c11",
          8155 => x"56567476",
          8156 => x"27843875",
          8157 => x"095c7b80",
          8158 => x"2e82f338",
          8159 => x"94180870",
          8160 => x"83ff0656",
          8161 => x"56748282",
          8162 => x"387e8a11",
          8163 => x"22ff0577",
          8164 => x"892a065c",
          8165 => x"557abf38",
          8166 => x"758c3888",
          8167 => x"18085574",
          8168 => x"9c387a52",
          8169 => x"85399818",
          8170 => x"08527751",
          8171 => x"c6ac3f82",
          8172 => x"e0980855",
          8173 => x"82e09808",
          8174 => x"802e82b2",
          8175 => x"3874812e",
          8176 => x"ff913874",
          8177 => x"ff2eff95",
          8178 => x"38749819",
          8179 => x"0c881808",
          8180 => x"85387488",
          8181 => x"190c7e55",
          8182 => x"b415089c",
          8183 => x"19082e09",
          8184 => x"81068e38",
          8185 => x"7451ffbd",
          8186 => x"853f82e0",
          8187 => x"9808feed",
          8188 => x"38981808",
          8189 => x"527e51ff",
          8190 => x"bfda3f82",
          8191 => x"e0980880",
          8192 => x"2efed038",
          8193 => x"82e09808",
          8194 => x"1b7c892a",
          8195 => x"5a577880",
          8196 => x"2e80d738",
          8197 => x"781b7f8a",
          8198 => x"1122585b",
          8199 => x"55757527",
          8200 => x"8538757b",
          8201 => x"31597854",
          8202 => x"76537c52",
          8203 => x"811a3351",
          8204 => x"ffb6c23f",
          8205 => x"82e09808",
          8206 => x"fea3387e",
          8207 => x"b4110878",
          8208 => x"31565674",
          8209 => x"79279c38",
          8210 => x"848053b4",
          8211 => x"16087731",
          8212 => x"892b7d05",
          8213 => x"52b81651",
          8214 => x"ffbab83f",
          8215 => x"7e55800b",
          8216 => x"83163478",
          8217 => x"892b5680",
          8218 => x"de398c18",
          8219 => x"08941908",
          8220 => x"2694387e",
          8221 => x"51ffbbf6",
          8222 => x"3f82e098",
          8223 => x"08fdde38",
          8224 => x"7e77b412",
          8225 => x"0c55769c",
          8226 => x"190c9418",
          8227 => x"0883ff06",
          8228 => x"84807131",
          8229 => x"57557b76",
          8230 => x"2783387b",
          8231 => x"569c1808",
          8232 => x"527e51ff",
          8233 => x"bcb83f82",
          8234 => x"e09808fd",
          8235 => x"b0387553",
          8236 => x"7c529418",
          8237 => x"0883ff06",
          8238 => x"1fb80551",
          8239 => x"ffb9d43f",
          8240 => x"7e55810b",
          8241 => x"8316347b",
          8242 => x"76317e08",
          8243 => x"177f0c76",
          8244 => x"1e941a08",
          8245 => x"1870941c",
          8246 => x"0c8c1b08",
          8247 => x"58585e5c",
          8248 => x"74762783",
          8249 => x"38755574",
          8250 => x"8c190cfd",
          8251 => x"89399018",
          8252 => x"3380c007",
          8253 => x"55749019",
          8254 => x"34805675",
          8255 => x"82e0980c",
          8256 => x"903d0d04",
          8257 => x"f83d0d7a",
          8258 => x"8b3dfc05",
          8259 => x"53705256",
          8260 => x"f2df3f82",
          8261 => x"e0980857",
          8262 => x"82e09808",
          8263 => x"81803890",
          8264 => x"16337086",
          8265 => x"2a708106",
          8266 => x"51555573",
          8267 => x"802e80ee",
          8268 => x"38a01608",
          8269 => x"527851ff",
          8270 => x"bba43f82",
          8271 => x"e0980857",
          8272 => x"82e09808",
          8273 => x"80d838a4",
          8274 => x"16088b11",
          8275 => x"33a00755",
          8276 => x"55738b16",
          8277 => x"34881608",
          8278 => x"53745275",
          8279 => x"0851cca5",
          8280 => x"3f8c1608",
          8281 => x"529c1551",
          8282 => x"ffb7f93f",
          8283 => x"8288b20a",
          8284 => x"52961551",
          8285 => x"ffb7ed3f",
          8286 => x"76529215",
          8287 => x"51ffb7c6",
          8288 => x"3f785481",
          8289 => x"0b831534",
          8290 => x"7851ffbb",
          8291 => x"983f82e0",
          8292 => x"98089017",
          8293 => x"3381bf06",
          8294 => x"55577390",
          8295 => x"17347682",
          8296 => x"e0980c8a",
          8297 => x"3d0d04fc",
          8298 => x"3d0d7670",
          8299 => x"5254fed4",
          8300 => x"3f82e098",
          8301 => x"085382e0",
          8302 => x"98089c38",
          8303 => x"863dfc05",
          8304 => x"527351f1",
          8305 => x"ac3f82e0",
          8306 => x"98085382",
          8307 => x"e0980887",
          8308 => x"3882e098",
          8309 => x"08740c72",
          8310 => x"82e0980c",
          8311 => x"863d0d04",
          8312 => x"ff3d0d84",
          8313 => x"3d51e689",
          8314 => x"3f8b5280",
          8315 => x"0b82e098",
          8316 => x"08248b38",
          8317 => x"82e09808",
          8318 => x"82f7f434",
          8319 => x"80527182",
          8320 => x"e0980c83",
          8321 => x"3d0d04ee",
          8322 => x"3d0d8053",
          8323 => x"943dcc05",
          8324 => x"52953d51",
          8325 => x"e8e63f82",
          8326 => x"e0980855",
          8327 => x"82e09808",
          8328 => x"80e03876",
          8329 => x"58645294",
          8330 => x"3dd00551",
          8331 => x"dce83f82",
          8332 => x"e0980855",
          8333 => x"82e09808",
          8334 => x"bc380280",
          8335 => x"c7053370",
          8336 => x"982b5556",
          8337 => x"73802589",
          8338 => x"38767a98",
          8339 => x"120c54b2",
          8340 => x"3902a205",
          8341 => x"3370842a",
          8342 => x"70810651",
          8343 => x"55567380",
          8344 => x"2e9e3876",
          8345 => x"7f537052",
          8346 => x"54c9e13f",
          8347 => x"82e09808",
          8348 => x"98150c8e",
          8349 => x"3982e098",
          8350 => x"08842e09",
          8351 => x"81068338",
          8352 => x"85557482",
          8353 => x"e0980c94",
          8354 => x"3d0d04ff",
          8355 => x"a33d0d80",
          8356 => x"e13d0880",
          8357 => x"e13d085b",
          8358 => x"5b807a34",
          8359 => x"805380df",
          8360 => x"3dfdb405",
          8361 => x"5280e03d",
          8362 => x"51e7d13f",
          8363 => x"82e09808",
          8364 => x"5782e098",
          8365 => x"0883a138",
          8366 => x"7b80d43d",
          8367 => x"0c7a7c98",
          8368 => x"110880d8",
          8369 => x"3d0c5558",
          8370 => x"80d53d08",
          8371 => x"5473802e",
          8372 => x"828338a0",
          8373 => x"5280d33d",
          8374 => x"705255c4",
          8375 => x"903f82e0",
          8376 => x"98085782",
          8377 => x"e0980882",
          8378 => x"ef3880d9",
          8379 => x"3d08527b",
          8380 => x"51ffb7ea",
          8381 => x"3f82e098",
          8382 => x"085782e0",
          8383 => x"980882d8",
          8384 => x"3880da3d",
          8385 => x"08527b51",
          8386 => x"c8c23f82",
          8387 => x"e0980880",
          8388 => x"d63d0c76",
          8389 => x"527451c3",
          8390 => x"d43f82e0",
          8391 => x"98085782",
          8392 => x"e0980882",
          8393 => x"b3388052",
          8394 => x"7451c9b6",
          8395 => x"3f82e098",
          8396 => x"085782e0",
          8397 => x"9808a738",
          8398 => x"80da3d08",
          8399 => x"527b51c8",
          8400 => x"8b3f7382",
          8401 => x"e098082e",
          8402 => x"a6387652",
          8403 => x"7451c4e8",
          8404 => x"3f82e098",
          8405 => x"085782e0",
          8406 => x"9808802e",
          8407 => x"c9387684",
          8408 => x"2e098106",
          8409 => x"86388257",
          8410 => x"81ee3976",
          8411 => x"81ea3880",
          8412 => x"df3dfdb8",
          8413 => x"05527451",
          8414 => x"d6a03f76",
          8415 => x"933d7811",
          8416 => x"82113351",
          8417 => x"565a5673",
          8418 => x"802e9238",
          8419 => x"0280c605",
          8420 => x"55811681",
          8421 => x"16703356",
          8422 => x"565673f5",
          8423 => x"38811654",
          8424 => x"73782681",
          8425 => x"99387580",
          8426 => x"2e9c3878",
          8427 => x"16820555",
          8428 => x"ff1880e1",
          8429 => x"3d0811ff",
          8430 => x"18ff1858",
          8431 => x"58555874",
          8432 => x"33743475",
          8433 => x"eb38ff18",
          8434 => x"80e13d08",
          8435 => x"115558af",
          8436 => x"7434fdf4",
          8437 => x"39777b2e",
          8438 => x"0981068d",
          8439 => x"38ff1880",
          8440 => x"e13d0811",
          8441 => x"5558af74",
          8442 => x"34800b82",
          8443 => x"f7f43370",
          8444 => x"842982d2",
          8445 => x"98057008",
          8446 => x"7033525c",
          8447 => x"56565673",
          8448 => x"762e8d38",
          8449 => x"8116701a",
          8450 => x"70335155",
          8451 => x"5673f538",
          8452 => x"82165473",
          8453 => x"7826a738",
          8454 => x"80557476",
          8455 => x"27913874",
          8456 => x"19547333",
          8457 => x"7a708105",
          8458 => x"5c348115",
          8459 => x"55ec39ba",
          8460 => x"7a708105",
          8461 => x"5c3474ff",
          8462 => x"2e098106",
          8463 => x"85389157",
          8464 => x"973980e0",
          8465 => x"3d081881",
          8466 => x"19595473",
          8467 => x"337a7081",
          8468 => x"055c347a",
          8469 => x"7826eb38",
          8470 => x"807a3476",
          8471 => x"82e0980c",
          8472 => x"80df3d0d",
          8473 => x"04f73d0d",
          8474 => x"7b7d8d3d",
          8475 => x"fc055471",
          8476 => x"535755eb",
          8477 => x"fc3f82e0",
          8478 => x"98085382",
          8479 => x"e0980882",
          8480 => x"fe389115",
          8481 => x"33537282",
          8482 => x"f6388c15",
          8483 => x"08547376",
          8484 => x"27923890",
          8485 => x"15337081",
          8486 => x"2a708106",
          8487 => x"51545772",
          8488 => x"83387356",
          8489 => x"94150854",
          8490 => x"80709417",
          8491 => x"0c587578",
          8492 => x"2e829b38",
          8493 => x"798a1122",
          8494 => x"70892b59",
          8495 => x"51537378",
          8496 => x"2eb73876",
          8497 => x"52ff1651",
          8498 => x"febc883f",
          8499 => x"82e09808",
          8500 => x"ff157854",
          8501 => x"70535553",
          8502 => x"febbf83f",
          8503 => x"82e09808",
          8504 => x"73269638",
          8505 => x"76307075",
          8506 => x"06709418",
          8507 => x"0c777131",
          8508 => x"98180857",
          8509 => x"585153b2",
          8510 => x"39881508",
          8511 => x"5473a738",
          8512 => x"73527451",
          8513 => x"ffbbd33f",
          8514 => x"82e09808",
          8515 => x"5482e098",
          8516 => x"08812e81",
          8517 => x"9d3882e0",
          8518 => x"9808ff2e",
          8519 => x"819e3882",
          8520 => x"e0980888",
          8521 => x"160c7398",
          8522 => x"160c7380",
          8523 => x"2e819f38",
          8524 => x"76762780",
          8525 => x"de387577",
          8526 => x"31941608",
          8527 => x"1894170c",
          8528 => x"90163370",
          8529 => x"812a7081",
          8530 => x"0651555a",
          8531 => x"5672802e",
          8532 => x"9b387352",
          8533 => x"7451ffbb",
          8534 => x"813f82e0",
          8535 => x"98085482",
          8536 => x"e0980895",
          8537 => x"3882e098",
          8538 => x"0856a839",
          8539 => x"73527451",
          8540 => x"ffb58b3f",
          8541 => x"82e09808",
          8542 => x"5473ff2e",
          8543 => x"bf388174",
          8544 => x"27b03879",
          8545 => x"53739c14",
          8546 => x"0827a738",
          8547 => x"7398160c",
          8548 => x"ff9e3994",
          8549 => x"15081694",
          8550 => x"160c7583",
          8551 => x"ff065372",
          8552 => x"802eab38",
          8553 => x"73527951",
          8554 => x"ffb4a93f",
          8555 => x"82e09808",
          8556 => x"9438820b",
          8557 => x"91163482",
          8558 => x"5380c439",
          8559 => x"810b9116",
          8560 => x"348153bb",
          8561 => x"3975892a",
          8562 => x"82e09808",
          8563 => x"05589415",
          8564 => x"08548c15",
          8565 => x"08742790",
          8566 => x"38738c16",
          8567 => x"0c901533",
          8568 => x"80c00753",
          8569 => x"72901634",
          8570 => x"7383ff06",
          8571 => x"5372802e",
          8572 => x"8c38779c",
          8573 => x"16082e85",
          8574 => x"38779c16",
          8575 => x"0c805372",
          8576 => x"82e0980c",
          8577 => x"8b3d0d04",
          8578 => x"f93d0d79",
          8579 => x"56895475",
          8580 => x"802e818b",
          8581 => x"38805389",
          8582 => x"3dfc0552",
          8583 => x"8a3d8405",
          8584 => x"51e0d93f",
          8585 => x"82e09808",
          8586 => x"5582e098",
          8587 => x"0880eb38",
          8588 => x"77760c7a",
          8589 => x"527551d4",
          8590 => x"dd3f82e0",
          8591 => x"98085582",
          8592 => x"e0980880",
          8593 => x"c438ab16",
          8594 => x"3370982b",
          8595 => x"55578074",
          8596 => x"24a23886",
          8597 => x"16337084",
          8598 => x"2a708106",
          8599 => x"51555773",
          8600 => x"802eae38",
          8601 => x"9c160852",
          8602 => x"7751c1e0",
          8603 => x"3f82e098",
          8604 => x"0888170c",
          8605 => x"77548614",
          8606 => x"22841723",
          8607 => x"74527551",
          8608 => x"ffbcea3f",
          8609 => x"82e09808",
          8610 => x"5574842e",
          8611 => x"09810685",
          8612 => x"38855586",
          8613 => x"3974802e",
          8614 => x"84388076",
          8615 => x"0c745473",
          8616 => x"82e0980c",
          8617 => x"893d0d04",
          8618 => x"fc3d0d76",
          8619 => x"873dfc05",
          8620 => x"53705253",
          8621 => x"e7bb3f82",
          8622 => x"e0980887",
          8623 => x"3882e098",
          8624 => x"08730c86",
          8625 => x"3d0d04fb",
          8626 => x"3d0d7779",
          8627 => x"893dfc05",
          8628 => x"54715356",
          8629 => x"54e79a3f",
          8630 => x"82e09808",
          8631 => x"5382e098",
          8632 => x"0880e138",
          8633 => x"74943882",
          8634 => x"e0980852",
          8635 => x"7351ffbb",
          8636 => x"fc3f82e0",
          8637 => x"98085380",
          8638 => x"cb3982e0",
          8639 => x"98085273",
          8640 => x"51c1df3f",
          8641 => x"82e09808",
          8642 => x"5382e098",
          8643 => x"08842e09",
          8644 => x"81068538",
          8645 => x"80538739",
          8646 => x"82e09808",
          8647 => x"a7387452",
          8648 => x"7351cef6",
          8649 => x"3f725273",
          8650 => x"51ffbd8c",
          8651 => x"3f82e098",
          8652 => x"08843270",
          8653 => x"30707207",
          8654 => x"9f2c7082",
          8655 => x"e0980806",
          8656 => x"51515454",
          8657 => x"7282e098",
          8658 => x"0c873d0d",
          8659 => x"04ed3d0d",
          8660 => x"66578053",
          8661 => x"893d7053",
          8662 => x"973d5256",
          8663 => x"de9e3f82",
          8664 => x"e0980855",
          8665 => x"82e09808",
          8666 => x"b2386552",
          8667 => x"7551d2a6",
          8668 => x"3f82e098",
          8669 => x"085582e0",
          8670 => x"9808a038",
          8671 => x"0280cb05",
          8672 => x"3370982b",
          8673 => x"55587380",
          8674 => x"25853886",
          8675 => x"558d3976",
          8676 => x"802e8838",
          8677 => x"76527551",
          8678 => x"ce803f74",
          8679 => x"82e0980c",
          8680 => x"953d0d04",
          8681 => x"f03d0d63",
          8682 => x"65555c80",
          8683 => x"53923dec",
          8684 => x"0552933d",
          8685 => x"51ddc53f",
          8686 => x"82e09808",
          8687 => x"5b82e098",
          8688 => x"08828238",
          8689 => x"7c740c73",
          8690 => x"089c1108",
          8691 => x"fe119413",
          8692 => x"08595658",
          8693 => x"55757426",
          8694 => x"9138757c",
          8695 => x"0c81e639",
          8696 => x"815b81ce",
          8697 => x"39825b81",
          8698 => x"c93982e0",
          8699 => x"98087533",
          8700 => x"55597381",
          8701 => x"2e098106",
          8702 => x"80c03882",
          8703 => x"755f5776",
          8704 => x"52923df0",
          8705 => x"0551ffaf",
          8706 => x"f53f82e0",
          8707 => x"9808ff2e",
          8708 => x"cf3882e0",
          8709 => x"9808812e",
          8710 => x"cc3882e0",
          8711 => x"98083070",
          8712 => x"82e09808",
          8713 => x"0780257a",
          8714 => x"0581197f",
          8715 => x"53595a54",
          8716 => x"9c140877",
          8717 => x"26c93880",
          8718 => x"f939a815",
          8719 => x"0882e098",
          8720 => x"08575875",
          8721 => x"98387752",
          8722 => x"81187d52",
          8723 => x"58ffad8e",
          8724 => x"3f82e098",
          8725 => x"085b82e0",
          8726 => x"980880d6",
          8727 => x"387c7033",
          8728 => x"7712ff1a",
          8729 => x"5d525654",
          8730 => x"74822e09",
          8731 => x"81069e38",
          8732 => x"b81451ff",
          8733 => x"a98e3f82",
          8734 => x"e0980883",
          8735 => x"ffff0670",
          8736 => x"30708025",
          8737 => x"1b821959",
          8738 => x"5b51549b",
          8739 => x"39b81451",
          8740 => x"ffa9883f",
          8741 => x"82e09808",
          8742 => x"f00a0670",
          8743 => x"30708025",
          8744 => x"1b841959",
          8745 => x"5b515475",
          8746 => x"83ff067a",
          8747 => x"585679ff",
          8748 => x"9238787c",
          8749 => x"0c7c7994",
          8750 => x"120c8411",
          8751 => x"33810756",
          8752 => x"54748415",
          8753 => x"347a82e0",
          8754 => x"980c923d",
          8755 => x"0d04f93d",
          8756 => x"0d798a3d",
          8757 => x"fc055370",
          8758 => x"5257e395",
          8759 => x"3f82e098",
          8760 => x"085682e0",
          8761 => x"980881aa",
          8762 => x"38911733",
          8763 => x"567581a2",
          8764 => x"38901733",
          8765 => x"70812a70",
          8766 => x"81065155",
          8767 => x"55875573",
          8768 => x"802e8190",
          8769 => x"38941708",
          8770 => x"54738c18",
          8771 => x"08278182",
          8772 => x"38739c38",
          8773 => x"82e09808",
          8774 => x"53881708",
          8775 => x"527651ff",
          8776 => x"b28c3f82",
          8777 => x"e0980874",
          8778 => x"88190c56",
          8779 => x"80ca3998",
          8780 => x"17085276",
          8781 => x"51ffadc6",
          8782 => x"3f82e098",
          8783 => x"08ff2e09",
          8784 => x"81068338",
          8785 => x"815682e0",
          8786 => x"9808812e",
          8787 => x"09810685",
          8788 => x"388256a4",
          8789 => x"3975a138",
          8790 => x"775482e0",
          8791 => x"98089c15",
          8792 => x"08279538",
          8793 => x"98170853",
          8794 => x"82e09808",
          8795 => x"527651ff",
          8796 => x"b1bc3f82",
          8797 => x"e0980856",
          8798 => x"9417088c",
          8799 => x"180c9017",
          8800 => x"3380c007",
          8801 => x"54739018",
          8802 => x"3475802e",
          8803 => x"85387591",
          8804 => x"18347555",
          8805 => x"7482e098",
          8806 => x"0c893d0d",
          8807 => x"04e03d0d",
          8808 => x"8253a23d",
          8809 => x"ff9c0552",
          8810 => x"a33d51d9",
          8811 => x"cf3f82e0",
          8812 => x"98085582",
          8813 => x"e0980881",
          8814 => x"f9387846",
          8815 => x"a33d0852",
          8816 => x"963d7052",
          8817 => x"58cdcf3f",
          8818 => x"82e09808",
          8819 => x"5582e098",
          8820 => x"0881df38",
          8821 => x"0280ff05",
          8822 => x"3370852a",
          8823 => x"70810651",
          8824 => x"55568655",
          8825 => x"7381cb38",
          8826 => x"75982b54",
          8827 => x"80742481",
          8828 => x"c1380280",
          8829 => x"da053370",
          8830 => x"81065854",
          8831 => x"87557681",
          8832 => x"b1386c52",
          8833 => x"7851ffba",
          8834 => x"c33f82e0",
          8835 => x"98087484",
          8836 => x"2a708106",
          8837 => x"51555673",
          8838 => x"802e80d6",
          8839 => x"38785482",
          8840 => x"e0980898",
          8841 => x"15082e81",
          8842 => x"8938735a",
          8843 => x"82e09808",
          8844 => x"5c76528a",
          8845 => x"3d705254",
          8846 => x"ffb5b23f",
          8847 => x"82e09808",
          8848 => x"5582e098",
          8849 => x"0880eb38",
          8850 => x"82e09808",
          8851 => x"527351ff",
          8852 => x"bb903f82",
          8853 => x"e0980855",
          8854 => x"82e09808",
          8855 => x"86388755",
          8856 => x"80d03982",
          8857 => x"e0980884",
          8858 => x"2e883882",
          8859 => x"e0980880",
          8860 => x"c1387751",
          8861 => x"c7ab3f82",
          8862 => x"e0980882",
          8863 => x"e0980830",
          8864 => x"7082e098",
          8865 => x"08078025",
          8866 => x"51555575",
          8867 => x"802e9538",
          8868 => x"73802e90",
          8869 => x"38805375",
          8870 => x"527751ff",
          8871 => x"af903f82",
          8872 => x"e0980855",
          8873 => x"748c3878",
          8874 => x"51ffa8f9",
          8875 => x"3f82e098",
          8876 => x"08557482",
          8877 => x"e0980ca2",
          8878 => x"3d0d04e8",
          8879 => x"3d0d8253",
          8880 => x"9a3dffbc",
          8881 => x"05529b3d",
          8882 => x"51d7b13f",
          8883 => x"82e09808",
          8884 => x"5482e098",
          8885 => x"0882b738",
          8886 => x"785e6a52",
          8887 => x"8e3d7052",
          8888 => x"58cbb33f",
          8889 => x"82e09808",
          8890 => x"5482e098",
          8891 => x"08863888",
          8892 => x"54829b39",
          8893 => x"82e09808",
          8894 => x"842e0981",
          8895 => x"06828f38",
          8896 => x"0280df05",
          8897 => x"3370852a",
          8898 => x"81065155",
          8899 => x"86547481",
          8900 => x"fd38785a",
          8901 => x"74528a3d",
          8902 => x"705257ff",
          8903 => x"afbc3f82",
          8904 => x"e0980875",
          8905 => x"555682e0",
          8906 => x"98088338",
          8907 => x"875482e0",
          8908 => x"9808812e",
          8909 => x"09810683",
          8910 => x"38825482",
          8911 => x"e09808ff",
          8912 => x"2e098106",
          8913 => x"86388154",
          8914 => x"81ba3973",
          8915 => x"81b63882",
          8916 => x"e0980852",
          8917 => x"7851ffb2",
          8918 => x"9c3f82e0",
          8919 => x"98085482",
          8920 => x"e0980881",
          8921 => x"9f388b53",
          8922 => x"a052b819",
          8923 => x"51ffa4c6",
          8924 => x"3f7854ae",
          8925 => x"0bb81534",
          8926 => x"7854900b",
          8927 => x"80c31534",
          8928 => x"8288b20a",
          8929 => x"5280ce19",
          8930 => x"51ffa3d8",
          8931 => x"3f755378",
          8932 => x"b8115351",
          8933 => x"ffb7ee3f",
          8934 => x"a05378b8",
          8935 => x"115380d8",
          8936 => x"0551ffa3",
          8937 => x"ee3f7854",
          8938 => x"ae0b80d9",
          8939 => x"15347f53",
          8940 => x"7880d811",
          8941 => x"5351ffb7",
          8942 => x"cc3f7854",
          8943 => x"810b8315",
          8944 => x"347751ff",
          8945 => x"bf893f82",
          8946 => x"e0980854",
          8947 => x"82e09808",
          8948 => x"b3388288",
          8949 => x"b20a5264",
          8950 => x"960551ff",
          8951 => x"a3863f75",
          8952 => x"53645278",
          8953 => x"51ffb79d",
          8954 => x"3f645490",
          8955 => x"0b8b1534",
          8956 => x"7854810b",
          8957 => x"83153478",
          8958 => x"51ffa6a9",
          8959 => x"3f82e098",
          8960 => x"08548b39",
          8961 => x"80537552",
          8962 => x"7651ffac",
          8963 => x"a13f7382",
          8964 => x"e0980c9a",
          8965 => x"3d0d04d8",
          8966 => x"3d0dab3d",
          8967 => x"840551d1",
          8968 => x"d03f8253",
          8969 => x"aa3dfefc",
          8970 => x"0552ab3d",
          8971 => x"51d4cd3f",
          8972 => x"82e09808",
          8973 => x"5582e098",
          8974 => x"0882d838",
          8975 => x"784eab3d",
          8976 => x"08529e3d",
          8977 => x"705258c8",
          8978 => x"cd3f82e0",
          8979 => x"98085582",
          8980 => x"e0980882",
          8981 => x"be380281",
          8982 => x"9f053381",
          8983 => x"a0065486",
          8984 => x"557382af",
          8985 => x"38a053a5",
          8986 => x"3d0852aa",
          8987 => x"3dff8005",
          8988 => x"51ffa29f",
          8989 => x"3fb05377",
          8990 => x"52923d70",
          8991 => x"5254ffa2",
          8992 => x"923fac3d",
          8993 => x"08527351",
          8994 => x"c88c3f82",
          8995 => x"e0980855",
          8996 => x"82e09808",
          8997 => x"973863a1",
          8998 => x"3d082e09",
          8999 => x"81068838",
          9000 => x"65a33d08",
          9001 => x"2e923888",
          9002 => x"5581e839",
          9003 => x"82e09808",
          9004 => x"842e0981",
          9005 => x"0681bb38",
          9006 => x"7351ffbd",
          9007 => x"923f82e0",
          9008 => x"98085582",
          9009 => x"e0980881",
          9010 => x"ca386856",
          9011 => x"9353aa3d",
          9012 => x"ff8d0552",
          9013 => x"8d1651ff",
          9014 => x"a1b93f02",
          9015 => x"af05338b",
          9016 => x"17348b16",
          9017 => x"3370842a",
          9018 => x"70810651",
          9019 => x"55557389",
          9020 => x"3874a007",
          9021 => x"54738b17",
          9022 => x"34785481",
          9023 => x"0b831534",
          9024 => x"8b163370",
          9025 => x"842a7081",
          9026 => x"06515555",
          9027 => x"73802e80",
          9028 => x"e7386f64",
          9029 => x"2e80e138",
          9030 => x"75527851",
          9031 => x"ffb4ad3f",
          9032 => x"82e09808",
          9033 => x"527851ff",
          9034 => x"a5aa3f82",
          9035 => x"5582e098",
          9036 => x"08802e80",
          9037 => x"de3882e0",
          9038 => x"98085278",
          9039 => x"51ffa39e",
          9040 => x"3f82e098",
          9041 => x"087980d8",
          9042 => x"11585855",
          9043 => x"82e09808",
          9044 => x"80c13881",
          9045 => x"16335473",
          9046 => x"ae2e0981",
          9047 => x"069a3863",
          9048 => x"53755276",
          9049 => x"51ffb49d",
          9050 => x"3f785481",
          9051 => x"0b831534",
          9052 => x"873982e0",
          9053 => x"98089c38",
          9054 => x"7751c1a5",
          9055 => x"3f82e098",
          9056 => x"085582e0",
          9057 => x"98088c38",
          9058 => x"7851ffa3",
          9059 => x"983f82e0",
          9060 => x"98085574",
          9061 => x"82e0980c",
          9062 => x"aa3d0d04",
          9063 => x"ec3d0d02",
          9064 => x"80df0533",
          9065 => x"02840580",
          9066 => x"e3053357",
          9067 => x"57825396",
          9068 => x"3dcc0552",
          9069 => x"973d51d1",
          9070 => x"c33f82e0",
          9071 => x"98085582",
          9072 => x"e0980880",
          9073 => x"cf38785a",
          9074 => x"6652963d",
          9075 => x"d00551c5",
          9076 => x"c53f82e0",
          9077 => x"98085582",
          9078 => x"e09808b8",
          9079 => x"380280cf",
          9080 => x"053381a0",
          9081 => x"06548655",
          9082 => x"73aa3875",
          9083 => x"a7066171",
          9084 => x"098b1233",
          9085 => x"71067a74",
          9086 => x"06075157",
          9087 => x"5556748b",
          9088 => x"15347854",
          9089 => x"810b8315",
          9090 => x"347851ff",
          9091 => x"a2973f82",
          9092 => x"e0980855",
          9093 => x"7482e098",
          9094 => x"0c963d0d",
          9095 => x"04ee3d0d",
          9096 => x"65568253",
          9097 => x"943dcc05",
          9098 => x"52953d51",
          9099 => x"d0ce3f82",
          9100 => x"e0980855",
          9101 => x"82e09808",
          9102 => x"80cb3876",
          9103 => x"58645294",
          9104 => x"3dd00551",
          9105 => x"c4d03f82",
          9106 => x"e0980855",
          9107 => x"82e09808",
          9108 => x"b4380280",
          9109 => x"c7053381",
          9110 => x"a0065486",
          9111 => x"5573a638",
          9112 => x"84162286",
          9113 => x"17227190",
          9114 => x"2b075354",
          9115 => x"961f51ff",
          9116 => x"9df23f76",
          9117 => x"54810b83",
          9118 => x"15347651",
          9119 => x"ffa1a63f",
          9120 => x"82e09808",
          9121 => x"557482e0",
          9122 => x"980c943d",
          9123 => x"0d04e93d",
          9124 => x"0d6a6c5c",
          9125 => x"5a805399",
          9126 => x"3dcc0552",
          9127 => x"9a3d51cf",
          9128 => x"db3f82e0",
          9129 => x"980882e0",
          9130 => x"98083070",
          9131 => x"82e09808",
          9132 => x"07802551",
          9133 => x"55577980",
          9134 => x"2e818638",
          9135 => x"81707506",
          9136 => x"55557380",
          9137 => x"2e80fa38",
          9138 => x"7b5d805f",
          9139 => x"80528d3d",
          9140 => x"705254ff",
          9141 => x"ac973f82",
          9142 => x"e0980857",
          9143 => x"82e09808",
          9144 => x"80d23874",
          9145 => x"527351ff",
          9146 => x"b1f83f82",
          9147 => x"e0980857",
          9148 => x"82e09808",
          9149 => x"bf3882e0",
          9150 => x"980882e0",
          9151 => x"9808655b",
          9152 => x"59567818",
          9153 => x"81197b18",
          9154 => x"56595574",
          9155 => x"33743481",
          9156 => x"16568a78",
          9157 => x"27ec388b",
          9158 => x"56751a54",
          9159 => x"80743475",
          9160 => x"802e9e38",
          9161 => x"ff16701b",
          9162 => x"70335155",
          9163 => x"5673a02e",
          9164 => x"e8388e39",
          9165 => x"76842e09",
          9166 => x"81068638",
          9167 => x"807a3480",
          9168 => x"57763070",
          9169 => x"78078025",
          9170 => x"51547a80",
          9171 => x"2e80c138",
          9172 => x"73802ebc",
          9173 => x"387ba411",
          9174 => x"085351ff",
          9175 => x"9f803f82",
          9176 => x"e0980857",
          9177 => x"82e09808",
          9178 => x"a7387b70",
          9179 => x"33555580",
          9180 => x"c3567383",
          9181 => x"2e8b3880",
          9182 => x"e4567384",
          9183 => x"2e8338a7",
          9184 => x"567515b8",
          9185 => x"0551ff9b",
          9186 => x"923f82e0",
          9187 => x"98087b0c",
          9188 => x"7682e098",
          9189 => x"0c993d0d",
          9190 => x"04e63d0d",
          9191 => x"82539c3d",
          9192 => x"ffb40552",
          9193 => x"9d3d51cd",
          9194 => x"d33f82e0",
          9195 => x"980882e0",
          9196 => x"98085654",
          9197 => x"82e09808",
          9198 => x"82dd388b",
          9199 => x"53a0528a",
          9200 => x"3d705258",
          9201 => x"ff9bef3f",
          9202 => x"736d7033",
          9203 => x"5155569f",
          9204 => x"74278186",
          9205 => x"3877579d",
          9206 => x"3d51ff9c",
          9207 => x"cc3f82e0",
          9208 => x"980883ff",
          9209 => x"ff2680c4",
          9210 => x"3882e098",
          9211 => x"085196c0",
          9212 => x"3f83b552",
          9213 => x"82e09808",
          9214 => x"5195903f",
          9215 => x"82e09808",
          9216 => x"83ffff06",
          9217 => x"5574802e",
          9218 => x"a3387452",
          9219 => x"82d3b851",
          9220 => x"ff9bee3f",
          9221 => x"82e09808",
          9222 => x"933881ff",
          9223 => x"75278838",
          9224 => x"75892688",
          9225 => x"388b398a",
          9226 => x"76278638",
          9227 => x"865581e7",
          9228 => x"3981ff75",
          9229 => x"278f3874",
          9230 => x"882a5473",
          9231 => x"77708105",
          9232 => x"59348116",
          9233 => x"56747770",
          9234 => x"81055934",
          9235 => x"81166d70",
          9236 => x"33515556",
          9237 => x"739f26fe",
          9238 => x"fe388a3d",
          9239 => x"33548655",
          9240 => x"7381e52e",
          9241 => x"81b13875",
          9242 => x"802e9938",
          9243 => x"02a30555",
          9244 => x"75157033",
          9245 => x"515473a0",
          9246 => x"2e098106",
          9247 => x"8738ff16",
          9248 => x"5675ed38",
          9249 => x"78408042",
          9250 => x"8052903d",
          9251 => x"705255ff",
          9252 => x"a8db3f82",
          9253 => x"e0980854",
          9254 => x"82e09808",
          9255 => x"80f73881",
          9256 => x"527451ff",
          9257 => x"aebc3f82",
          9258 => x"e0980854",
          9259 => x"82e09808",
          9260 => x"8d387580",
          9261 => x"c4386654",
          9262 => x"e5743480",
          9263 => x"c63982e0",
          9264 => x"9808842e",
          9265 => x"09810680",
          9266 => x"cc388054",
          9267 => x"75742e80",
          9268 => x"c4388152",
          9269 => x"7451ffab",
          9270 => x"d83f82e0",
          9271 => x"98085482",
          9272 => x"e09808b1",
          9273 => x"38a05382",
          9274 => x"e0980852",
          9275 => x"6651ff99",
          9276 => x"c53f6654",
          9277 => x"880b8b15",
          9278 => x"348b5377",
          9279 => x"526651ff",
          9280 => x"99913f78",
          9281 => x"54810b83",
          9282 => x"15347851",
          9283 => x"ff9c963f",
          9284 => x"82e09808",
          9285 => x"54735574",
          9286 => x"82e0980c",
          9287 => x"9c3d0d04",
          9288 => x"f23d0d60",
          9289 => x"62028805",
          9290 => x"80cb0533",
          9291 => x"933dfc05",
          9292 => x"55725440",
          9293 => x"5e5ad2b9",
          9294 => x"3f82e098",
          9295 => x"085882e0",
          9296 => x"980882bd",
          9297 => x"38911a33",
          9298 => x"587782b5",
          9299 => x"387c802e",
          9300 => x"97388c1a",
          9301 => x"08597890",
          9302 => x"38901a33",
          9303 => x"70812a70",
          9304 => x"81065155",
          9305 => x"55739038",
          9306 => x"87548297",
          9307 => x"39825882",
          9308 => x"90398158",
          9309 => x"828b397e",
          9310 => x"8a112270",
          9311 => x"892b7055",
          9312 => x"7f545656",
          9313 => x"56fea2cb",
          9314 => x"3fff147d",
          9315 => x"06703070",
          9316 => x"72079f2a",
          9317 => x"82e09808",
          9318 => x"05901908",
          9319 => x"7c405a5d",
          9320 => x"55558177",
          9321 => x"2788389c",
          9322 => x"16087726",
          9323 => x"83388257",
          9324 => x"76775659",
          9325 => x"80567452",
          9326 => x"7951ff9c",
          9327 => x"c13f8115",
          9328 => x"7f55559c",
          9329 => x"14087526",
          9330 => x"83388255",
          9331 => x"82e09808",
          9332 => x"812eff99",
          9333 => x"3882e098",
          9334 => x"08ff2eff",
          9335 => x"953882e0",
          9336 => x"98088e38",
          9337 => x"81165675",
          9338 => x"7b2e0981",
          9339 => x"06873893",
          9340 => x"39745980",
          9341 => x"5674772e",
          9342 => x"098106ff",
          9343 => x"b9388758",
          9344 => x"80ff397d",
          9345 => x"802eba38",
          9346 => x"787b5555",
          9347 => x"7a802eb4",
          9348 => x"38811556",
          9349 => x"73812e09",
          9350 => x"81068338",
          9351 => x"ff567553",
          9352 => x"74527e51",
          9353 => x"ff9dd03f",
          9354 => x"82e09808",
          9355 => x"5882e098",
          9356 => x"0880ce38",
          9357 => x"748116ff",
          9358 => x"1656565c",
          9359 => x"73d33884",
          9360 => x"39ff195c",
          9361 => x"7e7c9012",
          9362 => x"0c557d80",
          9363 => x"2eb33878",
          9364 => x"881b0c7c",
          9365 => x"8c1b0c90",
          9366 => x"1a3380c0",
          9367 => x"07547390",
          9368 => x"1b349c15",
          9369 => x"08fe0594",
          9370 => x"16085754",
          9371 => x"75742691",
          9372 => x"38757b31",
          9373 => x"94160c84",
          9374 => x"15338107",
          9375 => x"54738416",
          9376 => x"34775473",
          9377 => x"82e0980c",
          9378 => x"903d0d04",
          9379 => x"e83d0d6c",
          9380 => x"6e028805",
          9381 => x"80ef0533",
          9382 => x"9e3d5445",
          9383 => x"5c59c4d1",
          9384 => x"3f8b5680",
          9385 => x"0b82e098",
          9386 => x"08248da0",
          9387 => x"3882e098",
          9388 => x"08842982",
          9389 => x"f7e00570",
          9390 => x"08515574",
          9391 => x"802e8438",
          9392 => x"80753482",
          9393 => x"e0980882",
          9394 => x"e0980805",
          9395 => x"82e08c11",
          9396 => x"3382e08d",
          9397 => x"12334741",
          9398 => x"5581527f",
          9399 => x"51ff8eac",
          9400 => x"3f82e098",
          9401 => x"0881ff06",
          9402 => x"70810656",
          9403 => x"57835674",
          9404 => x"8cda3876",
          9405 => x"822a7081",
          9406 => x"0651558a",
          9407 => x"56748ccc",
          9408 => x"389a3dfc",
          9409 => x"05538352",
          9410 => x"7f51ff92",
          9411 => x"cc3f82e0",
          9412 => x"98089938",
          9413 => x"68557480",
          9414 => x"2e923874",
          9415 => x"82808026",
          9416 => x"8b38ff15",
          9417 => x"75065574",
          9418 => x"802e8338",
          9419 => x"81497880",
          9420 => x"2e873884",
          9421 => x"80792692",
          9422 => x"38788180",
          9423 => x"0a268b38",
          9424 => x"ff197906",
          9425 => x"5574802e",
          9426 => x"86389356",
          9427 => x"8bfe3978",
          9428 => x"892a6f89",
          9429 => x"2a70892b",
          9430 => x"77594943",
          9431 => x"597a8338",
          9432 => x"81566130",
          9433 => x"70802577",
          9434 => x"07515591",
          9435 => x"56748bdc",
          9436 => x"3864802e",
          9437 => x"80e03881",
          9438 => x"5474537a",
          9439 => x"527f51ff",
          9440 => x"8e893f81",
          9441 => x"5682e098",
          9442 => x"088bc138",
          9443 => x"83fe1b51",
          9444 => x"ff92f13f",
          9445 => x"82e09808",
          9446 => x"83ffff06",
          9447 => x"558e5674",
          9448 => x"82d4d52e",
          9449 => x"0981068b",
          9450 => x"a3386490",
          9451 => x"291b83b2",
          9452 => x"11335657",
          9453 => x"74802e8b",
          9454 => x"933883b6",
          9455 => x"1751ff92",
          9456 => x"da3f82e0",
          9457 => x"980883ba",
          9458 => x"18525fff",
          9459 => x"92cd3f82",
          9460 => x"e0980848",
          9461 => x"b7399a3d",
          9462 => x"f8055381",
          9463 => x"527f51ff",
          9464 => x"90f73f81",
          9465 => x"5682e098",
          9466 => x"088ae138",
          9467 => x"62832a70",
          9468 => x"770682e0",
          9469 => x"98084151",
          9470 => x"55748338",
          9471 => x"bf5f6755",
          9472 => x"8e567e75",
          9473 => x"268ac538",
          9474 => x"747f3148",
          9475 => x"8e5680ff",
          9476 => x"68278ab8",
          9477 => x"38935678",
          9478 => x"8180268a",
          9479 => x"af386281",
          9480 => x"2a708106",
          9481 => x"56447480",
          9482 => x"2e953862",
          9483 => x"87065574",
          9484 => x"822e838d",
          9485 => x"38628106",
          9486 => x"5574802e",
          9487 => x"83833862",
          9488 => x"81065593",
          9489 => x"56825e74",
          9490 => x"802e8a80",
          9491 => x"38785a7d",
          9492 => x"832e0981",
          9493 => x"0680e138",
          9494 => x"78ae3867",
          9495 => x"912a5781",
          9496 => x"0b82d3dc",
          9497 => x"22565a74",
          9498 => x"802e9d38",
          9499 => x"74772698",
          9500 => x"3882d3dc",
          9501 => x"56791082",
          9502 => x"17702257",
          9503 => x"575a7480",
          9504 => x"2e863876",
          9505 => x"7527ee38",
          9506 => x"79526751",
          9507 => x"fe9cc43f",
          9508 => x"82e09808",
          9509 => x"84298487",
          9510 => x"0570892a",
          9511 => x"5e55a05c",
          9512 => x"800b82e0",
          9513 => x"9808fc80",
          9514 => x"8a055646",
          9515 => x"fdfff00a",
          9516 => x"752780ec",
          9517 => x"38898839",
          9518 => x"78ae3867",
          9519 => x"8c2a5781",
          9520 => x"0b82d3cc",
          9521 => x"22565a74",
          9522 => x"802e9d38",
          9523 => x"74772698",
          9524 => x"3882d3cc",
          9525 => x"56791082",
          9526 => x"17702257",
          9527 => x"575a7480",
          9528 => x"2e863876",
          9529 => x"7527ee38",
          9530 => x"79526751",
          9531 => x"fe9be43f",
          9532 => x"82e09808",
          9533 => x"10840557",
          9534 => x"82e09808",
          9535 => x"9ff52696",
          9536 => x"38810b82",
          9537 => x"e0980810",
          9538 => x"82e09808",
          9539 => x"05711172",
          9540 => x"2a830559",
          9541 => x"565e83ff",
          9542 => x"17892a5d",
          9543 => x"815ca046",
          9544 => x"7b1f7d11",
          9545 => x"67056a70",
          9546 => x"12ff0571",
          9547 => x"30707206",
          9548 => x"74315c52",
          9549 => x"59575941",
          9550 => x"7d832e09",
          9551 => x"81068938",
          9552 => x"761c6118",
          9553 => x"425c8439",
          9554 => x"761d5d79",
          9555 => x"90291870",
          9556 => x"60316958",
          9557 => x"51557476",
          9558 => x"2687e438",
          9559 => x"757c317d",
          9560 => x"317a5370",
          9561 => x"67315255",
          9562 => x"fe9ae83f",
          9563 => x"82e09808",
          9564 => x"587d832e",
          9565 => x"0981069b",
          9566 => x"3882e098",
          9567 => x"0883fff5",
          9568 => x"2680dd38",
          9569 => x"7887b838",
          9570 => x"79812a59",
          9571 => x"78fdbe38",
          9572 => x"87ad397d",
          9573 => x"822e0981",
          9574 => x"0680c538",
          9575 => x"83fff50b",
          9576 => x"82e09808",
          9577 => x"27a03878",
          9578 => x"8f38791a",
          9579 => x"557480c0",
          9580 => x"26863874",
          9581 => x"59fd9639",
          9582 => x"63810655",
          9583 => x"74802e8f",
          9584 => x"38835efd",
          9585 => x"883982e0",
          9586 => x"98089ff5",
          9587 => x"26923878",
          9588 => x"86ed3879",
          9589 => x"1a598180",
          9590 => x"7927fcf1",
          9591 => x"3886e039",
          9592 => x"80557d81",
          9593 => x"2e098106",
          9594 => x"83387d55",
          9595 => x"9ff57827",
          9596 => x"8b387481",
          9597 => x"06558e56",
          9598 => x"7486d138",
          9599 => x"84805380",
          9600 => x"527a51ff",
          9601 => x"8fb03f8b",
          9602 => x"5382d1e4",
          9603 => x"527a51ff",
          9604 => x"8f813f84",
          9605 => x"80528b1b",
          9606 => x"51ff8eaa",
          9607 => x"3f798d1c",
          9608 => x"347b83ff",
          9609 => x"ff06528e",
          9610 => x"1b51ff8e",
          9611 => x"993f810b",
          9612 => x"901c347d",
          9613 => x"83327030",
          9614 => x"70962a84",
          9615 => x"80065451",
          9616 => x"55911b51",
          9617 => x"ff8dff3f",
          9618 => x"67557483",
          9619 => x"ffff2690",
          9620 => x"387483ff",
          9621 => x"ff065293",
          9622 => x"1b51ff8d",
          9623 => x"e93f8a39",
          9624 => x"7452a01b",
          9625 => x"51ff8dfc",
          9626 => x"3ff80b95",
          9627 => x"1c34bf52",
          9628 => x"981b51ff",
          9629 => x"8dd03f81",
          9630 => x"ff529a1b",
          9631 => x"51ff8dc6",
          9632 => x"3f7e529c",
          9633 => x"1b51ff8d",
          9634 => x"db3f7d83",
          9635 => x"2e098106",
          9636 => x"80cb3882",
          9637 => x"88b20a52",
          9638 => x"80c31b51",
          9639 => x"ff8dc53f",
          9640 => x"7c52a41b",
          9641 => x"51ff8dbc",
          9642 => x"3f8252ac",
          9643 => x"1b51ff8d",
          9644 => x"b33f8152",
          9645 => x"b01b51ff",
          9646 => x"8d8c3f86",
          9647 => x"52b21b51",
          9648 => x"ff8d833f",
          9649 => x"ff800b80",
          9650 => x"c01c34a9",
          9651 => x"0b80c21c",
          9652 => x"34935382",
          9653 => x"d1f05280",
          9654 => x"c71b51ae",
          9655 => x"398288b2",
          9656 => x"0a52a71b",
          9657 => x"51ff8cfc",
          9658 => x"3f7c83ff",
          9659 => x"ff065296",
          9660 => x"1b51ff8c",
          9661 => x"d13fff80",
          9662 => x"0ba41c34",
          9663 => x"a90ba61c",
          9664 => x"34935382",
          9665 => x"d28452ab",
          9666 => x"1b51ff8d",
          9667 => x"863f82d4",
          9668 => x"d55283fe",
          9669 => x"1b705259",
          9670 => x"ff8cab3f",
          9671 => x"81547e53",
          9672 => x"7a527f51",
          9673 => x"ff88ce3f",
          9674 => x"815682e0",
          9675 => x"9808849c",
          9676 => x"387d832e",
          9677 => x"09810680",
          9678 => x"ec387554",
          9679 => x"861f537a",
          9680 => x"527f51ff",
          9681 => x"88af3f84",
          9682 => x"80538052",
          9683 => x"7a51ff8c",
          9684 => x"e53f848b",
          9685 => x"85a4d252",
          9686 => x"7a51ff8c",
          9687 => x"873f868a",
          9688 => x"85e4f252",
          9689 => x"83e41b51",
          9690 => x"ff8bf93f",
          9691 => x"ff185283",
          9692 => x"e81b51ff",
          9693 => x"8bee3f82",
          9694 => x"5283ec1b",
          9695 => x"51ff8be4",
          9696 => x"3f82d4d5",
          9697 => x"527851ff",
          9698 => x"8bbc3f75",
          9699 => x"54871f53",
          9700 => x"7a527f51",
          9701 => x"ff87de3f",
          9702 => x"7554751f",
          9703 => x"537a527f",
          9704 => x"51ff87d1",
          9705 => x"3f665380",
          9706 => x"527a51ff",
          9707 => x"8c883f60",
          9708 => x"5680587d",
          9709 => x"832e0981",
          9710 => x"069a38f8",
          9711 => x"527a51ff",
          9712 => x"8ba23fff",
          9713 => x"52841b51",
          9714 => x"ff8b993f",
          9715 => x"f00a5288",
          9716 => x"1b519139",
          9717 => x"87fffff8",
          9718 => x"557d812e",
          9719 => x"8338f855",
          9720 => x"74527a51",
          9721 => x"ff8afd3f",
          9722 => x"7c556157",
          9723 => x"74622683",
          9724 => x"38745776",
          9725 => x"5475537a",
          9726 => x"527f51ff",
          9727 => x"86f73f82",
          9728 => x"e0980882",
          9729 => x"be388480",
          9730 => x"5382e098",
          9731 => x"08527a51",
          9732 => x"ff8ba33f",
          9733 => x"76167578",
          9734 => x"31565674",
          9735 => x"cd388118",
          9736 => x"5877802e",
          9737 => x"ff8d3879",
          9738 => x"557d832e",
          9739 => x"83386555",
          9740 => x"61577462",
          9741 => x"26833874",
          9742 => x"57765475",
          9743 => x"537a527f",
          9744 => x"51ff86b1",
          9745 => x"3f82e098",
          9746 => x"0881f838",
          9747 => x"76167578",
          9748 => x"31565674",
          9749 => x"db388c57",
          9750 => x"7d832e93",
          9751 => x"38865767",
          9752 => x"83ffff26",
          9753 => x"8a388457",
          9754 => x"7d822e83",
          9755 => x"38815764",
          9756 => x"802eb238",
          9757 => x"81548053",
          9758 => x"7a527f51",
          9759 => x"ff848c3f",
          9760 => x"815682e0",
          9761 => x"980881c4",
          9762 => x"38649029",
          9763 => x"1b557683",
          9764 => x"b2163475",
          9765 => x"5482e098",
          9766 => x"08537a52",
          9767 => x"7f51ff85",
          9768 => x"d43f8181",
          9769 => x"3962832a",
          9770 => x"81065877",
          9771 => x"80fd3884",
          9772 => x"80537752",
          9773 => x"7a51ff89",
          9774 => x"fd3f82d4",
          9775 => x"d5527851",
          9776 => x"ff89833f",
          9777 => x"83be1b55",
          9778 => x"77753481",
          9779 => x"0b811634",
          9780 => x"810b8216",
          9781 => x"34778316",
          9782 => x"34768416",
          9783 => x"34671f56",
          9784 => x"80fdc152",
          9785 => x"7551fe93",
          9786 => x"ea3ffe0b",
          9787 => x"85163482",
          9788 => x"e0980882",
          9789 => x"2abf0756",
          9790 => x"75861634",
          9791 => x"82e09808",
          9792 => x"8716347e",
          9793 => x"5283c61b",
          9794 => x"51ff88d8",
          9795 => x"3f675283",
          9796 => x"ca1b51ff",
          9797 => x"88ce3f81",
          9798 => x"5477537a",
          9799 => x"527f51ff",
          9800 => x"84d33f81",
          9801 => x"5682e098",
          9802 => x"08a23880",
          9803 => x"5380527f",
          9804 => x"51ff86a5",
          9805 => x"3f815682",
          9806 => x"e0980890",
          9807 => x"3889398e",
          9808 => x"568a3981",
          9809 => x"56863982",
          9810 => x"e0980856",
          9811 => x"7582e098",
          9812 => x"0c9a3d0d",
          9813 => x"04f53d0d",
          9814 => x"7d605b59",
          9815 => x"807960ff",
          9816 => x"055a5757",
          9817 => x"767825b4",
          9818 => x"388d3df8",
          9819 => x"11555581",
          9820 => x"53fc1552",
          9821 => x"7951c894",
          9822 => x"3f7a812e",
          9823 => x"0981069c",
          9824 => x"388c3d33",
          9825 => x"55748d2e",
          9826 => x"db387476",
          9827 => x"70810558",
          9828 => x"34811757",
          9829 => x"748a2e09",
          9830 => x"8106c938",
          9831 => x"80763478",
          9832 => x"55768338",
          9833 => x"76557482",
          9834 => x"e0980c8d",
          9835 => x"3d0d04f7",
          9836 => x"3d0d7b02",
          9837 => x"8405b305",
          9838 => x"33595777",
          9839 => x"8a2e0981",
          9840 => x"0687388d",
          9841 => x"527651e7",
          9842 => x"3f841708",
          9843 => x"56807624",
          9844 => x"be388817",
          9845 => x"0877178c",
          9846 => x"05565977",
          9847 => x"75348116",
          9848 => x"56bb7625",
          9849 => x"a1388b3d",
          9850 => x"fc055475",
          9851 => x"538c1752",
          9852 => x"760851ca",
          9853 => x"973f7976",
          9854 => x"32703070",
          9855 => x"72079f2a",
          9856 => x"70305351",
          9857 => x"56567584",
          9858 => x"180c8119",
          9859 => x"88180c8b",
          9860 => x"3d0d04f9",
          9861 => x"3d0d7984",
          9862 => x"11085656",
          9863 => x"807524a7",
          9864 => x"38893dfc",
          9865 => x"05547453",
          9866 => x"8c165275",
          9867 => x"0851c9dc",
          9868 => x"3f82e098",
          9869 => x"08913884",
          9870 => x"1608782e",
          9871 => x"09810687",
          9872 => x"38881608",
          9873 => x"558339ff",
          9874 => x"557482e0",
          9875 => x"980c893d",
          9876 => x"0d04fd3d",
          9877 => x"0d755480",
          9878 => x"cc538052",
          9879 => x"7351ff86",
          9880 => x"d53f7674",
          9881 => x"0c853d0d",
          9882 => x"04ea3d0d",
          9883 => x"0280e305",
          9884 => x"336a5386",
          9885 => x"3d705354",
          9886 => x"54d83f73",
          9887 => x"527251fe",
          9888 => x"ae3f7251",
          9889 => x"ff8d3f98",
          9890 => x"3d0d04fd",
          9891 => x"3d0d7502",
          9892 => x"84059a05",
          9893 => x"22555380",
          9894 => x"527280ff",
          9895 => x"268a3872",
          9896 => x"83ffff06",
          9897 => x"5280c339",
          9898 => x"83ffff73",
          9899 => x"27517383",
          9900 => x"b52e0981",
          9901 => x"06b43870",
          9902 => x"802eaf38",
          9903 => x"82d3ec22",
          9904 => x"5172712e",
          9905 => x"9c388112",
          9906 => x"7083ffff",
          9907 => x"06535171",
          9908 => x"80ff268d",
          9909 => x"38711082",
          9910 => x"d3ec0570",
          9911 => x"225151e1",
          9912 => x"39818012",
          9913 => x"7081ff06",
          9914 => x"53517182",
          9915 => x"e0980c85",
          9916 => x"3d0d04fe",
          9917 => x"3d0d0292",
          9918 => x"05220284",
          9919 => x"05960522",
          9920 => x"53518053",
          9921 => x"7080ff26",
          9922 => x"85387053",
          9923 => x"9a397183",
          9924 => x"b52e0981",
          9925 => x"06913870",
          9926 => x"81ff268b",
          9927 => x"38701082",
          9928 => x"d1ec0570",
          9929 => x"22545172",
          9930 => x"82e0980c",
          9931 => x"843d0d04",
          9932 => x"fb3d0d77",
          9933 => x"517083ff",
          9934 => x"ff2681a7",
          9935 => x"387083ff",
          9936 => x"ff0682d5",
          9937 => x"ec57529f",
          9938 => x"ff722785",
          9939 => x"3882d9e0",
          9940 => x"56757082",
          9941 => x"05572270",
          9942 => x"30708025",
          9943 => x"72752607",
          9944 => x"51525570",
          9945 => x"80fb3875",
          9946 => x"70820557",
          9947 => x"2270882a",
          9948 => x"7181ff06",
          9949 => x"70185452",
          9950 => x"55537171",
          9951 => x"2580d738",
          9952 => x"73882680",
          9953 => x"dc387384",
          9954 => x"2982b9b8",
          9955 => x"05517008",
          9956 => x"04717531",
          9957 => x"10761170",
          9958 => x"22545151",
          9959 => x"80c33971",
          9960 => x"75318106",
          9961 => x"72713151",
          9962 => x"51a439f0",
          9963 => x"12519f39",
          9964 => x"e012519a",
          9965 => x"39d01251",
          9966 => x"9539e612",
          9967 => x"51903988",
          9968 => x"12518b39",
          9969 => x"ffb01251",
          9970 => x"8539c7a0",
          9971 => x"12517083",
          9972 => x"ffff0652",
          9973 => x"8c3973fe",
          9974 => x"f8387210",
          9975 => x"1656fef1",
          9976 => x"39715170",
          9977 => x"82e0980c",
          9978 => x"873d0d04",
          9979 => x"00ffffff",
          9980 => x"ff00ffff",
          9981 => x"ffff00ff",
          9982 => x"ffffff00",
          9983 => x"00003101",
          9984 => x"00003085",
          9985 => x"0000308c",
          9986 => x"00003093",
          9987 => x"0000309a",
          9988 => x"000030a1",
          9989 => x"000030a8",
          9990 => x"000030af",
          9991 => x"000030b6",
          9992 => x"000030bd",
          9993 => x"000030c4",
          9994 => x"000030cb",
          9995 => x"000030d1",
          9996 => x"000030d7",
          9997 => x"000030dd",
          9998 => x"000030e3",
          9999 => x"000030e9",
         10000 => x"000030ef",
         10001 => x"000030f5",
         10002 => x"000030fb",
         10003 => x"00004781",
         10004 => x"00004787",
         10005 => x"0000478d",
         10006 => x"00004793",
         10007 => x"00004799",
         10008 => x"00004d79",
         10009 => x"00004e79",
         10010 => x"00004f8a",
         10011 => x"000051e2",
         10012 => x"00004e61",
         10013 => x"00004c4c",
         10014 => x"00005052",
         10015 => x"000051b3",
         10016 => x"00005095",
         10017 => x"0000512b",
         10018 => x"000050b1",
         10019 => x"00004f34",
         10020 => x"00004c4c",
         10021 => x"00004f8a",
         10022 => x"00004fb3",
         10023 => x"00005052",
         10024 => x"00004c4c",
         10025 => x"00004c4c",
         10026 => x"000050b1",
         10027 => x"0000512b",
         10028 => x"000051b3",
         10029 => x"000051e2",
         10030 => x"00009b91",
         10031 => x"00009b9f",
         10032 => x"00009bab",
         10033 => x"00009bb0",
         10034 => x"00009bb5",
         10035 => x"00009bba",
         10036 => x"00009bbf",
         10037 => x"00009bc4",
         10038 => x"00009bca",
         10039 => x"00000e65",
         10040 => x"0000174e",
         10041 => x"0000174e",
         10042 => x"00000e94",
         10043 => x"0000174e",
         10044 => x"0000174e",
         10045 => x"0000174e",
         10046 => x"0000174e",
         10047 => x"0000174e",
         10048 => x"0000174e",
         10049 => x"0000174e",
         10050 => x"00000e51",
         10051 => x"0000174e",
         10052 => x"00000e7c",
         10053 => x"00000eac",
         10054 => x"0000174e",
         10055 => x"0000174e",
         10056 => x"0000174e",
         10057 => x"0000174e",
         10058 => x"0000174e",
         10059 => x"0000174e",
         10060 => x"0000174e",
         10061 => x"0000174e",
         10062 => x"0000174e",
         10063 => x"0000174e",
         10064 => x"0000174e",
         10065 => x"0000174e",
         10066 => x"0000174e",
         10067 => x"0000174e",
         10068 => x"0000174e",
         10069 => x"0000174e",
         10070 => x"0000174e",
         10071 => x"0000174e",
         10072 => x"0000174e",
         10073 => x"0000174e",
         10074 => x"0000174e",
         10075 => x"0000174e",
         10076 => x"0000174e",
         10077 => x"0000174e",
         10078 => x"0000174e",
         10079 => x"0000174e",
         10080 => x"0000174e",
         10081 => x"0000174e",
         10082 => x"0000174e",
         10083 => x"0000174e",
         10084 => x"0000174e",
         10085 => x"0000174e",
         10086 => x"0000174e",
         10087 => x"0000174e",
         10088 => x"0000174e",
         10089 => x"0000174e",
         10090 => x"00000fdc",
         10091 => x"0000174e",
         10092 => x"0000174e",
         10093 => x"0000174e",
         10094 => x"0000174e",
         10095 => x"0000114a",
         10096 => x"0000174e",
         10097 => x"0000174e",
         10098 => x"0000174e",
         10099 => x"0000174e",
         10100 => x"0000174e",
         10101 => x"0000174e",
         10102 => x"0000174e",
         10103 => x"0000174e",
         10104 => x"0000174e",
         10105 => x"0000174e",
         10106 => x"00000f0c",
         10107 => x"00001073",
         10108 => x"00000ee3",
         10109 => x"00000ee3",
         10110 => x"00000ee3",
         10111 => x"0000174e",
         10112 => x"00001073",
         10113 => x"0000174e",
         10114 => x"0000174e",
         10115 => x"00000ecc",
         10116 => x"0000174e",
         10117 => x"0000174e",
         10118 => x"00001120",
         10119 => x"0000112b",
         10120 => x"0000174e",
         10121 => x"0000174e",
         10122 => x"00000f45",
         10123 => x"0000174e",
         10124 => x"00001153",
         10125 => x"0000174e",
         10126 => x"0000174e",
         10127 => x"0000114a",
         10128 => x"64696e69",
         10129 => x"74000000",
         10130 => x"64696f63",
         10131 => x"746c0000",
         10132 => x"66696e69",
         10133 => x"74000000",
         10134 => x"666c6f61",
         10135 => x"64000000",
         10136 => x"66657865",
         10137 => x"63000000",
         10138 => x"6d636c65",
         10139 => x"61720000",
         10140 => x"6d636f70",
         10141 => x"79000000",
         10142 => x"6d646966",
         10143 => x"66000000",
         10144 => x"6d64756d",
         10145 => x"70000000",
         10146 => x"6d656200",
         10147 => x"6d656800",
         10148 => x"6d657700",
         10149 => x"68696400",
         10150 => x"68696500",
         10151 => x"68666400",
         10152 => x"68666500",
         10153 => x"63616c6c",
         10154 => x"00000000",
         10155 => x"6a6d7000",
         10156 => x"72657374",
         10157 => x"61727400",
         10158 => x"72657365",
         10159 => x"74000000",
         10160 => x"696e666f",
         10161 => x"00000000",
         10162 => x"74626173",
         10163 => x"69630000",
         10164 => x"6d626173",
         10165 => x"69630000",
         10166 => x"6b696c6f",
         10167 => x"00000000",
         10168 => x"65640000",
         10169 => x"4469736b",
         10170 => x"20457272",
         10171 => x"6f720000",
         10172 => x"496e7465",
         10173 => x"726e616c",
         10174 => x"20657272",
         10175 => x"6f722e00",
         10176 => x"4469736b",
         10177 => x"206e6f74",
         10178 => x"20726561",
         10179 => x"64792e00",
         10180 => x"4e6f2066",
         10181 => x"696c6520",
         10182 => x"666f756e",
         10183 => x"642e0000",
         10184 => x"4e6f2070",
         10185 => x"61746820",
         10186 => x"666f756e",
         10187 => x"642e0000",
         10188 => x"496e7661",
         10189 => x"6c696420",
         10190 => x"66696c65",
         10191 => x"6e616d65",
         10192 => x"2e000000",
         10193 => x"41636365",
         10194 => x"73732064",
         10195 => x"656e6965",
         10196 => x"642e0000",
         10197 => x"46696c65",
         10198 => x"20616c72",
         10199 => x"65616479",
         10200 => x"20657869",
         10201 => x"7374732e",
         10202 => x"00000000",
         10203 => x"46696c65",
         10204 => x"2068616e",
         10205 => x"646c6520",
         10206 => x"696e7661",
         10207 => x"6c69642e",
         10208 => x"00000000",
         10209 => x"53442069",
         10210 => x"73207772",
         10211 => x"69746520",
         10212 => x"70726f74",
         10213 => x"65637465",
         10214 => x"642e0000",
         10215 => x"44726976",
         10216 => x"65206e75",
         10217 => x"6d626572",
         10218 => x"20697320",
         10219 => x"696e7661",
         10220 => x"6c69642e",
         10221 => x"00000000",
         10222 => x"4469736b",
         10223 => x"206e6f74",
         10224 => x"20656e61",
         10225 => x"626c6564",
         10226 => x"2e000000",
         10227 => x"4e6f2063",
         10228 => x"6f6d7061",
         10229 => x"7469626c",
         10230 => x"65206669",
         10231 => x"6c657379",
         10232 => x"7374656d",
         10233 => x"20666f75",
         10234 => x"6e64206f",
         10235 => x"6e206469",
         10236 => x"736b2e00",
         10237 => x"466f726d",
         10238 => x"61742061",
         10239 => x"626f7274",
         10240 => x"65642e00",
         10241 => x"54696d65",
         10242 => x"6f75742c",
         10243 => x"206f7065",
         10244 => x"72617469",
         10245 => x"6f6e2063",
         10246 => x"616e6365",
         10247 => x"6c6c6564",
         10248 => x"2e000000",
         10249 => x"46696c65",
         10250 => x"20697320",
         10251 => x"6c6f636b",
         10252 => x"65642e00",
         10253 => x"496e7375",
         10254 => x"66666963",
         10255 => x"69656e74",
         10256 => x"206d656d",
         10257 => x"6f72792e",
         10258 => x"00000000",
         10259 => x"546f6f20",
         10260 => x"6d616e79",
         10261 => x"206f7065",
         10262 => x"6e206669",
         10263 => x"6c65732e",
         10264 => x"00000000",
         10265 => x"50617261",
         10266 => x"6d657465",
         10267 => x"72732069",
         10268 => x"6e636f72",
         10269 => x"72656374",
         10270 => x"2e000000",
         10271 => x"53756363",
         10272 => x"6573732e",
         10273 => x"00000000",
         10274 => x"556e6b6e",
         10275 => x"6f776e20",
         10276 => x"6572726f",
         10277 => x"722e0000",
         10278 => x"0a256c75",
         10279 => x"20627974",
         10280 => x"65732025",
         10281 => x"73206174",
         10282 => x"20256c75",
         10283 => x"20627974",
         10284 => x"65732f73",
         10285 => x"65632e0a",
         10286 => x"00000000",
         10287 => x"72656164",
         10288 => x"00000000",
         10289 => x"2530386c",
         10290 => x"58000000",
         10291 => x"3a202000",
         10292 => x"25303458",
         10293 => x"00000000",
         10294 => x"20202020",
         10295 => x"20202020",
         10296 => x"00000000",
         10297 => x"25303258",
         10298 => x"00000000",
         10299 => x"20200000",
         10300 => x"207c0000",
         10301 => x"7c000000",
         10302 => x"7a4f5300",
         10303 => x"2a2a2025",
         10304 => x"73202800",
         10305 => x"31312f31",
         10306 => x"322f3230",
         10307 => x"32300000",
         10308 => x"76312e31",
         10309 => x"63000000",
         10310 => x"205a5055",
         10311 => x"2c207265",
         10312 => x"76202530",
         10313 => x"32782920",
         10314 => x"25732025",
         10315 => x"73202a2a",
         10316 => x"0a0a0000",
         10317 => x"5a505520",
         10318 => x"496e7465",
         10319 => x"72727570",
         10320 => x"74204861",
         10321 => x"6e646c65",
         10322 => x"72000000",
         10323 => x"54696d65",
         10324 => x"7220696e",
         10325 => x"74657272",
         10326 => x"75707400",
         10327 => x"50533220",
         10328 => x"696e7465",
         10329 => x"72727570",
         10330 => x"74000000",
         10331 => x"494f4354",
         10332 => x"4c205244",
         10333 => x"20696e74",
         10334 => x"65727275",
         10335 => x"70740000",
         10336 => x"494f4354",
         10337 => x"4c205752",
         10338 => x"20696e74",
         10339 => x"65727275",
         10340 => x"70740000",
         10341 => x"55415254",
         10342 => x"30205258",
         10343 => x"20696e74",
         10344 => x"65727275",
         10345 => x"70740000",
         10346 => x"55415254",
         10347 => x"30205458",
         10348 => x"20696e74",
         10349 => x"65727275",
         10350 => x"70740000",
         10351 => x"55415254",
         10352 => x"31205258",
         10353 => x"20696e74",
         10354 => x"65727275",
         10355 => x"70740000",
         10356 => x"55415254",
         10357 => x"31205458",
         10358 => x"20696e74",
         10359 => x"65727275",
         10360 => x"70740000",
         10361 => x"53657474",
         10362 => x"696e6720",
         10363 => x"75702074",
         10364 => x"696d6572",
         10365 => x"2e2e2e00",
         10366 => x"456e6162",
         10367 => x"6c696e67",
         10368 => x"2074696d",
         10369 => x"65722e2e",
         10370 => x"2e000000",
         10371 => x"6175746f",
         10372 => x"65786563",
         10373 => x"2e626174",
         10374 => x"00000000",
         10375 => x"7a4f535f",
         10376 => x"7a70752e",
         10377 => x"68737400",
         10378 => x"303a0000",
         10379 => x"4661696c",
         10380 => x"65642074",
         10381 => x"6f20696e",
         10382 => x"69746961",
         10383 => x"6c697365",
         10384 => x"20736420",
         10385 => x"63617264",
         10386 => x"20302c20",
         10387 => x"706c6561",
         10388 => x"73652069",
         10389 => x"6e697420",
         10390 => x"6d616e75",
         10391 => x"616c6c79",
         10392 => x"2e000000",
         10393 => x"2a200000",
         10394 => x"436c6561",
         10395 => x"72696e67",
         10396 => x"2e2e2e2e",
         10397 => x"00000000",
         10398 => x"436f7079",
         10399 => x"696e672e",
         10400 => x"2e2e0000",
         10401 => x"436f6d70",
         10402 => x"6172696e",
         10403 => x"672e2e2e",
         10404 => x"00000000",
         10405 => x"2530386c",
         10406 => x"78282530",
         10407 => x"3878292d",
         10408 => x"3e253038",
         10409 => x"6c782825",
         10410 => x"30387829",
         10411 => x"0a000000",
         10412 => x"44756d70",
         10413 => x"204d656d",
         10414 => x"6f727900",
         10415 => x"0a436f6d",
         10416 => x"706c6574",
         10417 => x"652e0000",
         10418 => x"2530386c",
         10419 => x"58202530",
         10420 => x"32582d00",
         10421 => x"3f3f3f00",
         10422 => x"2530386c",
         10423 => x"58202530",
         10424 => x"34582d00",
         10425 => x"2530386c",
         10426 => x"58202530",
         10427 => x"386c582d",
         10428 => x"00000000",
         10429 => x"45786563",
         10430 => x"7574696e",
         10431 => x"6720636f",
         10432 => x"64652040",
         10433 => x"20253038",
         10434 => x"6c78202e",
         10435 => x"2e2e0a00",
         10436 => x"43616c6c",
         10437 => x"696e6720",
         10438 => x"636f6465",
         10439 => x"20402025",
         10440 => x"30386c78",
         10441 => x"202e2e2e",
         10442 => x"0a000000",
         10443 => x"43616c6c",
         10444 => x"20726574",
         10445 => x"75726e65",
         10446 => x"6420636f",
         10447 => x"64652028",
         10448 => x"2564292e",
         10449 => x"0a000000",
         10450 => x"52657374",
         10451 => x"61727469",
         10452 => x"6e672061",
         10453 => x"70706c69",
         10454 => x"63617469",
         10455 => x"6f6e2e2e",
         10456 => x"2e000000",
         10457 => x"436f6c64",
         10458 => x"20726562",
         10459 => x"6f6f7469",
         10460 => x"6e672e2e",
         10461 => x"2e000000",
         10462 => x"5a505500",
         10463 => x"62696e00",
         10464 => x"25643a5c",
         10465 => x"25735c25",
         10466 => x"732e2573",
         10467 => x"00000000",
         10468 => x"25643a5c",
         10469 => x"25735c25",
         10470 => x"73000000",
         10471 => x"25643a5c",
         10472 => x"25730000",
         10473 => x"42616420",
         10474 => x"636f6d6d",
         10475 => x"616e642e",
         10476 => x"00000000",
         10477 => x"4d656d6f",
         10478 => x"72792065",
         10479 => x"78686175",
         10480 => x"73746564",
         10481 => x"2c206361",
         10482 => x"6e6e6f74",
         10483 => x"2070726f",
         10484 => x"63657373",
         10485 => x"20636f6d",
         10486 => x"6d616e64",
         10487 => x"2e000000",
         10488 => x"52756e6e",
         10489 => x"696e672e",
         10490 => x"2e2e0000",
         10491 => x"456e6162",
         10492 => x"6c696e67",
         10493 => x"20696e74",
         10494 => x"65727275",
         10495 => x"7074732e",
         10496 => x"2e2e0000",
         10497 => x"25642f25",
         10498 => x"642f2564",
         10499 => x"2025643a",
         10500 => x"25643a25",
         10501 => x"642e2564",
         10502 => x"25640a00",
         10503 => x"536f4320",
         10504 => x"436f6e66",
         10505 => x"69677572",
         10506 => x"6174696f",
         10507 => x"6e000000",
         10508 => x"20286672",
         10509 => x"6f6d2053",
         10510 => x"6f432063",
         10511 => x"6f6e6669",
         10512 => x"67290000",
         10513 => x"3a0a4465",
         10514 => x"76696365",
         10515 => x"7320696d",
         10516 => x"706c656d",
         10517 => x"656e7465",
         10518 => x"643a0000",
         10519 => x"20202020",
         10520 => x"57422053",
         10521 => x"4452414d",
         10522 => x"20202825",
         10523 => x"3038583a",
         10524 => x"25303858",
         10525 => x"292e0a00",
         10526 => x"20202020",
         10527 => x"53445241",
         10528 => x"4d202020",
         10529 => x"20202825",
         10530 => x"3038583a",
         10531 => x"25303858",
         10532 => x"292e0a00",
         10533 => x"20202020",
         10534 => x"494e534e",
         10535 => x"20425241",
         10536 => x"4d202825",
         10537 => x"3038583a",
         10538 => x"25303858",
         10539 => x"292e0a00",
         10540 => x"20202020",
         10541 => x"4252414d",
         10542 => x"20202020",
         10543 => x"20202825",
         10544 => x"3038583a",
         10545 => x"25303858",
         10546 => x"292e0a00",
         10547 => x"20202020",
         10548 => x"52414d20",
         10549 => x"20202020",
         10550 => x"20202825",
         10551 => x"3038583a",
         10552 => x"25303858",
         10553 => x"292e0a00",
         10554 => x"20202020",
         10555 => x"53442043",
         10556 => x"41524420",
         10557 => x"20202844",
         10558 => x"65766963",
         10559 => x"6573203d",
         10560 => x"25303264",
         10561 => x"292e0a00",
         10562 => x"20202020",
         10563 => x"54494d45",
         10564 => x"52312020",
         10565 => x"20202854",
         10566 => x"696d6572",
         10567 => x"7320203d",
         10568 => x"25303264",
         10569 => x"292e0a00",
         10570 => x"20202020",
         10571 => x"494e5452",
         10572 => x"20435452",
         10573 => x"4c202843",
         10574 => x"68616e6e",
         10575 => x"656c733d",
         10576 => x"25303264",
         10577 => x"292e0a00",
         10578 => x"20202020",
         10579 => x"57495348",
         10580 => x"424f4e45",
         10581 => x"20425553",
         10582 => x"00000000",
         10583 => x"20202020",
         10584 => x"57422049",
         10585 => x"32430000",
         10586 => x"20202020",
         10587 => x"494f4354",
         10588 => x"4c000000",
         10589 => x"20202020",
         10590 => x"50533200",
         10591 => x"20202020",
         10592 => x"53504900",
         10593 => x"41646472",
         10594 => x"65737365",
         10595 => x"733a0000",
         10596 => x"20202020",
         10597 => x"43505520",
         10598 => x"52657365",
         10599 => x"74205665",
         10600 => x"63746f72",
         10601 => x"20416464",
         10602 => x"72657373",
         10603 => x"203d2025",
         10604 => x"3038580a",
         10605 => x"00000000",
         10606 => x"20202020",
         10607 => x"43505520",
         10608 => x"4d656d6f",
         10609 => x"72792053",
         10610 => x"74617274",
         10611 => x"20416464",
         10612 => x"72657373",
         10613 => x"203d2025",
         10614 => x"3038580a",
         10615 => x"00000000",
         10616 => x"20202020",
         10617 => x"53746163",
         10618 => x"6b205374",
         10619 => x"61727420",
         10620 => x"41646472",
         10621 => x"65737320",
         10622 => x"20202020",
         10623 => x"203d2025",
         10624 => x"3038580a",
         10625 => x"00000000",
         10626 => x"4d697363",
         10627 => x"3a000000",
         10628 => x"20202020",
         10629 => x"5a505520",
         10630 => x"49642020",
         10631 => x"20202020",
         10632 => x"20202020",
         10633 => x"20202020",
         10634 => x"20202020",
         10635 => x"203d2025",
         10636 => x"3034580a",
         10637 => x"00000000",
         10638 => x"20202020",
         10639 => x"53797374",
         10640 => x"656d2043",
         10641 => x"6c6f636b",
         10642 => x"20467265",
         10643 => x"71202020",
         10644 => x"20202020",
         10645 => x"203d2025",
         10646 => x"642e2530",
         10647 => x"34644d48",
         10648 => x"7a0a0000",
         10649 => x"20202020",
         10650 => x"53445241",
         10651 => x"4d20436c",
         10652 => x"6f636b20",
         10653 => x"46726571",
         10654 => x"20202020",
         10655 => x"20202020",
         10656 => x"203d2025",
         10657 => x"642e2530",
         10658 => x"34644d48",
         10659 => x"7a0a0000",
         10660 => x"20202020",
         10661 => x"57697368",
         10662 => x"626f6e65",
         10663 => x"20534452",
         10664 => x"414d2043",
         10665 => x"6c6f636b",
         10666 => x"20467265",
         10667 => x"713d2025",
         10668 => x"642e2530",
         10669 => x"34644d48",
         10670 => x"7a0a0000",
         10671 => x"536d616c",
         10672 => x"6c000000",
         10673 => x"4d656469",
         10674 => x"756d0000",
         10675 => x"466c6578",
         10676 => x"00000000",
         10677 => x"45564f00",
         10678 => x"45564f6d",
         10679 => x"00000000",
         10680 => x"556e6b6e",
         10681 => x"6f776e00",
         10682 => x"0000a844",
         10683 => x"01000000",
         10684 => x"00000002",
         10685 => x"0000a840",
         10686 => x"01000000",
         10687 => x"00000003",
         10688 => x"0000a83c",
         10689 => x"01000000",
         10690 => x"00000004",
         10691 => x"0000a838",
         10692 => x"01000000",
         10693 => x"00000005",
         10694 => x"0000a834",
         10695 => x"01000000",
         10696 => x"00000006",
         10697 => x"0000a830",
         10698 => x"01000000",
         10699 => x"00000007",
         10700 => x"0000a82c",
         10701 => x"01000000",
         10702 => x"00000001",
         10703 => x"0000a828",
         10704 => x"01000000",
         10705 => x"00000008",
         10706 => x"0000a824",
         10707 => x"01000000",
         10708 => x"0000000b",
         10709 => x"0000a820",
         10710 => x"01000000",
         10711 => x"00000009",
         10712 => x"0000a81c",
         10713 => x"01000000",
         10714 => x"0000000a",
         10715 => x"0000a818",
         10716 => x"04000000",
         10717 => x"0000000d",
         10718 => x"0000a814",
         10719 => x"04000000",
         10720 => x"0000000c",
         10721 => x"0000a810",
         10722 => x"04000000",
         10723 => x"0000000e",
         10724 => x"0000a80c",
         10725 => x"03000000",
         10726 => x"0000000f",
         10727 => x"0000a808",
         10728 => x"04000000",
         10729 => x"0000000f",
         10730 => x"0000a804",
         10731 => x"04000000",
         10732 => x"00000010",
         10733 => x"0000a800",
         10734 => x"04000000",
         10735 => x"00000011",
         10736 => x"0000a7fc",
         10737 => x"03000000",
         10738 => x"00000012",
         10739 => x"0000a7f8",
         10740 => x"03000000",
         10741 => x"00000013",
         10742 => x"0000a7f4",
         10743 => x"03000000",
         10744 => x"00000014",
         10745 => x"0000a7f0",
         10746 => x"03000000",
         10747 => x"00000015",
         10748 => x"1b5b4400",
         10749 => x"1b5b4300",
         10750 => x"1b5b4200",
         10751 => x"1b5b4100",
         10752 => x"1b5b367e",
         10753 => x"1b5b357e",
         10754 => x"1b5b347e",
         10755 => x"1b304600",
         10756 => x"1b5b337e",
         10757 => x"1b5b327e",
         10758 => x"1b5b317e",
         10759 => x"10000000",
         10760 => x"0e000000",
         10761 => x"0d000000",
         10762 => x"0b000000",
         10763 => x"08000000",
         10764 => x"06000000",
         10765 => x"05000000",
         10766 => x"04000000",
         10767 => x"03000000",
         10768 => x"02000000",
         10769 => x"01000000",
         10770 => x"68697374",
         10771 => x"6f727900",
         10772 => x"68697374",
         10773 => x"00000000",
         10774 => x"21000000",
         10775 => x"2530346c",
         10776 => x"75202025",
         10777 => x"730a0000",
         10778 => x"4661696c",
         10779 => x"65642074",
         10780 => x"6f207265",
         10781 => x"73657420",
         10782 => x"74686520",
         10783 => x"68697374",
         10784 => x"6f727920",
         10785 => x"66696c65",
         10786 => x"20746f20",
         10787 => x"454f462e",
         10788 => x"00000000",
         10789 => x"43616e6e",
         10790 => x"6f74206f",
         10791 => x"70656e2f",
         10792 => x"63726561",
         10793 => x"74652068",
         10794 => x"6973746f",
         10795 => x"72792066",
         10796 => x"696c652c",
         10797 => x"20646973",
         10798 => x"61626c69",
         10799 => x"6e672e00",
         10800 => x"53440000",
         10801 => x"222a3a3c",
         10802 => x"3e3f7c7f",
         10803 => x"00000000",
         10804 => x"2b2c3b3d",
         10805 => x"5b5d0000",
         10806 => x"46415400",
         10807 => x"46415433",
         10808 => x"32000000",
         10809 => x"ebfe904d",
         10810 => x"53444f53",
         10811 => x"352e3000",
         10812 => x"4e4f204e",
         10813 => x"414d4520",
         10814 => x"20202046",
         10815 => x"41543332",
         10816 => x"20202000",
         10817 => x"4e4f204e",
         10818 => x"414d4520",
         10819 => x"20202046",
         10820 => x"41542020",
         10821 => x"20202000",
         10822 => x"0000a8c0",
         10823 => x"00000000",
         10824 => x"00000000",
         10825 => x"00000000",
         10826 => x"01030507",
         10827 => x"090e1012",
         10828 => x"1416181c",
         10829 => x"1e000000",
         10830 => x"809a4541",
         10831 => x"8e418f80",
         10832 => x"45454549",
         10833 => x"49498e8f",
         10834 => x"9092924f",
         10835 => x"994f5555",
         10836 => x"59999a9b",
         10837 => x"9c9d9e9f",
         10838 => x"41494f55",
         10839 => x"a5a5a6a7",
         10840 => x"a8a9aaab",
         10841 => x"acadaeaf",
         10842 => x"b0b1b2b3",
         10843 => x"b4b5b6b7",
         10844 => x"b8b9babb",
         10845 => x"bcbdbebf",
         10846 => x"c0c1c2c3",
         10847 => x"c4c5c6c7",
         10848 => x"c8c9cacb",
         10849 => x"cccdcecf",
         10850 => x"d0d1d2d3",
         10851 => x"d4d5d6d7",
         10852 => x"d8d9dadb",
         10853 => x"dcdddedf",
         10854 => x"e0e1e2e3",
         10855 => x"e4e5e6e7",
         10856 => x"e8e9eaeb",
         10857 => x"ecedeeef",
         10858 => x"f0f1f2f3",
         10859 => x"f4f5f6f7",
         10860 => x"f8f9fafb",
         10861 => x"fcfdfeff",
         10862 => x"2b2e2c3b",
         10863 => x"3d5b5d2f",
         10864 => x"5c222a3a",
         10865 => x"3c3e3f7c",
         10866 => x"7f000000",
         10867 => x"00010004",
         10868 => x"00100040",
         10869 => x"01000200",
         10870 => x"00000000",
         10871 => x"00010002",
         10872 => x"00040008",
         10873 => x"00100020",
         10874 => x"00000000",
         10875 => x"00c700fc",
         10876 => x"00e900e2",
         10877 => x"00e400e0",
         10878 => x"00e500e7",
         10879 => x"00ea00eb",
         10880 => x"00e800ef",
         10881 => x"00ee00ec",
         10882 => x"00c400c5",
         10883 => x"00c900e6",
         10884 => x"00c600f4",
         10885 => x"00f600f2",
         10886 => x"00fb00f9",
         10887 => x"00ff00d6",
         10888 => x"00dc00a2",
         10889 => x"00a300a5",
         10890 => x"20a70192",
         10891 => x"00e100ed",
         10892 => x"00f300fa",
         10893 => x"00f100d1",
         10894 => x"00aa00ba",
         10895 => x"00bf2310",
         10896 => x"00ac00bd",
         10897 => x"00bc00a1",
         10898 => x"00ab00bb",
         10899 => x"25912592",
         10900 => x"25932502",
         10901 => x"25242561",
         10902 => x"25622556",
         10903 => x"25552563",
         10904 => x"25512557",
         10905 => x"255d255c",
         10906 => x"255b2510",
         10907 => x"25142534",
         10908 => x"252c251c",
         10909 => x"2500253c",
         10910 => x"255e255f",
         10911 => x"255a2554",
         10912 => x"25692566",
         10913 => x"25602550",
         10914 => x"256c2567",
         10915 => x"25682564",
         10916 => x"25652559",
         10917 => x"25582552",
         10918 => x"2553256b",
         10919 => x"256a2518",
         10920 => x"250c2588",
         10921 => x"2584258c",
         10922 => x"25902580",
         10923 => x"03b100df",
         10924 => x"039303c0",
         10925 => x"03a303c3",
         10926 => x"00b503c4",
         10927 => x"03a60398",
         10928 => x"03a903b4",
         10929 => x"221e03c6",
         10930 => x"03b52229",
         10931 => x"226100b1",
         10932 => x"22652264",
         10933 => x"23202321",
         10934 => x"00f72248",
         10935 => x"00b02219",
         10936 => x"00b7221a",
         10937 => x"207f00b2",
         10938 => x"25a000a0",
         10939 => x"0061031a",
         10940 => x"00e00317",
         10941 => x"00f80307",
         10942 => x"00ff0001",
         10943 => x"01780100",
         10944 => x"01300132",
         10945 => x"01060139",
         10946 => x"0110014a",
         10947 => x"012e0179",
         10948 => x"01060180",
         10949 => x"004d0243",
         10950 => x"01810182",
         10951 => x"01820184",
         10952 => x"01840186",
         10953 => x"01870187",
         10954 => x"0189018a",
         10955 => x"018b018b",
         10956 => x"018d018e",
         10957 => x"018f0190",
         10958 => x"01910191",
         10959 => x"01930194",
         10960 => x"01f60196",
         10961 => x"01970198",
         10962 => x"0198023d",
         10963 => x"019b019c",
         10964 => x"019d0220",
         10965 => x"019f01a0",
         10966 => x"01a001a2",
         10967 => x"01a201a4",
         10968 => x"01a401a6",
         10969 => x"01a701a7",
         10970 => x"01a901aa",
         10971 => x"01ab01ac",
         10972 => x"01ac01ae",
         10973 => x"01af01af",
         10974 => x"01b101b2",
         10975 => x"01b301b3",
         10976 => x"01b501b5",
         10977 => x"01b701b8",
         10978 => x"01b801ba",
         10979 => x"01bb01bc",
         10980 => x"01bc01be",
         10981 => x"01f701c0",
         10982 => x"01c101c2",
         10983 => x"01c301c4",
         10984 => x"01c501c4",
         10985 => x"01c701c8",
         10986 => x"01c701ca",
         10987 => x"01cb01ca",
         10988 => x"01cd0110",
         10989 => x"01dd0001",
         10990 => x"018e01de",
         10991 => x"011201f3",
         10992 => x"000301f1",
         10993 => x"01f401f4",
         10994 => x"01f80128",
         10995 => x"02220112",
         10996 => x"023a0009",
         10997 => x"2c65023b",
         10998 => x"023b023d",
         10999 => x"2c66023f",
         11000 => x"02400241",
         11001 => x"02410246",
         11002 => x"010a0253",
         11003 => x"00400181",
         11004 => x"01860255",
         11005 => x"0189018a",
         11006 => x"0258018f",
         11007 => x"025a0190",
         11008 => x"025c025d",
         11009 => x"025e025f",
         11010 => x"01930261",
         11011 => x"02620194",
         11012 => x"02640265",
         11013 => x"02660267",
         11014 => x"01970196",
         11015 => x"026a2c62",
         11016 => x"026c026d",
         11017 => x"026e019c",
         11018 => x"02700271",
         11019 => x"019d0273",
         11020 => x"0274019f",
         11021 => x"02760277",
         11022 => x"02780279",
         11023 => x"027a027b",
         11024 => x"027c2c64",
         11025 => x"027e027f",
         11026 => x"01a60281",
         11027 => x"028201a9",
         11028 => x"02840285",
         11029 => x"02860287",
         11030 => x"01ae0244",
         11031 => x"01b101b2",
         11032 => x"0245028d",
         11033 => x"028e028f",
         11034 => x"02900291",
         11035 => x"01b7037b",
         11036 => x"000303fd",
         11037 => x"03fe03ff",
         11038 => x"03ac0004",
         11039 => x"03860388",
         11040 => x"0389038a",
         11041 => x"03b10311",
         11042 => x"03c20002",
         11043 => x"03a303a3",
         11044 => x"03c40308",
         11045 => x"03cc0003",
         11046 => x"038c038e",
         11047 => x"038f03d8",
         11048 => x"011803f2",
         11049 => x"000a03f9",
         11050 => x"03f303f4",
         11051 => x"03f503f6",
         11052 => x"03f703f7",
         11053 => x"03f903fa",
         11054 => x"03fa0430",
         11055 => x"03200450",
         11056 => x"07100460",
         11057 => x"0122048a",
         11058 => x"013604c1",
         11059 => x"010e04cf",
         11060 => x"000104c0",
         11061 => x"04d00144",
         11062 => x"05610426",
         11063 => x"00000000",
         11064 => x"1d7d0001",
         11065 => x"2c631e00",
         11066 => x"01961ea0",
         11067 => x"015a1f00",
         11068 => x"06081f10",
         11069 => x"06061f20",
         11070 => x"06081f30",
         11071 => x"06081f40",
         11072 => x"06061f51",
         11073 => x"00071f59",
         11074 => x"1f521f5b",
         11075 => x"1f541f5d",
         11076 => x"1f561f5f",
         11077 => x"1f600608",
         11078 => x"1f70000e",
         11079 => x"1fba1fbb",
         11080 => x"1fc81fc9",
         11081 => x"1fca1fcb",
         11082 => x"1fda1fdb",
         11083 => x"1ff81ff9",
         11084 => x"1fea1feb",
         11085 => x"1ffa1ffb",
         11086 => x"1f800608",
         11087 => x"1f900608",
         11088 => x"1fa00608",
         11089 => x"1fb00004",
         11090 => x"1fb81fb9",
         11091 => x"1fb21fbc",
         11092 => x"1fcc0001",
         11093 => x"1fc31fd0",
         11094 => x"06021fe0",
         11095 => x"06021fe5",
         11096 => x"00011fec",
         11097 => x"1ff30001",
         11098 => x"1ffc214e",
         11099 => x"00012132",
         11100 => x"21700210",
         11101 => x"21840001",
         11102 => x"218324d0",
         11103 => x"051a2c30",
         11104 => x"042f2c60",
         11105 => x"01022c67",
         11106 => x"01062c75",
         11107 => x"01022c80",
         11108 => x"01642d00",
         11109 => x"0826ff41",
         11110 => x"031a0000",
         11111 => x"00000000",
         11112 => x"00009e40",
         11113 => x"01020100",
         11114 => x"00000000",
         11115 => x"00000000",
         11116 => x"00009e48",
         11117 => x"01040100",
         11118 => x"00000000",
         11119 => x"00000000",
         11120 => x"00009e50",
         11121 => x"01140300",
         11122 => x"00000000",
         11123 => x"00000000",
         11124 => x"00009e58",
         11125 => x"012b0300",
         11126 => x"00000000",
         11127 => x"00000000",
         11128 => x"00009e60",
         11129 => x"01300300",
         11130 => x"00000000",
         11131 => x"00000000",
         11132 => x"00009e68",
         11133 => x"013c0400",
         11134 => x"00000000",
         11135 => x"00000000",
         11136 => x"00009e70",
         11137 => x"013d0400",
         11138 => x"00000000",
         11139 => x"00000000",
         11140 => x"00009e78",
         11141 => x"013f0400",
         11142 => x"00000000",
         11143 => x"00000000",
         11144 => x"00009e80",
         11145 => x"01400400",
         11146 => x"00000000",
         11147 => x"00000000",
         11148 => x"00009e88",
         11149 => x"01410400",
         11150 => x"00000000",
         11151 => x"00000000",
         11152 => x"00009e8c",
         11153 => x"01420400",
         11154 => x"00000000",
         11155 => x"00000000",
         11156 => x"00009e90",
         11157 => x"01430400",
         11158 => x"00000000",
         11159 => x"00000000",
         11160 => x"00009e94",
         11161 => x"01500500",
         11162 => x"00000000",
         11163 => x"00000000",
         11164 => x"00009e98",
         11165 => x"01510500",
         11166 => x"00000000",
         11167 => x"00000000",
         11168 => x"00009e9c",
         11169 => x"01540500",
         11170 => x"00000000",
         11171 => x"00000000",
         11172 => x"00009ea0",
         11173 => x"01550500",
         11174 => x"00000000",
         11175 => x"00000000",
         11176 => x"00009ea4",
         11177 => x"01790700",
         11178 => x"00000000",
         11179 => x"00000000",
         11180 => x"00009eac",
         11181 => x"01780700",
         11182 => x"00000000",
         11183 => x"00000000",
         11184 => x"00009eb0",
         11185 => x"01820800",
         11186 => x"00000000",
         11187 => x"00000000",
         11188 => x"00009eb8",
         11189 => x"01830800",
         11190 => x"00000000",
         11191 => x"00000000",
         11192 => x"00009ec0",
         11193 => x"01850800",
         11194 => x"00000000",
         11195 => x"00000000",
         11196 => x"00009ec8",
         11197 => x"018c0900",
         11198 => x"00000000",
         11199 => x"00000000",
         11200 => x"00009ed0",
         11201 => x"018d0900",
         11202 => x"00000000",
         11203 => x"00000000",
         11204 => x"00009ed8",
         11205 => x"018e0900",
         11206 => x"00000000",
         11207 => x"00000000",
         11208 => x"00009ee0",
         11209 => x"018f0900",
         11210 => x"00000000",
         11211 => x"00000000",
         11212 => x"00000000",
         11213 => x"00000000",
         11214 => x"00007fff",
         11215 => x"00000000",
         11216 => x"00007fff",
         11217 => x"00010000",
         11218 => x"00007fff",
         11219 => x"00010000",
         11220 => x"00810000",
         11221 => x"01000000",
         11222 => x"017fffff",
         11223 => x"00000000",
         11224 => x"00000000",
         11225 => x"00007800",
         11226 => x"00000000",
         11227 => x"05f5e100",
         11228 => x"05f5e100",
         11229 => x"05f5e100",
         11230 => x"00000000",
         11231 => x"01010101",
         11232 => x"01010101",
         11233 => x"01011001",
         11234 => x"01000000",
         11235 => x"00000000",
         11236 => x"00000000",
         11237 => x"00000000",
         11238 => x"00000000",
         11239 => x"00000000",
         11240 => x"00000000",
         11241 => x"00000000",
         11242 => x"00000000",
         11243 => x"00000000",
         11244 => x"00000000",
         11245 => x"00000000",
         11246 => x"00000000",
         11247 => x"00000000",
         11248 => x"00000000",
         11249 => x"00000000",
         11250 => x"00000000",
         11251 => x"00000000",
         11252 => x"00000000",
         11253 => x"00000000",
         11254 => x"00000000",
         11255 => x"00000000",
         11256 => x"00000000",
         11257 => x"00000000",
         11258 => x"00000000",
         11259 => x"0000a848",
         11260 => x"01000000",
         11261 => x"0000a850",
         11262 => x"01000000",
         11263 => x"0000a858",
         11264 => x"02000000",
         11265 => x"00000000",
         11266 => x"00000000",
         11267 => x"00010002",
         11268 => x"00030004",
         11269 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

