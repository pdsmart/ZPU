-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e9040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"cc738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8a",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"80040088",
           281 => x"e2040000",
           282 => x"009ff070",
           283 => x"a0a0278b",
           284 => x"38807170",
           285 => x"8405530c",
           286 => x"88eb0488",
           287 => x"e2519e99",
           288 => x"04940802",
           289 => x"940cfd3d",
           290 => x"0d805394",
           291 => x"088c0508",
           292 => x"52940888",
           293 => x"05085182",
           294 => x"de3f8808",
           295 => x"70880c54",
           296 => x"853d0d94",
           297 => x"0c049408",
           298 => x"02940cfd",
           299 => x"3d0d8153",
           300 => x"94088c05",
           301 => x"08529408",
           302 => x"88050851",
           303 => x"82b93f88",
           304 => x"0870880c",
           305 => x"54853d0d",
           306 => x"940c0494",
           307 => x"0802940c",
           308 => x"f93d0d80",
           309 => x"0b9408fc",
           310 => x"050c9408",
           311 => x"88050880",
           312 => x"25ab3894",
           313 => x"08880508",
           314 => x"30940888",
           315 => x"050c800b",
           316 => x"9408f405",
           317 => x"0c9408fc",
           318 => x"05088838",
           319 => x"810b9408",
           320 => x"f4050c94",
           321 => x"08f40508",
           322 => x"9408fc05",
           323 => x"0c94088c",
           324 => x"05088025",
           325 => x"ab389408",
           326 => x"8c050830",
           327 => x"94088c05",
           328 => x"0c800b94",
           329 => x"08f0050c",
           330 => x"9408fc05",
           331 => x"08883881",
           332 => x"0b9408f0",
           333 => x"050c9408",
           334 => x"f0050894",
           335 => x"08fc050c",
           336 => x"80539408",
           337 => x"8c050852",
           338 => x"94088805",
           339 => x"085181a7",
           340 => x"3f880870",
           341 => x"9408f805",
           342 => x"0c549408",
           343 => x"fc050880",
           344 => x"2e8c3894",
           345 => x"08f80508",
           346 => x"309408f8",
           347 => x"050c9408",
           348 => x"f8050870",
           349 => x"880c5489",
           350 => x"3d0d940c",
           351 => x"04940802",
           352 => x"940cfb3d",
           353 => x"0d800b94",
           354 => x"08fc050c",
           355 => x"94088805",
           356 => x"08802593",
           357 => x"38940888",
           358 => x"05083094",
           359 => x"0888050c",
           360 => x"810b9408",
           361 => x"fc050c94",
           362 => x"088c0508",
           363 => x"80258c38",
           364 => x"94088c05",
           365 => x"08309408",
           366 => x"8c050c81",
           367 => x"5394088c",
           368 => x"05085294",
           369 => x"08880508",
           370 => x"51ad3f88",
           371 => x"08709408",
           372 => x"f8050c54",
           373 => x"9408fc05",
           374 => x"08802e8c",
           375 => x"389408f8",
           376 => x"05083094",
           377 => x"08f8050c",
           378 => x"9408f805",
           379 => x"0870880c",
           380 => x"54873d0d",
           381 => x"940c0494",
           382 => x"0802940c",
           383 => x"fd3d0d81",
           384 => x"0b9408fc",
           385 => x"050c800b",
           386 => x"9408f805",
           387 => x"0c94088c",
           388 => x"05089408",
           389 => x"88050827",
           390 => x"ac389408",
           391 => x"fc050880",
           392 => x"2ea33880",
           393 => x"0b94088c",
           394 => x"05082499",
           395 => x"3894088c",
           396 => x"05081094",
           397 => x"088c050c",
           398 => x"9408fc05",
           399 => x"08109408",
           400 => x"fc050cc9",
           401 => x"399408fc",
           402 => x"0508802e",
           403 => x"80c93894",
           404 => x"088c0508",
           405 => x"94088805",
           406 => x"0826a138",
           407 => x"94088805",
           408 => x"0894088c",
           409 => x"05083194",
           410 => x"0888050c",
           411 => x"9408f805",
           412 => x"089408fc",
           413 => x"05080794",
           414 => x"08f8050c",
           415 => x"9408fc05",
           416 => x"08812a94",
           417 => x"08fc050c",
           418 => x"94088c05",
           419 => x"08812a94",
           420 => x"088c050c",
           421 => x"ffaf3994",
           422 => x"08900508",
           423 => x"802e8f38",
           424 => x"94088805",
           425 => x"08709408",
           426 => x"f4050c51",
           427 => x"8d399408",
           428 => x"f8050870",
           429 => x"9408f405",
           430 => x"0c519408",
           431 => x"f4050888",
           432 => x"0c853d0d",
           433 => x"940c04ff",
           434 => x"3d0d8188",
           435 => x"0b87c092",
           436 => x"8c0c810b",
           437 => x"87c0928c",
           438 => x"0c850b87",
           439 => x"c0988c0c",
           440 => x"87c0928c",
           441 => x"08708206",
           442 => x"51517080",
           443 => x"2e8a3887",
           444 => x"c0988c08",
           445 => x"5170e938",
           446 => x"87c0928c",
           447 => x"08fc8080",
           448 => x"06527193",
           449 => x"3887c098",
           450 => x"8c085170",
           451 => x"802e8838",
           452 => x"710b0b0b",
           453 => x"9fec340b",
           454 => x"0b0b9fec",
           455 => x"33880c83",
           456 => x"3d0d04fa",
           457 => x"3d0d787b",
           458 => x"7d565856",
           459 => x"800b0b0b",
           460 => x"0b9fec33",
           461 => x"81065255",
           462 => x"82527075",
           463 => x"2e098106",
           464 => x"819e3885",
           465 => x"0b87c098",
           466 => x"8c0c7987",
           467 => x"c092800c",
           468 => x"840b87c0",
           469 => x"928c0c87",
           470 => x"c0928c08",
           471 => x"70852a70",
           472 => x"81065152",
           473 => x"5370802e",
           474 => x"a73887c0",
           475 => x"92840870",
           476 => x"81ff0676",
           477 => x"79275253",
           478 => x"5173802e",
           479 => x"90387080",
           480 => x"2e8b3871",
           481 => x"76708105",
           482 => x"5834ff14",
           483 => x"54811555",
           484 => x"72a20651",
           485 => x"70802e8b",
           486 => x"3887c098",
           487 => x"8c085170",
           488 => x"ffb53887",
           489 => x"c0988c08",
           490 => x"51709538",
           491 => x"810b87c0",
           492 => x"928c0c87",
           493 => x"c0928c08",
           494 => x"70820651",
           495 => x"5170f438",
           496 => x"8073fc80",
           497 => x"80065252",
           498 => x"70722e09",
           499 => x"81068f38",
           500 => x"87c0988c",
           501 => x"08517072",
           502 => x"2e098106",
           503 => x"83388152",
           504 => x"71880c88",
           505 => x"3d0d04fe",
           506 => x"3d0d7481",
           507 => x"11337133",
           508 => x"71882b07",
           509 => x"880c5351",
           510 => x"843d0d04",
           511 => x"fd3d0d75",
           512 => x"83113382",
           513 => x"12337190",
           514 => x"2b71882b",
           515 => x"07811433",
           516 => x"70720788",
           517 => x"2b753371",
           518 => x"07880c52",
           519 => x"53545654",
           520 => x"52853d0d",
           521 => x"04f93d0d",
           522 => x"790b0b0b",
           523 => x"9ff00857",
           524 => x"57817727",
           525 => x"80ed3876",
           526 => x"88170827",
           527 => x"80e53875",
           528 => x"33557482",
           529 => x"2e893874",
           530 => x"832eae38",
           531 => x"80d53974",
           532 => x"54761083",
           533 => x"fe065376",
           534 => x"882a8c17",
           535 => x"08055288",
           536 => x"3d705255",
           537 => x"fdbd3f88",
           538 => x"08b93874",
           539 => x"51fef83f",
           540 => x"880883ff",
           541 => x"ff0655ad",
           542 => x"39845476",
           543 => x"822b83fc",
           544 => x"06537687",
           545 => x"2a8c1708",
           546 => x"0552883d",
           547 => x"705255fd",
           548 => x"923f8808",
           549 => x"8e387451",
           550 => x"fee23f88",
           551 => x"08f00a06",
           552 => x"55833981",
           553 => x"5574880c",
           554 => x"893d0d04",
           555 => x"fb3d0d0b",
           556 => x"0b0b9ff0",
           557 => x"08fe1988",
           558 => x"1208fe05",
           559 => x"55565480",
           560 => x"56747327",
           561 => x"8d388214",
           562 => x"33757129",
           563 => x"94160805",
           564 => x"57537588",
           565 => x"0c873d0d",
           566 => x"04fd3d0d",
           567 => x"7554800b",
           568 => x"0b0b0b9f",
           569 => x"f0087033",
           570 => x"51535371",
           571 => x"832e0981",
           572 => x"068c3894",
           573 => x"1451fdef",
           574 => x"3f880890",
           575 => x"2b539a14",
           576 => x"51fde43f",
           577 => x"880883ff",
           578 => x"ff067307",
           579 => x"880c853d",
           580 => x"0d04fc3d",
           581 => x"0d760b0b",
           582 => x"0b9ff008",
           583 => x"55558075",
           584 => x"23881508",
           585 => x"5372812e",
           586 => x"88388814",
           587 => x"08732685",
           588 => x"388152b0",
           589 => x"39729038",
           590 => x"73335271",
           591 => x"832e0981",
           592 => x"06853890",
           593 => x"14085372",
           594 => x"8c160c72",
           595 => x"802e8b38",
           596 => x"7251fed8",
           597 => x"3f880852",
           598 => x"85399014",
           599 => x"08527190",
           600 => x"160c8052",
           601 => x"71880c86",
           602 => x"3d0d04fa",
           603 => x"3d0d780b",
           604 => x"0b0b9ff0",
           605 => x"08712281",
           606 => x"057083ff",
           607 => x"ff065754",
           608 => x"57557380",
           609 => x"2e883890",
           610 => x"15085372",
           611 => x"86388352",
           612 => x"80dc3973",
           613 => x"8f065271",
           614 => x"80cf3881",
           615 => x"1390160c",
           616 => x"8c150853",
           617 => x"728f3883",
           618 => x"0b841722",
           619 => x"57527376",
           620 => x"27bc38b5",
           621 => x"39821633",
           622 => x"ff057484",
           623 => x"2a065271",
           624 => x"a8387251",
           625 => x"fcdf3f81",
           626 => x"52718808",
           627 => x"27a03883",
           628 => x"52880888",
           629 => x"17082796",
           630 => x"3888088c",
           631 => x"160c8808",
           632 => x"51fdc93f",
           633 => x"88089016",
           634 => x"0c737523",
           635 => x"80527188",
           636 => x"0c883d0d",
           637 => x"04f23d0d",
           638 => x"60626458",
           639 => x"5e5c7533",
           640 => x"5574a02e",
           641 => x"09810688",
           642 => x"38811670",
           643 => x"4456ef39",
           644 => x"62703356",
           645 => x"5674af2e",
           646 => x"09810684",
           647 => x"38811643",
           648 => x"800b881d",
           649 => x"0c627033",
           650 => x"5155749f",
           651 => x"268f387b",
           652 => x"51fddf3f",
           653 => x"88085680",
           654 => x"7d3482d3",
           655 => x"39933d84",
           656 => x"1d087058",
           657 => x"5a5f8a55",
           658 => x"a0767081",
           659 => x"055834ff",
           660 => x"155574ff",
           661 => x"2e098106",
           662 => x"ef388070",
           663 => x"595b887f",
           664 => x"085f5a7a",
           665 => x"811c7081",
           666 => x"ff066013",
           667 => x"703370af",
           668 => x"327030a0",
           669 => x"73277180",
           670 => x"25075151",
           671 => x"525b535d",
           672 => x"57557480",
           673 => x"c73876ae",
           674 => x"2e098106",
           675 => x"83388155",
           676 => x"777a2775",
           677 => x"07557480",
           678 => x"2e9f3879",
           679 => x"88327030",
           680 => x"78ae3270",
           681 => x"30707307",
           682 => x"9f2a5351",
           683 => x"57515675",
           684 => x"9b388858",
           685 => x"8b5affab",
           686 => x"39778119",
           687 => x"7081ff06",
           688 => x"721c535a",
           689 => x"57557675",
           690 => x"34ff9839",
           691 => x"7a1e7f0c",
           692 => x"805576a0",
           693 => x"26833881",
           694 => x"55748b1a",
           695 => x"347b51fc",
           696 => x"b13f8808",
           697 => x"80ef38a0",
           698 => x"547b2270",
           699 => x"852b83e0",
           700 => x"06545590",
           701 => x"1c08527c",
           702 => x"51f8a83f",
           703 => x"88085788",
           704 => x"0880fb38",
           705 => x"7c335574",
           706 => x"802e80ee",
           707 => x"388b1d33",
           708 => x"70832a70",
           709 => x"81065156",
           710 => x"5674b238",
           711 => x"8b7d841e",
           712 => x"08880859",
           713 => x"5b5b58ff",
           714 => x"185877ff",
           715 => x"2e9a3879",
           716 => x"7081055b",
           717 => x"33797081",
           718 => x"055b3371",
           719 => x"71315256",
           720 => x"5675802e",
           721 => x"e2388639",
           722 => x"75802e92",
           723 => x"387b51fc",
           724 => x"9a3fff8e",
           725 => x"39880856",
           726 => x"8808b438",
           727 => x"83397656",
           728 => x"841c088b",
           729 => x"11335155",
           730 => x"74a5388b",
           731 => x"1d337084",
           732 => x"2a708106",
           733 => x"51565674",
           734 => x"89388356",
           735 => x"92398156",
           736 => x"8e397c51",
           737 => x"fad33f88",
           738 => x"08881d0c",
           739 => x"fdaf3975",
           740 => x"880c903d",
           741 => x"0d04f93d",
           742 => x"0d797b59",
           743 => x"57825483",
           744 => x"fe537752",
           745 => x"7651f6fb",
           746 => x"3f835688",
           747 => x"0880e738",
           748 => x"7651f8b3",
           749 => x"3f880883",
           750 => x"ffff0655",
           751 => x"82567482",
           752 => x"d4d52e09",
           753 => x"810680ce",
           754 => x"387554b6",
           755 => x"53775276",
           756 => x"51f6d03f",
           757 => x"88085688",
           758 => x"08943876",
           759 => x"51f8883f",
           760 => x"880883ff",
           761 => x"ff065574",
           762 => x"8182c62e",
           763 => x"a9388254",
           764 => x"80d25377",
           765 => x"527651f6",
           766 => x"aa3f8808",
           767 => x"56880894",
           768 => x"387651f7",
           769 => x"e23f8808",
           770 => x"83ffff06",
           771 => x"55748182",
           772 => x"c62e8338",
           773 => x"81567588",
           774 => x"0c893d0d",
           775 => x"04ed3d0d",
           776 => x"6559800b",
           777 => x"0b0b0b9f",
           778 => x"f00cf59b",
           779 => x"3f880881",
           780 => x"06558256",
           781 => x"7482f238",
           782 => x"7475538d",
           783 => x"3d705357",
           784 => x"5afed33f",
           785 => x"880881ff",
           786 => x"06577681",
           787 => x"2e098106",
           788 => x"b3389054",
           789 => x"83be5374",
           790 => x"527551f5",
           791 => x"c63f8808",
           792 => x"ab388d3d",
           793 => x"33557480",
           794 => x"2eac3895",
           795 => x"3de40551",
           796 => x"f78a3f88",
           797 => x"08880853",
           798 => x"76525afe",
           799 => x"993f8808",
           800 => x"81ff0657",
           801 => x"76832e09",
           802 => x"81068638",
           803 => x"81568299",
           804 => x"3976802e",
           805 => x"86388656",
           806 => x"828f39a4",
           807 => x"548d5379",
           808 => x"527551f4",
           809 => x"fe3f8156",
           810 => x"880881fd",
           811 => x"38953de5",
           812 => x"0551f6b3",
           813 => x"3f880883",
           814 => x"ffff0658",
           815 => x"778c3895",
           816 => x"3df30551",
           817 => x"f6b63f88",
           818 => x"085802af",
           819 => x"05337871",
           820 => x"29028805",
           821 => x"ad057054",
           822 => x"52595bf6",
           823 => x"8a3f8808",
           824 => x"83ffff06",
           825 => x"7a058c1a",
           826 => x"0c8c3d33",
           827 => x"821a3495",
           828 => x"3de00551",
           829 => x"f5f13f88",
           830 => x"08841a23",
           831 => x"953de205",
           832 => x"51f5e43f",
           833 => x"880883ff",
           834 => x"ff065675",
           835 => x"8c38953d",
           836 => x"ef0551f5",
           837 => x"e73f8808",
           838 => x"567a51f5",
           839 => x"ca3f8808",
           840 => x"83ffff06",
           841 => x"76713179",
           842 => x"31841b22",
           843 => x"70842a82",
           844 => x"1d335672",
           845 => x"71315559",
           846 => x"5c5155ee",
           847 => x"c43f8808",
           848 => x"82057088",
           849 => x"1b0c8808",
           850 => x"e08a0556",
           851 => x"567483df",
           852 => x"fe268338",
           853 => x"825783ff",
           854 => x"f6762785",
           855 => x"38835789",
           856 => x"39865676",
           857 => x"802e80c1",
           858 => x"38767934",
           859 => x"76832e09",
           860 => x"81069038",
           861 => x"953dfb05",
           862 => x"51f5813f",
           863 => x"8808901a",
           864 => x"0c88398c",
           865 => x"19081890",
           866 => x"1a0c7983",
           867 => x"ffff068c",
           868 => x"1a081971",
           869 => x"842a0594",
           870 => x"1b0c5580",
           871 => x"0b811a34",
           872 => x"780b0b0b",
           873 => x"9ff00c80",
           874 => x"5675880c",
           875 => x"953d0d04",
           876 => x"ea3d0d0b",
           877 => x"0b0b9ff0",
           878 => x"08558554",
           879 => x"74802e80",
           880 => x"df38800b",
           881 => x"81163498",
           882 => x"3de01145",
           883 => x"6954893d",
           884 => x"705457ec",
           885 => x"0551f89d",
           886 => x"3f880854",
           887 => x"880880c0",
           888 => x"38883d33",
           889 => x"5473802e",
           890 => x"933802a7",
           891 => x"05337084",
           892 => x"2a708106",
           893 => x"51555773",
           894 => x"802e8538",
           895 => x"8354a139",
           896 => x"7551f5d5",
           897 => x"3f8808a0",
           898 => x"160c983d",
           899 => x"dc0551f3",
           900 => x"eb3f8808",
           901 => x"9c160c73",
           902 => x"98160c81",
           903 => x"0b811634",
           904 => x"73880c98",
           905 => x"3d0d04f6",
           906 => x"3d0d7d7f",
           907 => x"7e0b0b0b",
           908 => x"9ff00859",
           909 => x"5b5c5880",
           910 => x"7b0c8557",
           911 => x"75802e81",
           912 => x"d1388116",
           913 => x"33810655",
           914 => x"84577480",
           915 => x"2e81c338",
           916 => x"91397481",
           917 => x"17348639",
           918 => x"800b8117",
           919 => x"34815781",
           920 => x"b1399c16",
           921 => x"08981708",
           922 => x"31557478",
           923 => x"27833874",
           924 => x"5877802e",
           925 => x"819a3898",
           926 => x"16087083",
           927 => x"ff065657",
           928 => x"7480c738",
           929 => x"821633ff",
           930 => x"0577892a",
           931 => x"067081ff",
           932 => x"065b5579",
           933 => x"9e387687",
           934 => x"38a01608",
           935 => x"558b39a4",
           936 => x"160851f3",
           937 => x"803f8808",
           938 => x"55817527",
           939 => x"ffaa3874",
           940 => x"a4170ca4",
           941 => x"160851f3",
           942 => x"f33f8808",
           943 => x"55880880",
           944 => x"2eff8f38",
           945 => x"88081aa8",
           946 => x"170c9816",
           947 => x"0883ff06",
           948 => x"84807131",
           949 => x"51557775",
           950 => x"27833877",
           951 => x"55745498",
           952 => x"160883ff",
           953 => x"0653a816",
           954 => x"08527851",
           955 => x"f0b53f88",
           956 => x"08fee538",
           957 => x"98160815",
           958 => x"98170c77",
           959 => x"75317b08",
           960 => x"167c0c58",
           961 => x"78802efe",
           962 => x"e8387419",
           963 => x"59fee239",
           964 => x"80577688",
           965 => x"0c8c3d0d",
           966 => x"04fb3d0d",
           967 => x"87c0948c",
           968 => x"08548784",
           969 => x"80527351",
           970 => x"ead73f88",
           971 => x"08902b87",
           972 => x"c0948c08",
           973 => x"56548784",
           974 => x"80527451",
           975 => x"eac33f73",
           976 => x"88080787",
           977 => x"c0948c0c",
           978 => x"87c0949c",
           979 => x"08548784",
           980 => x"80527351",
           981 => x"eaab3f88",
           982 => x"08902b87",
           983 => x"c0949c08",
           984 => x"56548784",
           985 => x"80527451",
           986 => x"ea973f73",
           987 => x"88080787",
           988 => x"c0949c0c",
           989 => x"8c80830b",
           990 => x"87c09484",
           991 => x"0c8c8083",
           992 => x"0b87c094",
           993 => x"940c9ff4",
           994 => x"51f9923f",
           995 => x"8808b838",
           996 => x"9fdc51fc",
           997 => x"9b3f8808",
           998 => x"ae38a080",
           999 => x"0b880887",
          1000 => x"c098880c",
          1001 => x"55873dfc",
          1002 => x"05538480",
          1003 => x"527451fc",
          1004 => x"f63f8808",
          1005 => x"8d387554",
          1006 => x"73802e86",
          1007 => x"38731555",
          1008 => x"e439a080",
          1009 => x"54730480",
          1010 => x"54fb3900",
          1011 => x"00ffffff",
          1012 => x"ff00ffff",
          1013 => x"ffff00ff",
          1014 => x"ffffff00",
          1015 => x"424f4f54",
          1016 => x"54494e59",
          1017 => x"2e524f4d",
          1018 => x"00000000",
          1019 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

