-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use pkgs.config_pkg.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"84",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"84",
             9 => x"0b",
            10 => x"04",
            11 => x"84",
            12 => x"0b",
            13 => x"04",
            14 => x"84",
            15 => x"0b",
            16 => x"04",
            17 => x"84",
            18 => x"0b",
            19 => x"04",
            20 => x"84",
            21 => x"0b",
            22 => x"04",
            23 => x"85",
            24 => x"0b",
            25 => x"04",
            26 => x"85",
            27 => x"0b",
            28 => x"04",
            29 => x"85",
            30 => x"0b",
            31 => x"04",
            32 => x"85",
            33 => x"0b",
            34 => x"04",
            35 => x"86",
            36 => x"0b",
            37 => x"04",
            38 => x"86",
            39 => x"0b",
            40 => x"04",
            41 => x"86",
            42 => x"0b",
            43 => x"04",
            44 => x"86",
            45 => x"0b",
            46 => x"04",
            47 => x"87",
            48 => x"0b",
            49 => x"04",
            50 => x"87",
            51 => x"0b",
            52 => x"04",
            53 => x"87",
            54 => x"0b",
            55 => x"04",
            56 => x"87",
            57 => x"0b",
            58 => x"04",
            59 => x"88",
            60 => x"0b",
            61 => x"04",
            62 => x"88",
            63 => x"0b",
            64 => x"04",
            65 => x"88",
            66 => x"0b",
            67 => x"04",
            68 => x"88",
            69 => x"0b",
            70 => x"04",
            71 => x"89",
            72 => x"0b",
            73 => x"04",
            74 => x"89",
            75 => x"0b",
            76 => x"04",
            77 => x"89",
            78 => x"0b",
            79 => x"04",
            80 => x"89",
            81 => x"0b",
            82 => x"04",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"04",
           129 => x"0c",
           130 => x"81",
           131 => x"83",
           132 => x"81",
           133 => x"9f",
           134 => x"d3",
           135 => x"80",
           136 => x"d3",
           137 => x"ec",
           138 => x"b8",
           139 => x"90",
           140 => x"b8",
           141 => x"2d",
           142 => x"08",
           143 => x"04",
           144 => x"0c",
           145 => x"81",
           146 => x"83",
           147 => x"81",
           148 => x"a7",
           149 => x"d3",
           150 => x"80",
           151 => x"d3",
           152 => x"ab",
           153 => x"b8",
           154 => x"90",
           155 => x"b8",
           156 => x"2d",
           157 => x"08",
           158 => x"04",
           159 => x"0c",
           160 => x"81",
           161 => x"83",
           162 => x"81",
           163 => x"a6",
           164 => x"d3",
           165 => x"80",
           166 => x"d3",
           167 => x"9a",
           168 => x"b8",
           169 => x"90",
           170 => x"b8",
           171 => x"2d",
           172 => x"08",
           173 => x"04",
           174 => x"0c",
           175 => x"81",
           176 => x"83",
           177 => x"81",
           178 => x"97",
           179 => x"d3",
           180 => x"80",
           181 => x"d3",
           182 => x"bf",
           183 => x"b8",
           184 => x"90",
           185 => x"b8",
           186 => x"2d",
           187 => x"08",
           188 => x"04",
           189 => x"0c",
           190 => x"81",
           191 => x"83",
           192 => x"81",
           193 => x"80",
           194 => x"81",
           195 => x"83",
           196 => x"81",
           197 => x"80",
           198 => x"81",
           199 => x"83",
           200 => x"81",
           201 => x"80",
           202 => x"81",
           203 => x"83",
           204 => x"81",
           205 => x"80",
           206 => x"81",
           207 => x"83",
           208 => x"81",
           209 => x"80",
           210 => x"81",
           211 => x"83",
           212 => x"81",
           213 => x"80",
           214 => x"81",
           215 => x"83",
           216 => x"81",
           217 => x"80",
           218 => x"81",
           219 => x"83",
           220 => x"81",
           221 => x"80",
           222 => x"81",
           223 => x"83",
           224 => x"81",
           225 => x"80",
           226 => x"81",
           227 => x"83",
           228 => x"81",
           229 => x"80",
           230 => x"81",
           231 => x"83",
           232 => x"81",
           233 => x"81",
           234 => x"81",
           235 => x"83",
           236 => x"81",
           237 => x"80",
           238 => x"81",
           239 => x"83",
           240 => x"81",
           241 => x"81",
           242 => x"81",
           243 => x"83",
           244 => x"81",
           245 => x"80",
           246 => x"81",
           247 => x"83",
           248 => x"81",
           249 => x"81",
           250 => x"81",
           251 => x"83",
           252 => x"81",
           253 => x"81",
           254 => x"81",
           255 => x"83",
           256 => x"81",
           257 => x"80",
           258 => x"81",
           259 => x"83",
           260 => x"81",
           261 => x"80",
           262 => x"81",
           263 => x"83",
           264 => x"81",
           265 => x"80",
           266 => x"81",
           267 => x"83",
           268 => x"81",
           269 => x"80",
           270 => x"81",
           271 => x"83",
           272 => x"81",
           273 => x"81",
           274 => x"81",
           275 => x"83",
           276 => x"81",
           277 => x"81",
           278 => x"81",
           279 => x"83",
           280 => x"81",
           281 => x"81",
           282 => x"81",
           283 => x"83",
           284 => x"81",
           285 => x"80",
           286 => x"81",
           287 => x"83",
           288 => x"81",
           289 => x"81",
           290 => x"81",
           291 => x"83",
           292 => x"81",
           293 => x"ad",
           294 => x"d3",
           295 => x"80",
           296 => x"d3",
           297 => x"be",
           298 => x"b8",
           299 => x"90",
           300 => x"b8",
           301 => x"2d",
           302 => x"08",
           303 => x"04",
           304 => x"0c",
           305 => x"81",
           306 => x"83",
           307 => x"81",
           308 => x"90",
           309 => x"d3",
           310 => x"80",
           311 => x"d3",
           312 => x"da",
           313 => x"b8",
           314 => x"90",
           315 => x"b8",
           316 => x"c4",
           317 => x"b8",
           318 => x"90",
           319 => x"ac",
           320 => x"b0",
           321 => x"80",
           322 => x"05",
           323 => x"0b",
           324 => x"04",
           325 => x"81",
           326 => x"3c",
           327 => x"b8",
           328 => x"d3",
           329 => x"3d",
           330 => x"81",
           331 => x"8c",
           332 => x"81",
           333 => x"88",
           334 => x"80",
           335 => x"d3",
           336 => x"81",
           337 => x"54",
           338 => x"81",
           339 => x"04",
           340 => x"08",
           341 => x"b8",
           342 => x"0d",
           343 => x"d3",
           344 => x"05",
           345 => x"d3",
           346 => x"05",
           347 => x"3f",
           348 => x"08",
           349 => x"ac",
           350 => x"3d",
           351 => x"b8",
           352 => x"d3",
           353 => x"81",
           354 => x"fd",
           355 => x"0b",
           356 => x"08",
           357 => x"80",
           358 => x"b8",
           359 => x"0c",
           360 => x"08",
           361 => x"81",
           362 => x"88",
           363 => x"b9",
           364 => x"b8",
           365 => x"08",
           366 => x"38",
           367 => x"d3",
           368 => x"05",
           369 => x"38",
           370 => x"08",
           371 => x"10",
           372 => x"08",
           373 => x"81",
           374 => x"fc",
           375 => x"81",
           376 => x"fc",
           377 => x"b8",
           378 => x"b8",
           379 => x"08",
           380 => x"e1",
           381 => x"b8",
           382 => x"08",
           383 => x"08",
           384 => x"26",
           385 => x"d3",
           386 => x"05",
           387 => x"b8",
           388 => x"08",
           389 => x"b8",
           390 => x"0c",
           391 => x"08",
           392 => x"81",
           393 => x"fc",
           394 => x"81",
           395 => x"f8",
           396 => x"d3",
           397 => x"05",
           398 => x"81",
           399 => x"fc",
           400 => x"d3",
           401 => x"05",
           402 => x"81",
           403 => x"8c",
           404 => x"95",
           405 => x"b8",
           406 => x"08",
           407 => x"38",
           408 => x"08",
           409 => x"70",
           410 => x"08",
           411 => x"51",
           412 => x"d3",
           413 => x"05",
           414 => x"d3",
           415 => x"05",
           416 => x"d3",
           417 => x"05",
           418 => x"ac",
           419 => x"0d",
           420 => x"0c",
           421 => x"0d",
           422 => x"02",
           423 => x"05",
           424 => x"53",
           425 => x"27",
           426 => x"83",
           427 => x"80",
           428 => x"ff",
           429 => x"ff",
           430 => x"73",
           431 => x"05",
           432 => x"12",
           433 => x"2e",
           434 => x"ef",
           435 => x"d3",
           436 => x"3d",
           437 => x"74",
           438 => x"07",
           439 => x"2b",
           440 => x"51",
           441 => x"a5",
           442 => x"70",
           443 => x"0c",
           444 => x"84",
           445 => x"72",
           446 => x"05",
           447 => x"71",
           448 => x"53",
           449 => x"52",
           450 => x"dd",
           451 => x"27",
           452 => x"71",
           453 => x"53",
           454 => x"52",
           455 => x"f2",
           456 => x"ff",
           457 => x"3d",
           458 => x"70",
           459 => x"06",
           460 => x"70",
           461 => x"73",
           462 => x"56",
           463 => x"08",
           464 => x"38",
           465 => x"52",
           466 => x"81",
           467 => x"54",
           468 => x"9d",
           469 => x"55",
           470 => x"09",
           471 => x"38",
           472 => x"14",
           473 => x"81",
           474 => x"56",
           475 => x"e5",
           476 => x"55",
           477 => x"06",
           478 => x"06",
           479 => x"81",
           480 => x"52",
           481 => x"0d",
           482 => x"70",
           483 => x"ff",
           484 => x"f8",
           485 => x"80",
           486 => x"51",
           487 => x"84",
           488 => x"71",
           489 => x"54",
           490 => x"2e",
           491 => x"75",
           492 => x"94",
           493 => x"81",
           494 => x"87",
           495 => x"fe",
           496 => x"70",
           497 => x"88",
           498 => x"9b",
           499 => x"ac",
           500 => x"06",
           501 => x"14",
           502 => x"73",
           503 => x"71",
           504 => x"0c",
           505 => x"04",
           506 => x"76",
           507 => x"53",
           508 => x"80",
           509 => x"38",
           510 => x"70",
           511 => x"81",
           512 => x"81",
           513 => x"52",
           514 => x"2e",
           515 => x"52",
           516 => x"12",
           517 => x"33",
           518 => x"a0",
           519 => x"81",
           520 => x"70",
           521 => x"06",
           522 => x"e6",
           523 => x"51",
           524 => x"09",
           525 => x"38",
           526 => x"81",
           527 => x"71",
           528 => x"51",
           529 => x"ac",
           530 => x"0d",
           531 => x"0d",
           532 => x"08",
           533 => x"38",
           534 => x"05",
           535 => x"99",
           536 => x"d3",
           537 => x"38",
           538 => x"39",
           539 => x"81",
           540 => x"86",
           541 => x"f5",
           542 => x"82",
           543 => x"05",
           544 => x"5b",
           545 => x"81",
           546 => x"1c",
           547 => x"5a",
           548 => x"9e",
           549 => x"38",
           550 => x"5a",
           551 => x"97",
           552 => x"38",
           553 => x"5a",
           554 => x"bb",
           555 => x"38",
           556 => x"5a",
           557 => x"bb",
           558 => x"38",
           559 => x"5a",
           560 => x"87",
           561 => x"80",
           562 => x"22",
           563 => x"79",
           564 => x"80",
           565 => x"1c",
           566 => x"1c",
           567 => x"1c",
           568 => x"1c",
           569 => x"1c",
           570 => x"1c",
           571 => x"1c",
           572 => x"22",
           573 => x"8c",
           574 => x"3f",
           575 => x"9c",
           576 => x"0c",
           577 => x"c0",
           578 => x"82",
           579 => x"c0",
           580 => x"83",
           581 => x"c0",
           582 => x"84",
           583 => x"c0",
           584 => x"85",
           585 => x"c0",
           586 => x"86",
           587 => x"c0",
           588 => x"88",
           589 => x"c0",
           590 => x"8a",
           591 => x"c0",
           592 => x"80",
           593 => x"5b",
           594 => x"ac",
           595 => x"0d",
           596 => x"0d",
           597 => x"c0",
           598 => x"81",
           599 => x"c0",
           600 => x"5b",
           601 => x"87",
           602 => x"08",
           603 => x"1b",
           604 => x"98",
           605 => x"7a",
           606 => x"87",
           607 => x"08",
           608 => x"1b",
           609 => x"98",
           610 => x"7a",
           611 => x"87",
           612 => x"08",
           613 => x"1b",
           614 => x"98",
           615 => x"7a",
           616 => x"87",
           617 => x"08",
           618 => x"1b",
           619 => x"0c",
           620 => x"59",
           621 => x"58",
           622 => x"57",
           623 => x"56",
           624 => x"55",
           625 => x"54",
           626 => x"53",
           627 => x"81",
           628 => x"92",
           629 => x"3d",
           630 => x"3d",
           631 => x"05",
           632 => x"70",
           633 => x"51",
           634 => x"0b",
           635 => x"34",
           636 => x"04",
           637 => x"75",
           638 => x"cb",
           639 => x"54",
           640 => x"84",
           641 => x"2e",
           642 => x"c0",
           643 => x"70",
           644 => x"2a",
           645 => x"51",
           646 => x"80",
           647 => x"71",
           648 => x"81",
           649 => x"70",
           650 => x"96",
           651 => x"70",
           652 => x"51",
           653 => x"8d",
           654 => x"2a",
           655 => x"51",
           656 => x"bc",
           657 => x"81",
           658 => x"51",
           659 => x"80",
           660 => x"2e",
           661 => x"c0",
           662 => x"73",
           663 => x"81",
           664 => x"85",
           665 => x"fd",
           666 => x"97",
           667 => x"0b",
           668 => x"33",
           669 => x"c0",
           670 => x"72",
           671 => x"38",
           672 => x"94",
           673 => x"70",
           674 => x"81",
           675 => x"52",
           676 => x"8c",
           677 => x"2a",
           678 => x"51",
           679 => x"38",
           680 => x"81",
           681 => x"06",
           682 => x"80",
           683 => x"71",
           684 => x"81",
           685 => x"70",
           686 => x"0b",
           687 => x"a4",
           688 => x"c0",
           689 => x"70",
           690 => x"38",
           691 => x"90",
           692 => x"0c",
           693 => x"04",
           694 => x"77",
           695 => x"33",
           696 => x"76",
           697 => x"38",
           698 => x"05",
           699 => x"0b",
           700 => x"33",
           701 => x"c0",
           702 => x"72",
           703 => x"38",
           704 => x"94",
           705 => x"70",
           706 => x"81",
           707 => x"52",
           708 => x"8c",
           709 => x"2a",
           710 => x"51",
           711 => x"38",
           712 => x"81",
           713 => x"06",
           714 => x"80",
           715 => x"71",
           716 => x"81",
           717 => x"70",
           718 => x"0b",
           719 => x"a4",
           720 => x"c0",
           721 => x"70",
           722 => x"38",
           723 => x"90",
           724 => x"0c",
           725 => x"33",
           726 => x"ff",
           727 => x"81",
           728 => x"87",
           729 => x"ff",
           730 => x"0b",
           731 => x"33",
           732 => x"94",
           733 => x"80",
           734 => x"87",
           735 => x"51",
           736 => x"82",
           737 => x"06",
           738 => x"70",
           739 => x"38",
           740 => x"cb",
           741 => x"87",
           742 => x"52",
           743 => x"86",
           744 => x"94",
           745 => x"08",
           746 => x"06",
           747 => x"0c",
           748 => x"0d",
           749 => x"0d",
           750 => x"cb",
           751 => x"87",
           752 => x"52",
           753 => x"86",
           754 => x"94",
           755 => x"08",
           756 => x"70",
           757 => x"51",
           758 => x"70",
           759 => x"38",
           760 => x"cb",
           761 => x"87",
           762 => x"52",
           763 => x"86",
           764 => x"94",
           765 => x"08",
           766 => x"70",
           767 => x"53",
           768 => x"d3",
           769 => x"3d",
           770 => x"3d",
           771 => x"9e",
           772 => x"70",
           773 => x"06",
           774 => x"70",
           775 => x"9f",
           776 => x"a8",
           777 => x"9e",
           778 => x"0c",
           779 => x"c0",
           780 => x"71",
           781 => x"11",
           782 => x"8c",
           783 => x"52",
           784 => x"c0",
           785 => x"71",
           786 => x"11",
           787 => x"94",
           788 => x"52",
           789 => x"c0",
           790 => x"71",
           791 => x"11",
           792 => x"a4",
           793 => x"52",
           794 => x"c0",
           795 => x"71",
           796 => x"11",
           797 => x"ac",
           798 => x"52",
           799 => x"52",
           800 => x"23",
           801 => x"c0",
           802 => x"71",
           803 => x"0b",
           804 => x"ad",
           805 => x"0b",
           806 => x"88",
           807 => x"80",
           808 => x"53",
           809 => x"83",
           810 => x"72",
           811 => x"0b",
           812 => x"88",
           813 => x"80",
           814 => x"52",
           815 => x"2e",
           816 => x"52",
           817 => x"d6",
           818 => x"87",
           819 => x"08",
           820 => x"80",
           821 => x"52",
           822 => x"83",
           823 => x"71",
           824 => x"34",
           825 => x"c0",
           826 => x"70",
           827 => x"51",
           828 => x"80",
           829 => x"81",
           830 => x"cb",
           831 => x"0b",
           832 => x"88",
           833 => x"80",
           834 => x"52",
           835 => x"83",
           836 => x"71",
           837 => x"34",
           838 => x"c0",
           839 => x"70",
           840 => x"51",
           841 => x"80",
           842 => x"81",
           843 => x"cb",
           844 => x"0b",
           845 => x"88",
           846 => x"80",
           847 => x"52",
           848 => x"83",
           849 => x"71",
           850 => x"34",
           851 => x"c0",
           852 => x"70",
           853 => x"51",
           854 => x"80",
           855 => x"81",
           856 => x"cb",
           857 => x"cb",
           858 => x"c0",
           859 => x"08",
           860 => x"06",
           861 => x"51",
           862 => x"70",
           863 => x"05",
           864 => x"54",
           865 => x"70",
           866 => x"52",
           867 => x"2e",
           868 => x"52",
           869 => x"80",
           870 => x"9e",
           871 => x"88",
           872 => x"52",
           873 => x"83",
           874 => x"71",
           875 => x"34",
           876 => x"88",
           877 => x"06",
           878 => x"81",
           879 => x"85",
           880 => x"fc",
           881 => x"b6",
           882 => x"be",
           883 => x"d4",
           884 => x"80",
           885 => x"81",
           886 => x"84",
           887 => x"b6",
           888 => x"a6",
           889 => x"d5",
           890 => x"55",
           891 => x"91",
           892 => x"08",
           893 => x"a8",
           894 => x"b6",
           895 => x"84",
           896 => x"d6",
           897 => x"55",
           898 => x"90",
           899 => x"08",
           900 => x"08",
           901 => x"8c",
           902 => x"3f",
           903 => x"70",
           904 => x"73",
           905 => x"15",
           906 => x"80",
           907 => x"81",
           908 => x"08",
           909 => x"08",
           910 => x"b7",
           911 => x"c4",
           912 => x"d9",
           913 => x"80",
           914 => x"81",
           915 => x"83",
           916 => x"cb",
           917 => x"73",
           918 => x"38",
           919 => x"51",
           920 => x"81",
           921 => x"54",
           922 => x"88",
           923 => x"ec",
           924 => x"3f",
           925 => x"70",
           926 => x"73",
           927 => x"38",
           928 => x"52",
           929 => x"51",
           930 => x"81",
           931 => x"54",
           932 => x"88",
           933 => x"98",
           934 => x"3f",
           935 => x"70",
           936 => x"73",
           937 => x"38",
           938 => x"52",
           939 => x"51",
           940 => x"81",
           941 => x"82",
           942 => x"cb",
           943 => x"70",
           944 => x"08",
           945 => x"dc",
           946 => x"88",
           947 => x"08",
           948 => x"84",
           949 => x"3f",
           950 => x"52",
           951 => x"51",
           952 => x"8c",
           953 => x"81",
           954 => x"88",
           955 => x"15",
           956 => x"b9",
           957 => x"8c",
           958 => x"0d",
           959 => x"0d",
           960 => x"33",
           961 => x"26",
           962 => x"10",
           963 => x"81",
           964 => x"52",
           965 => x"81",
           966 => x"f7",
           967 => x"39",
           968 => x"51",
           969 => x"a3",
           970 => x"b4",
           971 => x"3f",
           972 => x"ba",
           973 => x"a0",
           974 => x"81",
           975 => x"f7",
           976 => x"39",
           977 => x"51",
           978 => x"83",
           979 => x"71",
           980 => x"04",
           981 => x"c0",
           982 => x"04",
           983 => x"87",
           984 => x"70",
           985 => x"80",
           986 => x"74",
           987 => x"cb",
           988 => x"0c",
           989 => x"04",
           990 => x"87",
           991 => x"70",
           992 => x"e4",
           993 => x"72",
           994 => x"70",
           995 => x"08",
           996 => x"cb",
           997 => x"0c",
           998 => x"0d",
           999 => x"e4",
          1000 => x"96",
          1001 => x"fe",
          1002 => x"93",
          1003 => x"72",
          1004 => x"81",
          1005 => x"8d",
          1006 => x"81",
          1007 => x"80",
          1008 => x"81",
          1009 => x"52",
          1010 => x"81",
          1011 => x"81",
          1012 => x"c4",
          1013 => x"81",
          1014 => x"80",
          1015 => x"72",
          1016 => x"bc",
          1017 => x"2d",
          1018 => x"04",
          1019 => x"02",
          1020 => x"81",
          1021 => x"76",
          1022 => x"0c",
          1023 => x"a7",
          1024 => x"d3",
          1025 => x"3d",
          1026 => x"3d",
          1027 => x"33",
          1028 => x"80",
          1029 => x"72",
          1030 => x"54",
          1031 => x"87",
          1032 => x"52",
          1033 => x"84",
          1034 => x"fd",
          1035 => x"81",
          1036 => x"77",
          1037 => x"0c",
          1038 => x"55",
          1039 => x"2e",
          1040 => x"70",
          1041 => x"33",
          1042 => x"3f",
          1043 => x"71",
          1044 => x"81",
          1045 => x"85",
          1046 => x"ec",
          1047 => x"68",
          1048 => x"70",
          1049 => x"33",
          1050 => x"2e",
          1051 => x"75",
          1052 => x"38",
          1053 => x"af",
          1054 => x"80",
          1055 => x"81",
          1056 => x"58",
          1057 => x"b0",
          1058 => x"06",
          1059 => x"79",
          1060 => x"5b",
          1061 => x"92",
          1062 => x"2e",
          1063 => x"8a",
          1064 => x"70",
          1065 => x"33",
          1066 => x"aa",
          1067 => x"06",
          1068 => x"84",
          1069 => x"7b",
          1070 => x"5d",
          1071 => x"5d",
          1072 => x"d0",
          1073 => x"89",
          1074 => x"79",
          1075 => x"d0",
          1076 => x"81",
          1077 => x"d0",
          1078 => x"5a",
          1079 => x"eb",
          1080 => x"ec",
          1081 => x"70",
          1082 => x"25",
          1083 => x"32",
          1084 => x"72",
          1085 => x"73",
          1086 => x"52",
          1087 => x"73",
          1088 => x"38",
          1089 => x"79",
          1090 => x"5b",
          1091 => x"75",
          1092 => x"ec",
          1093 => x"80",
          1094 => x"89",
          1095 => x"70",
          1096 => x"56",
          1097 => x"15",
          1098 => x"26",
          1099 => x"72",
          1100 => x"b0",
          1101 => x"72",
          1102 => x"84",
          1103 => x"57",
          1104 => x"75",
          1105 => x"72",
          1106 => x"38",
          1107 => x"16",
          1108 => x"54",
          1109 => x"38",
          1110 => x"70",
          1111 => x"53",
          1112 => x"73",
          1113 => x"53",
          1114 => x"99",
          1115 => x"2a",
          1116 => x"a0",
          1117 => x"3f",
          1118 => x"73",
          1119 => x"53",
          1120 => x"ef",
          1121 => x"fd",
          1122 => x"81",
          1123 => x"72",
          1124 => x"ce",
          1125 => x"fc",
          1126 => x"81",
          1127 => x"79",
          1128 => x"38",
          1129 => x"7b",
          1130 => x"12",
          1131 => x"53",
          1132 => x"fd",
          1133 => x"5b",
          1134 => x"5b",
          1135 => x"5b",
          1136 => x"5b",
          1137 => x"51",
          1138 => x"fd",
          1139 => x"82",
          1140 => x"06",
          1141 => x"80",
          1142 => x"7b",
          1143 => x"08",
          1144 => x"9c",
          1145 => x"c4",
          1146 => x"06",
          1147 => x"84",
          1148 => x"59",
          1149 => x"39",
          1150 => x"71",
          1151 => x"53",
          1152 => x"32",
          1153 => x"72",
          1154 => x"70",
          1155 => x"06",
          1156 => x"53",
          1157 => x"88",
          1158 => x"7d",
          1159 => x"57",
          1160 => x"52",
          1161 => x"a8",
          1162 => x"ac",
          1163 => x"06",
          1164 => x"52",
          1165 => x"3f",
          1166 => x"08",
          1167 => x"27",
          1168 => x"a7",
          1169 => x"ff",
          1170 => x"54",
          1171 => x"2e",
          1172 => x"14",
          1173 => x"06",
          1174 => x"3d",
          1175 => x"05",
          1176 => x"54",
          1177 => x"81",
          1178 => x"70",
          1179 => x"2a",
          1180 => x"27",
          1181 => x"54",
          1182 => x"a6",
          1183 => x"2a",
          1184 => x"51",
          1185 => x"2e",
          1186 => x"3d",
          1187 => x"05",
          1188 => x"34",
          1189 => x"77",
          1190 => x"54",
          1191 => x"72",
          1192 => x"55",
          1193 => x"70",
          1194 => x"53",
          1195 => x"73",
          1196 => x"53",
          1197 => x"99",
          1198 => x"2a",
          1199 => x"74",
          1200 => x"3f",
          1201 => x"73",
          1202 => x"53",
          1203 => x"ef",
          1204 => x"97",
          1205 => x"11",
          1206 => x"54",
          1207 => x"3f",
          1208 => x"73",
          1209 => x"53",
          1210 => x"fa",
          1211 => x"51",
          1212 => x"73",
          1213 => x"53",
          1214 => x"f2",
          1215 => x"39",
          1216 => x"04",
          1217 => x"86",
          1218 => x"84",
          1219 => x"55",
          1220 => x"fa",
          1221 => x"3d",
          1222 => x"3d",
          1223 => x"d3",
          1224 => x"3d",
          1225 => x"75",
          1226 => x"3f",
          1227 => x"08",
          1228 => x"34",
          1229 => x"d3",
          1230 => x"3d",
          1231 => x"3d",
          1232 => x"bc",
          1233 => x"d3",
          1234 => x"3d",
          1235 => x"77",
          1236 => x"87",
          1237 => x"d3",
          1238 => x"3d",
          1239 => x"3d",
          1240 => x"57",
          1241 => x"81",
          1242 => x"73",
          1243 => x"38",
          1244 => x"53",
          1245 => x"80",
          1246 => x"c0",
          1247 => x"2d",
          1248 => x"08",
          1249 => x"54",
          1250 => x"e6",
          1251 => x"2e",
          1252 => x"73",
          1253 => x"30",
          1254 => x"78",
          1255 => x"72",
          1256 => x"52",
          1257 => x"72",
          1258 => x"38",
          1259 => x"81",
          1260 => x"55",
          1261 => x"c1",
          1262 => x"25",
          1263 => x"ff",
          1264 => x"72",
          1265 => x"38",
          1266 => x"73",
          1267 => x"15",
          1268 => x"06",
          1269 => x"cf",
          1270 => x"39",
          1271 => x"80",
          1272 => x"51",
          1273 => x"81",
          1274 => x"d3",
          1275 => x"3d",
          1276 => x"3d",
          1277 => x"c0",
          1278 => x"d3",
          1279 => x"53",
          1280 => x"fe",
          1281 => x"81",
          1282 => x"84",
          1283 => x"f8",
          1284 => x"7c",
          1285 => x"70",
          1286 => x"08",
          1287 => x"54",
          1288 => x"2e",
          1289 => x"92",
          1290 => x"81",
          1291 => x"74",
          1292 => x"55",
          1293 => x"2e",
          1294 => x"ad",
          1295 => x"06",
          1296 => x"75",
          1297 => x"0c",
          1298 => x"33",
          1299 => x"73",
          1300 => x"81",
          1301 => x"38",
          1302 => x"05",
          1303 => x"08",
          1304 => x"53",
          1305 => x"2e",
          1306 => x"80",
          1307 => x"81",
          1308 => x"90",
          1309 => x"76",
          1310 => x"70",
          1311 => x"57",
          1312 => x"82",
          1313 => x"05",
          1314 => x"08",
          1315 => x"54",
          1316 => x"81",
          1317 => x"27",
          1318 => x"d0",
          1319 => x"56",
          1320 => x"73",
          1321 => x"80",
          1322 => x"14",
          1323 => x"72",
          1324 => x"e8",
          1325 => x"80",
          1326 => x"39",
          1327 => x"dc",
          1328 => x"80",
          1329 => x"27",
          1330 => x"80",
          1331 => x"89",
          1332 => x"70",
          1333 => x"55",
          1334 => x"70",
          1335 => x"55",
          1336 => x"27",
          1337 => x"14",
          1338 => x"06",
          1339 => x"74",
          1340 => x"73",
          1341 => x"38",
          1342 => x"14",
          1343 => x"05",
          1344 => x"08",
          1345 => x"54",
          1346 => x"26",
          1347 => x"77",
          1348 => x"38",
          1349 => x"75",
          1350 => x"56",
          1351 => x"ac",
          1352 => x"0d",
          1353 => x"0d",
          1354 => x"55",
          1355 => x"0c",
          1356 => x"33",
          1357 => x"73",
          1358 => x"81",
          1359 => x"74",
          1360 => x"75",
          1361 => x"70",
          1362 => x"73",
          1363 => x"38",
          1364 => x"09",
          1365 => x"38",
          1366 => x"11",
          1367 => x"08",
          1368 => x"54",
          1369 => x"2e",
          1370 => x"80",
          1371 => x"08",
          1372 => x"0c",
          1373 => x"33",
          1374 => x"80",
          1375 => x"38",
          1376 => x"2e",
          1377 => x"a1",
          1378 => x"81",
          1379 => x"75",
          1380 => x"56",
          1381 => x"c1",
          1382 => x"08",
          1383 => x"0c",
          1384 => x"33",
          1385 => x"b1",
          1386 => x"a0",
          1387 => x"82",
          1388 => x"53",
          1389 => x"57",
          1390 => x"9d",
          1391 => x"39",
          1392 => x"80",
          1393 => x"26",
          1394 => x"8b",
          1395 => x"80",
          1396 => x"56",
          1397 => x"8a",
          1398 => x"a0",
          1399 => x"c5",
          1400 => x"74",
          1401 => x"e0",
          1402 => x"ff",
          1403 => x"d0",
          1404 => x"ff",
          1405 => x"90",
          1406 => x"38",
          1407 => x"81",
          1408 => x"53",
          1409 => x"c5",
          1410 => x"27",
          1411 => x"76",
          1412 => x"08",
          1413 => x"0c",
          1414 => x"33",
          1415 => x"73",
          1416 => x"bd",
          1417 => x"2e",
          1418 => x"30",
          1419 => x"0c",
          1420 => x"81",
          1421 => x"8a",
          1422 => x"ff",
          1423 => x"8f",
          1424 => x"81",
          1425 => x"26",
          1426 => x"cb",
          1427 => x"52",
          1428 => x"ac",
          1429 => x"0d",
          1430 => x"0d",
          1431 => x"33",
          1432 => x"9b",
          1433 => x"53",
          1434 => x"81",
          1435 => x"38",
          1436 => x"87",
          1437 => x"05",
          1438 => x"73",
          1439 => x"38",
          1440 => x"71",
          1441 => x"90",
          1442 => x"92",
          1443 => x"81",
          1444 => x"0b",
          1445 => x"8c",
          1446 => x"87",
          1447 => x"54",
          1448 => x"82",
          1449 => x"70",
          1450 => x"38",
          1451 => x"70",
          1452 => x"90",
          1453 => x"92",
          1454 => x"08",
          1455 => x"06",
          1456 => x"92",
          1457 => x"98",
          1458 => x"70",
          1459 => x"38",
          1460 => x"e8",
          1461 => x"cb",
          1462 => x"51",
          1463 => x"ac",
          1464 => x"0d",
          1465 => x"0d",
          1466 => x"02",
          1467 => x"c3",
          1468 => x"41",
          1469 => x"73",
          1470 => x"bf",
          1471 => x"ac",
          1472 => x"7b",
          1473 => x"81",
          1474 => x"70",
          1475 => x"c0",
          1476 => x"84",
          1477 => x"92",
          1478 => x"c0",
          1479 => x"72",
          1480 => x"5b",
          1481 => x"0c",
          1482 => x"80",
          1483 => x"0c",
          1484 => x"0c",
          1485 => x"85",
          1486 => x"06",
          1487 => x"71",
          1488 => x"38",
          1489 => x"71",
          1490 => x"05",
          1491 => x"17",
          1492 => x"06",
          1493 => x"2e",
          1494 => x"08",
          1495 => x"38",
          1496 => x"71",
          1497 => x"38",
          1498 => x"2e",
          1499 => x"75",
          1500 => x"92",
          1501 => x"72",
          1502 => x"06",
          1503 => x"f7",
          1504 => x"5b",
          1505 => x"80",
          1506 => x"70",
          1507 => x"5f",
          1508 => x"80",
          1509 => x"73",
          1510 => x"06",
          1511 => x"38",
          1512 => x"ff",
          1513 => x"fc",
          1514 => x"52",
          1515 => x"83",
          1516 => x"71",
          1517 => x"d3",
          1518 => x"3d",
          1519 => x"3d",
          1520 => x"64",
          1521 => x"bf",
          1522 => x"40",
          1523 => x"73",
          1524 => x"e7",
          1525 => x"ac",
          1526 => x"7a",
          1527 => x"81",
          1528 => x"5c",
          1529 => x"8c",
          1530 => x"87",
          1531 => x"11",
          1532 => x"84",
          1533 => x"5b",
          1534 => x"85",
          1535 => x"c0",
          1536 => x"7b",
          1537 => x"82",
          1538 => x"53",
          1539 => x"84",
          1540 => x"06",
          1541 => x"71",
          1542 => x"38",
          1543 => x"05",
          1544 => x"0c",
          1545 => x"73",
          1546 => x"81",
          1547 => x"71",
          1548 => x"38",
          1549 => x"71",
          1550 => x"08",
          1551 => x"2e",
          1552 => x"84",
          1553 => x"38",
          1554 => x"87",
          1555 => x"1d",
          1556 => x"70",
          1557 => x"52",
          1558 => x"ff",
          1559 => x"39",
          1560 => x"81",
          1561 => x"80",
          1562 => x"52",
          1563 => x"90",
          1564 => x"80",
          1565 => x"71",
          1566 => x"7c",
          1567 => x"38",
          1568 => x"80",
          1569 => x"80",
          1570 => x"81",
          1571 => x"73",
          1572 => x"0c",
          1573 => x"04",
          1574 => x"7d",
          1575 => x"af",
          1576 => x"88",
          1577 => x"33",
          1578 => x"56",
          1579 => x"3f",
          1580 => x"08",
          1581 => x"83",
          1582 => x"38",
          1583 => x"74",
          1584 => x"72",
          1585 => x"38",
          1586 => x"8a",
          1587 => x"72",
          1588 => x"38",
          1589 => x"90",
          1590 => x"92",
          1591 => x"08",
          1592 => x"39",
          1593 => x"76",
          1594 => x"8b",
          1595 => x"76",
          1596 => x"83",
          1597 => x"73",
          1598 => x"0c",
          1599 => x"04",
          1600 => x"73",
          1601 => x"12",
          1602 => x"2b",
          1603 => x"d3",
          1604 => x"52",
          1605 => x"0d",
          1606 => x"0d",
          1607 => x"33",
          1608 => x"71",
          1609 => x"88",
          1610 => x"14",
          1611 => x"74",
          1612 => x"2b",
          1613 => x"ac",
          1614 => x"56",
          1615 => x"3d",
          1616 => x"3d",
          1617 => x"84",
          1618 => x"22",
          1619 => x"72",
          1620 => x"54",
          1621 => x"2a",
          1622 => x"34",
          1623 => x"04",
          1624 => x"73",
          1625 => x"70",
          1626 => x"05",
          1627 => x"88",
          1628 => x"72",
          1629 => x"54",
          1630 => x"2a",
          1631 => x"70",
          1632 => x"34",
          1633 => x"51",
          1634 => x"83",
          1635 => x"fe",
          1636 => x"75",
          1637 => x"51",
          1638 => x"93",
          1639 => x"81",
          1640 => x"73",
          1641 => x"55",
          1642 => x"51",
          1643 => x"84",
          1644 => x"fe",
          1645 => x"77",
          1646 => x"53",
          1647 => x"81",
          1648 => x"ff",
          1649 => x"f4",
          1650 => x"0d",
          1651 => x"0d",
          1652 => x"56",
          1653 => x"70",
          1654 => x"33",
          1655 => x"05",
          1656 => x"71",
          1657 => x"56",
          1658 => x"72",
          1659 => x"38",
          1660 => x"e2",
          1661 => x"d3",
          1662 => x"3d",
          1663 => x"3d",
          1664 => x"71",
          1665 => x"52",
          1666 => x"99",
          1667 => x"2e",
          1668 => x"12",
          1669 => x"52",
          1670 => x"89",
          1671 => x"2e",
          1672 => x"ee",
          1673 => x"81",
          1674 => x"84",
          1675 => x"80",
          1676 => x"ac",
          1677 => x"0b",
          1678 => x"0c",
          1679 => x"0d",
          1680 => x"0b",
          1681 => x"56",
          1682 => x"2e",
          1683 => x"81",
          1684 => x"08",
          1685 => x"70",
          1686 => x"33",
          1687 => x"de",
          1688 => x"ac",
          1689 => x"09",
          1690 => x"38",
          1691 => x"08",
          1692 => x"b0",
          1693 => x"17",
          1694 => x"74",
          1695 => x"27",
          1696 => x"16",
          1697 => x"82",
          1698 => x"06",
          1699 => x"54",
          1700 => x"9c",
          1701 => x"53",
          1702 => x"16",
          1703 => x"9e",
          1704 => x"81",
          1705 => x"d3",
          1706 => x"3d",
          1707 => x"3d",
          1708 => x"56",
          1709 => x"b0",
          1710 => x"2e",
          1711 => x"51",
          1712 => x"81",
          1713 => x"56",
          1714 => x"08",
          1715 => x"54",
          1716 => x"17",
          1717 => x"33",
          1718 => x"3f",
          1719 => x"08",
          1720 => x"38",
          1721 => x"56",
          1722 => x"0c",
          1723 => x"ac",
          1724 => x"0d",
          1725 => x"0d",
          1726 => x"57",
          1727 => x"81",
          1728 => x"58",
          1729 => x"08",
          1730 => x"76",
          1731 => x"83",
          1732 => x"06",
          1733 => x"84",
          1734 => x"78",
          1735 => x"81",
          1736 => x"38",
          1737 => x"81",
          1738 => x"52",
          1739 => x"52",
          1740 => x"3f",
          1741 => x"52",
          1742 => x"51",
          1743 => x"84",
          1744 => x"d2",
          1745 => x"fc",
          1746 => x"8a",
          1747 => x"52",
          1748 => x"51",
          1749 => x"90",
          1750 => x"84",
          1751 => x"fb",
          1752 => x"17",
          1753 => x"a0",
          1754 => x"f4",
          1755 => x"08",
          1756 => x"b0",
          1757 => x"55",
          1758 => x"81",
          1759 => x"f8",
          1760 => x"84",
          1761 => x"53",
          1762 => x"17",
          1763 => x"88",
          1764 => x"ac",
          1765 => x"83",
          1766 => x"77",
          1767 => x"0c",
          1768 => x"04",
          1769 => x"77",
          1770 => x"12",
          1771 => x"55",
          1772 => x"56",
          1773 => x"8d",
          1774 => x"22",
          1775 => x"ac",
          1776 => x"57",
          1777 => x"d3",
          1778 => x"3d",
          1779 => x"3d",
          1780 => x"70",
          1781 => x"55",
          1782 => x"88",
          1783 => x"08",
          1784 => x"38",
          1785 => x"d9",
          1786 => x"33",
          1787 => x"82",
          1788 => x"38",
          1789 => x"89",
          1790 => x"2e",
          1791 => x"bf",
          1792 => x"2e",
          1793 => x"81",
          1794 => x"81",
          1795 => x"89",
          1796 => x"08",
          1797 => x"52",
          1798 => x"3f",
          1799 => x"08",
          1800 => x"76",
          1801 => x"14",
          1802 => x"81",
          1803 => x"2a",
          1804 => x"05",
          1805 => x"59",
          1806 => x"f2",
          1807 => x"ac",
          1808 => x"38",
          1809 => x"06",
          1810 => x"33",
          1811 => x"7a",
          1812 => x"06",
          1813 => x"5a",
          1814 => x"53",
          1815 => x"38",
          1816 => x"06",
          1817 => x"39",
          1818 => x"a4",
          1819 => x"52",
          1820 => x"ba",
          1821 => x"ac",
          1822 => x"38",
          1823 => x"ff",
          1824 => x"b4",
          1825 => x"f8",
          1826 => x"ac",
          1827 => x"ff",
          1828 => x"39",
          1829 => x"a4",
          1830 => x"52",
          1831 => x"8e",
          1832 => x"ac",
          1833 => x"74",
          1834 => x"fc",
          1835 => x"b4",
          1836 => x"e5",
          1837 => x"ac",
          1838 => x"06",
          1839 => x"81",
          1840 => x"d3",
          1841 => x"3d",
          1842 => x"3d",
          1843 => x"7f",
          1844 => x"82",
          1845 => x"27",
          1846 => x"73",
          1847 => x"27",
          1848 => x"74",
          1849 => x"77",
          1850 => x"38",
          1851 => x"89",
          1852 => x"2e",
          1853 => x"91",
          1854 => x"2e",
          1855 => x"82",
          1856 => x"81",
          1857 => x"89",
          1858 => x"08",
          1859 => x"52",
          1860 => x"3f",
          1861 => x"08",
          1862 => x"ac",
          1863 => x"38",
          1864 => x"06",
          1865 => x"81",
          1866 => x"06",
          1867 => x"58",
          1868 => x"80",
          1869 => x"75",
          1870 => x"f0",
          1871 => x"8f",
          1872 => x"58",
          1873 => x"34",
          1874 => x"16",
          1875 => x"2a",
          1876 => x"05",
          1877 => x"fa",
          1878 => x"d3",
          1879 => x"81",
          1880 => x"81",
          1881 => x"83",
          1882 => x"b4",
          1883 => x"06",
          1884 => x"57",
          1885 => x"72",
          1886 => x"88",
          1887 => x"57",
          1888 => x"81",
          1889 => x"54",
          1890 => x"81",
          1891 => x"34",
          1892 => x"73",
          1893 => x"16",
          1894 => x"74",
          1895 => x"3f",
          1896 => x"08",
          1897 => x"ac",
          1898 => x"38",
          1899 => x"ff",
          1900 => x"14",
          1901 => x"75",
          1902 => x"51",
          1903 => x"81",
          1904 => x"34",
          1905 => x"73",
          1906 => x"16",
          1907 => x"74",
          1908 => x"3f",
          1909 => x"08",
          1910 => x"ac",
          1911 => x"75",
          1912 => x"74",
          1913 => x"fc",
          1914 => x"b4",
          1915 => x"51",
          1916 => x"a5",
          1917 => x"ac",
          1918 => x"06",
          1919 => x"72",
          1920 => x"3f",
          1921 => x"16",
          1922 => x"d3",
          1923 => x"3d",
          1924 => x"3d",
          1925 => x"7d",
          1926 => x"58",
          1927 => x"74",
          1928 => x"98",
          1929 => x"26",
          1930 => x"56",
          1931 => x"75",
          1932 => x"38",
          1933 => x"52",
          1934 => x"8e",
          1935 => x"ac",
          1936 => x"d3",
          1937 => x"f4",
          1938 => x"82",
          1939 => x"39",
          1940 => x"e8",
          1941 => x"ac",
          1942 => x"e0",
          1943 => x"76",
          1944 => x"3f",
          1945 => x"08",
          1946 => x"ac",
          1947 => x"80",
          1948 => x"d3",
          1949 => x"2e",
          1950 => x"d3",
          1951 => x"2e",
          1952 => x"53",
          1953 => x"51",
          1954 => x"81",
          1955 => x"c5",
          1956 => x"08",
          1957 => x"90",
          1958 => x"27",
          1959 => x"15",
          1960 => x"90",
          1961 => x"15",
          1962 => x"54",
          1963 => x"34",
          1964 => x"15",
          1965 => x"ff",
          1966 => x"56",
          1967 => x"ac",
          1968 => x"0d",
          1969 => x"0d",
          1970 => x"08",
          1971 => x"7a",
          1972 => x"19",
          1973 => x"80",
          1974 => x"98",
          1975 => x"26",
          1976 => x"58",
          1977 => x"52",
          1978 => x"e2",
          1979 => x"74",
          1980 => x"08",
          1981 => x"38",
          1982 => x"08",
          1983 => x"ac",
          1984 => x"82",
          1985 => x"d3",
          1986 => x"98",
          1987 => x"d3",
          1988 => x"82",
          1989 => x"58",
          1990 => x"19",
          1991 => x"82",
          1992 => x"57",
          1993 => x"09",
          1994 => x"db",
          1995 => x"57",
          1996 => x"77",
          1997 => x"82",
          1998 => x"7b",
          1999 => x"3f",
          2000 => x"08",
          2001 => x"81",
          2002 => x"81",
          2003 => x"06",
          2004 => x"d3",
          2005 => x"75",
          2006 => x"30",
          2007 => x"80",
          2008 => x"07",
          2009 => x"52",
          2010 => x"81",
          2011 => x"80",
          2012 => x"8c",
          2013 => x"81",
          2014 => x"38",
          2015 => x"08",
          2016 => x"75",
          2017 => x"76",
          2018 => x"77",
          2019 => x"57",
          2020 => x"77",
          2021 => x"82",
          2022 => x"26",
          2023 => x"76",
          2024 => x"f8",
          2025 => x"d3",
          2026 => x"81",
          2027 => x"80",
          2028 => x"80",
          2029 => x"ac",
          2030 => x"09",
          2031 => x"38",
          2032 => x"08",
          2033 => x"32",
          2034 => x"72",
          2035 => x"70",
          2036 => x"52",
          2037 => x"80",
          2038 => x"78",
          2039 => x"06",
          2040 => x"80",
          2041 => x"39",
          2042 => x"52",
          2043 => x"da",
          2044 => x"ac",
          2045 => x"ac",
          2046 => x"81",
          2047 => x"07",
          2048 => x"30",
          2049 => x"9f",
          2050 => x"52",
          2051 => x"56",
          2052 => x"8f",
          2053 => x"7a",
          2054 => x"f9",
          2055 => x"d3",
          2056 => x"75",
          2057 => x"8c",
          2058 => x"19",
          2059 => x"54",
          2060 => x"74",
          2061 => x"90",
          2062 => x"05",
          2063 => x"84",
          2064 => x"07",
          2065 => x"1a",
          2066 => x"ff",
          2067 => x"2e",
          2068 => x"39",
          2069 => x"39",
          2070 => x"39",
          2071 => x"55",
          2072 => x"ac",
          2073 => x"0d",
          2074 => x"0d",
          2075 => x"57",
          2076 => x"81",
          2077 => x"ac",
          2078 => x"38",
          2079 => x"51",
          2080 => x"81",
          2081 => x"81",
          2082 => x"b0",
          2083 => x"84",
          2084 => x"52",
          2085 => x"52",
          2086 => x"3f",
          2087 => x"58",
          2088 => x"39",
          2089 => x"8a",
          2090 => x"75",
          2091 => x"38",
          2092 => x"1a",
          2093 => x"81",
          2094 => x"ee",
          2095 => x"d3",
          2096 => x"2e",
          2097 => x"0b",
          2098 => x"56",
          2099 => x"2e",
          2100 => x"58",
          2101 => x"81",
          2102 => x"8b",
          2103 => x"f8",
          2104 => x"7c",
          2105 => x"56",
          2106 => x"80",
          2107 => x"38",
          2108 => x"53",
          2109 => x"86",
          2110 => x"81",
          2111 => x"90",
          2112 => x"17",
          2113 => x"aa",
          2114 => x"53",
          2115 => x"85",
          2116 => x"08",
          2117 => x"38",
          2118 => x"53",
          2119 => x"17",
          2120 => x"72",
          2121 => x"83",
          2122 => x"08",
          2123 => x"80",
          2124 => x"16",
          2125 => x"2b",
          2126 => x"75",
          2127 => x"73",
          2128 => x"f5",
          2129 => x"d3",
          2130 => x"81",
          2131 => x"ff",
          2132 => x"81",
          2133 => x"ac",
          2134 => x"38",
          2135 => x"81",
          2136 => x"26",
          2137 => x"58",
          2138 => x"74",
          2139 => x"74",
          2140 => x"38",
          2141 => x"51",
          2142 => x"81",
          2143 => x"98",
          2144 => x"94",
          2145 => x"58",
          2146 => x"80",
          2147 => x"85",
          2148 => x"97",
          2149 => x"2a",
          2150 => x"05",
          2151 => x"74",
          2152 => x"16",
          2153 => x"18",
          2154 => x"77",
          2155 => x"0c",
          2156 => x"04",
          2157 => x"79",
          2158 => x"90",
          2159 => x"05",
          2160 => x"55",
          2161 => x"76",
          2162 => x"80",
          2163 => x"0c",
          2164 => x"15",
          2165 => x"81",
          2166 => x"83",
          2167 => x"73",
          2168 => x"98",
          2169 => x"05",
          2170 => x"94",
          2171 => x"38",
          2172 => x"88",
          2173 => x"53",
          2174 => x"81",
          2175 => x"98",
          2176 => x"53",
          2177 => x"8a",
          2178 => x"11",
          2179 => x"06",
          2180 => x"81",
          2181 => x"15",
          2182 => x"51",
          2183 => x"81",
          2184 => x"54",
          2185 => x"0b",
          2186 => x"08",
          2187 => x"38",
          2188 => x"d3",
          2189 => x"2e",
          2190 => x"98",
          2191 => x"d3",
          2192 => x"80",
          2193 => x"8a",
          2194 => x"16",
          2195 => x"80",
          2196 => x"15",
          2197 => x"51",
          2198 => x"81",
          2199 => x"54",
          2200 => x"d3",
          2201 => x"2e",
          2202 => x"82",
          2203 => x"ac",
          2204 => x"bf",
          2205 => x"81",
          2206 => x"ff",
          2207 => x"81",
          2208 => x"52",
          2209 => x"e1",
          2210 => x"81",
          2211 => x"a3",
          2212 => x"16",
          2213 => x"76",
          2214 => x"3f",
          2215 => x"08",
          2216 => x"75",
          2217 => x"75",
          2218 => x"17",
          2219 => x"16",
          2220 => x"72",
          2221 => x"0c",
          2222 => x"04",
          2223 => x"7a",
          2224 => x"5a",
          2225 => x"52",
          2226 => x"93",
          2227 => x"ac",
          2228 => x"d3",
          2229 => x"e1",
          2230 => x"ac",
          2231 => x"16",
          2232 => x"51",
          2233 => x"81",
          2234 => x"54",
          2235 => x"08",
          2236 => x"81",
          2237 => x"9c",
          2238 => x"33",
          2239 => x"72",
          2240 => x"09",
          2241 => x"38",
          2242 => x"30",
          2243 => x"76",
          2244 => x"72",
          2245 => x"38",
          2246 => x"76",
          2247 => x"38",
          2248 => x"57",
          2249 => x"51",
          2250 => x"81",
          2251 => x"54",
          2252 => x"08",
          2253 => x"a6",
          2254 => x"2e",
          2255 => x"83",
          2256 => x"73",
          2257 => x"0c",
          2258 => x"04",
          2259 => x"76",
          2260 => x"54",
          2261 => x"81",
          2262 => x"83",
          2263 => x"76",
          2264 => x"53",
          2265 => x"2e",
          2266 => x"90",
          2267 => x"51",
          2268 => x"81",
          2269 => x"90",
          2270 => x"53",
          2271 => x"ac",
          2272 => x"0d",
          2273 => x"0d",
          2274 => x"83",
          2275 => x"54",
          2276 => x"55",
          2277 => x"3f",
          2278 => x"51",
          2279 => x"2e",
          2280 => x"8b",
          2281 => x"2a",
          2282 => x"51",
          2283 => x"86",
          2284 => x"f7",
          2285 => x"7d",
          2286 => x"76",
          2287 => x"98",
          2288 => x"2e",
          2289 => x"98",
          2290 => x"78",
          2291 => x"3f",
          2292 => x"08",
          2293 => x"ac",
          2294 => x"38",
          2295 => x"70",
          2296 => x"74",
          2297 => x"58",
          2298 => x"9c",
          2299 => x"11",
          2300 => x"06",
          2301 => x"06",
          2302 => x"53",
          2303 => x"34",
          2304 => x"32",
          2305 => x"ae",
          2306 => x"70",
          2307 => x"2a",
          2308 => x"51",
          2309 => x"2e",
          2310 => x"8f",
          2311 => x"80",
          2312 => x"54",
          2313 => x"2e",
          2314 => x"83",
          2315 => x"73",
          2316 => x"38",
          2317 => x"51",
          2318 => x"81",
          2319 => x"58",
          2320 => x"08",
          2321 => x"16",
          2322 => x"38",
          2323 => x"86",
          2324 => x"98",
          2325 => x"81",
          2326 => x"8b",
          2327 => x"f8",
          2328 => x"70",
          2329 => x"80",
          2330 => x"f8",
          2331 => x"d3",
          2332 => x"81",
          2333 => x"80",
          2334 => x"39",
          2335 => x"e6",
          2336 => x"08",
          2337 => x"ec",
          2338 => x"d3",
          2339 => x"81",
          2340 => x"80",
          2341 => x"16",
          2342 => x"51",
          2343 => x"2e",
          2344 => x"16",
          2345 => x"33",
          2346 => x"55",
          2347 => x"34",
          2348 => x"70",
          2349 => x"81",
          2350 => x"59",
          2351 => x"8b",
          2352 => x"52",
          2353 => x"85",
          2354 => x"ac",
          2355 => x"96",
          2356 => x"75",
          2357 => x"3f",
          2358 => x"08",
          2359 => x"ac",
          2360 => x"ff",
          2361 => x"54",
          2362 => x"ac",
          2363 => x"0d",
          2364 => x"0d",
          2365 => x"57",
          2366 => x"73",
          2367 => x"3f",
          2368 => x"08",
          2369 => x"ac",
          2370 => x"98",
          2371 => x"75",
          2372 => x"3f",
          2373 => x"08",
          2374 => x"ac",
          2375 => x"a0",
          2376 => x"ac",
          2377 => x"14",
          2378 => x"87",
          2379 => x"a0",
          2380 => x"14",
          2381 => x"d7",
          2382 => x"83",
          2383 => x"81",
          2384 => x"87",
          2385 => x"fc",
          2386 => x"70",
          2387 => x"08",
          2388 => x"56",
          2389 => x"3f",
          2390 => x"08",
          2391 => x"ac",
          2392 => x"9c",
          2393 => x"e5",
          2394 => x"0b",
          2395 => x"73",
          2396 => x"0c",
          2397 => x"04",
          2398 => x"78",
          2399 => x"80",
          2400 => x"34",
          2401 => x"80",
          2402 => x"38",
          2403 => x"55",
          2404 => x"14",
          2405 => x"16",
          2406 => x"72",
          2407 => x"38",
          2408 => x"09",
          2409 => x"38",
          2410 => x"73",
          2411 => x"81",
          2412 => x"75",
          2413 => x"52",
          2414 => x"13",
          2415 => x"55",
          2416 => x"05",
          2417 => x"13",
          2418 => x"55",
          2419 => x"c0",
          2420 => x"88",
          2421 => x"0b",
          2422 => x"9c",
          2423 => x"8b",
          2424 => x"17",
          2425 => x"08",
          2426 => x"e6",
          2427 => x"d3",
          2428 => x"0c",
          2429 => x"96",
          2430 => x"84",
          2431 => x"ac",
          2432 => x"23",
          2433 => x"98",
          2434 => x"f4",
          2435 => x"ac",
          2436 => x"23",
          2437 => x"04",
          2438 => x"7e",
          2439 => x"a0",
          2440 => x"5c",
          2441 => x"52",
          2442 => x"87",
          2443 => x"58",
          2444 => x"33",
          2445 => x"ae",
          2446 => x"06",
          2447 => x"78",
          2448 => x"81",
          2449 => x"32",
          2450 => x"9f",
          2451 => x"26",
          2452 => x"53",
          2453 => x"73",
          2454 => x"18",
          2455 => x"34",
          2456 => x"db",
          2457 => x"32",
          2458 => x"80",
          2459 => x"30",
          2460 => x"9f",
          2461 => x"56",
          2462 => x"80",
          2463 => x"86",
          2464 => x"26",
          2465 => x"76",
          2466 => x"a4",
          2467 => x"27",
          2468 => x"54",
          2469 => x"34",
          2470 => x"ce",
          2471 => x"70",
          2472 => x"59",
          2473 => x"76",
          2474 => x"38",
          2475 => x"70",
          2476 => x"dc",
          2477 => x"72",
          2478 => x"80",
          2479 => x"51",
          2480 => x"74",
          2481 => x"38",
          2482 => x"17",
          2483 => x"1a",
          2484 => x"55",
          2485 => x"2e",
          2486 => x"83",
          2487 => x"80",
          2488 => x"33",
          2489 => x"73",
          2490 => x"09",
          2491 => x"38",
          2492 => x"75",
          2493 => x"d2",
          2494 => x"39",
          2495 => x"70",
          2496 => x"25",
          2497 => x"07",
          2498 => x"73",
          2499 => x"38",
          2500 => x"70",
          2501 => x"32",
          2502 => x"80",
          2503 => x"2a",
          2504 => x"56",
          2505 => x"81",
          2506 => x"58",
          2507 => x"ed",
          2508 => x"2b",
          2509 => x"25",
          2510 => x"80",
          2511 => x"bb",
          2512 => x"57",
          2513 => x"e5",
          2514 => x"d3",
          2515 => x"2e",
          2516 => x"17",
          2517 => x"19",
          2518 => x"56",
          2519 => x"3f",
          2520 => x"08",
          2521 => x"38",
          2522 => x"73",
          2523 => x"38",
          2524 => x"f6",
          2525 => x"54",
          2526 => x"81",
          2527 => x"55",
          2528 => x"34",
          2529 => x"fe",
          2530 => x"52",
          2531 => x"51",
          2532 => x"81",
          2533 => x"80",
          2534 => x"9f",
          2535 => x"99",
          2536 => x"e0",
          2537 => x"ff",
          2538 => x"7a",
          2539 => x"74",
          2540 => x"58",
          2541 => x"76",
          2542 => x"86",
          2543 => x"2e",
          2544 => x"33",
          2545 => x"e5",
          2546 => x"06",
          2547 => x"7b",
          2548 => x"a0",
          2549 => x"38",
          2550 => x"54",
          2551 => x"54",
          2552 => x"54",
          2553 => x"34",
          2554 => x"81",
          2555 => x"8d",
          2556 => x"fa",
          2557 => x"70",
          2558 => x"80",
          2559 => x"51",
          2560 => x"af",
          2561 => x"81",
          2562 => x"70",
          2563 => x"54",
          2564 => x"2e",
          2565 => x"54",
          2566 => x"53",
          2567 => x"8c",
          2568 => x"08",
          2569 => x"b3",
          2570 => x"5a",
          2571 => x"33",
          2572 => x"72",
          2573 => x"81",
          2574 => x"81",
          2575 => x"70",
          2576 => x"54",
          2577 => x"2e",
          2578 => x"83",
          2579 => x"74",
          2580 => x"72",
          2581 => x"0b",
          2582 => x"79",
          2583 => x"53",
          2584 => x"9b",
          2585 => x"0b",
          2586 => x"80",
          2587 => x"f0",
          2588 => x"d3",
          2589 => x"81",
          2590 => x"55",
          2591 => x"89",
          2592 => x"52",
          2593 => x"90",
          2594 => x"ac",
          2595 => x"d3",
          2596 => x"8f",
          2597 => x"f7",
          2598 => x"d3",
          2599 => x"17",
          2600 => x"81",
          2601 => x"80",
          2602 => x"38",
          2603 => x"08",
          2604 => x"81",
          2605 => x"38",
          2606 => x"70",
          2607 => x"53",
          2608 => x"9a",
          2609 => x"2a",
          2610 => x"51",
          2611 => x"2e",
          2612 => x"ff",
          2613 => x"17",
          2614 => x"80",
          2615 => x"82",
          2616 => x"06",
          2617 => x"bb",
          2618 => x"b7",
          2619 => x"2a",
          2620 => x"51",
          2621 => x"38",
          2622 => x"70",
          2623 => x"81",
          2624 => x"54",
          2625 => x"fe",
          2626 => x"16",
          2627 => x"06",
          2628 => x"52",
          2629 => x"b4",
          2630 => x"ac",
          2631 => x"0c",
          2632 => x"74",
          2633 => x"0c",
          2634 => x"04",
          2635 => x"7c",
          2636 => x"08",
          2637 => x"59",
          2638 => x"80",
          2639 => x"38",
          2640 => x"05",
          2641 => x"ba",
          2642 => x"72",
          2643 => x"9f",
          2644 => x"51",
          2645 => x"e8",
          2646 => x"2e",
          2647 => x"81",
          2648 => x"33",
          2649 => x"52",
          2650 => x"92",
          2651 => x"72",
          2652 => x"d0",
          2653 => x"51",
          2654 => x"80",
          2655 => x"0b",
          2656 => x"5c",
          2657 => x"10",
          2658 => x"7a",
          2659 => x"51",
          2660 => x"05",
          2661 => x"70",
          2662 => x"33",
          2663 => x"53",
          2664 => x"99",
          2665 => x"e0",
          2666 => x"ff",
          2667 => x"ff",
          2668 => x"70",
          2669 => x"38",
          2670 => x"81",
          2671 => x"51",
          2672 => x"74",
          2673 => x"70",
          2674 => x"25",
          2675 => x"06",
          2676 => x"51",
          2677 => x"38",
          2678 => x"78",
          2679 => x"70",
          2680 => x"2a",
          2681 => x"07",
          2682 => x"51",
          2683 => x"8c",
          2684 => x"58",
          2685 => x"ff",
          2686 => x"39",
          2687 => x"86",
          2688 => x"7a",
          2689 => x"51",
          2690 => x"d3",
          2691 => x"70",
          2692 => x"0c",
          2693 => x"04",
          2694 => x"77",
          2695 => x"83",
          2696 => x"0b",
          2697 => x"78",
          2698 => x"e1",
          2699 => x"55",
          2700 => x"08",
          2701 => x"84",
          2702 => x"dd",
          2703 => x"d3",
          2704 => x"ff",
          2705 => x"83",
          2706 => x"d4",
          2707 => x"81",
          2708 => x"38",
          2709 => x"17",
          2710 => x"73",
          2711 => x"09",
          2712 => x"38",
          2713 => x"81",
          2714 => x"30",
          2715 => x"77",
          2716 => x"54",
          2717 => x"b4",
          2718 => x"73",
          2719 => x"09",
          2720 => x"38",
          2721 => x"ba",
          2722 => x"ea",
          2723 => x"bd",
          2724 => x"ac",
          2725 => x"d3",
          2726 => x"2e",
          2727 => x"53",
          2728 => x"52",
          2729 => x"51",
          2730 => x"81",
          2731 => x"55",
          2732 => x"08",
          2733 => x"38",
          2734 => x"81",
          2735 => x"87",
          2736 => x"f3",
          2737 => x"02",
          2738 => x"c7",
          2739 => x"54",
          2740 => x"7f",
          2741 => x"3f",
          2742 => x"08",
          2743 => x"80",
          2744 => x"ac",
          2745 => x"9e",
          2746 => x"ac",
          2747 => x"81",
          2748 => x"70",
          2749 => x"8c",
          2750 => x"2e",
          2751 => x"74",
          2752 => x"81",
          2753 => x"33",
          2754 => x"80",
          2755 => x"81",
          2756 => x"d6",
          2757 => x"d3",
          2758 => x"ff",
          2759 => x"06",
          2760 => x"99",
          2761 => x"2e",
          2762 => x"82",
          2763 => x"06",
          2764 => x"56",
          2765 => x"38",
          2766 => x"ca",
          2767 => x"34",
          2768 => x"34",
          2769 => x"15",
          2770 => x"8d",
          2771 => x"ac",
          2772 => x"06",
          2773 => x"54",
          2774 => x"72",
          2775 => x"76",
          2776 => x"38",
          2777 => x"70",
          2778 => x"53",
          2779 => x"86",
          2780 => x"70",
          2781 => x"5a",
          2782 => x"81",
          2783 => x"81",
          2784 => x"76",
          2785 => x"81",
          2786 => x"38",
          2787 => x"90",
          2788 => x"3d",
          2789 => x"05",
          2790 => x"f6",
          2791 => x"59",
          2792 => x"72",
          2793 => x"38",
          2794 => x"51",
          2795 => x"81",
          2796 => x"57",
          2797 => x"81",
          2798 => x"74",
          2799 => x"80",
          2800 => x"74",
          2801 => x"f0",
          2802 => x"53",
          2803 => x"80",
          2804 => x"79",
          2805 => x"fc",
          2806 => x"d3",
          2807 => x"ff",
          2808 => x"77",
          2809 => x"81",
          2810 => x"74",
          2811 => x"81",
          2812 => x"2e",
          2813 => x"8d",
          2814 => x"26",
          2815 => x"bf",
          2816 => x"fc",
          2817 => x"ac",
          2818 => x"ff",
          2819 => x"56",
          2820 => x"2e",
          2821 => x"84",
          2822 => x"ca",
          2823 => x"e0",
          2824 => x"ac",
          2825 => x"ff",
          2826 => x"8d",
          2827 => x"15",
          2828 => x"3f",
          2829 => x"08",
          2830 => x"16",
          2831 => x"15",
          2832 => x"34",
          2833 => x"33",
          2834 => x"8d",
          2835 => x"26",
          2836 => x"82",
          2837 => x"71",
          2838 => x"17",
          2839 => x"53",
          2840 => x"23",
          2841 => x"ff",
          2842 => x"80",
          2843 => x"ff",
          2844 => x"53",
          2845 => x"86",
          2846 => x"84",
          2847 => x"c5",
          2848 => x"fc",
          2849 => x"ac",
          2850 => x"23",
          2851 => x"08",
          2852 => x"06",
          2853 => x"8d",
          2854 => x"ea",
          2855 => x"15",
          2856 => x"3f",
          2857 => x"08",
          2858 => x"06",
          2859 => x"38",
          2860 => x"51",
          2861 => x"81",
          2862 => x"53",
          2863 => x"51",
          2864 => x"81",
          2865 => x"83",
          2866 => x"59",
          2867 => x"80",
          2868 => x"38",
          2869 => x"74",
          2870 => x"2a",
          2871 => x"8d",
          2872 => x"26",
          2873 => x"8a",
          2874 => x"72",
          2875 => x"ff",
          2876 => x"81",
          2877 => x"53",
          2878 => x"d3",
          2879 => x"2e",
          2880 => x"80",
          2881 => x"ac",
          2882 => x"ff",
          2883 => x"83",
          2884 => x"72",
          2885 => x"26",
          2886 => x"57",
          2887 => x"26",
          2888 => x"57",
          2889 => x"80",
          2890 => x"38",
          2891 => x"16",
          2892 => x"16",
          2893 => x"a4",
          2894 => x"1a",
          2895 => x"76",
          2896 => x"81",
          2897 => x"80",
          2898 => x"d7",
          2899 => x"d3",
          2900 => x"ff",
          2901 => x"8d",
          2902 => x"aa",
          2903 => x"22",
          2904 => x"72",
          2905 => x"80",
          2906 => x"d7",
          2907 => x"d3",
          2908 => x"16",
          2909 => x"08",
          2910 => x"b6",
          2911 => x"22",
          2912 => x"72",
          2913 => x"fe",
          2914 => x"08",
          2915 => x"0c",
          2916 => x"09",
          2917 => x"38",
          2918 => x"10",
          2919 => x"98",
          2920 => x"98",
          2921 => x"70",
          2922 => x"17",
          2923 => x"05",
          2924 => x"ff",
          2925 => x"53",
          2926 => x"9c",
          2927 => x"81",
          2928 => x"0b",
          2929 => x"ff",
          2930 => x"0c",
          2931 => x"84",
          2932 => x"83",
          2933 => x"06",
          2934 => x"80",
          2935 => x"d6",
          2936 => x"d3",
          2937 => x"ff",
          2938 => x"72",
          2939 => x"81",
          2940 => x"38",
          2941 => x"74",
          2942 => x"3f",
          2943 => x"08",
          2944 => x"81",
          2945 => x"84",
          2946 => x"b2",
          2947 => x"f0",
          2948 => x"ac",
          2949 => x"ff",
          2950 => x"82",
          2951 => x"09",
          2952 => x"c8",
          2953 => x"51",
          2954 => x"81",
          2955 => x"84",
          2956 => x"d2",
          2957 => x"06",
          2958 => x"98",
          2959 => x"d9",
          2960 => x"ac",
          2961 => x"85",
          2962 => x"09",
          2963 => x"38",
          2964 => x"51",
          2965 => x"81",
          2966 => x"90",
          2967 => x"a0",
          2968 => x"b5",
          2969 => x"ac",
          2970 => x"0c",
          2971 => x"81",
          2972 => x"81",
          2973 => x"81",
          2974 => x"72",
          2975 => x"80",
          2976 => x"0c",
          2977 => x"81",
          2978 => x"8f",
          2979 => x"fb",
          2980 => x"54",
          2981 => x"80",
          2982 => x"73",
          2983 => x"af",
          2984 => x"70",
          2985 => x"71",
          2986 => x"38",
          2987 => x"86",
          2988 => x"52",
          2989 => x"09",
          2990 => x"38",
          2991 => x"51",
          2992 => x"81",
          2993 => x"81",
          2994 => x"83",
          2995 => x"80",
          2996 => x"2e",
          2997 => x"84",
          2998 => x"53",
          2999 => x"0c",
          3000 => x"d3",
          3001 => x"3d",
          3002 => x"3d",
          3003 => x"05",
          3004 => x"89",
          3005 => x"52",
          3006 => x"3f",
          3007 => x"08",
          3008 => x"80",
          3009 => x"ac",
          3010 => x"c4",
          3011 => x"ac",
          3012 => x"81",
          3013 => x"70",
          3014 => x"73",
          3015 => x"38",
          3016 => x"78",
          3017 => x"38",
          3018 => x"74",
          3019 => x"10",
          3020 => x"05",
          3021 => x"54",
          3022 => x"80",
          3023 => x"80",
          3024 => x"70",
          3025 => x"51",
          3026 => x"81",
          3027 => x"54",
          3028 => x"ac",
          3029 => x"0d",
          3030 => x"0d",
          3031 => x"05",
          3032 => x"33",
          3033 => x"55",
          3034 => x"84",
          3035 => x"bf",
          3036 => x"98",
          3037 => x"53",
          3038 => x"05",
          3039 => x"c3",
          3040 => x"ac",
          3041 => x"d3",
          3042 => x"c5",
          3043 => x"68",
          3044 => x"d4",
          3045 => x"db",
          3046 => x"ac",
          3047 => x"d3",
          3048 => x"38",
          3049 => x"05",
          3050 => x"2b",
          3051 => x"80",
          3052 => x"86",
          3053 => x"06",
          3054 => x"2e",
          3055 => x"75",
          3056 => x"38",
          3057 => x"09",
          3058 => x"38",
          3059 => x"05",
          3060 => x"3f",
          3061 => x"08",
          3062 => x"07",
          3063 => x"02",
          3064 => x"91",
          3065 => x"80",
          3066 => x"87",
          3067 => x"76",
          3068 => x"81",
          3069 => x"74",
          3070 => x"38",
          3071 => x"83",
          3072 => x"83",
          3073 => x"06",
          3074 => x"80",
          3075 => x"38",
          3076 => x"51",
          3077 => x"81",
          3078 => x"59",
          3079 => x"0a",
          3080 => x"05",
          3081 => x"3f",
          3082 => x"0b",
          3083 => x"75",
          3084 => x"7a",
          3085 => x"3f",
          3086 => x"9c",
          3087 => x"a0",
          3088 => x"81",
          3089 => x"34",
          3090 => x"80",
          3091 => x"b0",
          3092 => x"55",
          3093 => x"3d",
          3094 => x"51",
          3095 => x"3f",
          3096 => x"08",
          3097 => x"ac",
          3098 => x"38",
          3099 => x"51",
          3100 => x"81",
          3101 => x"7b",
          3102 => x"12",
          3103 => x"b6",
          3104 => x"cd",
          3105 => x"05",
          3106 => x"2a",
          3107 => x"51",
          3108 => x"80",
          3109 => x"84",
          3110 => x"76",
          3111 => x"81",
          3112 => x"74",
          3113 => x"38",
          3114 => x"33",
          3115 => x"74",
          3116 => x"38",
          3117 => x"82",
          3118 => x"83",
          3119 => x"06",
          3120 => x"80",
          3121 => x"76",
          3122 => x"57",
          3123 => x"08",
          3124 => x"63",
          3125 => x"55",
          3126 => x"38",
          3127 => x"51",
          3128 => x"81",
          3129 => x"88",
          3130 => x"9c",
          3131 => x"a9",
          3132 => x"ac",
          3133 => x"0c",
          3134 => x"86",
          3135 => x"19",
          3136 => x"19",
          3137 => x"19",
          3138 => x"19",
          3139 => x"19",
          3140 => x"53",
          3141 => x"18",
          3142 => x"3f",
          3143 => x"70",
          3144 => x"55",
          3145 => x"81",
          3146 => x"18",
          3147 => x"81",
          3148 => x"18",
          3149 => x"0c",
          3150 => x"22",
          3151 => x"88",
          3152 => x"1c",
          3153 => x"5c",
          3154 => x"39",
          3155 => x"51",
          3156 => x"81",
          3157 => x"57",
          3158 => x"08",
          3159 => x"38",
          3160 => x"ff",
          3161 => x"06",
          3162 => x"56",
          3163 => x"59",
          3164 => x"77",
          3165 => x"70",
          3166 => x"06",
          3167 => x"74",
          3168 => x"98",
          3169 => x"80",
          3170 => x"83",
          3171 => x"74",
          3172 => x"38",
          3173 => x"51",
          3174 => x"81",
          3175 => x"85",
          3176 => x"a8",
          3177 => x"2a",
          3178 => x"08",
          3179 => x"1a",
          3180 => x"54",
          3181 => x"18",
          3182 => x"11",
          3183 => x"ca",
          3184 => x"d3",
          3185 => x"2e",
          3186 => x"56",
          3187 => x"84",
          3188 => x"0c",
          3189 => x"81",
          3190 => x"97",
          3191 => x"f3",
          3192 => x"62",
          3193 => x"5f",
          3194 => x"7d",
          3195 => x"fc",
          3196 => x"51",
          3197 => x"81",
          3198 => x"55",
          3199 => x"08",
          3200 => x"17",
          3201 => x"80",
          3202 => x"74",
          3203 => x"39",
          3204 => x"81",
          3205 => x"56",
          3206 => x"83",
          3207 => x"39",
          3208 => x"18",
          3209 => x"83",
          3210 => x"0b",
          3211 => x"81",
          3212 => x"39",
          3213 => x"18",
          3214 => x"83",
          3215 => x"0b",
          3216 => x"81",
          3217 => x"39",
          3218 => x"18",
          3219 => x"82",
          3220 => x"0b",
          3221 => x"81",
          3222 => x"39",
          3223 => x"94",
          3224 => x"55",
          3225 => x"83",
          3226 => x"78",
          3227 => x"cb",
          3228 => x"08",
          3229 => x"06",
          3230 => x"82",
          3231 => x"8a",
          3232 => x"05",
          3233 => x"06",
          3234 => x"a8",
          3235 => x"38",
          3236 => x"55",
          3237 => x"17",
          3238 => x"51",
          3239 => x"81",
          3240 => x"55",
          3241 => x"fe",
          3242 => x"ff",
          3243 => x"38",
          3244 => x"0c",
          3245 => x"52",
          3246 => x"e8",
          3247 => x"ac",
          3248 => x"fe",
          3249 => x"d3",
          3250 => x"79",
          3251 => x"58",
          3252 => x"80",
          3253 => x"1b",
          3254 => x"22",
          3255 => x"74",
          3256 => x"38",
          3257 => x"5a",
          3258 => x"53",
          3259 => x"81",
          3260 => x"55",
          3261 => x"81",
          3262 => x"fe",
          3263 => x"17",
          3264 => x"2b",
          3265 => x"80",
          3266 => x"9c",
          3267 => x"31",
          3268 => x"27",
          3269 => x"80",
          3270 => x"52",
          3271 => x"29",
          3272 => x"eb",
          3273 => x"2b",
          3274 => x"39",
          3275 => x"78",
          3276 => x"38",
          3277 => x"70",
          3278 => x"56",
          3279 => x"a5",
          3280 => x"9c",
          3281 => x"a8",
          3282 => x"81",
          3283 => x"55",
          3284 => x"81",
          3285 => x"fd",
          3286 => x"17",
          3287 => x"06",
          3288 => x"18",
          3289 => x"77",
          3290 => x"52",
          3291 => x"33",
          3292 => x"f1",
          3293 => x"ac",
          3294 => x"38",
          3295 => x"0c",
          3296 => x"83",
          3297 => x"80",
          3298 => x"55",
          3299 => x"83",
          3300 => x"75",
          3301 => x"08",
          3302 => x"17",
          3303 => x"7b",
          3304 => x"3f",
          3305 => x"7d",
          3306 => x"0c",
          3307 => x"19",
          3308 => x"1a",
          3309 => x"78",
          3310 => x"80",
          3311 => x"d3",
          3312 => x"3d",
          3313 => x"3d",
          3314 => x"64",
          3315 => x"5a",
          3316 => x"0c",
          3317 => x"05",
          3318 => x"f5",
          3319 => x"d3",
          3320 => x"81",
          3321 => x"8a",
          3322 => x"33",
          3323 => x"2e",
          3324 => x"56",
          3325 => x"90",
          3326 => x"81",
          3327 => x"06",
          3328 => x"87",
          3329 => x"2e",
          3330 => x"bd",
          3331 => x"91",
          3332 => x"56",
          3333 => x"81",
          3334 => x"34",
          3335 => x"d8",
          3336 => x"91",
          3337 => x"56",
          3338 => x"82",
          3339 => x"34",
          3340 => x"c4",
          3341 => x"91",
          3342 => x"56",
          3343 => x"81",
          3344 => x"34",
          3345 => x"b0",
          3346 => x"08",
          3347 => x"94",
          3348 => x"86",
          3349 => x"08",
          3350 => x"80",
          3351 => x"38",
          3352 => x"70",
          3353 => x"56",
          3354 => x"a8",
          3355 => x"11",
          3356 => x"77",
          3357 => x"5c",
          3358 => x"c6",
          3359 => x"38",
          3360 => x"55",
          3361 => x"7a",
          3362 => x"d4",
          3363 => x"d3",
          3364 => x"8f",
          3365 => x"08",
          3366 => x"d4",
          3367 => x"d3",
          3368 => x"74",
          3369 => x"c3",
          3370 => x"2e",
          3371 => x"74",
          3372 => x"e3",
          3373 => x"18",
          3374 => x"08",
          3375 => x"88",
          3376 => x"17",
          3377 => x"2b",
          3378 => x"80",
          3379 => x"81",
          3380 => x"08",
          3381 => x"52",
          3382 => x"33",
          3383 => x"de",
          3384 => x"ac",
          3385 => x"38",
          3386 => x"80",
          3387 => x"74",
          3388 => x"98",
          3389 => x"7d",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"a7",
          3393 => x"ac",
          3394 => x"89",
          3395 => x"79",
          3396 => x"d5",
          3397 => x"7e",
          3398 => x"51",
          3399 => x"76",
          3400 => x"74",
          3401 => x"79",
          3402 => x"7b",
          3403 => x"11",
          3404 => x"c5",
          3405 => x"d3",
          3406 => x"f9",
          3407 => x"08",
          3408 => x"74",
          3409 => x"38",
          3410 => x"74",
          3411 => x"1c",
          3412 => x"51",
          3413 => x"90",
          3414 => x"ff",
          3415 => x"90",
          3416 => x"89",
          3417 => x"db",
          3418 => x"08",
          3419 => x"38",
          3420 => x"8c",
          3421 => x"98",
          3422 => x"77",
          3423 => x"52",
          3424 => x"33",
          3425 => x"dd",
          3426 => x"ac",
          3427 => x"38",
          3428 => x"0c",
          3429 => x"83",
          3430 => x"80",
          3431 => x"55",
          3432 => x"83",
          3433 => x"75",
          3434 => x"94",
          3435 => x"ff",
          3436 => x"05",
          3437 => x"3f",
          3438 => x"ff",
          3439 => x"74",
          3440 => x"78",
          3441 => x"08",
          3442 => x"76",
          3443 => x"08",
          3444 => x"1b",
          3445 => x"08",
          3446 => x"59",
          3447 => x"83",
          3448 => x"74",
          3449 => x"78",
          3450 => x"90",
          3451 => x"c0",
          3452 => x"90",
          3453 => x"56",
          3454 => x"ac",
          3455 => x"0d",
          3456 => x"0d",
          3457 => x"fc",
          3458 => x"52",
          3459 => x"3f",
          3460 => x"08",
          3461 => x"ac",
          3462 => x"38",
          3463 => x"70",
          3464 => x"81",
          3465 => x"56",
          3466 => x"81",
          3467 => x"98",
          3468 => x"80",
          3469 => x"81",
          3470 => x"08",
          3471 => x"52",
          3472 => x"33",
          3473 => x"f6",
          3474 => x"81",
          3475 => x"80",
          3476 => x"18",
          3477 => x"06",
          3478 => x"19",
          3479 => x"08",
          3480 => x"c8",
          3481 => x"d3",
          3482 => x"81",
          3483 => x"80",
          3484 => x"18",
          3485 => x"33",
          3486 => x"56",
          3487 => x"34",
          3488 => x"53",
          3489 => x"08",
          3490 => x"3f",
          3491 => x"52",
          3492 => x"c5",
          3493 => x"88",
          3494 => x"96",
          3495 => x"c0",
          3496 => x"92",
          3497 => x"9a",
          3498 => x"81",
          3499 => x"34",
          3500 => x"c1",
          3501 => x"ac",
          3502 => x"33",
          3503 => x"56",
          3504 => x"19",
          3505 => x"74",
          3506 => x"0c",
          3507 => x"04",
          3508 => x"76",
          3509 => x"fe",
          3510 => x"d3",
          3511 => x"81",
          3512 => x"9c",
          3513 => x"fc",
          3514 => x"51",
          3515 => x"81",
          3516 => x"53",
          3517 => x"08",
          3518 => x"d3",
          3519 => x"0c",
          3520 => x"ac",
          3521 => x"0d",
          3522 => x"0d",
          3523 => x"e4",
          3524 => x"53",
          3525 => x"d3",
          3526 => x"8b",
          3527 => x"ac",
          3528 => x"dc",
          3529 => x"72",
          3530 => x"0c",
          3531 => x"04",
          3532 => x"80",
          3533 => x"d0",
          3534 => x"3d",
          3535 => x"3f",
          3536 => x"08",
          3537 => x"ac",
          3538 => x"38",
          3539 => x"52",
          3540 => x"05",
          3541 => x"3f",
          3542 => x"08",
          3543 => x"ac",
          3544 => x"02",
          3545 => x"33",
          3546 => x"55",
          3547 => x"25",
          3548 => x"7a",
          3549 => x"54",
          3550 => x"a2",
          3551 => x"84",
          3552 => x"06",
          3553 => x"73",
          3554 => x"38",
          3555 => x"70",
          3556 => x"b8",
          3557 => x"ac",
          3558 => x"0c",
          3559 => x"55",
          3560 => x"09",
          3561 => x"38",
          3562 => x"81",
          3563 => x"93",
          3564 => x"e1",
          3565 => x"3d",
          3566 => x"08",
          3567 => x"7a",
          3568 => x"a1",
          3569 => x"05",
          3570 => x"51",
          3571 => x"81",
          3572 => x"57",
          3573 => x"08",
          3574 => x"7e",
          3575 => x"94",
          3576 => x"55",
          3577 => x"74",
          3578 => x"f9",
          3579 => x"70",
          3580 => x"5e",
          3581 => x"7a",
          3582 => x"3f",
          3583 => x"08",
          3584 => x"ac",
          3585 => x"38",
          3586 => x"51",
          3587 => x"81",
          3588 => x"57",
          3589 => x"08",
          3590 => x"6c",
          3591 => x"d6",
          3592 => x"d3",
          3593 => x"76",
          3594 => x"d1",
          3595 => x"d3",
          3596 => x"81",
          3597 => x"81",
          3598 => x"54",
          3599 => x"51",
          3600 => x"81",
          3601 => x"57",
          3602 => x"08",
          3603 => x"52",
          3604 => x"f8",
          3605 => x"ac",
          3606 => x"95",
          3607 => x"73",
          3608 => x"3f",
          3609 => x"08",
          3610 => x"ac",
          3611 => x"cc",
          3612 => x"2e",
          3613 => x"83",
          3614 => x"76",
          3615 => x"a1",
          3616 => x"11",
          3617 => x"51",
          3618 => x"76",
          3619 => x"79",
          3620 => x"33",
          3621 => x"55",
          3622 => x"2e",
          3623 => x"16",
          3624 => x"11",
          3625 => x"56",
          3626 => x"81",
          3627 => x"74",
          3628 => x"91",
          3629 => x"75",
          3630 => x"38",
          3631 => x"19",
          3632 => x"11",
          3633 => x"1b",
          3634 => x"59",
          3635 => x"75",
          3636 => x"38",
          3637 => x"3d",
          3638 => x"59",
          3639 => x"67",
          3640 => x"91",
          3641 => x"85",
          3642 => x"2e",
          3643 => x"8c",
          3644 => x"a3",
          3645 => x"55",
          3646 => x"34",
          3647 => x"d3",
          3648 => x"10",
          3649 => x"cc",
          3650 => x"70",
          3651 => x"57",
          3652 => x"73",
          3653 => x"38",
          3654 => x"16",
          3655 => x"55",
          3656 => x"38",
          3657 => x"73",
          3658 => x"38",
          3659 => x"76",
          3660 => x"77",
          3661 => x"33",
          3662 => x"05",
          3663 => x"18",
          3664 => x"26",
          3665 => x"7a",
          3666 => x"5c",
          3667 => x"58",
          3668 => x"91",
          3669 => x"38",
          3670 => x"19",
          3671 => x"54",
          3672 => x"70",
          3673 => x"34",
          3674 => x"ec",
          3675 => x"34",
          3676 => x"ac",
          3677 => x"0d",
          3678 => x"0d",
          3679 => x"3d",
          3680 => x"71",
          3681 => x"ea",
          3682 => x"d3",
          3683 => x"81",
          3684 => x"8a",
          3685 => x"33",
          3686 => x"2e",
          3687 => x"55",
          3688 => x"8c",
          3689 => x"27",
          3690 => x"17",
          3691 => x"2a",
          3692 => x"51",
          3693 => x"85",
          3694 => x"08",
          3695 => x"08",
          3696 => x"94",
          3697 => x"77",
          3698 => x"b3",
          3699 => x"11",
          3700 => x"2b",
          3701 => x"75",
          3702 => x"38",
          3703 => x"18",
          3704 => x"b9",
          3705 => x"ac",
          3706 => x"7a",
          3707 => x"57",
          3708 => x"a9",
          3709 => x"ac",
          3710 => x"95",
          3711 => x"76",
          3712 => x"0c",
          3713 => x"08",
          3714 => x"08",
          3715 => x"c9",
          3716 => x"08",
          3717 => x"38",
          3718 => x"51",
          3719 => x"81",
          3720 => x"56",
          3721 => x"08",
          3722 => x"81",
          3723 => x"82",
          3724 => x"34",
          3725 => x"e3",
          3726 => x"ac",
          3727 => x"09",
          3728 => x"38",
          3729 => x"18",
          3730 => x"82",
          3731 => x"d3",
          3732 => x"18",
          3733 => x"18",
          3734 => x"2e",
          3735 => x"78",
          3736 => x"ea",
          3737 => x"31",
          3738 => x"1a",
          3739 => x"90",
          3740 => x"81",
          3741 => x"06",
          3742 => x"58",
          3743 => x"9a",
          3744 => x"76",
          3745 => x"3f",
          3746 => x"08",
          3747 => x"ac",
          3748 => x"81",
          3749 => x"58",
          3750 => x"52",
          3751 => x"ae",
          3752 => x"ac",
          3753 => x"ff",
          3754 => x"38",
          3755 => x"8a",
          3756 => x"98",
          3757 => x"26",
          3758 => x"0b",
          3759 => x"82",
          3760 => x"39",
          3761 => x"0c",
          3762 => x"ff",
          3763 => x"17",
          3764 => x"18",
          3765 => x"ff",
          3766 => x"80",
          3767 => x"75",
          3768 => x"c1",
          3769 => x"d3",
          3770 => x"38",
          3771 => x"18",
          3772 => x"81",
          3773 => x"89",
          3774 => x"ac",
          3775 => x"8c",
          3776 => x"18",
          3777 => x"38",
          3778 => x"8c",
          3779 => x"17",
          3780 => x"07",
          3781 => x"18",
          3782 => x"08",
          3783 => x"55",
          3784 => x"80",
          3785 => x"17",
          3786 => x"80",
          3787 => x"17",
          3788 => x"2b",
          3789 => x"80",
          3790 => x"81",
          3791 => x"08",
          3792 => x"52",
          3793 => x"33",
          3794 => x"b8",
          3795 => x"d3",
          3796 => x"2e",
          3797 => x"0b",
          3798 => x"81",
          3799 => x"90",
          3800 => x"ff",
          3801 => x"90",
          3802 => x"54",
          3803 => x"17",
          3804 => x"11",
          3805 => x"ff",
          3806 => x"81",
          3807 => x"80",
          3808 => x"81",
          3809 => x"34",
          3810 => x"39",
          3811 => x"18",
          3812 => x"87",
          3813 => x"18",
          3814 => x"74",
          3815 => x"0c",
          3816 => x"04",
          3817 => x"79",
          3818 => x"75",
          3819 => x"8f",
          3820 => x"89",
          3821 => x"52",
          3822 => x"05",
          3823 => x"3f",
          3824 => x"08",
          3825 => x"ac",
          3826 => x"38",
          3827 => x"7a",
          3828 => x"d8",
          3829 => x"d3",
          3830 => x"81",
          3831 => x"80",
          3832 => x"16",
          3833 => x"2b",
          3834 => x"74",
          3835 => x"86",
          3836 => x"84",
          3837 => x"06",
          3838 => x"73",
          3839 => x"38",
          3840 => x"52",
          3841 => x"c4",
          3842 => x"ac",
          3843 => x"0c",
          3844 => x"55",
          3845 => x"77",
          3846 => x"22",
          3847 => x"74",
          3848 => x"c9",
          3849 => x"d3",
          3850 => x"74",
          3851 => x"81",
          3852 => x"85",
          3853 => x"2e",
          3854 => x"76",
          3855 => x"73",
          3856 => x"0c",
          3857 => x"04",
          3858 => x"76",
          3859 => x"05",
          3860 => x"54",
          3861 => x"81",
          3862 => x"53",
          3863 => x"08",
          3864 => x"d3",
          3865 => x"0c",
          3866 => x"ac",
          3867 => x"0d",
          3868 => x"0d",
          3869 => x"3d",
          3870 => x"71",
          3871 => x"e4",
          3872 => x"d3",
          3873 => x"81",
          3874 => x"80",
          3875 => x"92",
          3876 => x"ac",
          3877 => x"51",
          3878 => x"81",
          3879 => x"53",
          3880 => x"52",
          3881 => x"8b",
          3882 => x"ac",
          3883 => x"d3",
          3884 => x"2e",
          3885 => x"83",
          3886 => x"72",
          3887 => x"52",
          3888 => x"b4",
          3889 => x"73",
          3890 => x"3f",
          3891 => x"08",
          3892 => x"ac",
          3893 => x"09",
          3894 => x"38",
          3895 => x"81",
          3896 => x"87",
          3897 => x"ef",
          3898 => x"56",
          3899 => x"3d",
          3900 => x"3d",
          3901 => x"cb",
          3902 => x"ac",
          3903 => x"d3",
          3904 => x"38",
          3905 => x"51",
          3906 => x"81",
          3907 => x"55",
          3908 => x"08",
          3909 => x"80",
          3910 => x"70",
          3911 => x"57",
          3912 => x"85",
          3913 => x"90",
          3914 => x"2e",
          3915 => x"52",
          3916 => x"05",
          3917 => x"3f",
          3918 => x"ac",
          3919 => x"0d",
          3920 => x"0d",
          3921 => x"5a",
          3922 => x"3d",
          3923 => x"91",
          3924 => x"ef",
          3925 => x"ac",
          3926 => x"d3",
          3927 => x"84",
          3928 => x"0c",
          3929 => x"11",
          3930 => x"55",
          3931 => x"08",
          3932 => x"38",
          3933 => x"7a",
          3934 => x"39",
          3935 => x"cf",
          3936 => x"81",
          3937 => x"7b",
          3938 => x"56",
          3939 => x"2e",
          3940 => x"80",
          3941 => x"75",
          3942 => x"52",
          3943 => x"05",
          3944 => x"aa",
          3945 => x"ac",
          3946 => x"d0",
          3947 => x"ac",
          3948 => x"cd",
          3949 => x"ac",
          3950 => x"81",
          3951 => x"07",
          3952 => x"05",
          3953 => x"53",
          3954 => x"98",
          3955 => x"26",
          3956 => x"fb",
          3957 => x"11",
          3958 => x"08",
          3959 => x"80",
          3960 => x"38",
          3961 => x"18",
          3962 => x"ff",
          3963 => x"81",
          3964 => x"59",
          3965 => x"08",
          3966 => x"7a",
          3967 => x"54",
          3968 => x"09",
          3969 => x"38",
          3970 => x"05",
          3971 => x"f0",
          3972 => x"ac",
          3973 => x"ff",
          3974 => x"70",
          3975 => x"82",
          3976 => x"51",
          3977 => x"7a",
          3978 => x"51",
          3979 => x"3f",
          3980 => x"08",
          3981 => x"70",
          3982 => x"25",
          3983 => x"58",
          3984 => x"74",
          3985 => x"ff",
          3986 => x"75",
          3987 => x"76",
          3988 => x"77",
          3989 => x"54",
          3990 => x"33",
          3991 => x"55",
          3992 => x"34",
          3993 => x"ac",
          3994 => x"0d",
          3995 => x"0d",
          3996 => x"fc",
          3997 => x"52",
          3998 => x"3f",
          3999 => x"08",
          4000 => x"ac",
          4001 => x"91",
          4002 => x"76",
          4003 => x"38",
          4004 => x"dc",
          4005 => x"33",
          4006 => x"70",
          4007 => x"56",
          4008 => x"74",
          4009 => x"c8",
          4010 => x"08",
          4011 => x"27",
          4012 => x"94",
          4013 => x"38",
          4014 => x"18",
          4015 => x"51",
          4016 => x"3f",
          4017 => x"08",
          4018 => x"88",
          4019 => x"ca",
          4020 => x"08",
          4021 => x"ff",
          4022 => x"81",
          4023 => x"81",
          4024 => x"ff",
          4025 => x"70",
          4026 => x"25",
          4027 => x"56",
          4028 => x"08",
          4029 => x"81",
          4030 => x"82",
          4031 => x"38",
          4032 => x"98",
          4033 => x"92",
          4034 => x"08",
          4035 => x"77",
          4036 => x"fe",
          4037 => x"ac",
          4038 => x"18",
          4039 => x"0c",
          4040 => x"80",
          4041 => x"74",
          4042 => x"76",
          4043 => x"98",
          4044 => x"80",
          4045 => x"81",
          4046 => x"08",
          4047 => x"52",
          4048 => x"33",
          4049 => x"b0",
          4050 => x"d3",
          4051 => x"2e",
          4052 => x"57",
          4053 => x"18",
          4054 => x"06",
          4055 => x"19",
          4056 => x"2e",
          4057 => x"91",
          4058 => x"56",
          4059 => x"56",
          4060 => x"ac",
          4061 => x"0d",
          4062 => x"0d",
          4063 => x"51",
          4064 => x"3f",
          4065 => x"3d",
          4066 => x"52",
          4067 => x"d6",
          4068 => x"d3",
          4069 => x"81",
          4070 => x"82",
          4071 => x"ba",
          4072 => x"96",
          4073 => x"44",
          4074 => x"3d",
          4075 => x"d0",
          4076 => x"d3",
          4077 => x"ba",
          4078 => x"ff",
          4079 => x"75",
          4080 => x"02",
          4081 => x"33",
          4082 => x"70",
          4083 => x"55",
          4084 => x"2e",
          4085 => x"56",
          4086 => x"38",
          4087 => x"51",
          4088 => x"3f",
          4089 => x"05",
          4090 => x"2b",
          4091 => x"80",
          4092 => x"86",
          4093 => x"02",
          4094 => x"33",
          4095 => x"73",
          4096 => x"38",
          4097 => x"81",
          4098 => x"52",
          4099 => x"bc",
          4100 => x"ac",
          4101 => x"05",
          4102 => x"33",
          4103 => x"70",
          4104 => x"56",
          4105 => x"80",
          4106 => x"38",
          4107 => x"51",
          4108 => x"3f",
          4109 => x"56",
          4110 => x"77",
          4111 => x"38",
          4112 => x"51",
          4113 => x"3f",
          4114 => x"5b",
          4115 => x"51",
          4116 => x"3f",
          4117 => x"3d",
          4118 => x"c1",
          4119 => x"d3",
          4120 => x"81",
          4121 => x"81",
          4122 => x"d3",
          4123 => x"73",
          4124 => x"3f",
          4125 => x"08",
          4126 => x"ac",
          4127 => x"87",
          4128 => x"32",
          4129 => x"72",
          4130 => x"78",
          4131 => x"54",
          4132 => x"38",
          4133 => x"51",
          4134 => x"3f",
          4135 => x"05",
          4136 => x"3f",
          4137 => x"08",
          4138 => x"08",
          4139 => x"d3",
          4140 => x"80",
          4141 => x"70",
          4142 => x"2a",
          4143 => x"57",
          4144 => x"74",
          4145 => x"38",
          4146 => x"51",
          4147 => x"3f",
          4148 => x"52",
          4149 => x"05",
          4150 => x"b6",
          4151 => x"ac",
          4152 => x"8c",
          4153 => x"ff",
          4154 => x"81",
          4155 => x"56",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"ac",
          4159 => x"0d",
          4160 => x"0d",
          4161 => x"3d",
          4162 => x"99",
          4163 => x"b3",
          4164 => x"ac",
          4165 => x"d3",
          4166 => x"b5",
          4167 => x"68",
          4168 => x"d4",
          4169 => x"cb",
          4170 => x"ac",
          4171 => x"d3",
          4172 => x"38",
          4173 => x"84",
          4174 => x"06",
          4175 => x"02",
          4176 => x"33",
          4177 => x"70",
          4178 => x"55",
          4179 => x"2e",
          4180 => x"55",
          4181 => x"09",
          4182 => x"f5",
          4183 => x"80",
          4184 => x"c4",
          4185 => x"ba",
          4186 => x"d3",
          4187 => x"80",
          4188 => x"ac",
          4189 => x"09",
          4190 => x"38",
          4191 => x"81",
          4192 => x"06",
          4193 => x"55",
          4194 => x"09",
          4195 => x"38",
          4196 => x"88",
          4197 => x"74",
          4198 => x"75",
          4199 => x"ff",
          4200 => x"81",
          4201 => x"55",
          4202 => x"08",
          4203 => x"8b",
          4204 => x"b4",
          4205 => x"af",
          4206 => x"54",
          4207 => x"15",
          4208 => x"90",
          4209 => x"34",
          4210 => x"ca",
          4211 => x"af",
          4212 => x"53",
          4213 => x"77",
          4214 => x"3f",
          4215 => x"18",
          4216 => x"18",
          4217 => x"a7",
          4218 => x"ae",
          4219 => x"15",
          4220 => x"80",
          4221 => x"77",
          4222 => x"3f",
          4223 => x"0b",
          4224 => x"98",
          4225 => x"51",
          4226 => x"81",
          4227 => x"55",
          4228 => x"08",
          4229 => x"52",
          4230 => x"51",
          4231 => x"3f",
          4232 => x"52",
          4233 => x"dd",
          4234 => x"90",
          4235 => x"34",
          4236 => x"0b",
          4237 => x"77",
          4238 => x"b9",
          4239 => x"ac",
          4240 => x"39",
          4241 => x"52",
          4242 => x"05",
          4243 => x"c2",
          4244 => x"d3",
          4245 => x"3d",
          4246 => x"3d",
          4247 => x"84",
          4248 => x"c8",
          4249 => x"a7",
          4250 => x"05",
          4251 => x"51",
          4252 => x"81",
          4253 => x"55",
          4254 => x"08",
          4255 => x"77",
          4256 => x"08",
          4257 => x"d4",
          4258 => x"e7",
          4259 => x"ac",
          4260 => x"d3",
          4261 => x"bd",
          4262 => x"97",
          4263 => x"a0",
          4264 => x"80",
          4265 => x"86",
          4266 => x"a9",
          4267 => x"a3",
          4268 => x"a7",
          4269 => x"05",
          4270 => x"d3",
          4271 => x"a7",
          4272 => x"52",
          4273 => x"52",
          4274 => x"c3",
          4275 => x"08",
          4276 => x"ca",
          4277 => x"d3",
          4278 => x"81",
          4279 => x"94",
          4280 => x"2e",
          4281 => x"8a",
          4282 => x"64",
          4283 => x"2e",
          4284 => x"55",
          4285 => x"09",
          4286 => x"b8",
          4287 => x"ff",
          4288 => x"c3",
          4289 => x"d3",
          4290 => x"81",
          4291 => x"81",
          4292 => x"56",
          4293 => x"3d",
          4294 => x"52",
          4295 => x"ff",
          4296 => x"02",
          4297 => x"8b",
          4298 => x"16",
          4299 => x"2a",
          4300 => x"51",
          4301 => x"89",
          4302 => x"07",
          4303 => x"17",
          4304 => x"81",
          4305 => x"34",
          4306 => x"70",
          4307 => x"81",
          4308 => x"57",
          4309 => x"80",
          4310 => x"63",
          4311 => x"38",
          4312 => x"51",
          4313 => x"3f",
          4314 => x"08",
          4315 => x"ff",
          4316 => x"82",
          4317 => x"ac",
          4318 => x"b8",
          4319 => x"ac",
          4320 => x"51",
          4321 => x"3f",
          4322 => x"08",
          4323 => x"57",
          4324 => x"ac",
          4325 => x"81",
          4326 => x"73",
          4327 => x"81",
          4328 => x"62",
          4329 => x"77",
          4330 => x"d9",
          4331 => x"81",
          4332 => x"34",
          4333 => x"a7",
          4334 => x"51",
          4335 => x"81",
          4336 => x"55",
          4337 => x"08",
          4338 => x"51",
          4339 => x"3f",
          4340 => x"08",
          4341 => x"d3",
          4342 => x"3d",
          4343 => x"3d",
          4344 => x"db",
          4345 => x"84",
          4346 => x"05",
          4347 => x"82",
          4348 => x"d0",
          4349 => x"3d",
          4350 => x"3f",
          4351 => x"08",
          4352 => x"ac",
          4353 => x"38",
          4354 => x"52",
          4355 => x"05",
          4356 => x"3f",
          4357 => x"08",
          4358 => x"ac",
          4359 => x"02",
          4360 => x"33",
          4361 => x"54",
          4362 => x"83",
          4363 => x"74",
          4364 => x"a7",
          4365 => x"09",
          4366 => x"71",
          4367 => x"06",
          4368 => x"55",
          4369 => x"15",
          4370 => x"81",
          4371 => x"34",
          4372 => x"ad",
          4373 => x"d3",
          4374 => x"74",
          4375 => x"0c",
          4376 => x"04",
          4377 => x"65",
          4378 => x"94",
          4379 => x"52",
          4380 => x"cc",
          4381 => x"d3",
          4382 => x"81",
          4383 => x"80",
          4384 => x"59",
          4385 => x"3d",
          4386 => x"c6",
          4387 => x"d3",
          4388 => x"81",
          4389 => x"bc",
          4390 => x"cb",
          4391 => x"a0",
          4392 => x"80",
          4393 => x"86",
          4394 => x"38",
          4395 => x"84",
          4396 => x"90",
          4397 => x"54",
          4398 => x"96",
          4399 => x"a9",
          4400 => x"54",
          4401 => x"15",
          4402 => x"ff",
          4403 => x"81",
          4404 => x"55",
          4405 => x"ac",
          4406 => x"0d",
          4407 => x"0d",
          4408 => x"59",
          4409 => x"3d",
          4410 => x"99",
          4411 => x"d3",
          4412 => x"ac",
          4413 => x"ac",
          4414 => x"81",
          4415 => x"07",
          4416 => x"30",
          4417 => x"9f",
          4418 => x"52",
          4419 => x"56",
          4420 => x"80",
          4421 => x"5d",
          4422 => x"52",
          4423 => x"52",
          4424 => x"bb",
          4425 => x"ac",
          4426 => x"d3",
          4427 => x"ce",
          4428 => x"73",
          4429 => x"fb",
          4430 => x"ac",
          4431 => x"d3",
          4432 => x"38",
          4433 => x"08",
          4434 => x"08",
          4435 => x"58",
          4436 => x"18",
          4437 => x"58",
          4438 => x"74",
          4439 => x"58",
          4440 => x"ec",
          4441 => x"54",
          4442 => x"77",
          4443 => x"38",
          4444 => x"11",
          4445 => x"55",
          4446 => x"2e",
          4447 => x"84",
          4448 => x"06",
          4449 => x"79",
          4450 => x"75",
          4451 => x"07",
          4452 => x"30",
          4453 => x"9f",
          4454 => x"52",
          4455 => x"74",
          4456 => x"38",
          4457 => x"08",
          4458 => x"aa",
          4459 => x"d3",
          4460 => x"81",
          4461 => x"a7",
          4462 => x"33",
          4463 => x"c3",
          4464 => x"2e",
          4465 => x"e4",
          4466 => x"2e",
          4467 => x"58",
          4468 => x"05",
          4469 => x"c1",
          4470 => x"ac",
          4471 => x"75",
          4472 => x"0c",
          4473 => x"04",
          4474 => x"82",
          4475 => x"ff",
          4476 => x"9b",
          4477 => x"cb",
          4478 => x"ac",
          4479 => x"d3",
          4480 => x"c8",
          4481 => x"a0",
          4482 => x"ff",
          4483 => x"ff",
          4484 => x"80",
          4485 => x"33",
          4486 => x"57",
          4487 => x"81",
          4488 => x"33",
          4489 => x"4c",
          4490 => x"06",
          4491 => x"a7",
          4492 => x"d3",
          4493 => x"2e",
          4494 => x"70",
          4495 => x"51",
          4496 => x"f2",
          4497 => x"ac",
          4498 => x"8d",
          4499 => x"2b",
          4500 => x"81",
          4501 => x"83",
          4502 => x"ff",
          4503 => x"73",
          4504 => x"38",
          4505 => x"83",
          4506 => x"57",
          4507 => x"76",
          4508 => x"81",
          4509 => x"33",
          4510 => x"2e",
          4511 => x"52",
          4512 => x"51",
          4513 => x"3f",
          4514 => x"08",
          4515 => x"ff",
          4516 => x"38",
          4517 => x"88",
          4518 => x"8a",
          4519 => x"38",
          4520 => x"a8",
          4521 => x"76",
          4522 => x"9a",
          4523 => x"ff",
          4524 => x"88",
          4525 => x"73",
          4526 => x"17",
          4527 => x"77",
          4528 => x"05",
          4529 => x"34",
          4530 => x"70",
          4531 => x"57",
          4532 => x"fe",
          4533 => x"3d",
          4534 => x"55",
          4535 => x"2e",
          4536 => x"76",
          4537 => x"38",
          4538 => x"70",
          4539 => x"33",
          4540 => x"54",
          4541 => x"09",
          4542 => x"38",
          4543 => x"76",
          4544 => x"38",
          4545 => x"33",
          4546 => x"a0",
          4547 => x"77",
          4548 => x"80",
          4549 => x"70",
          4550 => x"b3",
          4551 => x"d3",
          4552 => x"81",
          4553 => x"81",
          4554 => x"52",
          4555 => x"b9",
          4556 => x"d3",
          4557 => x"81",
          4558 => x"b0",
          4559 => x"2e",
          4560 => x"53",
          4561 => x"bc",
          4562 => x"51",
          4563 => x"3f",
          4564 => x"54",
          4565 => x"77",
          4566 => x"83",
          4567 => x"51",
          4568 => x"3f",
          4569 => x"08",
          4570 => x"39",
          4571 => x"08",
          4572 => x"81",
          4573 => x"38",
          4574 => x"74",
          4575 => x"38",
          4576 => x"3d",
          4577 => x"ff",
          4578 => x"81",
          4579 => x"54",
          4580 => x"08",
          4581 => x"53",
          4582 => x"08",
          4583 => x"ff",
          4584 => x"65",
          4585 => x"8b",
          4586 => x"53",
          4587 => x"bc",
          4588 => x"51",
          4589 => x"3f",
          4590 => x"0b",
          4591 => x"77",
          4592 => x"b1",
          4593 => x"ac",
          4594 => x"55",
          4595 => x"ac",
          4596 => x"0d",
          4597 => x"0d",
          4598 => x"88",
          4599 => x"05",
          4600 => x"fc",
          4601 => x"54",
          4602 => x"cd",
          4603 => x"d3",
          4604 => x"81",
          4605 => x"8a",
          4606 => x"33",
          4607 => x"2e",
          4608 => x"54",
          4609 => x"7a",
          4610 => x"38",
          4611 => x"90",
          4612 => x"33",
          4613 => x"70",
          4614 => x"55",
          4615 => x"38",
          4616 => x"99",
          4617 => x"81",
          4618 => x"57",
          4619 => x"7f",
          4620 => x"70",
          4621 => x"55",
          4622 => x"51",
          4623 => x"dd",
          4624 => x"7b",
          4625 => x"70",
          4626 => x"2a",
          4627 => x"08",
          4628 => x"11",
          4629 => x"40",
          4630 => x"5f",
          4631 => x"88",
          4632 => x"08",
          4633 => x"38",
          4634 => x"79",
          4635 => x"5a",
          4636 => x"51",
          4637 => x"3f",
          4638 => x"08",
          4639 => x"56",
          4640 => x"14",
          4641 => x"83",
          4642 => x"75",
          4643 => x"95",
          4644 => x"2e",
          4645 => x"75",
          4646 => x"1a",
          4647 => x"2e",
          4648 => x"39",
          4649 => x"5a",
          4650 => x"09",
          4651 => x"38",
          4652 => x"81",
          4653 => x"80",
          4654 => x"7c",
          4655 => x"7d",
          4656 => x"38",
          4657 => x"75",
          4658 => x"81",
          4659 => x"ff",
          4660 => x"74",
          4661 => x"ff",
          4662 => x"81",
          4663 => x"57",
          4664 => x"08",
          4665 => x"81",
          4666 => x"58",
          4667 => x"d4",
          4668 => x"ff",
          4669 => x"80",
          4670 => x"7f",
          4671 => x"54",
          4672 => x"b7",
          4673 => x"19",
          4674 => x"19",
          4675 => x"33",
          4676 => x"54",
          4677 => x"34",
          4678 => x"08",
          4679 => x"55",
          4680 => x"74",
          4681 => x"90",
          4682 => x"31",
          4683 => x"7f",
          4684 => x"81",
          4685 => x"73",
          4686 => x"76",
          4687 => x"d3",
          4688 => x"3d",
          4689 => x"3d",
          4690 => x"84",
          4691 => x"05",
          4692 => x"53",
          4693 => x"bf",
          4694 => x"d3",
          4695 => x"8b",
          4696 => x"81",
          4697 => x"24",
          4698 => x"81",
          4699 => x"10",
          4700 => x"c8",
          4701 => x"08",
          4702 => x"38",
          4703 => x"80",
          4704 => x"81",
          4705 => x"81",
          4706 => x"ff",
          4707 => x"81",
          4708 => x"81",
          4709 => x"81",
          4710 => x"83",
          4711 => x"9b",
          4712 => x"2a",
          4713 => x"51",
          4714 => x"74",
          4715 => x"98",
          4716 => x"53",
          4717 => x"51",
          4718 => x"3f",
          4719 => x"08",
          4720 => x"80",
          4721 => x"66",
          4722 => x"26",
          4723 => x"ff",
          4724 => x"55",
          4725 => x"83",
          4726 => x"84",
          4727 => x"80",
          4728 => x"7d",
          4729 => x"38",
          4730 => x"0a",
          4731 => x"ff",
          4732 => x"55",
          4733 => x"86",
          4734 => x"8b",
          4735 => x"52",
          4736 => x"f6",
          4737 => x"d3",
          4738 => x"7f",
          4739 => x"40",
          4740 => x"89",
          4741 => x"ac",
          4742 => x"d3",
          4743 => x"60",
          4744 => x"07",
          4745 => x"d3",
          4746 => x"70",
          4747 => x"08",
          4748 => x"72",
          4749 => x"51",
          4750 => x"91",
          4751 => x"fb",
          4752 => x"f8",
          4753 => x"52",
          4754 => x"9c",
          4755 => x"57",
          4756 => x"08",
          4757 => x"7c",
          4758 => x"81",
          4759 => x"80",
          4760 => x"2e",
          4761 => x"83",
          4762 => x"8e",
          4763 => x"26",
          4764 => x"65",
          4765 => x"8e",
          4766 => x"66",
          4767 => x"38",
          4768 => x"81",
          4769 => x"b3",
          4770 => x"2a",
          4771 => x"51",
          4772 => x"2e",
          4773 => x"87",
          4774 => x"82",
          4775 => x"7c",
          4776 => x"74",
          4777 => x"42",
          4778 => x"81",
          4779 => x"57",
          4780 => x"80",
          4781 => x"38",
          4782 => x"83",
          4783 => x"06",
          4784 => x"77",
          4785 => x"91",
          4786 => x"57",
          4787 => x"bd",
          4788 => x"22",
          4789 => x"59",
          4790 => x"9d",
          4791 => x"26",
          4792 => x"1b",
          4793 => x"10",
          4794 => x"51",
          4795 => x"74",
          4796 => x"38",
          4797 => x"ea",
          4798 => x"65",
          4799 => x"9d",
          4800 => x"ac",
          4801 => x"ac",
          4802 => x"1f",
          4803 => x"05",
          4804 => x"f4",
          4805 => x"d3",
          4806 => x"a0",
          4807 => x"fc",
          4808 => x"56",
          4809 => x"f0",
          4810 => x"81",
          4811 => x"57",
          4812 => x"77",
          4813 => x"8c",
          4814 => x"57",
          4815 => x"bc",
          4816 => x"22",
          4817 => x"59",
          4818 => x"9d",
          4819 => x"26",
          4820 => x"1b",
          4821 => x"10",
          4822 => x"51",
          4823 => x"74",
          4824 => x"38",
          4825 => x"ea",
          4826 => x"65",
          4827 => x"ad",
          4828 => x"ac",
          4829 => x"05",
          4830 => x"ac",
          4831 => x"26",
          4832 => x"0b",
          4833 => x"08",
          4834 => x"70",
          4835 => x"05",
          4836 => x"7d",
          4837 => x"ff",
          4838 => x"f3",
          4839 => x"d3",
          4840 => x"81",
          4841 => x"81",
          4842 => x"fe",
          4843 => x"81",
          4844 => x"83",
          4845 => x"43",
          4846 => x"11",
          4847 => x"11",
          4848 => x"30",
          4849 => x"73",
          4850 => x"59",
          4851 => x"83",
          4852 => x"06",
          4853 => x"1b",
          4854 => x"5b",
          4855 => x"1c",
          4856 => x"29",
          4857 => x"31",
          4858 => x"66",
          4859 => x"38",
          4860 => x"7c",
          4861 => x"70",
          4862 => x"56",
          4863 => x"3f",
          4864 => x"08",
          4865 => x"2e",
          4866 => x"9b",
          4867 => x"ac",
          4868 => x"f5",
          4869 => x"77",
          4870 => x"81",
          4871 => x"fd",
          4872 => x"57",
          4873 => x"61",
          4874 => x"81",
          4875 => x"38",
          4876 => x"76",
          4877 => x"77",
          4878 => x"19",
          4879 => x"c0",
          4880 => x"74",
          4881 => x"39",
          4882 => x"81",
          4883 => x"80",
          4884 => x"83",
          4885 => x"39",
          4886 => x"78",
          4887 => x"80",
          4888 => x"d4",
          4889 => x"86",
          4890 => x"9f",
          4891 => x"38",
          4892 => x"78",
          4893 => x"80",
          4894 => x"bc",
          4895 => x"86",
          4896 => x"55",
          4897 => x"09",
          4898 => x"38",
          4899 => x"9f",
          4900 => x"06",
          4901 => x"74",
          4902 => x"7d",
          4903 => x"7e",
          4904 => x"8f",
          4905 => x"81",
          4906 => x"7e",
          4907 => x"df",
          4908 => x"8b",
          4909 => x"99",
          4910 => x"7f",
          4911 => x"7a",
          4912 => x"06",
          4913 => x"51",
          4914 => x"3f",
          4915 => x"05",
          4916 => x"32",
          4917 => x"96",
          4918 => x"06",
          4919 => x"91",
          4920 => x"98",
          4921 => x"83",
          4922 => x"90",
          4923 => x"d6",
          4924 => x"93",
          4925 => x"98",
          4926 => x"39",
          4927 => x"1f",
          4928 => x"dc",
          4929 => x"95",
          4930 => x"52",
          4931 => x"ff",
          4932 => x"81",
          4933 => x"1f",
          4934 => x"a6",
          4935 => x"9c",
          4936 => x"98",
          4937 => x"83",
          4938 => x"06",
          4939 => x"82",
          4940 => x"52",
          4941 => x"51",
          4942 => x"3f",
          4943 => x"1f",
          4944 => x"9c",
          4945 => x"ac",
          4946 => x"98",
          4947 => x"52",
          4948 => x"ff",
          4949 => x"86",
          4950 => x"51",
          4951 => x"3f",
          4952 => x"80",
          4953 => x"a9",
          4954 => x"05",
          4955 => x"81",
          4956 => x"80",
          4957 => x"ff",
          4958 => x"b2",
          4959 => x"b2",
          4960 => x"1f",
          4961 => x"d8",
          4962 => x"ff",
          4963 => x"96",
          4964 => x"97",
          4965 => x"80",
          4966 => x"34",
          4967 => x"05",
          4968 => x"81",
          4969 => x"ab",
          4970 => x"97",
          4971 => x"d4",
          4972 => x"fe",
          4973 => x"97",
          4974 => x"54",
          4975 => x"52",
          4976 => x"93",
          4977 => x"57",
          4978 => x"08",
          4979 => x"61",
          4980 => x"81",
          4981 => x"38",
          4982 => x"86",
          4983 => x"52",
          4984 => x"93",
          4985 => x"53",
          4986 => x"51",
          4987 => x"3f",
          4988 => x"a4",
          4989 => x"51",
          4990 => x"3f",
          4991 => x"e4",
          4992 => x"e4",
          4993 => x"96",
          4994 => x"16",
          4995 => x"1f",
          4996 => x"cc",
          4997 => x"83",
          4998 => x"ff",
          4999 => x"82",
          5000 => x"83",
          5001 => x"ff",
          5002 => x"81",
          5003 => x"05",
          5004 => x"79",
          5005 => x"86",
          5006 => x"63",
          5007 => x"7e",
          5008 => x"ff",
          5009 => x"64",
          5010 => x"7e",
          5011 => x"e3",
          5012 => x"80",
          5013 => x"2e",
          5014 => x"9e",
          5015 => x"7e",
          5016 => x"fc",
          5017 => x"84",
          5018 => x"95",
          5019 => x"0a",
          5020 => x"51",
          5021 => x"3f",
          5022 => x"ff",
          5023 => x"61",
          5024 => x"38",
          5025 => x"52",
          5026 => x"95",
          5027 => x"55",
          5028 => x"61",
          5029 => x"74",
          5030 => x"75",
          5031 => x"79",
          5032 => x"9a",
          5033 => x"ac",
          5034 => x"38",
          5035 => x"52",
          5036 => x"95",
          5037 => x"16",
          5038 => x"56",
          5039 => x"38",
          5040 => x"7a",
          5041 => x"8d",
          5042 => x"61",
          5043 => x"38",
          5044 => x"57",
          5045 => x"83",
          5046 => x"76",
          5047 => x"7e",
          5048 => x"ff",
          5049 => x"81",
          5050 => x"81",
          5051 => x"16",
          5052 => x"56",
          5053 => x"38",
          5054 => x"83",
          5055 => x"86",
          5056 => x"ff",
          5057 => x"38",
          5058 => x"82",
          5059 => x"81",
          5060 => x"2a",
          5061 => x"77",
          5062 => x"7d",
          5063 => x"7e",
          5064 => x"8f",
          5065 => x"d5",
          5066 => x"1f",
          5067 => x"92",
          5068 => x"1f",
          5069 => x"34",
          5070 => x"17",
          5071 => x"82",
          5072 => x"83",
          5073 => x"84",
          5074 => x"66",
          5075 => x"fd",
          5076 => x"51",
          5077 => x"3f",
          5078 => x"17",
          5079 => x"ac",
          5080 => x"bf",
          5081 => x"86",
          5082 => x"d3",
          5083 => x"17",
          5084 => x"83",
          5085 => x"ff",
          5086 => x"65",
          5087 => x"1f",
          5088 => x"dc",
          5089 => x"77",
          5090 => x"79",
          5091 => x"ae",
          5092 => x"81",
          5093 => x"a3",
          5094 => x"80",
          5095 => x"ff",
          5096 => x"81",
          5097 => x"ac",
          5098 => x"8d",
          5099 => x"8b",
          5100 => x"87",
          5101 => x"83",
          5102 => x"76",
          5103 => x"0c",
          5104 => x"04",
          5105 => x"73",
          5106 => x"26",
          5107 => x"71",
          5108 => x"b1",
          5109 => x"71",
          5110 => x"c1",
          5111 => x"80",
          5112 => x"d4",
          5113 => x"e8",
          5114 => x"9e",
          5115 => x"39",
          5116 => x"51",
          5117 => x"3f",
          5118 => x"81",
          5119 => x"ff",
          5120 => x"81",
          5121 => x"c2",
          5122 => x"ff",
          5123 => x"a8",
          5124 => x"b0",
          5125 => x"f2",
          5126 => x"39",
          5127 => x"51",
          5128 => x"3f",
          5129 => x"81",
          5130 => x"fe",
          5131 => x"81",
          5132 => x"c2",
          5133 => x"ff",
          5134 => x"fc",
          5135 => x"84",
          5136 => x"c6",
          5137 => x"39",
          5138 => x"51",
          5139 => x"3f",
          5140 => x"81",
          5141 => x"fe",
          5142 => x"80",
          5143 => x"c3",
          5144 => x"ff",
          5145 => x"d0",
          5146 => x"f8",
          5147 => x"9a",
          5148 => x"39",
          5149 => x"51",
          5150 => x"3f",
          5151 => x"c4",
          5152 => x"ff",
          5153 => x"39",
          5154 => x"51",
          5155 => x"3f",
          5156 => x"c4",
          5157 => x"fe",
          5158 => x"39",
          5159 => x"51",
          5160 => x"3f",
          5161 => x"c5",
          5162 => x"fe",
          5163 => x"39",
          5164 => x"51",
          5165 => x"3f",
          5166 => x"04",
          5167 => x"77",
          5168 => x"74",
          5169 => x"93",
          5170 => x"75",
          5171 => x"51",
          5172 => x"3f",
          5173 => x"08",
          5174 => x"87",
          5175 => x"51",
          5176 => x"3f",
          5177 => x"08",
          5178 => x"fe",
          5179 => x"81",
          5180 => x"55",
          5181 => x"53",
          5182 => x"c5",
          5183 => x"84",
          5184 => x"3d",
          5185 => x"ec",
          5186 => x"97",
          5187 => x"99",
          5188 => x"88",
          5189 => x"05",
          5190 => x"30",
          5191 => x"80",
          5192 => x"75",
          5193 => x"59",
          5194 => x"58",
          5195 => x"81",
          5196 => x"53",
          5197 => x"96",
          5198 => x"05",
          5199 => x"99",
          5200 => x"ac",
          5201 => x"d3",
          5202 => x"38",
          5203 => x"08",
          5204 => x"88",
          5205 => x"ac",
          5206 => x"96",
          5207 => x"11",
          5208 => x"80",
          5209 => x"fb",
          5210 => x"c0",
          5211 => x"d3",
          5212 => x"81",
          5213 => x"8e",
          5214 => x"2e",
          5215 => x"19",
          5216 => x"59",
          5217 => x"96",
          5218 => x"05",
          5219 => x"3f",
          5220 => x"79",
          5221 => x"7b",
          5222 => x"2a",
          5223 => x"57",
          5224 => x"80",
          5225 => x"81",
          5226 => x"87",
          5227 => x"08",
          5228 => x"fe",
          5229 => x"55",
          5230 => x"ac",
          5231 => x"3d",
          5232 => x"3d",
          5233 => x"05",
          5234 => x"7d",
          5235 => x"53",
          5236 => x"51",
          5237 => x"81",
          5238 => x"a4",
          5239 => x"2e",
          5240 => x"81",
          5241 => x"98",
          5242 => x"60",
          5243 => x"ac",
          5244 => x"7e",
          5245 => x"81",
          5246 => x"59",
          5247 => x"04",
          5248 => x"ac",
          5249 => x"0d",
          5250 => x"0d",
          5251 => x"33",
          5252 => x"53",
          5253 => x"52",
          5254 => x"e8",
          5255 => x"cc",
          5256 => x"55",
          5257 => x"3f",
          5258 => x"54",
          5259 => x"53",
          5260 => x"52",
          5261 => x"51",
          5262 => x"3f",
          5263 => x"85",
          5264 => x"ff",
          5265 => x"0d",
          5266 => x"0d",
          5267 => x"80",
          5268 => x"f9",
          5269 => x"51",
          5270 => x"3f",
          5271 => x"51",
          5272 => x"3f",
          5273 => x"ee",
          5274 => x"81",
          5275 => x"06",
          5276 => x"80",
          5277 => x"81",
          5278 => x"de",
          5279 => x"b0",
          5280 => x"d4",
          5281 => x"fe",
          5282 => x"72",
          5283 => x"81",
          5284 => x"71",
          5285 => x"38",
          5286 => x"ee",
          5287 => x"c6",
          5288 => x"f0",
          5289 => x"51",
          5290 => x"3f",
          5291 => x"70",
          5292 => x"52",
          5293 => x"95",
          5294 => x"fe",
          5295 => x"81",
          5296 => x"fe",
          5297 => x"80",
          5298 => x"8e",
          5299 => x"2a",
          5300 => x"51",
          5301 => x"2e",
          5302 => x"51",
          5303 => x"3f",
          5304 => x"51",
          5305 => x"3f",
          5306 => x"ed",
          5307 => x"85",
          5308 => x"06",
          5309 => x"80",
          5310 => x"81",
          5311 => x"da",
          5312 => x"fc",
          5313 => x"d0",
          5314 => x"fe",
          5315 => x"72",
          5316 => x"81",
          5317 => x"71",
          5318 => x"38",
          5319 => x"ed",
          5320 => x"c7",
          5321 => x"ef",
          5322 => x"51",
          5323 => x"3f",
          5324 => x"70",
          5325 => x"52",
          5326 => x"95",
          5327 => x"fe",
          5328 => x"81",
          5329 => x"fe",
          5330 => x"80",
          5331 => x"8a",
          5332 => x"2a",
          5333 => x"51",
          5334 => x"2e",
          5335 => x"51",
          5336 => x"3f",
          5337 => x"51",
          5338 => x"3f",
          5339 => x"ec",
          5340 => x"f8",
          5341 => x"3d",
          5342 => x"3d",
          5343 => x"08",
          5344 => x"57",
          5345 => x"80",
          5346 => x"39",
          5347 => x"85",
          5348 => x"80",
          5349 => x"15",
          5350 => x"33",
          5351 => x"a0",
          5352 => x"81",
          5353 => x"70",
          5354 => x"06",
          5355 => x"e6",
          5356 => x"53",
          5357 => x"09",
          5358 => x"38",
          5359 => x"81",
          5360 => x"80",
          5361 => x"29",
          5362 => x"05",
          5363 => x"70",
          5364 => x"fe",
          5365 => x"81",
          5366 => x"8b",
          5367 => x"33",
          5368 => x"2e",
          5369 => x"81",
          5370 => x"ff",
          5371 => x"bb",
          5372 => x"38",
          5373 => x"81",
          5374 => x"88",
          5375 => x"ce",
          5376 => x"70",
          5377 => x"72",
          5378 => x"5e",
          5379 => x"81",
          5380 => x"ff",
          5381 => x"81",
          5382 => x"81",
          5383 => x"78",
          5384 => x"81",
          5385 => x"81",
          5386 => x"96",
          5387 => x"59",
          5388 => x"3f",
          5389 => x"52",
          5390 => x"51",
          5391 => x"3f",
          5392 => x"08",
          5393 => x"2e",
          5394 => x"c7",
          5395 => x"fd",
          5396 => x"39",
          5397 => x"5c",
          5398 => x"51",
          5399 => x"3f",
          5400 => x"43",
          5401 => x"70",
          5402 => x"52",
          5403 => x"e4",
          5404 => x"52",
          5405 => x"fd",
          5406 => x"3d",
          5407 => x"51",
          5408 => x"81",
          5409 => x"90",
          5410 => x"2c",
          5411 => x"81",
          5412 => x"af",
          5413 => x"10",
          5414 => x"05",
          5415 => x"04",
          5416 => x"f4",
          5417 => x"f8",
          5418 => x"fe",
          5419 => x"d3",
          5420 => x"38",
          5421 => x"51",
          5422 => x"3f",
          5423 => x"b4",
          5424 => x"11",
          5425 => x"05",
          5426 => x"c3",
          5427 => x"ac",
          5428 => x"88",
          5429 => x"25",
          5430 => x"40",
          5431 => x"33",
          5432 => x"c3",
          5433 => x"ff",
          5434 => x"81",
          5435 => x"81",
          5436 => x"78",
          5437 => x"c8",
          5438 => x"f6",
          5439 => x"5d",
          5440 => x"81",
          5441 => x"fe",
          5442 => x"fe",
          5443 => x"3d",
          5444 => x"53",
          5445 => x"51",
          5446 => x"3f",
          5447 => x"08",
          5448 => x"b4",
          5449 => x"80",
          5450 => x"c3",
          5451 => x"ff",
          5452 => x"81",
          5453 => x"52",
          5454 => x"51",
          5455 => x"3f",
          5456 => x"b4",
          5457 => x"11",
          5458 => x"05",
          5459 => x"bf",
          5460 => x"ac",
          5461 => x"87",
          5462 => x"26",
          5463 => x"b4",
          5464 => x"11",
          5465 => x"05",
          5466 => x"a3",
          5467 => x"ac",
          5468 => x"81",
          5469 => x"40",
          5470 => x"c8",
          5471 => x"3d",
          5472 => x"fe",
          5473 => x"02",
          5474 => x"53",
          5475 => x"84",
          5476 => x"e0",
          5477 => x"ff",
          5478 => x"81",
          5479 => x"80",
          5480 => x"81",
          5481 => x"51",
          5482 => x"fd",
          5483 => x"c8",
          5484 => x"f4",
          5485 => x"5c",
          5486 => x"b4",
          5487 => x"05",
          5488 => x"a4",
          5489 => x"ac",
          5490 => x"fe",
          5491 => x"5b",
          5492 => x"3f",
          5493 => x"d3",
          5494 => x"7a",
          5495 => x"3f",
          5496 => x"08",
          5497 => x"f0",
          5498 => x"ac",
          5499 => x"d4",
          5500 => x"39",
          5501 => x"f8",
          5502 => x"e3",
          5503 => x"d3",
          5504 => x"3d",
          5505 => x"52",
          5506 => x"c1",
          5507 => x"ac",
          5508 => x"fe",
          5509 => x"5a",
          5510 => x"3f",
          5511 => x"08",
          5512 => x"f8",
          5513 => x"fe",
          5514 => x"81",
          5515 => x"81",
          5516 => x"80",
          5517 => x"81",
          5518 => x"81",
          5519 => x"78",
          5520 => x"7a",
          5521 => x"3f",
          5522 => x"08",
          5523 => x"88",
          5524 => x"ac",
          5525 => x"ec",
          5526 => x"39",
          5527 => x"51",
          5528 => x"3f",
          5529 => x"f2",
          5530 => x"ec",
          5531 => x"94",
          5532 => x"96",
          5533 => x"fe",
          5534 => x"fb",
          5535 => x"80",
          5536 => x"c0",
          5537 => x"84",
          5538 => x"87",
          5539 => x"0c",
          5540 => x"51",
          5541 => x"3f",
          5542 => x"81",
          5543 => x"fe",
          5544 => x"8c",
          5545 => x"87",
          5546 => x"0c",
          5547 => x"0b",
          5548 => x"94",
          5549 => x"39",
          5550 => x"f4",
          5551 => x"f8",
          5552 => x"fa",
          5553 => x"d3",
          5554 => x"2e",
          5555 => x"60",
          5556 => x"d4",
          5557 => x"ac",
          5558 => x"78",
          5559 => x"fe",
          5560 => x"fe",
          5561 => x"fe",
          5562 => x"81",
          5563 => x"80",
          5564 => x"38",
          5565 => x"c9",
          5566 => x"f8",
          5567 => x"59",
          5568 => x"d3",
          5569 => x"81",
          5570 => x"80",
          5571 => x"38",
          5572 => x"08",
          5573 => x"8c",
          5574 => x"e8",
          5575 => x"39",
          5576 => x"51",
          5577 => x"3f",
          5578 => x"3f",
          5579 => x"81",
          5580 => x"fe",
          5581 => x"80",
          5582 => x"39",
          5583 => x"3f",
          5584 => x"61",
          5585 => x"59",
          5586 => x"fa",
          5587 => x"7c",
          5588 => x"80",
          5589 => x"38",
          5590 => x"f8",
          5591 => x"e1",
          5592 => x"ca",
          5593 => x"d3",
          5594 => x"81",
          5595 => x"80",
          5596 => x"e0",
          5597 => x"70",
          5598 => x"f7",
          5599 => x"cb",
          5600 => x"d3",
          5601 => x"56",
          5602 => x"42",
          5603 => x"54",
          5604 => x"53",
          5605 => x"52",
          5606 => x"a6",
          5607 => x"ac",
          5608 => x"81",
          5609 => x"32",
          5610 => x"8a",
          5611 => x"2e",
          5612 => x"f9",
          5613 => x"ca",
          5614 => x"f6",
          5615 => x"98",
          5616 => x"0d",
          5617 => x"d3",
          5618 => x"90",
          5619 => x"87",
          5620 => x"0c",
          5621 => x"e4",
          5622 => x"94",
          5623 => x"80",
          5624 => x"c0",
          5625 => x"8c",
          5626 => x"87",
          5627 => x"0c",
          5628 => x"81",
          5629 => x"96",
          5630 => x"d3",
          5631 => x"e8",
          5632 => x"ee",
          5633 => x"cb",
          5634 => x"e5",
          5635 => x"cb",
          5636 => x"ef",
          5637 => x"a4",
          5638 => x"ee",
          5639 => x"51",
          5640 => x"f7",
          5641 => x"04",
          5642 => x"44",
          5643 => x"17",
          5644 => x"20",
          5645 => x"29",
          5646 => x"32",
          5647 => x"3b",
          5648 => x"b6",
          5649 => x"a7",
          5650 => x"be",
          5651 => x"c6",
          5652 => x"c6",
          5653 => x"c6",
          5654 => x"c6",
          5655 => x"c6",
          5656 => x"c6",
          5657 => x"c6",
          5658 => x"c6",
          5659 => x"c6",
          5660 => x"c6",
          5661 => x"ba",
          5662 => x"c6",
          5663 => x"c6",
          5664 => x"c6",
          5665 => x"3a",
          5666 => x"c6",
          5667 => x"be",
          5668 => x"c6",
          5669 => x"c6",
          5670 => x"c2",
          5671 => x"a6",
          5672 => x"da",
          5673 => x"e5",
          5674 => x"f0",
          5675 => x"fb",
          5676 => x"06",
          5677 => x"11",
          5678 => x"1c",
          5679 => x"27",
          5680 => x"32",
          5681 => x"3d",
          5682 => x"48",
          5683 => x"53",
          5684 => x"5e",
          5685 => x"69",
          5686 => x"74",
          5687 => x"7e",
          5688 => x"88",
          5689 => x"92",
          5690 => x"9c",
          5691 => x"58",
          5692 => x"43",
          5693 => x"a0",
          5694 => x"43",
          5695 => x"0e",
          5696 => x"43",
          5697 => x"43",
          5698 => x"43",
          5699 => x"43",
          5700 => x"43",
          5701 => x"43",
          5702 => x"43",
          5703 => x"43",
          5704 => x"43",
          5705 => x"43",
          5706 => x"43",
          5707 => x"43",
          5708 => x"43",
          5709 => x"43",
          5710 => x"43",
          5711 => x"43",
          5712 => x"43",
          5713 => x"43",
          5714 => x"43",
          5715 => x"43",
          5716 => x"43",
          5717 => x"43",
          5718 => x"43",
          5719 => x"43",
          5720 => x"43",
          5721 => x"43",
          5722 => x"43",
          5723 => x"43",
          5724 => x"43",
          5725 => x"43",
          5726 => x"43",
          5727 => x"43",
          5728 => x"43",
          5729 => x"43",
          5730 => x"43",
          5731 => x"43",
          5732 => x"43",
          5733 => x"43",
          5734 => x"bb",
          5735 => x"43",
          5736 => x"43",
          5737 => x"43",
          5738 => x"43",
          5739 => x"f4",
          5740 => x"43",
          5741 => x"43",
          5742 => x"43",
          5743 => x"43",
          5744 => x"43",
          5745 => x"43",
          5746 => x"43",
          5747 => x"43",
          5748 => x"43",
          5749 => x"43",
          5750 => x"43",
          5751 => x"43",
          5752 => x"43",
          5753 => x"43",
          5754 => x"43",
          5755 => x"43",
          5756 => x"43",
          5757 => x"43",
          5758 => x"43",
          5759 => x"43",
          5760 => x"43",
          5761 => x"43",
          5762 => x"43",
          5763 => x"43",
          5764 => x"43",
          5765 => x"43",
          5766 => x"43",
          5767 => x"43",
          5768 => x"43",
          5769 => x"43",
          5770 => x"43",
          5771 => x"5c",
          5772 => x"6d",
          5773 => x"43",
          5774 => x"43",
          5775 => x"7e",
          5776 => x"9b",
          5777 => x"43",
          5778 => x"43",
          5779 => x"43",
          5780 => x"43",
          5781 => x"43",
          5782 => x"43",
          5783 => x"43",
          5784 => x"43",
          5785 => x"43",
          5786 => x"43",
          5787 => x"43",
          5788 => x"43",
          5789 => x"43",
          5790 => x"43",
          5791 => x"43",
          5792 => x"43",
          5793 => x"43",
          5794 => x"43",
          5795 => x"43",
          5796 => x"43",
          5797 => x"43",
          5798 => x"43",
          5799 => x"43",
          5800 => x"43",
          5801 => x"43",
          5802 => x"43",
          5803 => x"43",
          5804 => x"43",
          5805 => x"43",
          5806 => x"43",
          5807 => x"43",
          5808 => x"43",
          5809 => x"43",
          5810 => x"43",
          5811 => x"b8",
          5812 => x"dd",
          5813 => x"43",
          5814 => x"43",
          5815 => x"43",
          5816 => x"43",
          5817 => x"43",
          5818 => x"43",
          5819 => x"43",
          5820 => x"43",
          5821 => x"20",
          5822 => x"2f",
          5823 => x"43",
          5824 => x"3c",
          5825 => x"43",
          5826 => x"58",
          5827 => x"25",
          5828 => x"64",
          5829 => x"3a",
          5830 => x"25",
          5831 => x"64",
          5832 => x"00",
          5833 => x"20",
          5834 => x"66",
          5835 => x"72",
          5836 => x"6f",
          5837 => x"00",
          5838 => x"72",
          5839 => x"53",
          5840 => x"63",
          5841 => x"69",
          5842 => x"00",
          5843 => x"65",
          5844 => x"65",
          5845 => x"6d",
          5846 => x"6d",
          5847 => x"65",
          5848 => x"00",
          5849 => x"20",
          5850 => x"4e",
          5851 => x"41",
          5852 => x"53",
          5853 => x"74",
          5854 => x"38",
          5855 => x"53",
          5856 => x"3d",
          5857 => x"58",
          5858 => x"00",
          5859 => x"20",
          5860 => x"4d",
          5861 => x"74",
          5862 => x"3d",
          5863 => x"58",
          5864 => x"69",
          5865 => x"25",
          5866 => x"29",
          5867 => x"00",
          5868 => x"20",
          5869 => x"20",
          5870 => x"61",
          5871 => x"25",
          5872 => x"2c",
          5873 => x"7a",
          5874 => x"30",
          5875 => x"2e",
          5876 => x"00",
          5877 => x"20",
          5878 => x"54",
          5879 => x"00",
          5880 => x"20",
          5881 => x"0a",
          5882 => x"00",
          5883 => x"20",
          5884 => x"0a",
          5885 => x"00",
          5886 => x"20",
          5887 => x"43",
          5888 => x"20",
          5889 => x"76",
          5890 => x"73",
          5891 => x"32",
          5892 => x"0a",
          5893 => x"00",
          5894 => x"20",
          5895 => x"45",
          5896 => x"50",
          5897 => x"4f",
          5898 => x"4f",
          5899 => x"52",
          5900 => x"00",
          5901 => x"20",
          5902 => x"45",
          5903 => x"28",
          5904 => x"65",
          5905 => x"25",
          5906 => x"29",
          5907 => x"00",
          5908 => x"72",
          5909 => x"65",
          5910 => x"00",
          5911 => x"20",
          5912 => x"20",
          5913 => x"65",
          5914 => x"65",
          5915 => x"72",
          5916 => x"64",
          5917 => x"73",
          5918 => x"25",
          5919 => x"0a",
          5920 => x"00",
          5921 => x"20",
          5922 => x"20",
          5923 => x"6f",
          5924 => x"53",
          5925 => x"74",
          5926 => x"64",
          5927 => x"73",
          5928 => x"25",
          5929 => x"0a",
          5930 => x"00",
          5931 => x"20",
          5932 => x"63",
          5933 => x"74",
          5934 => x"20",
          5935 => x"72",
          5936 => x"20",
          5937 => x"20",
          5938 => x"25",
          5939 => x"0a",
          5940 => x"00",
          5941 => x"20",
          5942 => x"20",
          5943 => x"20",
          5944 => x"20",
          5945 => x"20",
          5946 => x"20",
          5947 => x"20",
          5948 => x"25",
          5949 => x"0a",
          5950 => x"00",
          5951 => x"20",
          5952 => x"74",
          5953 => x"43",
          5954 => x"6b",
          5955 => x"65",
          5956 => x"20",
          5957 => x"20",
          5958 => x"25",
          5959 => x"0a",
          5960 => x"00",
          5961 => x"6c",
          5962 => x"00",
          5963 => x"69",
          5964 => x"00",
          5965 => x"78",
          5966 => x"00",
          5967 => x"00",
          5968 => x"6d",
          5969 => x"00",
          5970 => x"6e",
          5971 => x"00",
          5972 => x"00",
          5973 => x"2c",
          5974 => x"3d",
          5975 => x"5d",
          5976 => x"00",
          5977 => x"00",
          5978 => x"33",
          5979 => x"00",
          5980 => x"00",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"00",
          5985 => x"00",
          5986 => x"00",
          5987 => x"00",
          5988 => x"00",
          5989 => x"00",
          5990 => x"4d",
          5991 => x"53",
          5992 => x"00",
          5993 => x"4e",
          5994 => x"20",
          5995 => x"46",
          5996 => x"32",
          5997 => x"00",
          5998 => x"4e",
          5999 => x"20",
          6000 => x"46",
          6001 => x"20",
          6002 => x"00",
          6003 => x"50",
          6004 => x"00",
          6005 => x"00",
          6006 => x"00",
          6007 => x"41",
          6008 => x"80",
          6009 => x"49",
          6010 => x"8f",
          6011 => x"4f",
          6012 => x"55",
          6013 => x"9b",
          6014 => x"9f",
          6015 => x"55",
          6016 => x"a7",
          6017 => x"ab",
          6018 => x"af",
          6019 => x"b3",
          6020 => x"b7",
          6021 => x"bb",
          6022 => x"bf",
          6023 => x"c3",
          6024 => x"c7",
          6025 => x"cb",
          6026 => x"cf",
          6027 => x"d3",
          6028 => x"d7",
          6029 => x"db",
          6030 => x"df",
          6031 => x"e3",
          6032 => x"e7",
          6033 => x"eb",
          6034 => x"ef",
          6035 => x"f3",
          6036 => x"f7",
          6037 => x"fb",
          6038 => x"ff",
          6039 => x"3b",
          6040 => x"2f",
          6041 => x"3a",
          6042 => x"7c",
          6043 => x"00",
          6044 => x"04",
          6045 => x"40",
          6046 => x"00",
          6047 => x"00",
          6048 => x"02",
          6049 => x"08",
          6050 => x"20",
          6051 => x"00",
          6052 => x"31",
          6053 => x"00",
          6054 => x"31",
          6055 => x"00",
          6056 => x"41",
          6057 => x"00",
          6058 => x"4b",
          6059 => x"20",
          6060 => x"54",
          6061 => x"53",
          6062 => x"00",
          6063 => x"4b",
          6064 => x"46",
          6065 => x"20",
          6066 => x"54",
          6067 => x"53",
          6068 => x"00",
          6069 => x"45",
          6070 => x"54",
          6071 => x"43",
          6072 => x"52",
          6073 => x"00",
          6074 => x"4f",
          6075 => x"00",
          6076 => x"44",
          6077 => x"45",
          6078 => x"00",
          6079 => x"54",
          6080 => x"00",
          6081 => x"43",
          6082 => x"4f",
          6083 => x"00",
          6084 => x"43",
          6085 => x"4d",
          6086 => x"44",
          6087 => x"00",
          6088 => x"6d",
          6089 => x"00",
          6090 => x"69",
          6091 => x"00",
          6092 => x"61",
          6093 => x"00",
          6094 => x"63",
          6095 => x"00",
          6096 => x"6d",
          6097 => x"00",
          6098 => x"69",
          6099 => x"00",
          6100 => x"61",
          6101 => x"00",
          6102 => x"69",
          6103 => x"00",
          6104 => x"6c",
          6105 => x"00",
          6106 => x"6e",
          6107 => x"00",
          6108 => x"69",
          6109 => x"00",
          6110 => x"65",
          6111 => x"00",
          6112 => x"6f",
          6113 => x"00",
          6114 => x"65",
          6115 => x"00",
          6116 => x"61",
          6117 => x"00",
          6118 => x"73",
          6119 => x"74",
          6120 => x"00",
          6121 => x"69",
          6122 => x"00",
          6123 => x"75",
          6124 => x"00",
          6125 => x"6c",
          6126 => x"00",
          6127 => x"74",
          6128 => x"00",
          6129 => x"6d",
          6130 => x"00",
          6131 => x"6e",
          6132 => x"00",
          6133 => x"6c",
          6134 => x"00",
          6135 => x"64",
          6136 => x"00",
          6137 => x"61",
          6138 => x"00",
          6139 => x"72",
          6140 => x"00",
          6141 => x"74",
          6142 => x"00",
          6143 => x"00",
          6144 => x"6e",
          6145 => x"00",
          6146 => x"72",
          6147 => x"00",
          6148 => x"61",
          6149 => x"00",
          6150 => x"65",
          6151 => x"00",
          6152 => x"76",
          6153 => x"00",
          6154 => x"6d",
          6155 => x"00",
          6156 => x"00",
          6157 => x"69",
          6158 => x"00",
          6159 => x"6f",
          6160 => x"72",
          6161 => x"00",
          6162 => x"62",
          6163 => x"00",
          6164 => x"66",
          6165 => x"00",
          6166 => x"72",
          6167 => x"00",
          6168 => x"6d",
          6169 => x"00",
          6170 => x"00",
          6171 => x"00",
          6172 => x"00",
          6173 => x"00",
          6174 => x"00",
          6175 => x"00",
          6176 => x"00",
          6177 => x"00",
          6178 => x"00",
          6179 => x"79",
          6180 => x"00",
          6181 => x"65",
          6182 => x"6b",
          6183 => x"00",
          6184 => x"6c",
          6185 => x"00",
          6186 => x"00",
          6187 => x"74",
          6188 => x"00",
          6189 => x"65",
          6190 => x"00",
          6191 => x"70",
          6192 => x"00",
          6193 => x"6f",
          6194 => x"00",
          6195 => x"65",
          6196 => x"00",
          6197 => x"74",
          6198 => x"00",
          6199 => x"6b",
          6200 => x"72",
          6201 => x"00",
          6202 => x"65",
          6203 => x"6c",
          6204 => x"72",
          6205 => x"0a",
          6206 => x"00",
          6207 => x"6b",
          6208 => x"74",
          6209 => x"61",
          6210 => x"0a",
          6211 => x"00",
          6212 => x"66",
          6213 => x"20",
          6214 => x"6e",
          6215 => x"00",
          6216 => x"70",
          6217 => x"20",
          6218 => x"6e",
          6219 => x"00",
          6220 => x"61",
          6221 => x"20",
          6222 => x"65",
          6223 => x"65",
          6224 => x"00",
          6225 => x"65",
          6226 => x"64",
          6227 => x"65",
          6228 => x"00",
          6229 => x"65",
          6230 => x"72",
          6231 => x"79",
          6232 => x"69",
          6233 => x"2e",
          6234 => x"00",
          6235 => x"65",
          6236 => x"6e",
          6237 => x"20",
          6238 => x"61",
          6239 => x"2e",
          6240 => x"00",
          6241 => x"69",
          6242 => x"72",
          6243 => x"20",
          6244 => x"74",
          6245 => x"65",
          6246 => x"00",
          6247 => x"76",
          6248 => x"75",
          6249 => x"72",
          6250 => x"20",
          6251 => x"61",
          6252 => x"2e",
          6253 => x"00",
          6254 => x"6b",
          6255 => x"74",
          6256 => x"61",
          6257 => x"64",
          6258 => x"00",
          6259 => x"63",
          6260 => x"61",
          6261 => x"6c",
          6262 => x"69",
          6263 => x"79",
          6264 => x"6d",
          6265 => x"75",
          6266 => x"6f",
          6267 => x"69",
          6268 => x"0a",
          6269 => x"00",
          6270 => x"6d",
          6271 => x"61",
          6272 => x"74",
          6273 => x"0a",
          6274 => x"00",
          6275 => x"65",
          6276 => x"2c",
          6277 => x"65",
          6278 => x"69",
          6279 => x"63",
          6280 => x"65",
          6281 => x"64",
          6282 => x"00",
          6283 => x"65",
          6284 => x"20",
          6285 => x"6b",
          6286 => x"0a",
          6287 => x"00",
          6288 => x"75",
          6289 => x"63",
          6290 => x"74",
          6291 => x"6d",
          6292 => x"2e",
          6293 => x"00",
          6294 => x"20",
          6295 => x"79",
          6296 => x"65",
          6297 => x"69",
          6298 => x"2e",
          6299 => x"00",
          6300 => x"61",
          6301 => x"65",
          6302 => x"69",
          6303 => x"72",
          6304 => x"74",
          6305 => x"00",
          6306 => x"63",
          6307 => x"2e",
          6308 => x"00",
          6309 => x"6e",
          6310 => x"20",
          6311 => x"6f",
          6312 => x"00",
          6313 => x"75",
          6314 => x"74",
          6315 => x"25",
          6316 => x"74",
          6317 => x"75",
          6318 => x"74",
          6319 => x"73",
          6320 => x"0a",
          6321 => x"00",
          6322 => x"64",
          6323 => x"00",
          6324 => x"54",
          6325 => x"00",
          6326 => x"20",
          6327 => x"28",
          6328 => x"00",
          6329 => x"30",
          6330 => x"30",
          6331 => x"00",
          6332 => x"33",
          6333 => x"00",
          6334 => x"55",
          6335 => x"65",
          6336 => x"30",
          6337 => x"20",
          6338 => x"25",
          6339 => x"2a",
          6340 => x"00",
          6341 => x"54",
          6342 => x"6e",
          6343 => x"72",
          6344 => x"20",
          6345 => x"64",
          6346 => x"0a",
          6347 => x"00",
          6348 => x"65",
          6349 => x"6e",
          6350 => x"72",
          6351 => x"0a",
          6352 => x"00",
          6353 => x"20",
          6354 => x"65",
          6355 => x"70",
          6356 => x"00",
          6357 => x"54",
          6358 => x"44",
          6359 => x"74",
          6360 => x"75",
          6361 => x"00",
          6362 => x"54",
          6363 => x"52",
          6364 => x"74",
          6365 => x"75",
          6366 => x"00",
          6367 => x"54",
          6368 => x"58",
          6369 => x"74",
          6370 => x"75",
          6371 => x"00",
          6372 => x"54",
          6373 => x"58",
          6374 => x"74",
          6375 => x"75",
          6376 => x"00",
          6377 => x"54",
          6378 => x"58",
          6379 => x"74",
          6380 => x"75",
          6381 => x"00",
          6382 => x"54",
          6383 => x"58",
          6384 => x"74",
          6385 => x"75",
          6386 => x"00",
          6387 => x"74",
          6388 => x"20",
          6389 => x"74",
          6390 => x"72",
          6391 => x"0a",
          6392 => x"00",
          6393 => x"62",
          6394 => x"67",
          6395 => x"6d",
          6396 => x"2e",
          6397 => x"00",
          6398 => x"00",
          6399 => x"6c",
          6400 => x"74",
          6401 => x"6e",
          6402 => x"61",
          6403 => x"65",
          6404 => x"20",
          6405 => x"64",
          6406 => x"20",
          6407 => x"61",
          6408 => x"69",
          6409 => x"20",
          6410 => x"75",
          6411 => x"79",
          6412 => x"00",
          6413 => x"00",
          6414 => x"20",
          6415 => x"6b",
          6416 => x"21",
          6417 => x"00",
          6418 => x"74",
          6419 => x"69",
          6420 => x"2e",
          6421 => x"00",
          6422 => x"6c",
          6423 => x"74",
          6424 => x"6e",
          6425 => x"61",
          6426 => x"65",
          6427 => x"00",
          6428 => x"25",
          6429 => x"00",
          6430 => x"00",
          6431 => x"61",
          6432 => x"6e",
          6433 => x"6e",
          6434 => x"72",
          6435 => x"73",
          6436 => x"00",
          6437 => x"62",
          6438 => x"67",
          6439 => x"74",
          6440 => x"75",
          6441 => x"0a",
          6442 => x"00",
          6443 => x"61",
          6444 => x"64",
          6445 => x"72",
          6446 => x"69",
          6447 => x"00",
          6448 => x"62",
          6449 => x"67",
          6450 => x"72",
          6451 => x"69",
          6452 => x"00",
          6453 => x"63",
          6454 => x"6e",
          6455 => x"6f",
          6456 => x"40",
          6457 => x"38",
          6458 => x"2e",
          6459 => x"00",
          6460 => x"6c",
          6461 => x"20",
          6462 => x"65",
          6463 => x"25",
          6464 => x"20",
          6465 => x"0a",
          6466 => x"00",
          6467 => x"6c",
          6468 => x"74",
          6469 => x"65",
          6470 => x"6f",
          6471 => x"28",
          6472 => x"2e",
          6473 => x"00",
          6474 => x"74",
          6475 => x"69",
          6476 => x"61",
          6477 => x"69",
          6478 => x"69",
          6479 => x"2e",
          6480 => x"00",
          6481 => x"64",
          6482 => x"62",
          6483 => x"69",
          6484 => x"2e",
          6485 => x"00",
          6486 => x"00",
          6487 => x"00",
          6488 => x"5c",
          6489 => x"25",
          6490 => x"73",
          6491 => x"00",
          6492 => x"20",
          6493 => x"6d",
          6494 => x"2e",
          6495 => x"00",
          6496 => x"6e",
          6497 => x"2e",
          6498 => x"00",
          6499 => x"62",
          6500 => x"67",
          6501 => x"74",
          6502 => x"75",
          6503 => x"2e",
          6504 => x"00",
          6505 => x"00",
          6506 => x"00",
          6507 => x"ff",
          6508 => x"00",
          6509 => x"ff",
          6510 => x"00",
          6511 => x"ff",
          6512 => x"00",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"00",
          6517 => x"01",
          6518 => x"01",
          6519 => x"01",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"20",
          6524 => x"00",
          6525 => x"00",
          6526 => x"00",
          6527 => x"28",
          6528 => x"00",
          6529 => x"00",
          6530 => x"00",
          6531 => x"30",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"38",
          6536 => x"00",
          6537 => x"00",
          6538 => x"00",
          6539 => x"40",
          6540 => x"00",
          6541 => x"00",
          6542 => x"00",
          6543 => x"48",
          6544 => x"00",
          6545 => x"00",
          6546 => x"00",
          6547 => x"50",
          6548 => x"00",
          6549 => x"00",
          6550 => x"00",
          6551 => x"58",
          6552 => x"00",
          6553 => x"00",
          6554 => x"00",
          6555 => x"60",
          6556 => x"00",
          6557 => x"00",
          6558 => x"00",
          6559 => x"68",
          6560 => x"00",
          6561 => x"00",
          6562 => x"00",
          6563 => x"70",
          6564 => x"00",
          6565 => x"00",
          6566 => x"00",
          6567 => x"78",
          6568 => x"00",
          6569 => x"00",
          6570 => x"00",
          6571 => x"80",
          6572 => x"00",
          6573 => x"00",
          6574 => x"00",
          6575 => x"88",
          6576 => x"00",
          6577 => x"00",
          6578 => x"00",
          6579 => x"90",
          6580 => x"00",
          6581 => x"00",
          6582 => x"00",
          6583 => x"98",
          6584 => x"00",
          6585 => x"00",
          6586 => x"00",
          6587 => x"a4",
          6588 => x"00",
          6589 => x"00",
          6590 => x"00",
          6591 => x"ac",
          6592 => x"00",
          6593 => x"00",
          6594 => x"00",
          6595 => x"b4",
          6596 => x"00",
          6597 => x"00",
          6598 => x"00",
          6599 => x"bc",
          6600 => x"00",
          6601 => x"00",
          6602 => x"00",
          6603 => x"c4",
          6604 => x"00",
          6605 => x"00",
          6606 => x"00",
          6607 => x"cc",
          6608 => x"00",
          6609 => x"00",
          6610 => x"00",
          6611 => x"d4",
          6612 => x"00",
          6613 => x"00",
          6614 => x"00",
          6615 => x"dc",
          6616 => x"00",
          6617 => x"00",
          6618 => x"00",
          6619 => x"e4",
          6620 => x"00",
          6621 => x"00",
          6622 => x"00",
          6623 => x"ec",
          6624 => x"00",
          6625 => x"00",
          6626 => x"00",
          6627 => x"f4",
          6628 => x"00",
          6629 => x"00",
          6630 => x"00",
          6631 => x"fc",
          6632 => x"00",
          6633 => x"00",
          6634 => x"00",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"00",
          6639 => x"08",
          6640 => x"00",
          6641 => x"00",
          6642 => x"00",
          6643 => x"10",
          6644 => x"00",
          6645 => x"00",
          6646 => x"00",
          6647 => x"18",
          6648 => x"00",
          6649 => x"00",
          6650 => x"00",
          6651 => x"20",
          6652 => x"00",
          6653 => x"00",
          6654 => x"00",
          6655 => x"28",
          6656 => x"00",
          6657 => x"00",
          6658 => x"00",
          6659 => x"30",
          6660 => x"00",
          6661 => x"00",
          6662 => x"00",
          6663 => x"34",
          6664 => x"00",
          6665 => x"00",
          6666 => x"00",
          6667 => x"3c",
          6668 => x"00",
          6669 => x"00",
          6670 => x"00",
          6671 => x"48",
          6672 => x"00",
          6673 => x"00",
          6674 => x"00",
          6675 => x"50",
          6676 => x"00",
          6677 => x"00",
          6678 => x"00",
          6679 => x"58",
          6680 => x"00",
          6681 => x"00",
          6682 => x"00",
          6683 => x"60",
          6684 => x"00",
          6685 => x"00",
          6686 => x"00",
          6687 => x"68",
          6688 => x"00",
          6689 => x"00",
          6690 => x"00",
          6691 => x"6c",
          6692 => x"00",
          6693 => x"00",
          6694 => x"00",
          6695 => x"70",
          6696 => x"00",
          6697 => x"00",
          6698 => x"00",
          6699 => x"74",
          6700 => x"00",
          6701 => x"00",
          6702 => x"00",
          6703 => x"78",
          6704 => x"00",
          6705 => x"00",
          6706 => x"00",
          6707 => x"7c",
          6708 => x"00",
          6709 => x"00",
          6710 => x"00",
          6711 => x"80",
          6712 => x"00",
          6713 => x"00",
          6714 => x"00",
          6715 => x"84",
          6716 => x"00",
          6717 => x"00",
          6718 => x"00",
          6719 => x"88",
          6720 => x"00",
          6721 => x"00",
          6722 => x"00",
          6723 => x"8c",
          6724 => x"00",
          6725 => x"00",
          6726 => x"00",
          6727 => x"94",
          6728 => x"00",
          6729 => x"00",
          6730 => x"00",
          6731 => x"a0",
          6732 => x"00",
          6733 => x"00",
          6734 => x"00",
          6735 => x"a8",
          6736 => x"00",
          6737 => x"00",
          6738 => x"00",
          6739 => x"ac",
          6740 => x"00",
          6741 => x"00",
          6742 => x"00",
          6743 => x"b4",
          6744 => x"00",
          6745 => x"00",
          6746 => x"00",
          6747 => x"bc",
          6748 => x"00",
          6749 => x"00",
          6750 => x"00",
          6751 => x"c4",
          6752 => x"00",
          6753 => x"00",
          6754 => x"00",
          6755 => x"cc",
          6756 => x"00",
          6757 => x"00",
          6758 => x"00",
          6759 => x"d4",
          6760 => x"00",
          6761 => x"00",
          6762 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"fd",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"0b",
            10 => x"84",
            11 => x"0b",
            12 => x"0b",
            13 => x"a2",
            14 => x"0b",
            15 => x"0b",
            16 => x"c0",
            17 => x"0b",
            18 => x"0b",
            19 => x"de",
            20 => x"0b",
            21 => x"0b",
            22 => x"fc",
            23 => x"0b",
            24 => x"0b",
            25 => x"9a",
            26 => x"0b",
            27 => x"0b",
            28 => x"b8",
            29 => x"0b",
            30 => x"0b",
            31 => x"d6",
            32 => x"0b",
            33 => x"0b",
            34 => x"f4",
            35 => x"0b",
            36 => x"0b",
            37 => x"93",
            38 => x"0b",
            39 => x"0b",
            40 => x"b3",
            41 => x"0b",
            42 => x"0b",
            43 => x"d3",
            44 => x"0b",
            45 => x"0b",
            46 => x"f3",
            47 => x"0b",
            48 => x"0b",
            49 => x"93",
            50 => x"0b",
            51 => x"0b",
            52 => x"b3",
            53 => x"0b",
            54 => x"0b",
            55 => x"d3",
            56 => x"0b",
            57 => x"0b",
            58 => x"f3",
            59 => x"0b",
            60 => x"0b",
            61 => x"93",
            62 => x"0b",
            63 => x"0b",
            64 => x"b3",
            65 => x"0b",
            66 => x"0b",
            67 => x"d3",
            68 => x"0b",
            69 => x"0b",
            70 => x"f3",
            71 => x"0b",
            72 => x"0b",
            73 => x"93",
            74 => x"0b",
            75 => x"0b",
            76 => x"b1",
            77 => x"0b",
            78 => x"0b",
            79 => x"cf",
            80 => x"0b",
            81 => x"0b",
            82 => x"ed",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"80",
           129 => x"b8",
           130 => x"2d",
           131 => x"08",
           132 => x"04",
           133 => x"0c",
           134 => x"81",
           135 => x"83",
           136 => x"81",
           137 => x"9f",
           138 => x"d3",
           139 => x"80",
           140 => x"d3",
           141 => x"8a",
           142 => x"b8",
           143 => x"90",
           144 => x"b8",
           145 => x"2d",
           146 => x"08",
           147 => x"04",
           148 => x"0c",
           149 => x"81",
           150 => x"83",
           151 => x"81",
           152 => x"a0",
           153 => x"d3",
           154 => x"80",
           155 => x"d3",
           156 => x"8f",
           157 => x"b8",
           158 => x"90",
           159 => x"b8",
           160 => x"2d",
           161 => x"08",
           162 => x"04",
           163 => x"0c",
           164 => x"81",
           165 => x"83",
           166 => x"81",
           167 => x"a6",
           168 => x"d3",
           169 => x"80",
           170 => x"d3",
           171 => x"be",
           172 => x"b8",
           173 => x"90",
           174 => x"b8",
           175 => x"2d",
           176 => x"08",
           177 => x"04",
           178 => x"0c",
           179 => x"81",
           180 => x"83",
           181 => x"81",
           182 => x"8f",
           183 => x"d3",
           184 => x"80",
           185 => x"d3",
           186 => x"f7",
           187 => x"b8",
           188 => x"90",
           189 => x"b8",
           190 => x"2d",
           191 => x"08",
           192 => x"04",
           193 => x"0c",
           194 => x"2d",
           195 => x"08",
           196 => x"04",
           197 => x"0c",
           198 => x"2d",
           199 => x"08",
           200 => x"04",
           201 => x"0c",
           202 => x"2d",
           203 => x"08",
           204 => x"04",
           205 => x"0c",
           206 => x"2d",
           207 => x"08",
           208 => x"04",
           209 => x"0c",
           210 => x"2d",
           211 => x"08",
           212 => x"04",
           213 => x"0c",
           214 => x"2d",
           215 => x"08",
           216 => x"04",
           217 => x"0c",
           218 => x"2d",
           219 => x"08",
           220 => x"04",
           221 => x"0c",
           222 => x"2d",
           223 => x"08",
           224 => x"04",
           225 => x"0c",
           226 => x"2d",
           227 => x"08",
           228 => x"04",
           229 => x"0c",
           230 => x"2d",
           231 => x"08",
           232 => x"04",
           233 => x"0c",
           234 => x"2d",
           235 => x"08",
           236 => x"04",
           237 => x"0c",
           238 => x"2d",
           239 => x"08",
           240 => x"04",
           241 => x"0c",
           242 => x"2d",
           243 => x"08",
           244 => x"04",
           245 => x"0c",
           246 => x"2d",
           247 => x"08",
           248 => x"04",
           249 => x"0c",
           250 => x"2d",
           251 => x"08",
           252 => x"04",
           253 => x"0c",
           254 => x"2d",
           255 => x"08",
           256 => x"04",
           257 => x"0c",
           258 => x"2d",
           259 => x"08",
           260 => x"04",
           261 => x"0c",
           262 => x"2d",
           263 => x"08",
           264 => x"04",
           265 => x"0c",
           266 => x"2d",
           267 => x"08",
           268 => x"04",
           269 => x"0c",
           270 => x"2d",
           271 => x"08",
           272 => x"04",
           273 => x"0c",
           274 => x"2d",
           275 => x"08",
           276 => x"04",
           277 => x"0c",
           278 => x"2d",
           279 => x"08",
           280 => x"04",
           281 => x"0c",
           282 => x"2d",
           283 => x"08",
           284 => x"04",
           285 => x"0c",
           286 => x"2d",
           287 => x"08",
           288 => x"04",
           289 => x"0c",
           290 => x"2d",
           291 => x"08",
           292 => x"04",
           293 => x"0c",
           294 => x"81",
           295 => x"83",
           296 => x"81",
           297 => x"af",
           298 => x"d3",
           299 => x"80",
           300 => x"d3",
           301 => x"98",
           302 => x"b8",
           303 => x"90",
           304 => x"b8",
           305 => x"2d",
           306 => x"08",
           307 => x"04",
           308 => x"0c",
           309 => x"81",
           310 => x"83",
           311 => x"81",
           312 => x"93",
           313 => x"d3",
           314 => x"80",
           315 => x"d3",
           316 => x"9f",
           317 => x"d3",
           318 => x"80",
           319 => x"d3",
           320 => x"f6",
           321 => x"38",
           322 => x"84",
           323 => x"0b",
           324 => x"80",
           325 => x"51",
           326 => x"04",
           327 => x"d3",
           328 => x"81",
           329 => x"fd",
           330 => x"53",
           331 => x"08",
           332 => x"52",
           333 => x"08",
           334 => x"51",
           335 => x"81",
           336 => x"70",
           337 => x"0c",
           338 => x"0d",
           339 => x"0c",
           340 => x"b8",
           341 => x"d3",
           342 => x"3d",
           343 => x"81",
           344 => x"8c",
           345 => x"81",
           346 => x"88",
           347 => x"93",
           348 => x"ac",
           349 => x"d3",
           350 => x"85",
           351 => x"d3",
           352 => x"81",
           353 => x"02",
           354 => x"0c",
           355 => x"81",
           356 => x"b8",
           357 => x"0c",
           358 => x"d3",
           359 => x"05",
           360 => x"b8",
           361 => x"08",
           362 => x"08",
           363 => x"27",
           364 => x"d3",
           365 => x"05",
           366 => x"ae",
           367 => x"81",
           368 => x"8c",
           369 => x"a2",
           370 => x"b8",
           371 => x"08",
           372 => x"b8",
           373 => x"0c",
           374 => x"08",
           375 => x"10",
           376 => x"08",
           377 => x"ff",
           378 => x"d3",
           379 => x"05",
           380 => x"80",
           381 => x"d3",
           382 => x"05",
           383 => x"b8",
           384 => x"08",
           385 => x"81",
           386 => x"88",
           387 => x"d3",
           388 => x"05",
           389 => x"d3",
           390 => x"05",
           391 => x"b8",
           392 => x"08",
           393 => x"08",
           394 => x"07",
           395 => x"08",
           396 => x"81",
           397 => x"fc",
           398 => x"2a",
           399 => x"08",
           400 => x"81",
           401 => x"8c",
           402 => x"2a",
           403 => x"08",
           404 => x"ff",
           405 => x"d3",
           406 => x"05",
           407 => x"93",
           408 => x"b8",
           409 => x"08",
           410 => x"b8",
           411 => x"0c",
           412 => x"81",
           413 => x"f8",
           414 => x"81",
           415 => x"f4",
           416 => x"81",
           417 => x"f4",
           418 => x"d3",
           419 => x"3d",
           420 => x"b8",
           421 => x"3d",
           422 => x"71",
           423 => x"9f",
           424 => x"55",
           425 => x"72",
           426 => x"74",
           427 => x"70",
           428 => x"38",
           429 => x"71",
           430 => x"38",
           431 => x"81",
           432 => x"ff",
           433 => x"ff",
           434 => x"06",
           435 => x"81",
           436 => x"86",
           437 => x"74",
           438 => x"75",
           439 => x"90",
           440 => x"54",
           441 => x"27",
           442 => x"71",
           443 => x"53",
           444 => x"70",
           445 => x"0c",
           446 => x"84",
           447 => x"72",
           448 => x"05",
           449 => x"12",
           450 => x"26",
           451 => x"72",
           452 => x"72",
           453 => x"05",
           454 => x"12",
           455 => x"26",
           456 => x"53",
           457 => x"fb",
           458 => x"79",
           459 => x"83",
           460 => x"52",
           461 => x"71",
           462 => x"54",
           463 => x"73",
           464 => x"c6",
           465 => x"54",
           466 => x"70",
           467 => x"52",
           468 => x"2e",
           469 => x"33",
           470 => x"2e",
           471 => x"95",
           472 => x"81",
           473 => x"70",
           474 => x"54",
           475 => x"70",
           476 => x"33",
           477 => x"ff",
           478 => x"ff",
           479 => x"31",
           480 => x"0c",
           481 => x"3d",
           482 => x"09",
           483 => x"fd",
           484 => x"70",
           485 => x"81",
           486 => x"51",
           487 => x"38",
           488 => x"16",
           489 => x"56",
           490 => x"08",
           491 => x"73",
           492 => x"ff",
           493 => x"0b",
           494 => x"0c",
           495 => x"04",
           496 => x"80",
           497 => x"71",
           498 => x"87",
           499 => x"d3",
           500 => x"ff",
           501 => x"81",
           502 => x"83",
           503 => x"38",
           504 => x"ac",
           505 => x"0d",
           506 => x"0d",
           507 => x"70",
           508 => x"73",
           509 => x"cd",
           510 => x"51",
           511 => x"09",
           512 => x"38",
           513 => x"33",
           514 => x"a0",
           515 => x"73",
           516 => x"81",
           517 => x"72",
           518 => x"70",
           519 => x"38",
           520 => x"30",
           521 => x"74",
           522 => x"70",
           523 => x"33",
           524 => x"2e",
           525 => x"88",
           526 => x"70",
           527 => x"34",
           528 => x"73",
           529 => x"d3",
           530 => x"3d",
           531 => x"3d",
           532 => x"72",
           533 => x"91",
           534 => x"fc",
           535 => x"51",
           536 => x"81",
           537 => x"85",
           538 => x"83",
           539 => x"72",
           540 => x"0c",
           541 => x"04",
           542 => x"7d",
           543 => x"ff",
           544 => x"81",
           545 => x"26",
           546 => x"83",
           547 => x"05",
           548 => x"79",
           549 => x"b1",
           550 => x"33",
           551 => x"79",
           552 => x"a5",
           553 => x"33",
           554 => x"79",
           555 => x"99",
           556 => x"33",
           557 => x"79",
           558 => x"8d",
           559 => x"22",
           560 => x"79",
           561 => x"81",
           562 => x"1c",
           563 => x"5b",
           564 => x"26",
           565 => x"8a",
           566 => x"88",
           567 => x"86",
           568 => x"85",
           569 => x"84",
           570 => x"83",
           571 => x"82",
           572 => x"7b",
           573 => x"b6",
           574 => x"89",
           575 => x"98",
           576 => x"7b",
           577 => x"87",
           578 => x"0c",
           579 => x"87",
           580 => x"0c",
           581 => x"87",
           582 => x"0c",
           583 => x"87",
           584 => x"0c",
           585 => x"87",
           586 => x"0c",
           587 => x"87",
           588 => x"0c",
           589 => x"87",
           590 => x"0c",
           591 => x"87",
           592 => x"0c",
           593 => x"80",
           594 => x"d3",
           595 => x"3d",
           596 => x"3d",
           597 => x"87",
           598 => x"5c",
           599 => x"87",
           600 => x"08",
           601 => x"23",
           602 => x"b8",
           603 => x"82",
           604 => x"c0",
           605 => x"5b",
           606 => x"34",
           607 => x"b0",
           608 => x"84",
           609 => x"c0",
           610 => x"5b",
           611 => x"34",
           612 => x"a8",
           613 => x"86",
           614 => x"c0",
           615 => x"5b",
           616 => x"23",
           617 => x"a0",
           618 => x"8a",
           619 => x"7c",
           620 => x"22",
           621 => x"22",
           622 => x"33",
           623 => x"33",
           624 => x"33",
           625 => x"33",
           626 => x"33",
           627 => x"52",
           628 => x"51",
           629 => x"8d",
           630 => x"80",
           631 => x"8b",
           632 => x"30",
           633 => x"51",
           634 => x"0b",
           635 => x"a4",
           636 => x"0d",
           637 => x"0d",
           638 => x"81",
           639 => x"54",
           640 => x"94",
           641 => x"80",
           642 => x"87",
           643 => x"51",
           644 => x"96",
           645 => x"06",
           646 => x"70",
           647 => x"38",
           648 => x"70",
           649 => x"51",
           650 => x"71",
           651 => x"32",
           652 => x"51",
           653 => x"2e",
           654 => x"93",
           655 => x"06",
           656 => x"ff",
           657 => x"0b",
           658 => x"33",
           659 => x"94",
           660 => x"80",
           661 => x"87",
           662 => x"52",
           663 => x"73",
           664 => x"0c",
           665 => x"04",
           666 => x"02",
           667 => x"0b",
           668 => x"a4",
           669 => x"87",
           670 => x"51",
           671 => x"86",
           672 => x"94",
           673 => x"08",
           674 => x"70",
           675 => x"52",
           676 => x"2e",
           677 => x"91",
           678 => x"06",
           679 => x"d7",
           680 => x"2a",
           681 => x"81",
           682 => x"70",
           683 => x"38",
           684 => x"70",
           685 => x"51",
           686 => x"38",
           687 => x"cb",
           688 => x"87",
           689 => x"52",
           690 => x"86",
           691 => x"94",
           692 => x"72",
           693 => x"0d",
           694 => x"0d",
           695 => x"74",
           696 => x"70",
           697 => x"f7",
           698 => x"81",
           699 => x"0b",
           700 => x"a4",
           701 => x"87",
           702 => x"51",
           703 => x"86",
           704 => x"94",
           705 => x"08",
           706 => x"70",
           707 => x"52",
           708 => x"2e",
           709 => x"91",
           710 => x"06",
           711 => x"d7",
           712 => x"2a",
           713 => x"81",
           714 => x"70",
           715 => x"38",
           716 => x"70",
           717 => x"51",
           718 => x"38",
           719 => x"cb",
           720 => x"87",
           721 => x"52",
           722 => x"86",
           723 => x"94",
           724 => x"72",
           725 => x"74",
           726 => x"70",
           727 => x"75",
           728 => x"0c",
           729 => x"04",
           730 => x"0b",
           731 => x"a4",
           732 => x"c0",
           733 => x"71",
           734 => x"38",
           735 => x"94",
           736 => x"70",
           737 => x"81",
           738 => x"51",
           739 => x"e2",
           740 => x"81",
           741 => x"51",
           742 => x"80",
           743 => x"2e",
           744 => x"c0",
           745 => x"71",
           746 => x"ff",
           747 => x"ac",
           748 => x"3d",
           749 => x"3d",
           750 => x"81",
           751 => x"51",
           752 => x"84",
           753 => x"2e",
           754 => x"c0",
           755 => x"71",
           756 => x"2a",
           757 => x"51",
           758 => x"52",
           759 => x"a2",
           760 => x"81",
           761 => x"51",
           762 => x"80",
           763 => x"2e",
           764 => x"c0",
           765 => x"71",
           766 => x"2b",
           767 => x"51",
           768 => x"81",
           769 => x"83",
           770 => x"fd",
           771 => x"c0",
           772 => x"08",
           773 => x"8a",
           774 => x"53",
           775 => x"83",
           776 => x"cb",
           777 => x"c0",
           778 => x"71",
           779 => x"87",
           780 => x"08",
           781 => x"88",
           782 => x"9e",
           783 => x"0c",
           784 => x"87",
           785 => x"08",
           786 => x"90",
           787 => x"9e",
           788 => x"0c",
           789 => x"87",
           790 => x"08",
           791 => x"98",
           792 => x"9e",
           793 => x"0c",
           794 => x"87",
           795 => x"08",
           796 => x"a0",
           797 => x"9e",
           798 => x"0c",
           799 => x"52",
           800 => x"13",
           801 => x"87",
           802 => x"08",
           803 => x"81",
           804 => x"34",
           805 => x"80",
           806 => x"9e",
           807 => x"a0",
           808 => x"52",
           809 => x"2e",
           810 => x"53",
           811 => x"80",
           812 => x"9e",
           813 => x"81",
           814 => x"51",
           815 => x"80",
           816 => x"81",
           817 => x"cb",
           818 => x"0b",
           819 => x"88",
           820 => x"c0",
           821 => x"52",
           822 => x"2e",
           823 => x"52",
           824 => x"d7",
           825 => x"87",
           826 => x"08",
           827 => x"06",
           828 => x"70",
           829 => x"38",
           830 => x"81",
           831 => x"80",
           832 => x"9e",
           833 => x"88",
           834 => x"52",
           835 => x"2e",
           836 => x"52",
           837 => x"d9",
           838 => x"87",
           839 => x"08",
           840 => x"06",
           841 => x"70",
           842 => x"38",
           843 => x"81",
           844 => x"80",
           845 => x"9e",
           846 => x"82",
           847 => x"52",
           848 => x"2e",
           849 => x"52",
           850 => x"db",
           851 => x"87",
           852 => x"08",
           853 => x"06",
           854 => x"70",
           855 => x"38",
           856 => x"81",
           857 => x"81",
           858 => x"87",
           859 => x"70",
           860 => x"e0",
           861 => x"2c",
           862 => x"53",
           863 => x"81",
           864 => x"71",
           865 => x"08",
           866 => x"51",
           867 => x"80",
           868 => x"81",
           869 => x"34",
           870 => x"c0",
           871 => x"70",
           872 => x"52",
           873 => x"2e",
           874 => x"52",
           875 => x"df",
           876 => x"9e",
           877 => x"87",
           878 => x"70",
           879 => x"34",
           880 => x"04",
           881 => x"81",
           882 => x"84",
           883 => x"cb",
           884 => x"73",
           885 => x"38",
           886 => x"51",
           887 => x"81",
           888 => x"84",
           889 => x"cb",
           890 => x"55",
           891 => x"2e",
           892 => x"15",
           893 => x"cb",
           894 => x"81",
           895 => x"8a",
           896 => x"cb",
           897 => x"55",
           898 => x"2e",
           899 => x"15",
           900 => x"15",
           901 => x"b7",
           902 => x"e9",
           903 => x"d7",
           904 => x"55",
           905 => x"81",
           906 => x"73",
           907 => x"38",
           908 => x"70",
           909 => x"11",
           910 => x"81",
           911 => x"89",
           912 => x"cb",
           913 => x"73",
           914 => x"38",
           915 => x"51",
           916 => x"81",
           917 => x"54",
           918 => x"88",
           919 => x"e0",
           920 => x"3f",
           921 => x"33",
           922 => x"2e",
           923 => x"b7",
           924 => x"97",
           925 => x"dc",
           926 => x"55",
           927 => x"8c",
           928 => x"33",
           929 => x"f8",
           930 => x"3f",
           931 => x"33",
           932 => x"2e",
           933 => x"b8",
           934 => x"ef",
           935 => x"df",
           936 => x"55",
           937 => x"8c",
           938 => x"33",
           939 => x"b4",
           940 => x"3f",
           941 => x"51",
           942 => x"81",
           943 => x"70",
           944 => x"52",
           945 => x"b8",
           946 => x"55",
           947 => x"73",
           948 => x"b9",
           949 => x"ad",
           950 => x"08",
           951 => x"ac",
           952 => x"3f",
           953 => x"52",
           954 => x"51",
           955 => x"90",
           956 => x"81",
           957 => x"88",
           958 => x"3d",
           959 => x"3d",
           960 => x"05",
           961 => x"85",
           962 => x"71",
           963 => x"0b",
           964 => x"05",
           965 => x"04",
           966 => x"51",
           967 => x"ac",
           968 => x"ac",
           969 => x"3f",
           970 => x"ba",
           971 => x"a9",
           972 => x"81",
           973 => x"f7",
           974 => x"39",
           975 => x"51",
           976 => x"88",
           977 => x"c8",
           978 => x"3f",
           979 => x"04",
           980 => x"0c",
           981 => x"87",
           982 => x"0c",
           983 => x"0d",
           984 => x"84",
           985 => x"52",
           986 => x"70",
           987 => x"81",
           988 => x"72",
           989 => x"0d",
           990 => x"0d",
           991 => x"84",
           992 => x"cb",
           993 => x"80",
           994 => x"09",
           995 => x"e4",
           996 => x"81",
           997 => x"73",
           998 => x"3d",
           999 => x"cb",
          1000 => x"c0",
          1001 => x"04",
          1002 => x"02",
          1003 => x"53",
          1004 => x"09",
          1005 => x"38",
          1006 => x"3f",
          1007 => x"08",
          1008 => x"38",
          1009 => x"08",
          1010 => x"34",
          1011 => x"08",
          1012 => x"d3",
          1013 => x"39",
          1014 => x"08",
          1015 => x"38",
          1016 => x"d3",
          1017 => x"71",
          1018 => x"0d",
          1019 => x"0d",
          1020 => x"33",
          1021 => x"08",
          1022 => x"bc",
          1023 => x"ff",
          1024 => x"81",
          1025 => x"84",
          1026 => x"fe",
          1027 => x"70",
          1028 => x"71",
          1029 => x"38",
          1030 => x"05",
          1031 => x"ff",
          1032 => x"33",
          1033 => x"38",
          1034 => x"04",
          1035 => x"76",
          1036 => x"08",
          1037 => x"bc",
          1038 => x"54",
          1039 => x"80",
          1040 => x"72",
          1041 => x"54",
          1042 => x"dc",
          1043 => x"52",
          1044 => x"73",
          1045 => x"0c",
          1046 => x"04",
          1047 => x"66",
          1048 => x"78",
          1049 => x"5a",
          1050 => x"80",
          1051 => x"38",
          1052 => x"88",
          1053 => x"fe",
          1054 => x"39",
          1055 => x"70",
          1056 => x"33",
          1057 => x"75",
          1058 => x"81",
          1059 => x"81",
          1060 => x"05",
          1061 => x"5d",
          1062 => x"ad",
          1063 => x"06",
          1064 => x"79",
          1065 => x"5b",
          1066 => x"75",
          1067 => x"81",
          1068 => x"7b",
          1069 => x"08",
          1070 => x"05",
          1071 => x"5c",
          1072 => x"39",
          1073 => x"72",
          1074 => x"38",
          1075 => x"16",
          1076 => x"70",
          1077 => x"33",
          1078 => x"57",
          1079 => x"27",
          1080 => x"80",
          1081 => x"30",
          1082 => x"80",
          1083 => x"cc",
          1084 => x"70",
          1085 => x"25",
          1086 => x"59",
          1087 => x"54",
          1088 => x"8c",
          1089 => x"07",
          1090 => x"05",
          1091 => x"5d",
          1092 => x"83",
          1093 => x"55",
          1094 => x"27",
          1095 => x"16",
          1096 => x"06",
          1097 => x"be",
          1098 => x"96",
          1099 => x"38",
          1100 => x"81",
          1101 => x"53",
          1102 => x"7b",
          1103 => x"08",
          1104 => x"80",
          1105 => x"54",
          1106 => x"8d",
          1107 => x"70",
          1108 => x"51",
          1109 => x"f5",
          1110 => x"2a",
          1111 => x"51",
          1112 => x"38",
          1113 => x"55",
          1114 => x"27",
          1115 => x"81",
          1116 => x"56",
          1117 => x"b0",
          1118 => x"38",
          1119 => x"55",
          1120 => x"26",
          1121 => x"51",
          1122 => x"73",
          1123 => x"53",
          1124 => x"fd",
          1125 => x"51",
          1126 => x"73",
          1127 => x"53",
          1128 => x"f2",
          1129 => x"39",
          1130 => x"83",
          1131 => x"5d",
          1132 => x"3f",
          1133 => x"82",
          1134 => x"88",
          1135 => x"8a",
          1136 => x"90",
          1137 => x"75",
          1138 => x"3f",
          1139 => x"7c",
          1140 => x"81",
          1141 => x"72",
          1142 => x"38",
          1143 => x"71",
          1144 => x"53",
          1145 => x"80",
          1146 => x"81",
          1147 => x"7b",
          1148 => x"08",
          1149 => x"89",
          1150 => x"1d",
          1151 => x"5d",
          1152 => x"c4",
          1153 => x"70",
          1154 => x"25",
          1155 => x"24",
          1156 => x"55",
          1157 => x"2e",
          1158 => x"30",
          1159 => x"5e",
          1160 => x"7a",
          1161 => x"e6",
          1162 => x"d3",
          1163 => x"ff",
          1164 => x"77",
          1165 => x"e6",
          1166 => x"ac",
          1167 => x"75",
          1168 => x"74",
          1169 => x"81",
          1170 => x"54",
          1171 => x"f8",
          1172 => x"87",
          1173 => x"ff",
          1174 => x"96",
          1175 => x"e0",
          1176 => x"54",
          1177 => x"34",
          1178 => x"30",
          1179 => x"9f",
          1180 => x"74",
          1181 => x"51",
          1182 => x"ff",
          1183 => x"84",
          1184 => x"06",
          1185 => x"80",
          1186 => x"96",
          1187 => x"e0",
          1188 => x"73",
          1189 => x"58",
          1190 => x"06",
          1191 => x"55",
          1192 => x"a0",
          1193 => x"2a",
          1194 => x"51",
          1195 => x"38",
          1196 => x"55",
          1197 => x"27",
          1198 => x"81",
          1199 => x"56",
          1200 => x"e4",
          1201 => x"38",
          1202 => x"55",
          1203 => x"26",
          1204 => x"18",
          1205 => x"05",
          1206 => x"53",
          1207 => x"c8",
          1208 => x"38",
          1209 => x"55",
          1210 => x"27",
          1211 => x"a0",
          1212 => x"3f",
          1213 => x"55",
          1214 => x"26",
          1215 => x"e3",
          1216 => x"0d",
          1217 => x"0d",
          1218 => x"70",
          1219 => x"08",
          1220 => x"51",
          1221 => x"85",
          1222 => x"fe",
          1223 => x"81",
          1224 => x"85",
          1225 => x"52",
          1226 => x"b0",
          1227 => x"c4",
          1228 => x"73",
          1229 => x"81",
          1230 => x"84",
          1231 => x"fd",
          1232 => x"d3",
          1233 => x"81",
          1234 => x"87",
          1235 => x"53",
          1236 => x"fa",
          1237 => x"81",
          1238 => x"85",
          1239 => x"fa",
          1240 => x"7a",
          1241 => x"53",
          1242 => x"08",
          1243 => x"fa",
          1244 => x"73",
          1245 => x"39",
          1246 => x"d3",
          1247 => x"71",
          1248 => x"ac",
          1249 => x"06",
          1250 => x"2e",
          1251 => x"8d",
          1252 => x"38",
          1253 => x"70",
          1254 => x"70",
          1255 => x"2a",
          1256 => x"06",
          1257 => x"53",
          1258 => x"8e",
          1259 => x"74",
          1260 => x"52",
          1261 => x"3f",
          1262 => x"74",
          1263 => x"38",
          1264 => x"74",
          1265 => x"b2",
          1266 => x"52",
          1267 => x"81",
          1268 => x"ff",
          1269 => x"f7",
          1270 => x"9e",
          1271 => x"52",
          1272 => x"8a",
          1273 => x"3f",
          1274 => x"81",
          1275 => x"88",
          1276 => x"fe",
          1277 => x"d3",
          1278 => x"81",
          1279 => x"77",
          1280 => x"53",
          1281 => x"72",
          1282 => x"0c",
          1283 => x"04",
          1284 => x"7a",
          1285 => x"80",
          1286 => x"75",
          1287 => x"56",
          1288 => x"a0",
          1289 => x"06",
          1290 => x"08",
          1291 => x"0c",
          1292 => x"33",
          1293 => x"a0",
          1294 => x"73",
          1295 => x"81",
          1296 => x"81",
          1297 => x"76",
          1298 => x"70",
          1299 => x"58",
          1300 => x"09",
          1301 => x"d3",
          1302 => x"81",
          1303 => x"74",
          1304 => x"55",
          1305 => x"e2",
          1306 => x"73",
          1307 => x"09",
          1308 => x"38",
          1309 => x"14",
          1310 => x"08",
          1311 => x"54",
          1312 => x"39",
          1313 => x"81",
          1314 => x"75",
          1315 => x"56",
          1316 => x"39",
          1317 => x"74",
          1318 => x"38",
          1319 => x"80",
          1320 => x"89",
          1321 => x"38",
          1322 => x"d0",
          1323 => x"56",
          1324 => x"80",
          1325 => x"39",
          1326 => x"e1",
          1327 => x"80",
          1328 => x"57",
          1329 => x"74",
          1330 => x"38",
          1331 => x"27",
          1332 => x"14",
          1333 => x"06",
          1334 => x"14",
          1335 => x"06",
          1336 => x"74",
          1337 => x"f9",
          1338 => x"ff",
          1339 => x"89",
          1340 => x"38",
          1341 => x"c5",
          1342 => x"29",
          1343 => x"81",
          1344 => x"75",
          1345 => x"56",
          1346 => x"a0",
          1347 => x"38",
          1348 => x"84",
          1349 => x"56",
          1350 => x"81",
          1351 => x"d3",
          1352 => x"3d",
          1353 => x"3d",
          1354 => x"5a",
          1355 => x"7a",
          1356 => x"70",
          1357 => x"58",
          1358 => x"09",
          1359 => x"38",
          1360 => x"05",
          1361 => x"08",
          1362 => x"53",
          1363 => x"f0",
          1364 => x"2e",
          1365 => x"8e",
          1366 => x"08",
          1367 => x"75",
          1368 => x"56",
          1369 => x"b0",
          1370 => x"06",
          1371 => x"74",
          1372 => x"75",
          1373 => x"70",
          1374 => x"73",
          1375 => x"9a",
          1376 => x"f8",
          1377 => x"06",
          1378 => x"0b",
          1379 => x"0c",
          1380 => x"33",
          1381 => x"80",
          1382 => x"75",
          1383 => x"76",
          1384 => x"70",
          1385 => x"57",
          1386 => x"56",
          1387 => x"81",
          1388 => x"14",
          1389 => x"88",
          1390 => x"27",
          1391 => x"f3",
          1392 => x"53",
          1393 => x"89",
          1394 => x"38",
          1395 => x"56",
          1396 => x"80",
          1397 => x"39",
          1398 => x"56",
          1399 => x"80",
          1400 => x"e0",
          1401 => x"38",
          1402 => x"81",
          1403 => x"53",
          1404 => x"81",
          1405 => x"53",
          1406 => x"8e",
          1407 => x"70",
          1408 => x"55",
          1409 => x"27",
          1410 => x"77",
          1411 => x"76",
          1412 => x"75",
          1413 => x"76",
          1414 => x"70",
          1415 => x"56",
          1416 => x"ff",
          1417 => x"80",
          1418 => x"75",
          1419 => x"79",
          1420 => x"75",
          1421 => x"0c",
          1422 => x"04",
          1423 => x"02",
          1424 => x"51",
          1425 => x"72",
          1426 => x"81",
          1427 => x"33",
          1428 => x"d3",
          1429 => x"3d",
          1430 => x"3d",
          1431 => x"05",
          1432 => x"05",
          1433 => x"55",
          1434 => x"72",
          1435 => x"ed",
          1436 => x"29",
          1437 => x"8c",
          1438 => x"52",
          1439 => x"84",
          1440 => x"52",
          1441 => x"72",
          1442 => x"c0",
          1443 => x"51",
          1444 => x"85",
          1445 => x"98",
          1446 => x"52",
          1447 => x"8c",
          1448 => x"70",
          1449 => x"51",
          1450 => x"87",
          1451 => x"51",
          1452 => x"72",
          1453 => x"c0",
          1454 => x"70",
          1455 => x"80",
          1456 => x"71",
          1457 => x"c0",
          1458 => x"51",
          1459 => x"87",
          1460 => x"cb",
          1461 => x"81",
          1462 => x"33",
          1463 => x"d3",
          1464 => x"3d",
          1465 => x"3d",
          1466 => x"65",
          1467 => x"80",
          1468 => x"56",
          1469 => x"83",
          1470 => x"fe",
          1471 => x"d3",
          1472 => x"06",
          1473 => x"71",
          1474 => x"80",
          1475 => x"87",
          1476 => x"73",
          1477 => x"c0",
          1478 => x"87",
          1479 => x"12",
          1480 => x"57",
          1481 => x"76",
          1482 => x"92",
          1483 => x"71",
          1484 => x"75",
          1485 => x"70",
          1486 => x"81",
          1487 => x"54",
          1488 => x"8e",
          1489 => x"52",
          1490 => x"81",
          1491 => x"81",
          1492 => x"a2",
          1493 => x"80",
          1494 => x"75",
          1495 => x"d5",
          1496 => x"52",
          1497 => x"87",
          1498 => x"80",
          1499 => x"81",
          1500 => x"c0",
          1501 => x"53",
          1502 => x"82",
          1503 => x"71",
          1504 => x"1b",
          1505 => x"84",
          1506 => x"1e",
          1507 => x"06",
          1508 => x"7a",
          1509 => x"38",
          1510 => x"80",
          1511 => x"87",
          1512 => x"26",
          1513 => x"73",
          1514 => x"06",
          1515 => x"2e",
          1516 => x"52",
          1517 => x"81",
          1518 => x"90",
          1519 => x"f3",
          1520 => x"62",
          1521 => x"05",
          1522 => x"56",
          1523 => x"83",
          1524 => x"fc",
          1525 => x"d3",
          1526 => x"06",
          1527 => x"71",
          1528 => x"80",
          1529 => x"98",
          1530 => x"2b",
          1531 => x"8c",
          1532 => x"92",
          1533 => x"41",
          1534 => x"56",
          1535 => x"87",
          1536 => x"19",
          1537 => x"52",
          1538 => x"80",
          1539 => x"70",
          1540 => x"81",
          1541 => x"54",
          1542 => x"8c",
          1543 => x"81",
          1544 => x"78",
          1545 => x"53",
          1546 => x"70",
          1547 => x"52",
          1548 => x"87",
          1549 => x"52",
          1550 => x"75",
          1551 => x"80",
          1552 => x"72",
          1553 => x"99",
          1554 => x"0c",
          1555 => x"8c",
          1556 => x"08",
          1557 => x"51",
          1558 => x"38",
          1559 => x"8d",
          1560 => x"70",
          1561 => x"84",
          1562 => x"5d",
          1563 => x"2e",
          1564 => x"fc",
          1565 => x"52",
          1566 => x"7d",
          1567 => x"fc",
          1568 => x"80",
          1569 => x"71",
          1570 => x"38",
          1571 => x"54",
          1572 => x"ac",
          1573 => x"0d",
          1574 => x"0d",
          1575 => x"05",
          1576 => x"02",
          1577 => x"05",
          1578 => x"55",
          1579 => x"8c",
          1580 => x"ac",
          1581 => x"52",
          1582 => x"bc",
          1583 => x"72",
          1584 => x"38",
          1585 => x"88",
          1586 => x"2e",
          1587 => x"39",
          1588 => x"9a",
          1589 => x"74",
          1590 => x"c0",
          1591 => x"70",
          1592 => x"94",
          1593 => x"0a",
          1594 => x"54",
          1595 => x"80",
          1596 => x"54",
          1597 => x"54",
          1598 => x"ac",
          1599 => x"0d",
          1600 => x"0d",
          1601 => x"81",
          1602 => x"88",
          1603 => x"81",
          1604 => x"52",
          1605 => x"3d",
          1606 => x"3d",
          1607 => x"11",
          1608 => x"33",
          1609 => x"71",
          1610 => x"81",
          1611 => x"07",
          1612 => x"88",
          1613 => x"d3",
          1614 => x"54",
          1615 => x"85",
          1616 => x"ff",
          1617 => x"02",
          1618 => x"05",
          1619 => x"70",
          1620 => x"05",
          1621 => x"88",
          1622 => x"72",
          1623 => x"0d",
          1624 => x"0d",
          1625 => x"52",
          1626 => x"81",
          1627 => x"70",
          1628 => x"70",
          1629 => x"05",
          1630 => x"88",
          1631 => x"72",
          1632 => x"54",
          1633 => x"2a",
          1634 => x"34",
          1635 => x"04",
          1636 => x"76",
          1637 => x"54",
          1638 => x"2e",
          1639 => x"70",
          1640 => x"33",
          1641 => x"05",
          1642 => x"11",
          1643 => x"38",
          1644 => x"04",
          1645 => x"75",
          1646 => x"52",
          1647 => x"70",
          1648 => x"34",
          1649 => x"70",
          1650 => x"3d",
          1651 => x"3d",
          1652 => x"79",
          1653 => x"74",
          1654 => x"56",
          1655 => x"81",
          1656 => x"71",
          1657 => x"16",
          1658 => x"52",
          1659 => x"86",
          1660 => x"2e",
          1661 => x"81",
          1662 => x"86",
          1663 => x"fe",
          1664 => x"76",
          1665 => x"54",
          1666 => x"2e",
          1667 => x"73",
          1668 => x"81",
          1669 => x"52",
          1670 => x"2e",
          1671 => x"73",
          1672 => x"06",
          1673 => x"33",
          1674 => x"0c",
          1675 => x"04",
          1676 => x"d3",
          1677 => x"80",
          1678 => x"ac",
          1679 => x"3d",
          1680 => x"80",
          1681 => x"33",
          1682 => x"78",
          1683 => x"38",
          1684 => x"16",
          1685 => x"16",
          1686 => x"17",
          1687 => x"fa",
          1688 => x"d3",
          1689 => x"2e",
          1690 => x"b8",
          1691 => x"ac",
          1692 => x"34",
          1693 => x"a4",
          1694 => x"55",
          1695 => x"08",
          1696 => x"82",
          1697 => x"74",
          1698 => x"81",
          1699 => x"81",
          1700 => x"08",
          1701 => x"05",
          1702 => x"81",
          1703 => x"fa",
          1704 => x"39",
          1705 => x"81",
          1706 => x"89",
          1707 => x"fa",
          1708 => x"7a",
          1709 => x"56",
          1710 => x"75",
          1711 => x"76",
          1712 => x"3f",
          1713 => x"08",
          1714 => x"ac",
          1715 => x"81",
          1716 => x"b4",
          1717 => x"17",
          1718 => x"8a",
          1719 => x"ac",
          1720 => x"85",
          1721 => x"81",
          1722 => x"18",
          1723 => x"d3",
          1724 => x"3d",
          1725 => x"3d",
          1726 => x"52",
          1727 => x"3f",
          1728 => x"08",
          1729 => x"ac",
          1730 => x"38",
          1731 => x"74",
          1732 => x"81",
          1733 => x"38",
          1734 => x"59",
          1735 => x"09",
          1736 => x"e3",
          1737 => x"53",
          1738 => x"08",
          1739 => x"70",
          1740 => x"80",
          1741 => x"d5",
          1742 => x"17",
          1743 => x"3f",
          1744 => x"a4",
          1745 => x"51",
          1746 => x"86",
          1747 => x"f2",
          1748 => x"17",
          1749 => x"3f",
          1750 => x"52",
          1751 => x"51",
          1752 => x"8c",
          1753 => x"84",
          1754 => x"fb",
          1755 => x"17",
          1756 => x"70",
          1757 => x"79",
          1758 => x"52",
          1759 => x"51",
          1760 => x"77",
          1761 => x"80",
          1762 => x"81",
          1763 => x"fa",
          1764 => x"d3",
          1765 => x"2e",
          1766 => x"58",
          1767 => x"ac",
          1768 => x"0d",
          1769 => x"0d",
          1770 => x"98",
          1771 => x"05",
          1772 => x"80",
          1773 => x"27",
          1774 => x"14",
          1775 => x"29",
          1776 => x"05",
          1777 => x"81",
          1778 => x"87",
          1779 => x"f9",
          1780 => x"7a",
          1781 => x"54",
          1782 => x"27",
          1783 => x"14",
          1784 => x"86",
          1785 => x"81",
          1786 => x"74",
          1787 => x"72",
          1788 => x"f5",
          1789 => x"24",
          1790 => x"81",
          1791 => x"81",
          1792 => x"83",
          1793 => x"38",
          1794 => x"74",
          1795 => x"70",
          1796 => x"16",
          1797 => x"74",
          1798 => x"93",
          1799 => x"ac",
          1800 => x"38",
          1801 => x"06",
          1802 => x"33",
          1803 => x"89",
          1804 => x"08",
          1805 => x"54",
          1806 => x"fc",
          1807 => x"d3",
          1808 => x"fe",
          1809 => x"ff",
          1810 => x"11",
          1811 => x"2b",
          1812 => x"81",
          1813 => x"2a",
          1814 => x"51",
          1815 => x"e2",
          1816 => x"ff",
          1817 => x"da",
          1818 => x"2a",
          1819 => x"05",
          1820 => x"fc",
          1821 => x"d3",
          1822 => x"c6",
          1823 => x"83",
          1824 => x"05",
          1825 => x"f8",
          1826 => x"d3",
          1827 => x"ff",
          1828 => x"ae",
          1829 => x"2a",
          1830 => x"05",
          1831 => x"fc",
          1832 => x"d3",
          1833 => x"38",
          1834 => x"83",
          1835 => x"05",
          1836 => x"f8",
          1837 => x"d3",
          1838 => x"0a",
          1839 => x"39",
          1840 => x"81",
          1841 => x"89",
          1842 => x"f7",
          1843 => x"7d",
          1844 => x"55",
          1845 => x"74",
          1846 => x"38",
          1847 => x"08",
          1848 => x"38",
          1849 => x"72",
          1850 => x"a8",
          1851 => x"24",
          1852 => x"81",
          1853 => x"82",
          1854 => x"83",
          1855 => x"38",
          1856 => x"73",
          1857 => x"70",
          1858 => x"17",
          1859 => x"75",
          1860 => x"9b",
          1861 => x"ac",
          1862 => x"d3",
          1863 => x"ea",
          1864 => x"ff",
          1865 => x"11",
          1866 => x"81",
          1867 => x"51",
          1868 => x"72",
          1869 => x"38",
          1870 => x"9f",
          1871 => x"33",
          1872 => x"07",
          1873 => x"78",
          1874 => x"83",
          1875 => x"89",
          1876 => x"08",
          1877 => x"51",
          1878 => x"81",
          1879 => x"57",
          1880 => x"08",
          1881 => x"78",
          1882 => x"15",
          1883 => x"81",
          1884 => x"2a",
          1885 => x"58",
          1886 => x"75",
          1887 => x"33",
          1888 => x"76",
          1889 => x"07",
          1890 => x"34",
          1891 => x"16",
          1892 => x"39",
          1893 => x"a4",
          1894 => x"52",
          1895 => x"8f",
          1896 => x"ac",
          1897 => x"d3",
          1898 => x"de",
          1899 => x"ff",
          1900 => x"73",
          1901 => x"06",
          1902 => x"05",
          1903 => x"3f",
          1904 => x"16",
          1905 => x"39",
          1906 => x"a4",
          1907 => x"52",
          1908 => x"db",
          1909 => x"ac",
          1910 => x"d3",
          1911 => x"38",
          1912 => x"06",
          1913 => x"83",
          1914 => x"11",
          1915 => x"54",
          1916 => x"f6",
          1917 => x"d3",
          1918 => x"0a",
          1919 => x"52",
          1920 => x"dd",
          1921 => x"83",
          1922 => x"81",
          1923 => x"8b",
          1924 => x"f9",
          1925 => x"7b",
          1926 => x"58",
          1927 => x"81",
          1928 => x"38",
          1929 => x"74",
          1930 => x"82",
          1931 => x"39",
          1932 => x"aa",
          1933 => x"75",
          1934 => x"fd",
          1935 => x"d3",
          1936 => x"81",
          1937 => x"80",
          1938 => x"39",
          1939 => x"ed",
          1940 => x"80",
          1941 => x"d3",
          1942 => x"80",
          1943 => x"52",
          1944 => x"eb",
          1945 => x"ac",
          1946 => x"d3",
          1947 => x"2e",
          1948 => x"81",
          1949 => x"81",
          1950 => x"81",
          1951 => x"ff",
          1952 => x"80",
          1953 => x"74",
          1954 => x"3f",
          1955 => x"08",
          1956 => x"15",
          1957 => x"54",
          1958 => x"74",
          1959 => x"90",
          1960 => x"05",
          1961 => x"84",
          1962 => x"07",
          1963 => x"16",
          1964 => x"98",
          1965 => x"26",
          1966 => x"80",
          1967 => x"d3",
          1968 => x"3d",
          1969 => x"3d",
          1970 => x"71",
          1971 => x"5c",
          1972 => x"8c",
          1973 => x"77",
          1974 => x"38",
          1975 => x"78",
          1976 => x"81",
          1977 => x"7a",
          1978 => x"f9",
          1979 => x"55",
          1980 => x"ac",
          1981 => x"e9",
          1982 => x"ac",
          1983 => x"d3",
          1984 => x"2e",
          1985 => x"81",
          1986 => x"55",
          1987 => x"81",
          1988 => x"26",
          1989 => x"7a",
          1990 => x"90",
          1991 => x"2e",
          1992 => x"80",
          1993 => x"2e",
          1994 => x"80",
          1995 => x"1b",
          1996 => x"08",
          1997 => x"38",
          1998 => x"52",
          1999 => x"8f",
          2000 => x"ac",
          2001 => x"5a",
          2002 => x"08",
          2003 => x"81",
          2004 => x"81",
          2005 => x"5a",
          2006 => x"70",
          2007 => x"07",
          2008 => x"7d",
          2009 => x"51",
          2010 => x"73",
          2011 => x"75",
          2012 => x"38",
          2013 => x"56",
          2014 => x"8a",
          2015 => x"1a",
          2016 => x"38",
          2017 => x"57",
          2018 => x"38",
          2019 => x"17",
          2020 => x"08",
          2021 => x"38",
          2022 => x"78",
          2023 => x"38",
          2024 => x"51",
          2025 => x"81",
          2026 => x"56",
          2027 => x"08",
          2028 => x"38",
          2029 => x"d3",
          2030 => x"2e",
          2031 => x"86",
          2032 => x"ac",
          2033 => x"ff",
          2034 => x"70",
          2035 => x"25",
          2036 => x"51",
          2037 => x"73",
          2038 => x"76",
          2039 => x"81",
          2040 => x"38",
          2041 => x"f9",
          2042 => x"76",
          2043 => x"f9",
          2044 => x"d3",
          2045 => x"d3",
          2046 => x"70",
          2047 => x"08",
          2048 => x"7d",
          2049 => x"07",
          2050 => x"06",
          2051 => x"56",
          2052 => x"2e",
          2053 => x"53",
          2054 => x"51",
          2055 => x"81",
          2056 => x"56",
          2057 => x"76",
          2058 => x"98",
          2059 => x"05",
          2060 => x"08",
          2061 => x"38",
          2062 => x"ff",
          2063 => x"0c",
          2064 => x"81",
          2065 => x"84",
          2066 => x"39",
          2067 => x"81",
          2068 => x"89",
          2069 => x"89",
          2070 => x"85",
          2071 => x"76",
          2072 => x"d3",
          2073 => x"3d",
          2074 => x"3d",
          2075 => x"52",
          2076 => x"3f",
          2077 => x"d3",
          2078 => x"db",
          2079 => x"76",
          2080 => x"3f",
          2081 => x"08",
          2082 => x"08",
          2083 => x"5a",
          2084 => x"80",
          2085 => x"70",
          2086 => x"98",
          2087 => x"81",
          2088 => x"84",
          2089 => x"56",
          2090 => x"55",
          2091 => x"97",
          2092 => x"75",
          2093 => x"52",
          2094 => x"51",
          2095 => x"81",
          2096 => x"80",
          2097 => x"80",
          2098 => x"22",
          2099 => x"76",
          2100 => x"81",
          2101 => x"74",
          2102 => x"0c",
          2103 => x"04",
          2104 => x"7a",
          2105 => x"58",
          2106 => x"f0",
          2107 => x"8a",
          2108 => x"06",
          2109 => x"2e",
          2110 => x"58",
          2111 => x"74",
          2112 => x"88",
          2113 => x"73",
          2114 => x"33",
          2115 => x"27",
          2116 => x"16",
          2117 => x"9b",
          2118 => x"2a",
          2119 => x"88",
          2120 => x"58",
          2121 => x"81",
          2122 => x"16",
          2123 => x"0c",
          2124 => x"8a",
          2125 => x"89",
          2126 => x"72",
          2127 => x"38",
          2128 => x"51",
          2129 => x"81",
          2130 => x"54",
          2131 => x"08",
          2132 => x"38",
          2133 => x"d3",
          2134 => x"8b",
          2135 => x"08",
          2136 => x"08",
          2137 => x"82",
          2138 => x"39",
          2139 => x"55",
          2140 => x"cc",
          2141 => x"75",
          2142 => x"3f",
          2143 => x"08",
          2144 => x"73",
          2145 => x"82",
          2146 => x"08",
          2147 => x"38",
          2148 => x"58",
          2149 => x"89",
          2150 => x"08",
          2151 => x"0c",
          2152 => x"06",
          2153 => x"9c",
          2154 => x"58",
          2155 => x"ac",
          2156 => x"0d",
          2157 => x"0d",
          2158 => x"08",
          2159 => x"a0",
          2160 => x"59",
          2161 => x"0a",
          2162 => x"38",
          2163 => x"16",
          2164 => x"98",
          2165 => x"2e",
          2166 => x"75",
          2167 => x"54",
          2168 => x"38",
          2169 => x"81",
          2170 => x"0c",
          2171 => x"98",
          2172 => x"2a",
          2173 => x"59",
          2174 => x"26",
          2175 => x"73",
          2176 => x"84",
          2177 => x"39",
          2178 => x"ff",
          2179 => x"2a",
          2180 => x"72",
          2181 => x"94",
          2182 => x"74",
          2183 => x"3f",
          2184 => x"08",
          2185 => x"81",
          2186 => x"ac",
          2187 => x"84",
          2188 => x"81",
          2189 => x"ff",
          2190 => x"38",
          2191 => x"81",
          2192 => x"26",
          2193 => x"77",
          2194 => x"98",
          2195 => x"53",
          2196 => x"94",
          2197 => x"74",
          2198 => x"3f",
          2199 => x"08",
          2200 => x"81",
          2201 => x"80",
          2202 => x"38",
          2203 => x"d3",
          2204 => x"2e",
          2205 => x"53",
          2206 => x"08",
          2207 => x"38",
          2208 => x"08",
          2209 => x"fb",
          2210 => x"53",
          2211 => x"08",
          2212 => x"94",
          2213 => x"52",
          2214 => x"89",
          2215 => x"ac",
          2216 => x"0c",
          2217 => x"0c",
          2218 => x"06",
          2219 => x"9c",
          2220 => x"53",
          2221 => x"ac",
          2222 => x"0d",
          2223 => x"0d",
          2224 => x"08",
          2225 => x"80",
          2226 => x"fc",
          2227 => x"d3",
          2228 => x"81",
          2229 => x"80",
          2230 => x"d3",
          2231 => x"98",
          2232 => x"77",
          2233 => x"3f",
          2234 => x"08",
          2235 => x"ac",
          2236 => x"38",
          2237 => x"08",
          2238 => x"70",
          2239 => x"55",
          2240 => x"2e",
          2241 => x"83",
          2242 => x"72",
          2243 => x"25",
          2244 => x"53",
          2245 => x"8b",
          2246 => x"57",
          2247 => x"9a",
          2248 => x"80",
          2249 => x"75",
          2250 => x"3f",
          2251 => x"08",
          2252 => x"ac",
          2253 => x"ff",
          2254 => x"84",
          2255 => x"06",
          2256 => x"54",
          2257 => x"ac",
          2258 => x"0d",
          2259 => x"0d",
          2260 => x"52",
          2261 => x"3f",
          2262 => x"08",
          2263 => x"06",
          2264 => x"51",
          2265 => x"83",
          2266 => x"06",
          2267 => x"14",
          2268 => x"3f",
          2269 => x"08",
          2270 => x"07",
          2271 => x"d3",
          2272 => x"3d",
          2273 => x"3d",
          2274 => x"70",
          2275 => x"06",
          2276 => x"53",
          2277 => x"ab",
          2278 => x"33",
          2279 => x"83",
          2280 => x"06",
          2281 => x"90",
          2282 => x"15",
          2283 => x"3f",
          2284 => x"04",
          2285 => x"7b",
          2286 => x"84",
          2287 => x"58",
          2288 => x"80",
          2289 => x"38",
          2290 => x"52",
          2291 => x"df",
          2292 => x"ac",
          2293 => x"d3",
          2294 => x"f1",
          2295 => x"08",
          2296 => x"53",
          2297 => x"84",
          2298 => x"39",
          2299 => x"8b",
          2300 => x"bf",
          2301 => x"ff",
          2302 => x"51",
          2303 => x"17",
          2304 => x"e5",
          2305 => x"76",
          2306 => x"30",
          2307 => x"9f",
          2308 => x"55",
          2309 => x"80",
          2310 => x"76",
          2311 => x"38",
          2312 => x"06",
          2313 => x"88",
          2314 => x"06",
          2315 => x"54",
          2316 => x"99",
          2317 => x"75",
          2318 => x"3f",
          2319 => x"08",
          2320 => x"ac",
          2321 => x"98",
          2322 => x"fc",
          2323 => x"2e",
          2324 => x"0b",
          2325 => x"77",
          2326 => x"0c",
          2327 => x"04",
          2328 => x"7a",
          2329 => x"56",
          2330 => x"51",
          2331 => x"81",
          2332 => x"54",
          2333 => x"08",
          2334 => x"86",
          2335 => x"80",
          2336 => x"16",
          2337 => x"51",
          2338 => x"81",
          2339 => x"57",
          2340 => x"08",
          2341 => x"9c",
          2342 => x"33",
          2343 => x"80",
          2344 => x"9c",
          2345 => x"11",
          2346 => x"55",
          2347 => x"17",
          2348 => x"33",
          2349 => x"70",
          2350 => x"55",
          2351 => x"38",
          2352 => x"16",
          2353 => x"ea",
          2354 => x"d3",
          2355 => x"2e",
          2356 => x"52",
          2357 => x"dd",
          2358 => x"ac",
          2359 => x"d3",
          2360 => x"2e",
          2361 => x"76",
          2362 => x"d3",
          2363 => x"3d",
          2364 => x"3d",
          2365 => x"08",
          2366 => x"52",
          2367 => x"bd",
          2368 => x"ac",
          2369 => x"d3",
          2370 => x"38",
          2371 => x"52",
          2372 => x"9b",
          2373 => x"ac",
          2374 => x"d3",
          2375 => x"38",
          2376 => x"d3",
          2377 => x"9c",
          2378 => x"e9",
          2379 => x"53",
          2380 => x"9c",
          2381 => x"e8",
          2382 => x"0b",
          2383 => x"74",
          2384 => x"0c",
          2385 => x"04",
          2386 => x"76",
          2387 => x"12",
          2388 => x"53",
          2389 => x"d7",
          2390 => x"ac",
          2391 => x"d3",
          2392 => x"38",
          2393 => x"53",
          2394 => x"81",
          2395 => x"34",
          2396 => x"ac",
          2397 => x"0d",
          2398 => x"0d",
          2399 => x"57",
          2400 => x"17",
          2401 => x"08",
          2402 => x"89",
          2403 => x"55",
          2404 => x"08",
          2405 => x"81",
          2406 => x"52",
          2407 => x"ad",
          2408 => x"2e",
          2409 => x"84",
          2410 => x"53",
          2411 => x"09",
          2412 => x"38",
          2413 => x"05",
          2414 => x"81",
          2415 => x"15",
          2416 => x"88",
          2417 => x"81",
          2418 => x"15",
          2419 => x"27",
          2420 => x"15",
          2421 => x"80",
          2422 => x"34",
          2423 => x"52",
          2424 => x"88",
          2425 => x"17",
          2426 => x"51",
          2427 => x"81",
          2428 => x"76",
          2429 => x"08",
          2430 => x"e6",
          2431 => x"d3",
          2432 => x"17",
          2433 => x"08",
          2434 => x"e5",
          2435 => x"d3",
          2436 => x"17",
          2437 => x"0d",
          2438 => x"0d",
          2439 => x"7f",
          2440 => x"5a",
          2441 => x"a0",
          2442 => x"e7",
          2443 => x"70",
          2444 => x"79",
          2445 => x"73",
          2446 => x"81",
          2447 => x"38",
          2448 => x"33",
          2449 => x"ae",
          2450 => x"70",
          2451 => x"82",
          2452 => x"51",
          2453 => x"54",
          2454 => x"7a",
          2455 => x"74",
          2456 => x"58",
          2457 => x"af",
          2458 => x"77",
          2459 => x"70",
          2460 => x"06",
          2461 => x"51",
          2462 => x"74",
          2463 => x"38",
          2464 => x"a0",
          2465 => x"38",
          2466 => x"0c",
          2467 => x"76",
          2468 => x"a0",
          2469 => x"1c",
          2470 => x"82",
          2471 => x"17",
          2472 => x"19",
          2473 => x"a0",
          2474 => x"8c",
          2475 => x"32",
          2476 => x"80",
          2477 => x"30",
          2478 => x"71",
          2479 => x"53",
          2480 => x"55",
          2481 => x"b5",
          2482 => x"81",
          2483 => x"77",
          2484 => x"51",
          2485 => x"af",
          2486 => x"06",
          2487 => x"5a",
          2488 => x"70",
          2489 => x"55",
          2490 => x"2e",
          2491 => x"83",
          2492 => x"79",
          2493 => x"73",
          2494 => x"bc",
          2495 => x"32",
          2496 => x"80",
          2497 => x"27",
          2498 => x"54",
          2499 => x"a2",
          2500 => x"32",
          2501 => x"ae",
          2502 => x"72",
          2503 => x"9f",
          2504 => x"51",
          2505 => x"74",
          2506 => x"88",
          2507 => x"fe",
          2508 => x"98",
          2509 => x"80",
          2510 => x"75",
          2511 => x"81",
          2512 => x"33",
          2513 => x"51",
          2514 => x"81",
          2515 => x"80",
          2516 => x"78",
          2517 => x"81",
          2518 => x"59",
          2519 => x"d7",
          2520 => x"ac",
          2521 => x"89",
          2522 => x"54",
          2523 => x"86",
          2524 => x"80",
          2525 => x"18",
          2526 => x"34",
          2527 => x"11",
          2528 => x"74",
          2529 => x"58",
          2530 => x"75",
          2531 => x"d4",
          2532 => x"3f",
          2533 => x"08",
          2534 => x"ff",
          2535 => x"73",
          2536 => x"38",
          2537 => x"81",
          2538 => x"54",
          2539 => x"75",
          2540 => x"18",
          2541 => x"39",
          2542 => x"0c",
          2543 => x"80",
          2544 => x"7a",
          2545 => x"81",
          2546 => x"81",
          2547 => x"85",
          2548 => x"54",
          2549 => x"8d",
          2550 => x"86",
          2551 => x"86",
          2552 => x"80",
          2553 => x"1c",
          2554 => x"73",
          2555 => x"0c",
          2556 => x"04",
          2557 => x"78",
          2558 => x"56",
          2559 => x"33",
          2560 => x"72",
          2561 => x"38",
          2562 => x"7a",
          2563 => x"54",
          2564 => x"dc",
          2565 => x"81",
          2566 => x"06",
          2567 => x"2e",
          2568 => x"17",
          2569 => x"0c",
          2570 => x"1a",
          2571 => x"70",
          2572 => x"55",
          2573 => x"09",
          2574 => x"38",
          2575 => x"7a",
          2576 => x"54",
          2577 => x"dc",
          2578 => x"06",
          2579 => x"54",
          2580 => x"53",
          2581 => x"80",
          2582 => x"0c",
          2583 => x"51",
          2584 => x"26",
          2585 => x"80",
          2586 => x"34",
          2587 => x"51",
          2588 => x"81",
          2589 => x"55",
          2590 => x"85",
          2591 => x"39",
          2592 => x"05",
          2593 => x"fb",
          2594 => x"d3",
          2595 => x"81",
          2596 => x"81",
          2597 => x"51",
          2598 => x"81",
          2599 => x"ab",
          2600 => x"55",
          2601 => x"08",
          2602 => x"c2",
          2603 => x"ac",
          2604 => x"09",
          2605 => x"ec",
          2606 => x"2a",
          2607 => x"51",
          2608 => x"2e",
          2609 => x"82",
          2610 => x"06",
          2611 => x"80",
          2612 => x"38",
          2613 => x"ab",
          2614 => x"55",
          2615 => x"73",
          2616 => x"81",
          2617 => x"72",
          2618 => x"55",
          2619 => x"82",
          2620 => x"06",
          2621 => x"ac",
          2622 => x"33",
          2623 => x"70",
          2624 => x"54",
          2625 => x"2e",
          2626 => x"90",
          2627 => x"ff",
          2628 => x"05",
          2629 => x"f4",
          2630 => x"d3",
          2631 => x"17",
          2632 => x"39",
          2633 => x"ac",
          2634 => x"0d",
          2635 => x"0d",
          2636 => x"79",
          2637 => x"54",
          2638 => x"74",
          2639 => x"d0",
          2640 => x"81",
          2641 => x"70",
          2642 => x"30",
          2643 => x"71",
          2644 => x"51",
          2645 => x"70",
          2646 => x"ba",
          2647 => x"06",
          2648 => x"74",
          2649 => x"52",
          2650 => x"26",
          2651 => x"15",
          2652 => x"06",
          2653 => x"59",
          2654 => x"2e",
          2655 => x"80",
          2656 => x"cc",
          2657 => x"10",
          2658 => x"08",
          2659 => x"57",
          2660 => x"81",
          2661 => x"75",
          2662 => x"57",
          2663 => x"12",
          2664 => x"70",
          2665 => x"38",
          2666 => x"81",
          2667 => x"51",
          2668 => x"51",
          2669 => x"89",
          2670 => x"70",
          2671 => x"54",
          2672 => x"74",
          2673 => x"30",
          2674 => x"80",
          2675 => x"2a",
          2676 => x"53",
          2677 => x"b9",
          2678 => x"75",
          2679 => x"30",
          2680 => x"9f",
          2681 => x"2a",
          2682 => x"53",
          2683 => x"2e",
          2684 => x"18",
          2685 => x"25",
          2686 => x"8b",
          2687 => x"24",
          2688 => x"77",
          2689 => x"79",
          2690 => x"81",
          2691 => x"51",
          2692 => x"ac",
          2693 => x"0d",
          2694 => x"0d",
          2695 => x"0b",
          2696 => x"ff",
          2697 => x"0c",
          2698 => x"51",
          2699 => x"84",
          2700 => x"ac",
          2701 => x"38",
          2702 => x"51",
          2703 => x"81",
          2704 => x"83",
          2705 => x"54",
          2706 => x"82",
          2707 => x"09",
          2708 => x"e7",
          2709 => x"b4",
          2710 => x"55",
          2711 => x"2e",
          2712 => x"83",
          2713 => x"73",
          2714 => x"70",
          2715 => x"25",
          2716 => x"51",
          2717 => x"38",
          2718 => x"54",
          2719 => x"2e",
          2720 => x"b5",
          2721 => x"81",
          2722 => x"80",
          2723 => x"de",
          2724 => x"d3",
          2725 => x"81",
          2726 => x"80",
          2727 => x"85",
          2728 => x"e8",
          2729 => x"16",
          2730 => x"3f",
          2731 => x"08",
          2732 => x"ac",
          2733 => x"83",
          2734 => x"74",
          2735 => x"0c",
          2736 => x"04",
          2737 => x"60",
          2738 => x"80",
          2739 => x"58",
          2740 => x"0c",
          2741 => x"d5",
          2742 => x"ac",
          2743 => x"56",
          2744 => x"d3",
          2745 => x"87",
          2746 => x"d3",
          2747 => x"10",
          2748 => x"05",
          2749 => x"53",
          2750 => x"80",
          2751 => x"38",
          2752 => x"76",
          2753 => x"75",
          2754 => x"72",
          2755 => x"38",
          2756 => x"51",
          2757 => x"81",
          2758 => x"81",
          2759 => x"81",
          2760 => x"72",
          2761 => x"80",
          2762 => x"73",
          2763 => x"81",
          2764 => x"8a",
          2765 => x"cf",
          2766 => x"86",
          2767 => x"75",
          2768 => x"16",
          2769 => x"81",
          2770 => x"d6",
          2771 => x"d3",
          2772 => x"ff",
          2773 => x"06",
          2774 => x"56",
          2775 => x"38",
          2776 => x"8f",
          2777 => x"2a",
          2778 => x"51",
          2779 => x"72",
          2780 => x"80",
          2781 => x"52",
          2782 => x"3f",
          2783 => x"08",
          2784 => x"57",
          2785 => x"09",
          2786 => x"e4",
          2787 => x"73",
          2788 => x"90",
          2789 => x"10",
          2790 => x"83",
          2791 => x"55",
          2792 => x"57",
          2793 => x"8d",
          2794 => x"16",
          2795 => x"3f",
          2796 => x"08",
          2797 => x"0c",
          2798 => x"83",
          2799 => x"38",
          2800 => x"3d",
          2801 => x"05",
          2802 => x"5b",
          2803 => x"79",
          2804 => x"38",
          2805 => x"51",
          2806 => x"81",
          2807 => x"81",
          2808 => x"81",
          2809 => x"38",
          2810 => x"83",
          2811 => x"38",
          2812 => x"84",
          2813 => x"38",
          2814 => x"81",
          2815 => x"38",
          2816 => x"d9",
          2817 => x"d3",
          2818 => x"ff",
          2819 => x"8d",
          2820 => x"80",
          2821 => x"06",
          2822 => x"80",
          2823 => x"d9",
          2824 => x"d3",
          2825 => x"ff",
          2826 => x"73",
          2827 => x"d8",
          2828 => x"e6",
          2829 => x"ac",
          2830 => x"9c",
          2831 => x"c4",
          2832 => x"16",
          2833 => x"15",
          2834 => x"53",
          2835 => x"81",
          2836 => x"38",
          2837 => x"74",
          2838 => x"c1",
          2839 => x"55",
          2840 => x"16",
          2841 => x"ff",
          2842 => x"72",
          2843 => x"38",
          2844 => x"06",
          2845 => x"2e",
          2846 => x"56",
          2847 => x"80",
          2848 => x"d8",
          2849 => x"d3",
          2850 => x"16",
          2851 => x"ac",
          2852 => x"ff",
          2853 => x"53",
          2854 => x"83",
          2855 => x"c7",
          2856 => x"dd",
          2857 => x"ac",
          2858 => x"ff",
          2859 => x"8d",
          2860 => x"15",
          2861 => x"3f",
          2862 => x"08",
          2863 => x"15",
          2864 => x"3f",
          2865 => x"08",
          2866 => x"06",
          2867 => x"78",
          2868 => x"b3",
          2869 => x"22",
          2870 => x"84",
          2871 => x"56",
          2872 => x"73",
          2873 => x"38",
          2874 => x"52",
          2875 => x"51",
          2876 => x"3f",
          2877 => x"08",
          2878 => x"81",
          2879 => x"80",
          2880 => x"38",
          2881 => x"d3",
          2882 => x"ff",
          2883 => x"26",
          2884 => x"57",
          2885 => x"f5",
          2886 => x"82",
          2887 => x"f5",
          2888 => x"81",
          2889 => x"76",
          2890 => x"db",
          2891 => x"98",
          2892 => x"a0",
          2893 => x"19",
          2894 => x"77",
          2895 => x"0c",
          2896 => x"09",
          2897 => x"38",
          2898 => x"51",
          2899 => x"81",
          2900 => x"83",
          2901 => x"53",
          2902 => x"82",
          2903 => x"15",
          2904 => x"56",
          2905 => x"38",
          2906 => x"51",
          2907 => x"81",
          2908 => x"a8",
          2909 => x"15",
          2910 => x"53",
          2911 => x"15",
          2912 => x"56",
          2913 => x"81",
          2914 => x"15",
          2915 => x"16",
          2916 => x"2e",
          2917 => x"88",
          2918 => x"08",
          2919 => x"39",
          2920 => x"10",
          2921 => x"05",
          2922 => x"98",
          2923 => x"06",
          2924 => x"83",
          2925 => x"2a",
          2926 => x"72",
          2927 => x"26",
          2928 => x"ff",
          2929 => x"0c",
          2930 => x"16",
          2931 => x"0b",
          2932 => x"76",
          2933 => x"81",
          2934 => x"38",
          2935 => x"51",
          2936 => x"81",
          2937 => x"83",
          2938 => x"53",
          2939 => x"09",
          2940 => x"f9",
          2941 => x"52",
          2942 => x"b3",
          2943 => x"ac",
          2944 => x"38",
          2945 => x"08",
          2946 => x"84",
          2947 => x"d5",
          2948 => x"d3",
          2949 => x"ff",
          2950 => x"72",
          2951 => x"2e",
          2952 => x"80",
          2953 => x"15",
          2954 => x"3f",
          2955 => x"08",
          2956 => x"a4",
          2957 => x"81",
          2958 => x"84",
          2959 => x"d5",
          2960 => x"d3",
          2961 => x"8a",
          2962 => x"2e",
          2963 => x"9d",
          2964 => x"15",
          2965 => x"3f",
          2966 => x"08",
          2967 => x"84",
          2968 => x"d5",
          2969 => x"d3",
          2970 => x"16",
          2971 => x"34",
          2972 => x"22",
          2973 => x"72",
          2974 => x"23",
          2975 => x"23",
          2976 => x"16",
          2977 => x"75",
          2978 => x"0c",
          2979 => x"04",
          2980 => x"77",
          2981 => x"73",
          2982 => x"38",
          2983 => x"2e",
          2984 => x"08",
          2985 => x"53",
          2986 => x"a4",
          2987 => x"22",
          2988 => x"57",
          2989 => x"2e",
          2990 => x"94",
          2991 => x"33",
          2992 => x"3f",
          2993 => x"08",
          2994 => x"71",
          2995 => x"55",
          2996 => x"73",
          2997 => x"06",
          2998 => x"08",
          2999 => x"71",
          3000 => x"81",
          3001 => x"87",
          3002 => x"fa",
          3003 => x"ab",
          3004 => x"58",
          3005 => x"05",
          3006 => x"b1",
          3007 => x"ac",
          3008 => x"54",
          3009 => x"d3",
          3010 => x"80",
          3011 => x"d3",
          3012 => x"10",
          3013 => x"05",
          3014 => x"54",
          3015 => x"84",
          3016 => x"34",
          3017 => x"86",
          3018 => x"80",
          3019 => x"10",
          3020 => x"c8",
          3021 => x"0c",
          3022 => x"75",
          3023 => x"38",
          3024 => x"3d",
          3025 => x"05",
          3026 => x"3f",
          3027 => x"08",
          3028 => x"d3",
          3029 => x"3d",
          3030 => x"3d",
          3031 => x"84",
          3032 => x"05",
          3033 => x"89",
          3034 => x"2e",
          3035 => x"76",
          3036 => x"54",
          3037 => x"05",
          3038 => x"84",
          3039 => x"f6",
          3040 => x"d3",
          3041 => x"81",
          3042 => x"84",
          3043 => x"5c",
          3044 => x"3d",
          3045 => x"f0",
          3046 => x"d3",
          3047 => x"81",
          3048 => x"92",
          3049 => x"d7",
          3050 => x"98",
          3051 => x"74",
          3052 => x"38",
          3053 => x"9c",
          3054 => x"80",
          3055 => x"38",
          3056 => x"9c",
          3057 => x"2e",
          3058 => x"8e",
          3059 => x"d4",
          3060 => x"9e",
          3061 => x"ac",
          3062 => x"88",
          3063 => x"39",
          3064 => x"33",
          3065 => x"74",
          3066 => x"38",
          3067 => x"39",
          3068 => x"70",
          3069 => x"55",
          3070 => x"83",
          3071 => x"75",
          3072 => x"76",
          3073 => x"81",
          3074 => x"74",
          3075 => x"a7",
          3076 => x"7a",
          3077 => x"3f",
          3078 => x"08",
          3079 => x"b2",
          3080 => x"8e",
          3081 => x"b9",
          3082 => x"a0",
          3083 => x"34",
          3084 => x"52",
          3085 => x"ce",
          3086 => x"62",
          3087 => x"d2",
          3088 => x"55",
          3089 => x"16",
          3090 => x"2e",
          3091 => x"7a",
          3092 => x"77",
          3093 => x"99",
          3094 => x"53",
          3095 => x"b3",
          3096 => x"ac",
          3097 => x"d3",
          3098 => x"e6",
          3099 => x"7a",
          3100 => x"3f",
          3101 => x"08",
          3102 => x"8c",
          3103 => x"56",
          3104 => x"82",
          3105 => x"b2",
          3106 => x"84",
          3107 => x"06",
          3108 => x"74",
          3109 => x"38",
          3110 => x"39",
          3111 => x"70",
          3112 => x"55",
          3113 => x"8f",
          3114 => x"05",
          3115 => x"55",
          3116 => x"83",
          3117 => x"75",
          3118 => x"76",
          3119 => x"81",
          3120 => x"74",
          3121 => x"38",
          3122 => x"07",
          3123 => x"11",
          3124 => x"0c",
          3125 => x"0c",
          3126 => x"f6",
          3127 => x"74",
          3128 => x"3f",
          3129 => x"08",
          3130 => x"62",
          3131 => x"d0",
          3132 => x"d3",
          3133 => x"19",
          3134 => x"0c",
          3135 => x"84",
          3136 => x"90",
          3137 => x"91",
          3138 => x"9c",
          3139 => x"94",
          3140 => x"80",
          3141 => x"a8",
          3142 => x"98",
          3143 => x"2a",
          3144 => x"51",
          3145 => x"2e",
          3146 => x"8c",
          3147 => x"2e",
          3148 => x"8c",
          3149 => x"19",
          3150 => x"11",
          3151 => x"2b",
          3152 => x"8c",
          3153 => x"5a",
          3154 => x"a5",
          3155 => x"77",
          3156 => x"3f",
          3157 => x"08",
          3158 => x"ac",
          3159 => x"83",
          3160 => x"76",
          3161 => x"81",
          3162 => x"81",
          3163 => x"31",
          3164 => x"70",
          3165 => x"25",
          3166 => x"26",
          3167 => x"55",
          3168 => x"76",
          3169 => x"75",
          3170 => x"78",
          3171 => x"55",
          3172 => x"b9",
          3173 => x"7a",
          3174 => x"3f",
          3175 => x"08",
          3176 => x"56",
          3177 => x"89",
          3178 => x"ac",
          3179 => x"9c",
          3180 => x"81",
          3181 => x"a8",
          3182 => x"81",
          3183 => x"55",
          3184 => x"81",
          3185 => x"80",
          3186 => x"81",
          3187 => x"2e",
          3188 => x"78",
          3189 => x"74",
          3190 => x"0c",
          3191 => x"04",
          3192 => x"7f",
          3193 => x"5f",
          3194 => x"80",
          3195 => x"3d",
          3196 => x"76",
          3197 => x"3f",
          3198 => x"08",
          3199 => x"ac",
          3200 => x"91",
          3201 => x"74",
          3202 => x"38",
          3203 => x"ae",
          3204 => x"33",
          3205 => x"87",
          3206 => x"2e",
          3207 => x"bd",
          3208 => x"91",
          3209 => x"56",
          3210 => x"81",
          3211 => x"34",
          3212 => x"8a",
          3213 => x"91",
          3214 => x"56",
          3215 => x"81",
          3216 => x"34",
          3217 => x"f6",
          3218 => x"91",
          3219 => x"56",
          3220 => x"81",
          3221 => x"34",
          3222 => x"e2",
          3223 => x"08",
          3224 => x"31",
          3225 => x"27",
          3226 => x"59",
          3227 => x"82",
          3228 => x"17",
          3229 => x"ff",
          3230 => x"74",
          3231 => x"7d",
          3232 => x"ff",
          3233 => x"2a",
          3234 => x"7a",
          3235 => x"87",
          3236 => x"08",
          3237 => x"98",
          3238 => x"76",
          3239 => x"3f",
          3240 => x"08",
          3241 => x"27",
          3242 => x"74",
          3243 => x"fb",
          3244 => x"18",
          3245 => x"08",
          3246 => x"d1",
          3247 => x"d3",
          3248 => x"2e",
          3249 => x"81",
          3250 => x"1b",
          3251 => x"5b",
          3252 => x"2e",
          3253 => x"79",
          3254 => x"11",
          3255 => x"56",
          3256 => x"85",
          3257 => x"31",
          3258 => x"77",
          3259 => x"7d",
          3260 => x"52",
          3261 => x"3f",
          3262 => x"08",
          3263 => x"90",
          3264 => x"98",
          3265 => x"74",
          3266 => x"38",
          3267 => x"78",
          3268 => x"7a",
          3269 => x"84",
          3270 => x"17",
          3271 => x"80",
          3272 => x"cc",
          3273 => x"89",
          3274 => x"f9",
          3275 => x"08",
          3276 => x"c9",
          3277 => x"33",
          3278 => x"56",
          3279 => x"25",
          3280 => x"54",
          3281 => x"53",
          3282 => x"7d",
          3283 => x"52",
          3284 => x"3f",
          3285 => x"08",
          3286 => x"90",
          3287 => x"ff",
          3288 => x"90",
          3289 => x"54",
          3290 => x"17",
          3291 => x"11",
          3292 => x"c6",
          3293 => x"d3",
          3294 => x"d7",
          3295 => x"18",
          3296 => x"08",
          3297 => x"84",
          3298 => x"57",
          3299 => x"27",
          3300 => x"56",
          3301 => x"17",
          3302 => x"06",
          3303 => x"52",
          3304 => x"ec",
          3305 => x"31",
          3306 => x"7e",
          3307 => x"94",
          3308 => x"94",
          3309 => x"59",
          3310 => x"38",
          3311 => x"81",
          3312 => x"8f",
          3313 => x"f3",
          3314 => x"62",
          3315 => x"5f",
          3316 => x"7d",
          3317 => x"fc",
          3318 => x"51",
          3319 => x"81",
          3320 => x"55",
          3321 => x"08",
          3322 => x"17",
          3323 => x"80",
          3324 => x"74",
          3325 => x"39",
          3326 => x"70",
          3327 => x"81",
          3328 => x"56",
          3329 => x"80",
          3330 => x"38",
          3331 => x"0b",
          3332 => x"82",
          3333 => x"39",
          3334 => x"18",
          3335 => x"83",
          3336 => x"0b",
          3337 => x"81",
          3338 => x"39",
          3339 => x"18",
          3340 => x"83",
          3341 => x"0b",
          3342 => x"81",
          3343 => x"39",
          3344 => x"18",
          3345 => x"83",
          3346 => x"17",
          3347 => x"74",
          3348 => x"27",
          3349 => x"17",
          3350 => x"78",
          3351 => x"8c",
          3352 => x"08",
          3353 => x"06",
          3354 => x"82",
          3355 => x"8a",
          3356 => x"05",
          3357 => x"06",
          3358 => x"80",
          3359 => x"96",
          3360 => x"08",
          3361 => x"38",
          3362 => x"51",
          3363 => x"81",
          3364 => x"55",
          3365 => x"17",
          3366 => x"51",
          3367 => x"81",
          3368 => x"55",
          3369 => x"82",
          3370 => x"81",
          3371 => x"38",
          3372 => x"fe",
          3373 => x"98",
          3374 => x"17",
          3375 => x"74",
          3376 => x"90",
          3377 => x"98",
          3378 => x"74",
          3379 => x"38",
          3380 => x"17",
          3381 => x"17",
          3382 => x"11",
          3383 => x"c5",
          3384 => x"d3",
          3385 => x"ba",
          3386 => x"33",
          3387 => x"55",
          3388 => x"34",
          3389 => x"52",
          3390 => x"a9",
          3391 => x"ac",
          3392 => x"fe",
          3393 => x"d3",
          3394 => x"79",
          3395 => x"58",
          3396 => x"80",
          3397 => x"1b",
          3398 => x"22",
          3399 => x"74",
          3400 => x"38",
          3401 => x"5a",
          3402 => x"53",
          3403 => x"81",
          3404 => x"55",
          3405 => x"81",
          3406 => x"fd",
          3407 => x"17",
          3408 => x"55",
          3409 => x"9b",
          3410 => x"53",
          3411 => x"29",
          3412 => x"17",
          3413 => x"3f",
          3414 => x"80",
          3415 => x"74",
          3416 => x"79",
          3417 => x"80",
          3418 => x"17",
          3419 => x"a1",
          3420 => x"08",
          3421 => x"27",
          3422 => x"54",
          3423 => x"17",
          3424 => x"11",
          3425 => x"c2",
          3426 => x"d3",
          3427 => x"b0",
          3428 => x"18",
          3429 => x"08",
          3430 => x"84",
          3431 => x"57",
          3432 => x"27",
          3433 => x"56",
          3434 => x"52",
          3435 => x"83",
          3436 => x"a8",
          3437 => x"d8",
          3438 => x"33",
          3439 => x"55",
          3440 => x"34",
          3441 => x"7d",
          3442 => x"0c",
          3443 => x"19",
          3444 => x"94",
          3445 => x"1a",
          3446 => x"5d",
          3447 => x"27",
          3448 => x"55",
          3449 => x"0c",
          3450 => x"38",
          3451 => x"80",
          3452 => x"74",
          3453 => x"80",
          3454 => x"d3",
          3455 => x"3d",
          3456 => x"3d",
          3457 => x"3d",
          3458 => x"70",
          3459 => x"80",
          3460 => x"ac",
          3461 => x"d3",
          3462 => x"aa",
          3463 => x"33",
          3464 => x"70",
          3465 => x"56",
          3466 => x"2e",
          3467 => x"75",
          3468 => x"74",
          3469 => x"38",
          3470 => x"18",
          3471 => x"18",
          3472 => x"11",
          3473 => x"c2",
          3474 => x"55",
          3475 => x"08",
          3476 => x"90",
          3477 => x"ff",
          3478 => x"90",
          3479 => x"18",
          3480 => x"51",
          3481 => x"81",
          3482 => x"57",
          3483 => x"08",
          3484 => x"a4",
          3485 => x"11",
          3486 => x"56",
          3487 => x"17",
          3488 => x"08",
          3489 => x"77",
          3490 => x"fa",
          3491 => x"08",
          3492 => x"51",
          3493 => x"82",
          3494 => x"52",
          3495 => x"c5",
          3496 => x"52",
          3497 => x"c5",
          3498 => x"55",
          3499 => x"16",
          3500 => x"c8",
          3501 => x"d3",
          3502 => x"19",
          3503 => x"06",
          3504 => x"90",
          3505 => x"55",
          3506 => x"ac",
          3507 => x"0d",
          3508 => x"0d",
          3509 => x"54",
          3510 => x"81",
          3511 => x"53",
          3512 => x"08",
          3513 => x"3d",
          3514 => x"73",
          3515 => x"3f",
          3516 => x"08",
          3517 => x"ac",
          3518 => x"81",
          3519 => x"74",
          3520 => x"d3",
          3521 => x"3d",
          3522 => x"3d",
          3523 => x"51",
          3524 => x"8b",
          3525 => x"81",
          3526 => x"24",
          3527 => x"d3",
          3528 => x"d3",
          3529 => x"53",
          3530 => x"ac",
          3531 => x"0d",
          3532 => x"0d",
          3533 => x"3d",
          3534 => x"94",
          3535 => x"84",
          3536 => x"ac",
          3537 => x"d3",
          3538 => x"df",
          3539 => x"63",
          3540 => x"d4",
          3541 => x"9c",
          3542 => x"ac",
          3543 => x"d3",
          3544 => x"38",
          3545 => x"05",
          3546 => x"2b",
          3547 => x"80",
          3548 => x"76",
          3549 => x"0c",
          3550 => x"02",
          3551 => x"70",
          3552 => x"81",
          3553 => x"56",
          3554 => x"93",
          3555 => x"53",
          3556 => x"d7",
          3557 => x"d3",
          3558 => x"15",
          3559 => x"85",
          3560 => x"2e",
          3561 => x"83",
          3562 => x"74",
          3563 => x"0c",
          3564 => x"04",
          3565 => x"a3",
          3566 => x"3d",
          3567 => x"80",
          3568 => x"53",
          3569 => x"b8",
          3570 => x"3d",
          3571 => x"3f",
          3572 => x"08",
          3573 => x"ac",
          3574 => x"38",
          3575 => x"7f",
          3576 => x"4a",
          3577 => x"59",
          3578 => x"81",
          3579 => x"3d",
          3580 => x"40",
          3581 => x"52",
          3582 => x"e4",
          3583 => x"ac",
          3584 => x"d3",
          3585 => x"de",
          3586 => x"7e",
          3587 => x"3f",
          3588 => x"08",
          3589 => x"ac",
          3590 => x"38",
          3591 => x"51",
          3592 => x"81",
          3593 => x"48",
          3594 => x"51",
          3595 => x"81",
          3596 => x"57",
          3597 => x"08",
          3598 => x"7c",
          3599 => x"73",
          3600 => x"3f",
          3601 => x"08",
          3602 => x"ac",
          3603 => x"6c",
          3604 => x"d5",
          3605 => x"d3",
          3606 => x"2e",
          3607 => x"52",
          3608 => x"d1",
          3609 => x"ac",
          3610 => x"d3",
          3611 => x"2e",
          3612 => x"84",
          3613 => x"06",
          3614 => x"57",
          3615 => x"38",
          3616 => x"bc",
          3617 => x"05",
          3618 => x"3f",
          3619 => x"70",
          3620 => x"11",
          3621 => x"57",
          3622 => x"80",
          3623 => x"81",
          3624 => x"81",
          3625 => x"55",
          3626 => x"38",
          3627 => x"78",
          3628 => x"38",
          3629 => x"39",
          3630 => x"99",
          3631 => x"ff",
          3632 => x"08",
          3633 => x"70",
          3634 => x"56",
          3635 => x"33",
          3636 => x"eb",
          3637 => x"a3",
          3638 => x"55",
          3639 => x"34",
          3640 => x"fe",
          3641 => x"81",
          3642 => x"7c",
          3643 => x"06",
          3644 => x"19",
          3645 => x"11",
          3646 => x"74",
          3647 => x"81",
          3648 => x"70",
          3649 => x"bb",
          3650 => x"08",
          3651 => x"52",
          3652 => x"58",
          3653 => x"8d",
          3654 => x"70",
          3655 => x"51",
          3656 => x"f5",
          3657 => x"54",
          3658 => x"a5",
          3659 => x"77",
          3660 => x"38",
          3661 => x"73",
          3662 => x"81",
          3663 => x"81",
          3664 => x"78",
          3665 => x"ba",
          3666 => x"05",
          3667 => x"18",
          3668 => x"38",
          3669 => x"96",
          3670 => x"08",
          3671 => x"5a",
          3672 => x"7a",
          3673 => x"5c",
          3674 => x"26",
          3675 => x"7a",
          3676 => x"d3",
          3677 => x"3d",
          3678 => x"3d",
          3679 => x"90",
          3680 => x"54",
          3681 => x"57",
          3682 => x"81",
          3683 => x"5a",
          3684 => x"08",
          3685 => x"17",
          3686 => x"80",
          3687 => x"79",
          3688 => x"39",
          3689 => x"78",
          3690 => x"90",
          3691 => x"81",
          3692 => x"06",
          3693 => x"74",
          3694 => x"17",
          3695 => x"17",
          3696 => x"70",
          3697 => x"5b",
          3698 => x"82",
          3699 => x"8a",
          3700 => x"89",
          3701 => x"55",
          3702 => x"b6",
          3703 => x"ff",
          3704 => x"96",
          3705 => x"d3",
          3706 => x"17",
          3707 => x"53",
          3708 => x"96",
          3709 => x"d3",
          3710 => x"26",
          3711 => x"30",
          3712 => x"18",
          3713 => x"18",
          3714 => x"18",
          3715 => x"80",
          3716 => x"17",
          3717 => x"be",
          3718 => x"76",
          3719 => x"3f",
          3720 => x"08",
          3721 => x"ac",
          3722 => x"09",
          3723 => x"38",
          3724 => x"18",
          3725 => x"82",
          3726 => x"d3",
          3727 => x"2e",
          3728 => x"8b",
          3729 => x"91",
          3730 => x"55",
          3731 => x"81",
          3732 => x"88",
          3733 => x"98",
          3734 => x"80",
          3735 => x"38",
          3736 => x"80",
          3737 => x"79",
          3738 => x"08",
          3739 => x"0c",
          3740 => x"70",
          3741 => x"81",
          3742 => x"5d",
          3743 => x"2e",
          3744 => x"52",
          3745 => x"be",
          3746 => x"ac",
          3747 => x"d3",
          3748 => x"38",
          3749 => x"08",
          3750 => x"75",
          3751 => x"c2",
          3752 => x"d3",
          3753 => x"75",
          3754 => x"e1",
          3755 => x"27",
          3756 => x"55",
          3757 => x"76",
          3758 => x"82",
          3759 => x"34",
          3760 => x"d8",
          3761 => x"18",
          3762 => x"26",
          3763 => x"94",
          3764 => x"94",
          3765 => x"83",
          3766 => x"74",
          3767 => x"38",
          3768 => x"51",
          3769 => x"81",
          3770 => x"8b",
          3771 => x"91",
          3772 => x"55",
          3773 => x"77",
          3774 => x"d3",
          3775 => x"5b",
          3776 => x"94",
          3777 => x"92",
          3778 => x"08",
          3779 => x"90",
          3780 => x"c0",
          3781 => x"90",
          3782 => x"17",
          3783 => x"06",
          3784 => x"2e",
          3785 => x"9c",
          3786 => x"2e",
          3787 => x"90",
          3788 => x"98",
          3789 => x"74",
          3790 => x"38",
          3791 => x"17",
          3792 => x"17",
          3793 => x"11",
          3794 => x"ff",
          3795 => x"81",
          3796 => x"80",
          3797 => x"81",
          3798 => x"34",
          3799 => x"39",
          3800 => x"80",
          3801 => x"74",
          3802 => x"81",
          3803 => x"a8",
          3804 => x"81",
          3805 => x"55",
          3806 => x"3f",
          3807 => x"08",
          3808 => x"38",
          3809 => x"18",
          3810 => x"90",
          3811 => x"91",
          3812 => x"55",
          3813 => x"9c",
          3814 => x"55",
          3815 => x"ac",
          3816 => x"0d",
          3817 => x"0d",
          3818 => x"54",
          3819 => x"81",
          3820 => x"53",
          3821 => x"05",
          3822 => x"84",
          3823 => x"84",
          3824 => x"ac",
          3825 => x"d3",
          3826 => x"ef",
          3827 => x"0c",
          3828 => x"51",
          3829 => x"81",
          3830 => x"55",
          3831 => x"08",
          3832 => x"ab",
          3833 => x"98",
          3834 => x"80",
          3835 => x"38",
          3836 => x"70",
          3837 => x"81",
          3838 => x"57",
          3839 => x"93",
          3840 => x"08",
          3841 => x"ce",
          3842 => x"d3",
          3843 => x"17",
          3844 => x"85",
          3845 => x"38",
          3846 => x"14",
          3847 => x"23",
          3848 => x"51",
          3849 => x"81",
          3850 => x"55",
          3851 => x"09",
          3852 => x"38",
          3853 => x"80",
          3854 => x"80",
          3855 => x"54",
          3856 => x"ac",
          3857 => x"0d",
          3858 => x"0d",
          3859 => x"fc",
          3860 => x"52",
          3861 => x"3f",
          3862 => x"08",
          3863 => x"ac",
          3864 => x"81",
          3865 => x"74",
          3866 => x"d3",
          3867 => x"3d",
          3868 => x"3d",
          3869 => x"89",
          3870 => x"54",
          3871 => x"54",
          3872 => x"81",
          3873 => x"53",
          3874 => x"08",
          3875 => x"74",
          3876 => x"d3",
          3877 => x"73",
          3878 => x"3f",
          3879 => x"08",
          3880 => x"80",
          3881 => x"ce",
          3882 => x"d3",
          3883 => x"81",
          3884 => x"84",
          3885 => x"06",
          3886 => x"53",
          3887 => x"74",
          3888 => x"d1",
          3889 => x"52",
          3890 => x"e9",
          3891 => x"ac",
          3892 => x"d3",
          3893 => x"2e",
          3894 => x"83",
          3895 => x"72",
          3896 => x"0c",
          3897 => x"04",
          3898 => x"64",
          3899 => x"88",
          3900 => x"95",
          3901 => x"db",
          3902 => x"d3",
          3903 => x"81",
          3904 => x"b5",
          3905 => x"73",
          3906 => x"3f",
          3907 => x"08",
          3908 => x"ac",
          3909 => x"02",
          3910 => x"33",
          3911 => x"55",
          3912 => x"25",
          3913 => x"55",
          3914 => x"80",
          3915 => x"75",
          3916 => x"d4",
          3917 => x"c1",
          3918 => x"d3",
          3919 => x"3d",
          3920 => x"3d",
          3921 => x"55",
          3922 => x"90",
          3923 => x"52",
          3924 => x"da",
          3925 => x"d3",
          3926 => x"81",
          3927 => x"82",
          3928 => x"74",
          3929 => x"98",
          3930 => x"05",
          3931 => x"15",
          3932 => x"93",
          3933 => x"08",
          3934 => x"e9",
          3935 => x"81",
          3936 => x"59",
          3937 => x"80",
          3938 => x"56",
          3939 => x"81",
          3940 => x"06",
          3941 => x"82",
          3942 => x"75",
          3943 => x"f0",
          3944 => x"bc",
          3945 => x"d3",
          3946 => x"2e",
          3947 => x"d3",
          3948 => x"2e",
          3949 => x"d3",
          3950 => x"70",
          3951 => x"08",
          3952 => x"78",
          3953 => x"7d",
          3954 => x"54",
          3955 => x"76",
          3956 => x"80",
          3957 => x"98",
          3958 => x"12",
          3959 => x"54",
          3960 => x"98",
          3961 => x"81",
          3962 => x"58",
          3963 => x"3f",
          3964 => x"08",
          3965 => x"ac",
          3966 => x"38",
          3967 => x"51",
          3968 => x"2e",
          3969 => x"a0",
          3970 => x"b4",
          3971 => x"b5",
          3972 => x"d3",
          3973 => x"ff",
          3974 => x"30",
          3975 => x"19",
          3976 => x"59",
          3977 => x"39",
          3978 => x"05",
          3979 => x"ea",
          3980 => x"ac",
          3981 => x"06",
          3982 => x"80",
          3983 => x"18",
          3984 => x"54",
          3985 => x"06",
          3986 => x"55",
          3987 => x"38",
          3988 => x"7a",
          3989 => x"0c",
          3990 => x"11",
          3991 => x"55",
          3992 => x"16",
          3993 => x"d3",
          3994 => x"3d",
          3995 => x"3d",
          3996 => x"3d",
          3997 => x"70",
          3998 => x"94",
          3999 => x"ac",
          4000 => x"d3",
          4001 => x"38",
          4002 => x"57",
          4003 => x"86",
          4004 => x"81",
          4005 => x"18",
          4006 => x"2a",
          4007 => x"51",
          4008 => x"56",
          4009 => x"81",
          4010 => x"18",
          4011 => x"08",
          4012 => x"38",
          4013 => x"9a",
          4014 => x"88",
          4015 => x"77",
          4016 => x"cf",
          4017 => x"ac",
          4018 => x"0b",
          4019 => x"80",
          4020 => x"18",
          4021 => x"51",
          4022 => x"3f",
          4023 => x"08",
          4024 => x"08",
          4025 => x"30",
          4026 => x"80",
          4027 => x"58",
          4028 => x"ac",
          4029 => x"09",
          4030 => x"38",
          4031 => x"9b",
          4032 => x"75",
          4033 => x"27",
          4034 => x"18",
          4035 => x"52",
          4036 => x"bd",
          4037 => x"d3",
          4038 => x"94",
          4039 => x"19",
          4040 => x"33",
          4041 => x"55",
          4042 => x"34",
          4043 => x"74",
          4044 => x"74",
          4045 => x"38",
          4046 => x"18",
          4047 => x"18",
          4048 => x"11",
          4049 => x"ff",
          4050 => x"81",
          4051 => x"80",
          4052 => x"81",
          4053 => x"90",
          4054 => x"ff",
          4055 => x"90",
          4056 => x"80",
          4057 => x"76",
          4058 => x"76",
          4059 => x"76",
          4060 => x"d3",
          4061 => x"3d",
          4062 => x"3d",
          4063 => x"f0",
          4064 => x"d5",
          4065 => x"9f",
          4066 => x"05",
          4067 => x"51",
          4068 => x"81",
          4069 => x"56",
          4070 => x"08",
          4071 => x"81",
          4072 => x"ff",
          4073 => x"77",
          4074 => x"9f",
          4075 => x"51",
          4076 => x"81",
          4077 => x"81",
          4078 => x"56",
          4079 => x"3f",
          4080 => x"38",
          4081 => x"05",
          4082 => x"2a",
          4083 => x"51",
          4084 => x"80",
          4085 => x"86",
          4086 => x"95",
          4087 => x"fc",
          4088 => x"f5",
          4089 => x"f7",
          4090 => x"98",
          4091 => x"73",
          4092 => x"38",
          4093 => x"39",
          4094 => x"05",
          4095 => x"54",
          4096 => x"83",
          4097 => x"75",
          4098 => x"6a",
          4099 => x"c6",
          4100 => x"d3",
          4101 => x"84",
          4102 => x"05",
          4103 => x"2a",
          4104 => x"51",
          4105 => x"73",
          4106 => x"e5",
          4107 => x"80",
          4108 => x"a5",
          4109 => x"55",
          4110 => x"08",
          4111 => x"d1",
          4112 => x"84",
          4113 => x"91",
          4114 => x"76",
          4115 => x"88",
          4116 => x"85",
          4117 => x"89",
          4118 => x"54",
          4119 => x"81",
          4120 => x"56",
          4121 => x"08",
          4122 => x"81",
          4123 => x"52",
          4124 => x"c0",
          4125 => x"ac",
          4126 => x"d3",
          4127 => x"38",
          4128 => x"84",
          4129 => x"70",
          4130 => x"2c",
          4131 => x"56",
          4132 => x"dd",
          4133 => x"8c",
          4134 => x"bd",
          4135 => x"d4",
          4136 => x"a4",
          4137 => x"ac",
          4138 => x"ac",
          4139 => x"81",
          4140 => x"07",
          4141 => x"30",
          4142 => x"9f",
          4143 => x"52",
          4144 => x"56",
          4145 => x"9b",
          4146 => x"90",
          4147 => x"89",
          4148 => x"76",
          4149 => x"d4",
          4150 => x"ba",
          4151 => x"d3",
          4152 => x"75",
          4153 => x"51",
          4154 => x"3f",
          4155 => x"08",
          4156 => x"94",
          4157 => x"e1",
          4158 => x"d3",
          4159 => x"3d",
          4160 => x"3d",
          4161 => x"98",
          4162 => x"52",
          4163 => x"d3",
          4164 => x"d3",
          4165 => x"81",
          4166 => x"82",
          4167 => x"5d",
          4168 => x"3d",
          4169 => x"cd",
          4170 => x"d3",
          4171 => x"81",
          4172 => x"83",
          4173 => x"74",
          4174 => x"81",
          4175 => x"38",
          4176 => x"05",
          4177 => x"2a",
          4178 => x"51",
          4179 => x"80",
          4180 => x"86",
          4181 => x"2e",
          4182 => x"81",
          4183 => x"59",
          4184 => x"3d",
          4185 => x"ff",
          4186 => x"81",
          4187 => x"56",
          4188 => x"d3",
          4189 => x"2e",
          4190 => x"83",
          4191 => x"75",
          4192 => x"81",
          4193 => x"82",
          4194 => x"2e",
          4195 => x"83",
          4196 => x"82",
          4197 => x"57",
          4198 => x"38",
          4199 => x"51",
          4200 => x"3f",
          4201 => x"08",
          4202 => x"ac",
          4203 => x"38",
          4204 => x"52",
          4205 => x"ff",
          4206 => x"77",
          4207 => x"b4",
          4208 => x"54",
          4209 => x"15",
          4210 => x"80",
          4211 => x"ff",
          4212 => x"75",
          4213 => x"52",
          4214 => x"aa",
          4215 => x"b4",
          4216 => x"d4",
          4217 => x"af",
          4218 => x"54",
          4219 => x"d5",
          4220 => x"53",
          4221 => x"52",
          4222 => x"8a",
          4223 => x"81",
          4224 => x"34",
          4225 => x"05",
          4226 => x"3f",
          4227 => x"08",
          4228 => x"ac",
          4229 => x"76",
          4230 => x"05",
          4231 => x"c1",
          4232 => x"63",
          4233 => x"c2",
          4234 => x"54",
          4235 => x"15",
          4236 => x"81",
          4237 => x"34",
          4238 => x"b1",
          4239 => x"d3",
          4240 => x"8e",
          4241 => x"75",
          4242 => x"c4",
          4243 => x"b7",
          4244 => x"81",
          4245 => x"98",
          4246 => x"db",
          4247 => x"3d",
          4248 => x"cd",
          4249 => x"53",
          4250 => x"84",
          4251 => x"3d",
          4252 => x"3f",
          4253 => x"08",
          4254 => x"ac",
          4255 => x"38",
          4256 => x"3d",
          4257 => x"3d",
          4258 => x"ca",
          4259 => x"d3",
          4260 => x"81",
          4261 => x"82",
          4262 => x"81",
          4263 => x"81",
          4264 => x"73",
          4265 => x"38",
          4266 => x"82",
          4267 => x"53",
          4268 => x"52",
          4269 => x"88",
          4270 => x"ad",
          4271 => x"53",
          4272 => x"05",
          4273 => x"70",
          4274 => x"ad",
          4275 => x"3d",
          4276 => x"51",
          4277 => x"81",
          4278 => x"55",
          4279 => x"08",
          4280 => x"6e",
          4281 => x"06",
          4282 => x"55",
          4283 => x"08",
          4284 => x"88",
          4285 => x"2e",
          4286 => x"81",
          4287 => x"3d",
          4288 => x"51",
          4289 => x"81",
          4290 => x"55",
          4291 => x"08",
          4292 => x"67",
          4293 => x"a7",
          4294 => x"05",
          4295 => x"51",
          4296 => x"3f",
          4297 => x"33",
          4298 => x"8b",
          4299 => x"84",
          4300 => x"06",
          4301 => x"73",
          4302 => x"a0",
          4303 => x"8b",
          4304 => x"54",
          4305 => x"15",
          4306 => x"33",
          4307 => x"70",
          4308 => x"55",
          4309 => x"2e",
          4310 => x"6d",
          4311 => x"d5",
          4312 => x"77",
          4313 => x"e5",
          4314 => x"ac",
          4315 => x"51",
          4316 => x"3f",
          4317 => x"d3",
          4318 => x"2e",
          4319 => x"d3",
          4320 => x"77",
          4321 => x"a7",
          4322 => x"ac",
          4323 => x"19",
          4324 => x"d3",
          4325 => x"38",
          4326 => x"54",
          4327 => x"09",
          4328 => x"38",
          4329 => x"52",
          4330 => x"bf",
          4331 => x"54",
          4332 => x"15",
          4333 => x"38",
          4334 => x"05",
          4335 => x"3f",
          4336 => x"08",
          4337 => x"ac",
          4338 => x"77",
          4339 => x"a6",
          4340 => x"ac",
          4341 => x"81",
          4342 => x"a7",
          4343 => x"ed",
          4344 => x"80",
          4345 => x"02",
          4346 => x"df",
          4347 => x"57",
          4348 => x"3d",
          4349 => x"96",
          4350 => x"c8",
          4351 => x"ac",
          4352 => x"d3",
          4353 => x"d4",
          4354 => x"65",
          4355 => x"d4",
          4356 => x"e0",
          4357 => x"ac",
          4358 => x"d3",
          4359 => x"38",
          4360 => x"05",
          4361 => x"06",
          4362 => x"2e",
          4363 => x"55",
          4364 => x"75",
          4365 => x"71",
          4366 => x"33",
          4367 => x"74",
          4368 => x"57",
          4369 => x"8b",
          4370 => x"54",
          4371 => x"15",
          4372 => x"ff",
          4373 => x"81",
          4374 => x"55",
          4375 => x"ac",
          4376 => x"0d",
          4377 => x"0d",
          4378 => x"53",
          4379 => x"05",
          4380 => x"51",
          4381 => x"81",
          4382 => x"55",
          4383 => x"08",
          4384 => x"77",
          4385 => x"94",
          4386 => x"51",
          4387 => x"81",
          4388 => x"55",
          4389 => x"08",
          4390 => x"80",
          4391 => x"81",
          4392 => x"73",
          4393 => x"38",
          4394 => x"a9",
          4395 => x"22",
          4396 => x"70",
          4397 => x"07",
          4398 => x"7f",
          4399 => x"ff",
          4400 => x"77",
          4401 => x"83",
          4402 => x"51",
          4403 => x"3f",
          4404 => x"08",
          4405 => x"d3",
          4406 => x"3d",
          4407 => x"3d",
          4408 => x"5c",
          4409 => x"98",
          4410 => x"52",
          4411 => x"cb",
          4412 => x"d3",
          4413 => x"d3",
          4414 => x"70",
          4415 => x"08",
          4416 => x"7b",
          4417 => x"07",
          4418 => x"06",
          4419 => x"56",
          4420 => x"2e",
          4421 => x"7b",
          4422 => x"80",
          4423 => x"70",
          4424 => x"b7",
          4425 => x"d3",
          4426 => x"81",
          4427 => x"80",
          4428 => x"52",
          4429 => x"bc",
          4430 => x"d3",
          4431 => x"81",
          4432 => x"bb",
          4433 => x"ac",
          4434 => x"ac",
          4435 => x"58",
          4436 => x"81",
          4437 => x"56",
          4438 => x"33",
          4439 => x"18",
          4440 => x"27",
          4441 => x"19",
          4442 => x"34",
          4443 => x"8f",
          4444 => x"79",
          4445 => x"51",
          4446 => x"a0",
          4447 => x"75",
          4448 => x"81",
          4449 => x"80",
          4450 => x"56",
          4451 => x"77",
          4452 => x"7c",
          4453 => x"07",
          4454 => x"06",
          4455 => x"55",
          4456 => x"bc",
          4457 => x"11",
          4458 => x"ff",
          4459 => x"81",
          4460 => x"56",
          4461 => x"08",
          4462 => x"70",
          4463 => x"80",
          4464 => x"83",
          4465 => x"80",
          4466 => x"84",
          4467 => x"a7",
          4468 => x"b4",
          4469 => x"a6",
          4470 => x"d3",
          4471 => x"0c",
          4472 => x"ac",
          4473 => x"0d",
          4474 => x"0d",
          4475 => x"3d",
          4476 => x"52",
          4477 => x"c9",
          4478 => x"d3",
          4479 => x"81",
          4480 => x"83",
          4481 => x"53",
          4482 => x"3d",
          4483 => x"51",
          4484 => x"3f",
          4485 => x"71",
          4486 => x"55",
          4487 => x"27",
          4488 => x"74",
          4489 => x"05",
          4490 => x"ff",
          4491 => x"ff",
          4492 => x"81",
          4493 => x"80",
          4494 => x"6a",
          4495 => x"53",
          4496 => x"a7",
          4497 => x"d3",
          4498 => x"2e",
          4499 => x"88",
          4500 => x"6b",
          4501 => x"56",
          4502 => x"56",
          4503 => x"54",
          4504 => x"8a",
          4505 => x"70",
          4506 => x"06",
          4507 => x"ff",
          4508 => x"38",
          4509 => x"16",
          4510 => x"80",
          4511 => x"75",
          4512 => x"dc",
          4513 => x"f7",
          4514 => x"ac",
          4515 => x"81",
          4516 => x"88",
          4517 => x"26",
          4518 => x"39",
          4519 => x"86",
          4520 => x"82",
          4521 => x"ff",
          4522 => x"38",
          4523 => x"05",
          4524 => x"76",
          4525 => x"55",
          4526 => x"81",
          4527 => x"3d",
          4528 => x"bc",
          4529 => x"74",
          4530 => x"6b",
          4531 => x"56",
          4532 => x"26",
          4533 => x"89",
          4534 => x"86",
          4535 => x"e5",
          4536 => x"38",
          4537 => x"a8",
          4538 => x"05",
          4539 => x"70",
          4540 => x"56",
          4541 => x"2e",
          4542 => x"94",
          4543 => x"57",
          4544 => x"8c",
          4545 => x"70",
          4546 => x"73",
          4547 => x"38",
          4548 => x"41",
          4549 => x"3d",
          4550 => x"ff",
          4551 => x"81",
          4552 => x"54",
          4553 => x"08",
          4554 => x"81",
          4555 => x"ff",
          4556 => x"81",
          4557 => x"54",
          4558 => x"08",
          4559 => x"80",
          4560 => x"8b",
          4561 => x"ff",
          4562 => x"65",
          4563 => x"c0",
          4564 => x"65",
          4565 => x"34",
          4566 => x"0b",
          4567 => x"77",
          4568 => x"92",
          4569 => x"ac",
          4570 => x"df",
          4571 => x"ac",
          4572 => x"09",
          4573 => x"d3",
          4574 => x"76",
          4575 => x"cb",
          4576 => x"9a",
          4577 => x"51",
          4578 => x"3f",
          4579 => x"08",
          4580 => x"ac",
          4581 => x"a0",
          4582 => x"ac",
          4583 => x"51",
          4584 => x"3f",
          4585 => x"0b",
          4586 => x"8b",
          4587 => x"ff",
          4588 => x"65",
          4589 => x"d8",
          4590 => x"81",
          4591 => x"34",
          4592 => x"a6",
          4593 => x"d3",
          4594 => x"73",
          4595 => x"d3",
          4596 => x"3d",
          4597 => x"3d",
          4598 => x"02",
          4599 => x"cf",
          4600 => x"3d",
          4601 => x"72",
          4602 => x"58",
          4603 => x"81",
          4604 => x"57",
          4605 => x"08",
          4606 => x"18",
          4607 => x"80",
          4608 => x"76",
          4609 => x"39",
          4610 => x"95",
          4611 => x"08",
          4612 => x"18",
          4613 => x"2a",
          4614 => x"51",
          4615 => x"90",
          4616 => x"82",
          4617 => x"57",
          4618 => x"81",
          4619 => x"39",
          4620 => x"22",
          4621 => x"70",
          4622 => x"58",
          4623 => x"f9",
          4624 => x"16",
          4625 => x"30",
          4626 => x"9f",
          4627 => x"ac",
          4628 => x"8c",
          4629 => x"52",
          4630 => x"80",
          4631 => x"27",
          4632 => x"14",
          4633 => x"83",
          4634 => x"78",
          4635 => x"80",
          4636 => x"77",
          4637 => x"d7",
          4638 => x"ac",
          4639 => x"61",
          4640 => x"98",
          4641 => x"26",
          4642 => x"55",
          4643 => x"ff",
          4644 => x"ff",
          4645 => x"38",
          4646 => x"81",
          4647 => x"7e",
          4648 => x"85",
          4649 => x"80",
          4650 => x"2e",
          4651 => x"c1",
          4652 => x"76",
          4653 => x"7b",
          4654 => x"38",
          4655 => x"55",
          4656 => x"b3",
          4657 => x"54",
          4658 => x"09",
          4659 => x"38",
          4660 => x"53",
          4661 => x"51",
          4662 => x"3f",
          4663 => x"08",
          4664 => x"ac",
          4665 => x"74",
          4666 => x"18",
          4667 => x"75",
          4668 => x"39",
          4669 => x"76",
          4670 => x"7f",
          4671 => x"0c",
          4672 => x"2e",
          4673 => x"88",
          4674 => x"8c",
          4675 => x"18",
          4676 => x"07",
          4677 => x"19",
          4678 => x"11",
          4679 => x"55",
          4680 => x"08",
          4681 => x"38",
          4682 => x"7e",
          4683 => x"0c",
          4684 => x"33",
          4685 => x"55",
          4686 => x"34",
          4687 => x"81",
          4688 => x"91",
          4689 => x"ea",
          4690 => x"02",
          4691 => x"e7",
          4692 => x"3d",
          4693 => x"ff",
          4694 => x"81",
          4695 => x"56",
          4696 => x"0b",
          4697 => x"08",
          4698 => x"38",
          4699 => x"08",
          4700 => x"d3",
          4701 => x"74",
          4702 => x"87",
          4703 => x"55",
          4704 => x"75",
          4705 => x"5a",
          4706 => x"51",
          4707 => x"3f",
          4708 => x"08",
          4709 => x"70",
          4710 => x"56",
          4711 => x"8c",
          4712 => x"82",
          4713 => x"06",
          4714 => x"57",
          4715 => x"38",
          4716 => x"05",
          4717 => x"79",
          4718 => x"dd",
          4719 => x"ac",
          4720 => x"66",
          4721 => x"38",
          4722 => x"80",
          4723 => x"66",
          4724 => x"06",
          4725 => x"2e",
          4726 => x"47",
          4727 => x"77",
          4728 => x"38",
          4729 => x"92",
          4730 => x"80",
          4731 => x"38",
          4732 => x"06",
          4733 => x"2e",
          4734 => x"57",
          4735 => x"7d",
          4736 => x"fe",
          4737 => x"81",
          4738 => x"6c",
          4739 => x"53",
          4740 => x"f6",
          4741 => x"d3",
          4742 => x"81",
          4743 => x"29",
          4744 => x"62",
          4745 => x"81",
          4746 => x"30",
          4747 => x"ac",
          4748 => x"25",
          4749 => x"59",
          4750 => x"41",
          4751 => x"8a",
          4752 => x"3d",
          4753 => x"81",
          4754 => x"ff",
          4755 => x"81",
          4756 => x"ac",
          4757 => x"38",
          4758 => x"70",
          4759 => x"55",
          4760 => x"64",
          4761 => x"06",
          4762 => x"44",
          4763 => x"66",
          4764 => x"38",
          4765 => x"46",
          4766 => x"ff",
          4767 => x"bc",
          4768 => x"77",
          4769 => x"8a",
          4770 => x"81",
          4771 => x"06",
          4772 => x"80",
          4773 => x"7c",
          4774 => x"74",
          4775 => x"38",
          4776 => x"55",
          4777 => x"83",
          4778 => x"7c",
          4779 => x"93",
          4780 => x"74",
          4781 => x"84",
          4782 => x"61",
          4783 => x"81",
          4784 => x"38",
          4785 => x"65",
          4786 => x"5c",
          4787 => x"81",
          4788 => x"71",
          4789 => x"56",
          4790 => x"2e",
          4791 => x"77",
          4792 => x"81",
          4793 => x"71",
          4794 => x"22",
          4795 => x"5b",
          4796 => x"86",
          4797 => x"27",
          4798 => x"52",
          4799 => x"f4",
          4800 => x"d3",
          4801 => x"d3",
          4802 => x"10",
          4803 => x"87",
          4804 => x"fe",
          4805 => x"81",
          4806 => x"5c",
          4807 => x"0b",
          4808 => x"17",
          4809 => x"ff",
          4810 => x"27",
          4811 => x"8e",
          4812 => x"39",
          4813 => x"65",
          4814 => x"5c",
          4815 => x"81",
          4816 => x"71",
          4817 => x"56",
          4818 => x"2e",
          4819 => x"77",
          4820 => x"81",
          4821 => x"71",
          4822 => x"22",
          4823 => x"5b",
          4824 => x"86",
          4825 => x"27",
          4826 => x"52",
          4827 => x"f3",
          4828 => x"d3",
          4829 => x"84",
          4830 => x"d3",
          4831 => x"f5",
          4832 => x"81",
          4833 => x"ac",
          4834 => x"11",
          4835 => x"83",
          4836 => x"42",
          4837 => x"1e",
          4838 => x"fe",
          4839 => x"81",
          4840 => x"5c",
          4841 => x"5b",
          4842 => x"51",
          4843 => x"3f",
          4844 => x"08",
          4845 => x"06",
          4846 => x"7c",
          4847 => x"68",
          4848 => x"69",
          4849 => x"06",
          4850 => x"58",
          4851 => x"61",
          4852 => x"81",
          4853 => x"76",
          4854 => x"41",
          4855 => x"76",
          4856 => x"90",
          4857 => x"65",
          4858 => x"74",
          4859 => x"be",
          4860 => x"31",
          4861 => x"53",
          4862 => x"52",
          4863 => x"9e",
          4864 => x"ac",
          4865 => x"83",
          4866 => x"06",
          4867 => x"d3",
          4868 => x"ff",
          4869 => x"38",
          4870 => x"78",
          4871 => x"77",
          4872 => x"8e",
          4873 => x"39",
          4874 => x"09",
          4875 => x"d3",
          4876 => x"f5",
          4877 => x"38",
          4878 => x"78",
          4879 => x"80",
          4880 => x"38",
          4881 => x"f1",
          4882 => x"2a",
          4883 => x"74",
          4884 => x"38",
          4885 => x"e1",
          4886 => x"38",
          4887 => x"81",
          4888 => x"fc",
          4889 => x"57",
          4890 => x"75",
          4891 => x"93",
          4892 => x"38",
          4893 => x"81",
          4894 => x"fc",
          4895 => x"57",
          4896 => x"80",
          4897 => x"2e",
          4898 => x"83",
          4899 => x"75",
          4900 => x"75",
          4901 => x"57",
          4902 => x"38",
          4903 => x"52",
          4904 => x"9a",
          4905 => x"53",
          4906 => x"52",
          4907 => x"99",
          4908 => x"52",
          4909 => x"ff",
          4910 => x"78",
          4911 => x"34",
          4912 => x"ff",
          4913 => x"1f",
          4914 => x"f7",
          4915 => x"90",
          4916 => x"83",
          4917 => x"70",
          4918 => x"80",
          4919 => x"55",
          4920 => x"ff",
          4921 => x"65",
          4922 => x"26",
          4923 => x"80",
          4924 => x"52",
          4925 => x"ff",
          4926 => x"8a",
          4927 => x"a0",
          4928 => x"98",
          4929 => x"7f",
          4930 => x"bf",
          4931 => x"51",
          4932 => x"3f",
          4933 => x"9a",
          4934 => x"98",
          4935 => x"52",
          4936 => x"ff",
          4937 => x"61",
          4938 => x"81",
          4939 => x"38",
          4940 => x"0a",
          4941 => x"1f",
          4942 => x"a5",
          4943 => x"a4",
          4944 => x"98",
          4945 => x"52",
          4946 => x"ff",
          4947 => x"81",
          4948 => x"51",
          4949 => x"3f",
          4950 => x"1f",
          4951 => x"e3",
          4952 => x"7f",
          4953 => x"34",
          4954 => x"c2",
          4955 => x"53",
          4956 => x"52",
          4957 => x"51",
          4958 => x"3f",
          4959 => x"88",
          4960 => x"a7",
          4961 => x"97",
          4962 => x"83",
          4963 => x"52",
          4964 => x"ff",
          4965 => x"ff",
          4966 => x"05",
          4967 => x"a6",
          4968 => x"53",
          4969 => x"52",
          4970 => x"ff",
          4971 => x"82",
          4972 => x"83",
          4973 => x"ff",
          4974 => x"81",
          4975 => x"7e",
          4976 => x"ff",
          4977 => x"81",
          4978 => x"ac",
          4979 => x"38",
          4980 => x"09",
          4981 => x"f0",
          4982 => x"63",
          4983 => x"7e",
          4984 => x"ff",
          4985 => x"7d",
          4986 => x"7e",
          4987 => x"c4",
          4988 => x"85",
          4989 => x"7e",
          4990 => x"e5",
          4991 => x"85",
          4992 => x"83",
          4993 => x"ff",
          4994 => x"ff",
          4995 => x"e8",
          4996 => x"96",
          4997 => x"52",
          4998 => x"51",
          4999 => x"3f",
          5000 => x"52",
          5001 => x"51",
          5002 => x"3f",
          5003 => x"87",
          5004 => x"52",
          5005 => x"93",
          5006 => x"54",
          5007 => x"53",
          5008 => x"51",
          5009 => x"3f",
          5010 => x"52",
          5011 => x"96",
          5012 => x"56",
          5013 => x"83",
          5014 => x"06",
          5015 => x"52",
          5016 => x"95",
          5017 => x"52",
          5018 => x"ff",
          5019 => x"f0",
          5020 => x"1f",
          5021 => x"e9",
          5022 => x"87",
          5023 => x"55",
          5024 => x"83",
          5025 => x"74",
          5026 => x"ff",
          5027 => x"7b",
          5028 => x"74",
          5029 => x"38",
          5030 => x"54",
          5031 => x"52",
          5032 => x"92",
          5033 => x"d3",
          5034 => x"86",
          5035 => x"80",
          5036 => x"ff",
          5037 => x"76",
          5038 => x"31",
          5039 => x"d1",
          5040 => x"5b",
          5041 => x"ff",
          5042 => x"55",
          5043 => x"83",
          5044 => x"60",
          5045 => x"26",
          5046 => x"57",
          5047 => x"53",
          5048 => x"51",
          5049 => x"3f",
          5050 => x"08",
          5051 => x"76",
          5052 => x"31",
          5053 => x"db",
          5054 => x"61",
          5055 => x"38",
          5056 => x"83",
          5057 => x"8a",
          5058 => x"61",
          5059 => x"38",
          5060 => x"83",
          5061 => x"58",
          5062 => x"38",
          5063 => x"52",
          5064 => x"95",
          5065 => x"d4",
          5066 => x"fe",
          5067 => x"94",
          5068 => x"be",
          5069 => x"76",
          5070 => x"81",
          5071 => x"0b",
          5072 => x"77",
          5073 => x"76",
          5074 => x"63",
          5075 => x"80",
          5076 => x"76",
          5077 => x"c6",
          5078 => x"85",
          5079 => x"d3",
          5080 => x"2a",
          5081 => x"74",
          5082 => x"81",
          5083 => x"87",
          5084 => x"52",
          5085 => x"51",
          5086 => x"3f",
          5087 => x"ca",
          5088 => x"93",
          5089 => x"54",
          5090 => x"52",
          5091 => x"90",
          5092 => x"57",
          5093 => x"08",
          5094 => x"53",
          5095 => x"51",
          5096 => x"3f",
          5097 => x"d3",
          5098 => x"38",
          5099 => x"57",
          5100 => x"57",
          5101 => x"57",
          5102 => x"57",
          5103 => x"ac",
          5104 => x"0d",
          5105 => x"0d",
          5106 => x"93",
          5107 => x"38",
          5108 => x"81",
          5109 => x"52",
          5110 => x"81",
          5111 => x"ff",
          5112 => x"81",
          5113 => x"c1",
          5114 => x"80",
          5115 => x"c9",
          5116 => x"fc",
          5117 => x"93",
          5118 => x"39",
          5119 => x"51",
          5120 => x"3f",
          5121 => x"81",
          5122 => x"fe",
          5123 => x"81",
          5124 => x"c2",
          5125 => x"ff",
          5126 => x"9d",
          5127 => x"c4",
          5128 => x"e7",
          5129 => x"39",
          5130 => x"51",
          5131 => x"3f",
          5132 => x"81",
          5133 => x"fe",
          5134 => x"80",
          5135 => x"c3",
          5136 => x"ff",
          5137 => x"f1",
          5138 => x"9c",
          5139 => x"bb",
          5140 => x"39",
          5141 => x"51",
          5142 => x"3f",
          5143 => x"81",
          5144 => x"fe",
          5145 => x"80",
          5146 => x"c3",
          5147 => x"ff",
          5148 => x"c5",
          5149 => x"8c",
          5150 => x"8f",
          5151 => x"81",
          5152 => x"fe",
          5153 => x"b1",
          5154 => x"c0",
          5155 => x"fb",
          5156 => x"81",
          5157 => x"fe",
          5158 => x"9d",
          5159 => x"f0",
          5160 => x"e7",
          5161 => x"81",
          5162 => x"fe",
          5163 => x"89",
          5164 => x"94",
          5165 => x"d3",
          5166 => x"0d",
          5167 => x"0d",
          5168 => x"56",
          5169 => x"26",
          5170 => x"52",
          5171 => x"29",
          5172 => x"ca",
          5173 => x"ac",
          5174 => x"39",
          5175 => x"74",
          5176 => x"ba",
          5177 => x"ac",
          5178 => x"51",
          5179 => x"3f",
          5180 => x"08",
          5181 => x"79",
          5182 => x"81",
          5183 => x"ff",
          5184 => x"87",
          5185 => x"fe",
          5186 => x"81",
          5187 => x"81",
          5188 => x"02",
          5189 => x"e3",
          5190 => x"73",
          5191 => x"07",
          5192 => x"ff",
          5193 => x"54",
          5194 => x"57",
          5195 => x"75",
          5196 => x"81",
          5197 => x"81",
          5198 => x"d8",
          5199 => x"bc",
          5200 => x"d3",
          5201 => x"81",
          5202 => x"bb",
          5203 => x"ac",
          5204 => x"98",
          5205 => x"d3",
          5206 => x"81",
          5207 => x"d4",
          5208 => x"84",
          5209 => x"52",
          5210 => x"51",
          5211 => x"81",
          5212 => x"58",
          5213 => x"08",
          5214 => x"80",
          5215 => x"7a",
          5216 => x"58",
          5217 => x"81",
          5218 => x"d8",
          5219 => x"c1",
          5220 => x"70",
          5221 => x"25",
          5222 => x"9f",
          5223 => x"51",
          5224 => x"74",
          5225 => x"38",
          5226 => x"53",
          5227 => x"88",
          5228 => x"51",
          5229 => x"77",
          5230 => x"d3",
          5231 => x"96",
          5232 => x"f8",
          5233 => x"b7",
          5234 => x"ff",
          5235 => x"80",
          5236 => x"7a",
          5237 => x"3f",
          5238 => x"08",
          5239 => x"80",
          5240 => x"76",
          5241 => x"38",
          5242 => x"55",
          5243 => x"d3",
          5244 => x"52",
          5245 => x"2d",
          5246 => x"08",
          5247 => x"75",
          5248 => x"d3",
          5249 => x"3d",
          5250 => x"3d",
          5251 => x"05",
          5252 => x"d0",
          5253 => x"d8",
          5254 => x"81",
          5255 => x"cb",
          5256 => x"52",
          5257 => x"d6",
          5258 => x"e4",
          5259 => x"f0",
          5260 => x"33",
          5261 => x"f8",
          5262 => x"c9",
          5263 => x"2e",
          5264 => x"f6",
          5265 => x"3d",
          5266 => x"3d",
          5267 => x"96",
          5268 => x"fe",
          5269 => x"81",
          5270 => x"ff",
          5271 => x"94",
          5272 => x"f5",
          5273 => x"fe",
          5274 => x"72",
          5275 => x"81",
          5276 => x"71",
          5277 => x"38",
          5278 => x"ee",
          5279 => x"c6",
          5280 => x"f0",
          5281 => x"51",
          5282 => x"3f",
          5283 => x"70",
          5284 => x"52",
          5285 => x"95",
          5286 => x"fe",
          5287 => x"81",
          5288 => x"fe",
          5289 => x"80",
          5290 => x"af",
          5291 => x"2a",
          5292 => x"51",
          5293 => x"2e",
          5294 => x"51",
          5295 => x"3f",
          5296 => x"51",
          5297 => x"3f",
          5298 => x"ee",
          5299 => x"84",
          5300 => x"06",
          5301 => x"80",
          5302 => x"81",
          5303 => x"fb",
          5304 => x"e8",
          5305 => x"f1",
          5306 => x"fe",
          5307 => x"72",
          5308 => x"81",
          5309 => x"71",
          5310 => x"38",
          5311 => x"ed",
          5312 => x"c6",
          5313 => x"ef",
          5314 => x"51",
          5315 => x"3f",
          5316 => x"70",
          5317 => x"52",
          5318 => x"95",
          5319 => x"fe",
          5320 => x"81",
          5321 => x"fe",
          5322 => x"80",
          5323 => x"ab",
          5324 => x"2a",
          5325 => x"51",
          5326 => x"2e",
          5327 => x"51",
          5328 => x"3f",
          5329 => x"51",
          5330 => x"3f",
          5331 => x"ed",
          5332 => x"88",
          5333 => x"06",
          5334 => x"80",
          5335 => x"81",
          5336 => x"f7",
          5337 => x"b8",
          5338 => x"ed",
          5339 => x"fe",
          5340 => x"fe",
          5341 => x"84",
          5342 => x"fa",
          5343 => x"70",
          5344 => x"56",
          5345 => x"2e",
          5346 => x"8e",
          5347 => x"0c",
          5348 => x"53",
          5349 => x"81",
          5350 => x"75",
          5351 => x"72",
          5352 => x"38",
          5353 => x"30",
          5354 => x"75",
          5355 => x"72",
          5356 => x"33",
          5357 => x"2e",
          5358 => x"88",
          5359 => x"70",
          5360 => x"34",
          5361 => x"90",
          5362 => x"ec",
          5363 => x"53",
          5364 => x"54",
          5365 => x"3f",
          5366 => x"08",
          5367 => x"14",
          5368 => x"81",
          5369 => x"38",
          5370 => x"81",
          5371 => x"53",
          5372 => x"d2",
          5373 => x"72",
          5374 => x"0c",
          5375 => x"04",
          5376 => x"80",
          5377 => x"ac",
          5378 => x"5d",
          5379 => x"5a",
          5380 => x"51",
          5381 => x"3f",
          5382 => x"08",
          5383 => x"59",
          5384 => x"09",
          5385 => x"38",
          5386 => x"52",
          5387 => x"52",
          5388 => x"e7",
          5389 => x"78",
          5390 => x"1b",
          5391 => x"ab",
          5392 => x"ac",
          5393 => x"80",
          5394 => x"81",
          5395 => x"fe",
          5396 => x"85",
          5397 => x"5e",
          5398 => x"b4",
          5399 => x"ab",
          5400 => x"70",
          5401 => x"f8",
          5402 => x"80",
          5403 => x"fe",
          5404 => x"79",
          5405 => x"fe",
          5406 => x"b4",
          5407 => x"05",
          5408 => x"3f",
          5409 => x"08",
          5410 => x"90",
          5411 => x"78",
          5412 => x"85",
          5413 => x"10",
          5414 => x"ec",
          5415 => x"08",
          5416 => x"fe",
          5417 => x"fe",
          5418 => x"fe",
          5419 => x"81",
          5420 => x"8c",
          5421 => x"b8",
          5422 => x"c9",
          5423 => x"39",
          5424 => x"f0",
          5425 => x"f8",
          5426 => x"fe",
          5427 => x"d3",
          5428 => x"2e",
          5429 => x"60",
          5430 => x"80",
          5431 => x"05",
          5432 => x"80",
          5433 => x"51",
          5434 => x"3f",
          5435 => x"08",
          5436 => x"59",
          5437 => x"81",
          5438 => x"fe",
          5439 => x"81",
          5440 => x"39",
          5441 => x"51",
          5442 => x"3f",
          5443 => x"b4",
          5444 => x"11",
          5445 => x"05",
          5446 => x"f4",
          5447 => x"ac",
          5448 => x"fe",
          5449 => x"53",
          5450 => x"80",
          5451 => x"51",
          5452 => x"3f",
          5453 => x"08",
          5454 => x"f0",
          5455 => x"c5",
          5456 => x"39",
          5457 => x"f4",
          5458 => x"f8",
          5459 => x"fd",
          5460 => x"d3",
          5461 => x"2e",
          5462 => x"89",
          5463 => x"38",
          5464 => x"f0",
          5465 => x"f8",
          5466 => x"fd",
          5467 => x"d3",
          5468 => x"38",
          5469 => x"08",
          5470 => x"81",
          5471 => x"96",
          5472 => x"59",
          5473 => x"3f",
          5474 => x"33",
          5475 => x"60",
          5476 => x"81",
          5477 => x"51",
          5478 => x"3f",
          5479 => x"08",
          5480 => x"38",
          5481 => x"08",
          5482 => x"3f",
          5483 => x"81",
          5484 => x"fe",
          5485 => x"81",
          5486 => x"39",
          5487 => x"f8",
          5488 => x"e4",
          5489 => x"d3",
          5490 => x"3d",
          5491 => x"52",
          5492 => x"fa",
          5493 => x"81",
          5494 => x"52",
          5495 => x"a7",
          5496 => x"ac",
          5497 => x"fc",
          5498 => x"d3",
          5499 => x"f3",
          5500 => x"e5",
          5501 => x"fe",
          5502 => x"fe",
          5503 => x"81",
          5504 => x"b5",
          5505 => x"05",
          5506 => x"e4",
          5507 => x"d3",
          5508 => x"3d",
          5509 => x"52",
          5510 => x"b2",
          5511 => x"ac",
          5512 => x"fe",
          5513 => x"59",
          5514 => x"3f",
          5515 => x"58",
          5516 => x"57",
          5517 => x"55",
          5518 => x"08",
          5519 => x"54",
          5520 => x"52",
          5521 => x"fb",
          5522 => x"ac",
          5523 => x"fc",
          5524 => x"d3",
          5525 => x"f2",
          5526 => x"fd",
          5527 => x"fc",
          5528 => x"a7",
          5529 => x"fe",
          5530 => x"fb",
          5531 => x"c9",
          5532 => x"f3",
          5533 => x"51",
          5534 => x"3f",
          5535 => x"84",
          5536 => x"87",
          5537 => x"0c",
          5538 => x"0b",
          5539 => x"94",
          5540 => x"ac",
          5541 => x"f3",
          5542 => x"39",
          5543 => x"51",
          5544 => x"3f",
          5545 => x"0b",
          5546 => x"84",
          5547 => x"83",
          5548 => x"94",
          5549 => x"a1",
          5550 => x"fe",
          5551 => x"fe",
          5552 => x"fe",
          5553 => x"81",
          5554 => x"80",
          5555 => x"38",
          5556 => x"c9",
          5557 => x"f8",
          5558 => x"59",
          5559 => x"3d",
          5560 => x"53",
          5561 => x"51",
          5562 => x"3f",
          5563 => x"08",
          5564 => x"e5",
          5565 => x"81",
          5566 => x"fe",
          5567 => x"60",
          5568 => x"81",
          5569 => x"5e",
          5570 => x"08",
          5571 => x"c9",
          5572 => x"ac",
          5573 => x"ca",
          5574 => x"f7",
          5575 => x"b9",
          5576 => x"a8",
          5577 => x"e3",
          5578 => x"d5",
          5579 => x"39",
          5580 => x"51",
          5581 => x"3f",
          5582 => x"a0",
          5583 => x"84",
          5584 => x"39",
          5585 => x"51",
          5586 => x"2e",
          5587 => x"7c",
          5588 => x"78",
          5589 => x"cb",
          5590 => x"fe",
          5591 => x"fe",
          5592 => x"81",
          5593 => x"81",
          5594 => x"55",
          5595 => x"54",
          5596 => x"ca",
          5597 => x"3d",
          5598 => x"fe",
          5599 => x"81",
          5600 => x"81",
          5601 => x"80",
          5602 => x"05",
          5603 => x"80",
          5604 => x"80",
          5605 => x"80",
          5606 => x"f4",
          5607 => x"d3",
          5608 => x"7c",
          5609 => x"81",
          5610 => x"78",
          5611 => x"ff",
          5612 => x"06",
          5613 => x"81",
          5614 => x"fe",
          5615 => x"f9",
          5616 => x"3d",
          5617 => x"81",
          5618 => x"9b",
          5619 => x"0b",
          5620 => x"8c",
          5621 => x"86",
          5622 => x"c0",
          5623 => x"8c",
          5624 => x"87",
          5625 => x"0c",
          5626 => x"0b",
          5627 => x"94",
          5628 => x"0b",
          5629 => x"0c",
          5630 => x"81",
          5631 => x"fe",
          5632 => x"fe",
          5633 => x"81",
          5634 => x"fe",
          5635 => x"81",
          5636 => x"fe",
          5637 => x"81",
          5638 => x"fe",
          5639 => x"81",
          5640 => x"3f",
          5641 => x"80",
          5642 => x"0f",
          5643 => x"0f",
          5644 => x"0f",
          5645 => x"0f",
          5646 => x"0f",
          5647 => x"0f",
          5648 => x"11",
          5649 => x"11",
          5650 => x"11",
          5651 => x"11",
          5652 => x"11",
          5653 => x"11",
          5654 => x"11",
          5655 => x"11",
          5656 => x"11",
          5657 => x"11",
          5658 => x"11",
          5659 => x"11",
          5660 => x"11",
          5661 => x"11",
          5662 => x"11",
          5663 => x"11",
          5664 => x"11",
          5665 => x"11",
          5666 => x"11",
          5667 => x"11",
          5668 => x"11",
          5669 => x"11",
          5670 => x"11",
          5671 => x"50",
          5672 => x"4f",
          5673 => x"4f",
          5674 => x"4f",
          5675 => x"4f",
          5676 => x"50",
          5677 => x"50",
          5678 => x"50",
          5679 => x"50",
          5680 => x"50",
          5681 => x"50",
          5682 => x"50",
          5683 => x"50",
          5684 => x"50",
          5685 => x"50",
          5686 => x"50",
          5687 => x"50",
          5688 => x"50",
          5689 => x"50",
          5690 => x"50",
          5691 => x"54",
          5692 => x"57",
          5693 => x"54",
          5694 => x"57",
          5695 => x"55",
          5696 => x"57",
          5697 => x"57",
          5698 => x"57",
          5699 => x"57",
          5700 => x"57",
          5701 => x"57",
          5702 => x"57",
          5703 => x"57",
          5704 => x"57",
          5705 => x"57",
          5706 => x"57",
          5707 => x"57",
          5708 => x"57",
          5709 => x"57",
          5710 => x"57",
          5711 => x"55",
          5712 => x"57",
          5713 => x"57",
          5714 => x"57",
          5715 => x"57",
          5716 => x"57",
          5717 => x"57",
          5718 => x"57",
          5719 => x"57",
          5720 => x"57",
          5721 => x"57",
          5722 => x"57",
          5723 => x"57",
          5724 => x"57",
          5725 => x"57",
          5726 => x"57",
          5727 => x"57",
          5728 => x"57",
          5729 => x"57",
          5730 => x"57",
          5731 => x"57",
          5732 => x"57",
          5733 => x"57",
          5734 => x"55",
          5735 => x"57",
          5736 => x"57",
          5737 => x"57",
          5738 => x"57",
          5739 => x"55",
          5740 => x"57",
          5741 => x"57",
          5742 => x"57",
          5743 => x"57",
          5744 => x"57",
          5745 => x"57",
          5746 => x"57",
          5747 => x"57",
          5748 => x"57",
          5749 => x"57",
          5750 => x"57",
          5751 => x"57",
          5752 => x"57",
          5753 => x"57",
          5754 => x"57",
          5755 => x"57",
          5756 => x"57",
          5757 => x"57",
          5758 => x"57",
          5759 => x"57",
          5760 => x"57",
          5761 => x"57",
          5762 => x"57",
          5763 => x"57",
          5764 => x"57",
          5765 => x"57",
          5766 => x"57",
          5767 => x"57",
          5768 => x"57",
          5769 => x"57",
          5770 => x"57",
          5771 => x"56",
          5772 => x"56",
          5773 => x"57",
          5774 => x"57",
          5775 => x"56",
          5776 => x"56",
          5777 => x"57",
          5778 => x"57",
          5779 => x"57",
          5780 => x"57",
          5781 => x"57",
          5782 => x"57",
          5783 => x"57",
          5784 => x"57",
          5785 => x"57",
          5786 => x"57",
          5787 => x"57",
          5788 => x"57",
          5789 => x"57",
          5790 => x"57",
          5791 => x"57",
          5792 => x"57",
          5793 => x"57",
          5794 => x"57",
          5795 => x"57",
          5796 => x"57",
          5797 => x"57",
          5798 => x"57",
          5799 => x"57",
          5800 => x"57",
          5801 => x"57",
          5802 => x"57",
          5803 => x"57",
          5804 => x"57",
          5805 => x"57",
          5806 => x"57",
          5807 => x"57",
          5808 => x"57",
          5809 => x"57",
          5810 => x"57",
          5811 => x"56",
          5812 => x"56",
          5813 => x"57",
          5814 => x"57",
          5815 => x"57",
          5816 => x"57",
          5817 => x"57",
          5818 => x"57",
          5819 => x"57",
          5820 => x"57",
          5821 => x"57",
          5822 => x"57",
          5823 => x"57",
          5824 => x"57",
          5825 => x"57",
          5826 => x"54",
          5827 => x"2f",
          5828 => x"25",
          5829 => x"64",
          5830 => x"3a",
          5831 => x"25",
          5832 => x"0a",
          5833 => x"43",
          5834 => x"6e",
          5835 => x"75",
          5836 => x"69",
          5837 => x"00",
          5838 => x"66",
          5839 => x"20",
          5840 => x"20",
          5841 => x"66",
          5842 => x"00",
          5843 => x"44",
          5844 => x"63",
          5845 => x"69",
          5846 => x"65",
          5847 => x"74",
          5848 => x"0a",
          5849 => x"20",
          5850 => x"53",
          5851 => x"52",
          5852 => x"28",
          5853 => x"72",
          5854 => x"30",
          5855 => x"20",
          5856 => x"65",
          5857 => x"38",
          5858 => x"0a",
          5859 => x"20",
          5860 => x"41",
          5861 => x"53",
          5862 => x"74",
          5863 => x"38",
          5864 => x"53",
          5865 => x"3d",
          5866 => x"58",
          5867 => x"00",
          5868 => x"20",
          5869 => x"4d",
          5870 => x"74",
          5871 => x"3d",
          5872 => x"58",
          5873 => x"69",
          5874 => x"25",
          5875 => x"29",
          5876 => x"00",
          5877 => x"20",
          5878 => x"43",
          5879 => x"00",
          5880 => x"20",
          5881 => x"32",
          5882 => x"00",
          5883 => x"20",
          5884 => x"49",
          5885 => x"00",
          5886 => x"20",
          5887 => x"20",
          5888 => x"64",
          5889 => x"65",
          5890 => x"65",
          5891 => x"30",
          5892 => x"2e",
          5893 => x"00",
          5894 => x"20",
          5895 => x"54",
          5896 => x"55",
          5897 => x"43",
          5898 => x"52",
          5899 => x"45",
          5900 => x"00",
          5901 => x"20",
          5902 => x"4d",
          5903 => x"20",
          5904 => x"6d",
          5905 => x"3d",
          5906 => x"58",
          5907 => x"00",
          5908 => x"64",
          5909 => x"73",
          5910 => x"0a",
          5911 => x"20",
          5912 => x"55",
          5913 => x"73",
          5914 => x"56",
          5915 => x"6f",
          5916 => x"64",
          5917 => x"73",
          5918 => x"20",
          5919 => x"58",
          5920 => x"00",
          5921 => x"20",
          5922 => x"55",
          5923 => x"6d",
          5924 => x"20",
          5925 => x"72",
          5926 => x"64",
          5927 => x"73",
          5928 => x"20",
          5929 => x"58",
          5930 => x"00",
          5931 => x"20",
          5932 => x"61",
          5933 => x"53",
          5934 => x"74",
          5935 => x"64",
          5936 => x"73",
          5937 => x"20",
          5938 => x"20",
          5939 => x"58",
          5940 => x"00",
          5941 => x"20",
          5942 => x"55",
          5943 => x"20",
          5944 => x"20",
          5945 => x"20",
          5946 => x"20",
          5947 => x"20",
          5948 => x"20",
          5949 => x"58",
          5950 => x"00",
          5951 => x"20",
          5952 => x"73",
          5953 => x"20",
          5954 => x"63",
          5955 => x"72",
          5956 => x"20",
          5957 => x"20",
          5958 => x"20",
          5959 => x"58",
          5960 => x"00",
          5961 => x"61",
          5962 => x"00",
          5963 => x"64",
          5964 => x"00",
          5965 => x"65",
          5966 => x"00",
          5967 => x"4f",
          5968 => x"4f",
          5969 => x"00",
          5970 => x"6b",
          5971 => x"6e",
          5972 => x"00",
          5973 => x"2b",
          5974 => x"3c",
          5975 => x"5b",
          5976 => x"00",
          5977 => x"54",
          5978 => x"54",
          5979 => x"00",
          5980 => x"00",
          5981 => x"00",
          5982 => x"00",
          5983 => x"00",
          5984 => x"00",
          5985 => x"00",
          5986 => x"00",
          5987 => x"00",
          5988 => x"00",
          5989 => x"0a",
          5990 => x"90",
          5991 => x"4f",
          5992 => x"30",
          5993 => x"20",
          5994 => x"45",
          5995 => x"20",
          5996 => x"33",
          5997 => x"20",
          5998 => x"20",
          5999 => x"45",
          6000 => x"20",
          6001 => x"20",
          6002 => x"20",
          6003 => x"5d",
          6004 => x"00",
          6005 => x"00",
          6006 => x"00",
          6007 => x"45",
          6008 => x"8f",
          6009 => x"45",
          6010 => x"8e",
          6011 => x"92",
          6012 => x"55",
          6013 => x"9a",
          6014 => x"9e",
          6015 => x"4f",
          6016 => x"a6",
          6017 => x"aa",
          6018 => x"ae",
          6019 => x"b2",
          6020 => x"b6",
          6021 => x"ba",
          6022 => x"be",
          6023 => x"c2",
          6024 => x"c6",
          6025 => x"ca",
          6026 => x"ce",
          6027 => x"d2",
          6028 => x"d6",
          6029 => x"da",
          6030 => x"de",
          6031 => x"e2",
          6032 => x"e6",
          6033 => x"ea",
          6034 => x"ee",
          6035 => x"f2",
          6036 => x"f6",
          6037 => x"fa",
          6038 => x"fe",
          6039 => x"2c",
          6040 => x"5d",
          6041 => x"2a",
          6042 => x"3f",
          6043 => x"00",
          6044 => x"00",
          6045 => x"00",
          6046 => x"02",
          6047 => x"00",
          6048 => x"00",
          6049 => x"00",
          6050 => x"00",
          6051 => x"00",
          6052 => x"54",
          6053 => x"00",
          6054 => x"54",
          6055 => x"00",
          6056 => x"46",
          6057 => x"00",
          6058 => x"53",
          6059 => x"4f",
          6060 => x"4e",
          6061 => x"4c",
          6062 => x"00",
          6063 => x"53",
          6064 => x"55",
          6065 => x"52",
          6066 => x"4e",
          6067 => x"4c",
          6068 => x"00",
          6069 => x"4c",
          6070 => x"53",
          6071 => x"20",
          6072 => x"54",
          6073 => x"53",
          6074 => x"4d",
          6075 => x"00",
          6076 => x"52",
          6077 => x"52",
          6078 => x"00",
          6079 => x"53",
          6080 => x"47",
          6081 => x"45",
          6082 => x"49",
          6083 => x"00",
          6084 => x"53",
          6085 => x"4f",
          6086 => x"4e",
          6087 => x"00",
          6088 => x"75",
          6089 => x"00",
          6090 => x"6e",
          6091 => x"00",
          6092 => x"74",
          6093 => x"00",
          6094 => x"6f",
          6095 => x"00",
          6096 => x"75",
          6097 => x"00",
          6098 => x"64",
          6099 => x"00",
          6100 => x"65",
          6101 => x"00",
          6102 => x"72",
          6103 => x"00",
          6104 => x"69",
          6105 => x"00",
          6106 => x"65",
          6107 => x"00",
          6108 => x"6e",
          6109 => x"00",
          6110 => x"70",
          6111 => x"00",
          6112 => x"6c",
          6113 => x"00",
          6114 => x"65",
          6115 => x"00",
          6116 => x"65",
          6117 => x"00",
          6118 => x"6e",
          6119 => x"63",
          6120 => x"00",
          6121 => x"72",
          6122 => x"00",
          6123 => x"72",
          6124 => x"00",
          6125 => x"6c",
          6126 => x"00",
          6127 => x"74",
          6128 => x"00",
          6129 => x"69",
          6130 => x"00",
          6131 => x"65",
          6132 => x"65",
          6133 => x"65",
          6134 => x"00",
          6135 => x"6b",
          6136 => x"00",
          6137 => x"74",
          6138 => x"00",
          6139 => x"69",
          6140 => x"00",
          6141 => x"61",
          6142 => x"00",
          6143 => x"70",
          6144 => x"6f",
          6145 => x"74",
          6146 => x"74",
          6147 => x"74",
          6148 => x"6f",
          6149 => x"00",
          6150 => x"78",
          6151 => x"00",
          6152 => x"61",
          6153 => x"00",
          6154 => x"75",
          6155 => x"00",
          6156 => x"64",
          6157 => x"72",
          6158 => x"00",
          6159 => x"68",
          6160 => x"69",
          6161 => x"00",
          6162 => x"61",
          6163 => x"00",
          6164 => x"6b",
          6165 => x"00",
          6166 => x"6c",
          6167 => x"00",
          6168 => x"75",
          6169 => x"00",
          6170 => x"62",
          6171 => x"68",
          6172 => x"77",
          6173 => x"64",
          6174 => x"65",
          6175 => x"00",
          6176 => x"00",
          6177 => x"64",
          6178 => x"65",
          6179 => x"72",
          6180 => x"00",
          6181 => x"72",
          6182 => x"72",
          6183 => x"00",
          6184 => x"6c",
          6185 => x"00",
          6186 => x"70",
          6187 => x"73",
          6188 => x"74",
          6189 => x"73",
          6190 => x"00",
          6191 => x"6c",
          6192 => x"00",
          6193 => x"66",
          6194 => x"00",
          6195 => x"6d",
          6196 => x"00",
          6197 => x"73",
          6198 => x"00",
          6199 => x"73",
          6200 => x"72",
          6201 => x"0a",
          6202 => x"74",
          6203 => x"61",
          6204 => x"72",
          6205 => x"2e",
          6206 => x"00",
          6207 => x"73",
          6208 => x"6f",
          6209 => x"65",
          6210 => x"2e",
          6211 => x"00",
          6212 => x"20",
          6213 => x"65",
          6214 => x"75",
          6215 => x"0a",
          6216 => x"20",
          6217 => x"68",
          6218 => x"75",
          6219 => x"0a",
          6220 => x"76",
          6221 => x"64",
          6222 => x"6c",
          6223 => x"6d",
          6224 => x"00",
          6225 => x"63",
          6226 => x"20",
          6227 => x"69",
          6228 => x"0a",
          6229 => x"6c",
          6230 => x"6c",
          6231 => x"64",
          6232 => x"78",
          6233 => x"73",
          6234 => x"00",
          6235 => x"6c",
          6236 => x"61",
          6237 => x"65",
          6238 => x"76",
          6239 => x"64",
          6240 => x"00",
          6241 => x"20",
          6242 => x"77",
          6243 => x"65",
          6244 => x"6f",
          6245 => x"74",
          6246 => x"0a",
          6247 => x"69",
          6248 => x"6e",
          6249 => x"65",
          6250 => x"73",
          6251 => x"76",
          6252 => x"64",
          6253 => x"00",
          6254 => x"73",
          6255 => x"6f",
          6256 => x"6e",
          6257 => x"65",
          6258 => x"00",
          6259 => x"20",
          6260 => x"70",
          6261 => x"62",
          6262 => x"66",
          6263 => x"73",
          6264 => x"65",
          6265 => x"6f",
          6266 => x"20",
          6267 => x"64",
          6268 => x"2e",
          6269 => x"00",
          6270 => x"72",
          6271 => x"20",
          6272 => x"72",
          6273 => x"2e",
          6274 => x"00",
          6275 => x"6d",
          6276 => x"74",
          6277 => x"70",
          6278 => x"74",
          6279 => x"20",
          6280 => x"63",
          6281 => x"65",
          6282 => x"00",
          6283 => x"6c",
          6284 => x"73",
          6285 => x"63",
          6286 => x"2e",
          6287 => x"00",
          6288 => x"73",
          6289 => x"69",
          6290 => x"6e",
          6291 => x"65",
          6292 => x"79",
          6293 => x"00",
          6294 => x"6f",
          6295 => x"6e",
          6296 => x"70",
          6297 => x"66",
          6298 => x"73",
          6299 => x"00",
          6300 => x"72",
          6301 => x"74",
          6302 => x"20",
          6303 => x"6f",
          6304 => x"63",
          6305 => x"00",
          6306 => x"63",
          6307 => x"73",
          6308 => x"00",
          6309 => x"6b",
          6310 => x"6e",
          6311 => x"72",
          6312 => x"0a",
          6313 => x"6c",
          6314 => x"79",
          6315 => x"20",
          6316 => x"61",
          6317 => x"6c",
          6318 => x"79",
          6319 => x"2f",
          6320 => x"2e",
          6321 => x"00",
          6322 => x"61",
          6323 => x"00",
          6324 => x"55",
          6325 => x"00",
          6326 => x"2a",
          6327 => x"20",
          6328 => x"00",
          6329 => x"2f",
          6330 => x"32",
          6331 => x"00",
          6332 => x"2e",
          6333 => x"00",
          6334 => x"50",
          6335 => x"72",
          6336 => x"25",
          6337 => x"29",
          6338 => x"20",
          6339 => x"2a",
          6340 => x"00",
          6341 => x"55",
          6342 => x"49",
          6343 => x"72",
          6344 => x"74",
          6345 => x"6e",
          6346 => x"72",
          6347 => x"00",
          6348 => x"6d",
          6349 => x"69",
          6350 => x"72",
          6351 => x"74",
          6352 => x"00",
          6353 => x"32",
          6354 => x"74",
          6355 => x"75",
          6356 => x"00",
          6357 => x"43",
          6358 => x"52",
          6359 => x"6e",
          6360 => x"72",
          6361 => x"0a",
          6362 => x"43",
          6363 => x"57",
          6364 => x"6e",
          6365 => x"72",
          6366 => x"0a",
          6367 => x"52",
          6368 => x"52",
          6369 => x"6e",
          6370 => x"72",
          6371 => x"0a",
          6372 => x"52",
          6373 => x"54",
          6374 => x"6e",
          6375 => x"72",
          6376 => x"0a",
          6377 => x"52",
          6378 => x"52",
          6379 => x"6e",
          6380 => x"72",
          6381 => x"0a",
          6382 => x"52",
          6383 => x"54",
          6384 => x"6e",
          6385 => x"72",
          6386 => x"0a",
          6387 => x"74",
          6388 => x"67",
          6389 => x"20",
          6390 => x"65",
          6391 => x"2e",
          6392 => x"00",
          6393 => x"61",
          6394 => x"6e",
          6395 => x"69",
          6396 => x"2e",
          6397 => x"00",
          6398 => x"00",
          6399 => x"69",
          6400 => x"20",
          6401 => x"69",
          6402 => x"69",
          6403 => x"73",
          6404 => x"64",
          6405 => x"72",
          6406 => x"2c",
          6407 => x"65",
          6408 => x"20",
          6409 => x"74",
          6410 => x"6e",
          6411 => x"6c",
          6412 => x"00",
          6413 => x"00",
          6414 => x"64",
          6415 => x"73",
          6416 => x"64",
          6417 => x"00",
          6418 => x"69",
          6419 => x"6c",
          6420 => x"64",
          6421 => x"00",
          6422 => x"69",
          6423 => x"20",
          6424 => x"69",
          6425 => x"69",
          6426 => x"73",
          6427 => x"00",
          6428 => x"3d",
          6429 => x"00",
          6430 => x"3a",
          6431 => x"73",
          6432 => x"69",
          6433 => x"69",
          6434 => x"72",
          6435 => x"74",
          6436 => x"00",
          6437 => x"61",
          6438 => x"6e",
          6439 => x"6e",
          6440 => x"72",
          6441 => x"73",
          6442 => x"00",
          6443 => x"73",
          6444 => x"65",
          6445 => x"61",
          6446 => x"66",
          6447 => x"0a",
          6448 => x"61",
          6449 => x"6e",
          6450 => x"61",
          6451 => x"66",
          6452 => x"0a",
          6453 => x"65",
          6454 => x"69",
          6455 => x"63",
          6456 => x"20",
          6457 => x"30",
          6458 => x"2e",
          6459 => x"00",
          6460 => x"6c",
          6461 => x"67",
          6462 => x"64",
          6463 => x"20",
          6464 => x"78",
          6465 => x"2e",
          6466 => x"00",
          6467 => x"6c",
          6468 => x"65",
          6469 => x"6e",
          6470 => x"63",
          6471 => x"20",
          6472 => x"29",
          6473 => x"00",
          6474 => x"73",
          6475 => x"74",
          6476 => x"20",
          6477 => x"6c",
          6478 => x"74",
          6479 => x"2e",
          6480 => x"00",
          6481 => x"6c",
          6482 => x"65",
          6483 => x"74",
          6484 => x"2e",
          6485 => x"00",
          6486 => x"55",
          6487 => x"6e",
          6488 => x"3a",
          6489 => x"5c",
          6490 => x"25",
          6491 => x"00",
          6492 => x"64",
          6493 => x"6d",
          6494 => x"64",
          6495 => x"00",
          6496 => x"6e",
          6497 => x"67",
          6498 => x"0a",
          6499 => x"61",
          6500 => x"6e",
          6501 => x"6e",
          6502 => x"72",
          6503 => x"73",
          6504 => x"0a",
          6505 => x"00",
          6506 => x"00",
          6507 => x"7f",
          6508 => x"00",
          6509 => x"7f",
          6510 => x"00",
          6511 => x"7f",
          6512 => x"00",
          6513 => x"00",
          6514 => x"78",
          6515 => x"00",
          6516 => x"e1",
          6517 => x"01",
          6518 => x"01",
          6519 => x"01",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"5f",
          6524 => x"01",
          6525 => x"00",
          6526 => x"00",
          6527 => x"5f",
          6528 => x"01",
          6529 => x"00",
          6530 => x"00",
          6531 => x"5f",
          6532 => x"01",
          6533 => x"00",
          6534 => x"00",
          6535 => x"5f",
          6536 => x"01",
          6537 => x"00",
          6538 => x"00",
          6539 => x"5f",
          6540 => x"02",
          6541 => x"00",
          6542 => x"00",
          6543 => x"5f",
          6544 => x"02",
          6545 => x"00",
          6546 => x"00",
          6547 => x"5f",
          6548 => x"02",
          6549 => x"00",
          6550 => x"00",
          6551 => x"5f",
          6552 => x"02",
          6553 => x"00",
          6554 => x"00",
          6555 => x"5f",
          6556 => x"02",
          6557 => x"00",
          6558 => x"00",
          6559 => x"5f",
          6560 => x"02",
          6561 => x"00",
          6562 => x"00",
          6563 => x"5f",
          6564 => x"03",
          6565 => x"00",
          6566 => x"00",
          6567 => x"5f",
          6568 => x"03",
          6569 => x"00",
          6570 => x"00",
          6571 => x"5f",
          6572 => x"03",
          6573 => x"00",
          6574 => x"00",
          6575 => x"5f",
          6576 => x"03",
          6577 => x"00",
          6578 => x"00",
          6579 => x"5f",
          6580 => x"03",
          6581 => x"00",
          6582 => x"00",
          6583 => x"5f",
          6584 => x"03",
          6585 => x"00",
          6586 => x"00",
          6587 => x"5f",
          6588 => x"03",
          6589 => x"00",
          6590 => x"00",
          6591 => x"5f",
          6592 => x"03",
          6593 => x"00",
          6594 => x"00",
          6595 => x"5f",
          6596 => x"03",
          6597 => x"00",
          6598 => x"00",
          6599 => x"5f",
          6600 => x"03",
          6601 => x"00",
          6602 => x"00",
          6603 => x"5f",
          6604 => x"03",
          6605 => x"00",
          6606 => x"00",
          6607 => x"5f",
          6608 => x"03",
          6609 => x"00",
          6610 => x"00",
          6611 => x"5f",
          6612 => x"03",
          6613 => x"00",
          6614 => x"00",
          6615 => x"5f",
          6616 => x"03",
          6617 => x"00",
          6618 => x"00",
          6619 => x"5f",
          6620 => x"03",
          6621 => x"00",
          6622 => x"00",
          6623 => x"5f",
          6624 => x"03",
          6625 => x"00",
          6626 => x"00",
          6627 => x"5f",
          6628 => x"03",
          6629 => x"00",
          6630 => x"00",
          6631 => x"5f",
          6632 => x"03",
          6633 => x"00",
          6634 => x"00",
          6635 => x"60",
          6636 => x"03",
          6637 => x"00",
          6638 => x"00",
          6639 => x"60",
          6640 => x"03",
          6641 => x"00",
          6642 => x"00",
          6643 => x"60",
          6644 => x"03",
          6645 => x"00",
          6646 => x"00",
          6647 => x"60",
          6648 => x"03",
          6649 => x"00",
          6650 => x"00",
          6651 => x"60",
          6652 => x"03",
          6653 => x"00",
          6654 => x"00",
          6655 => x"60",
          6656 => x"03",
          6657 => x"00",
          6658 => x"00",
          6659 => x"60",
          6660 => x"03",
          6661 => x"00",
          6662 => x"00",
          6663 => x"60",
          6664 => x"03",
          6665 => x"00",
          6666 => x"00",
          6667 => x"60",
          6668 => x"03",
          6669 => x"00",
          6670 => x"00",
          6671 => x"60",
          6672 => x"03",
          6673 => x"00",
          6674 => x"00",
          6675 => x"60",
          6676 => x"03",
          6677 => x"00",
          6678 => x"00",
          6679 => x"60",
          6680 => x"04",
          6681 => x"00",
          6682 => x"00",
          6683 => x"60",
          6684 => x"04",
          6685 => x"00",
          6686 => x"00",
          6687 => x"60",
          6688 => x"04",
          6689 => x"00",
          6690 => x"00",
          6691 => x"60",
          6692 => x"04",
          6693 => x"00",
          6694 => x"00",
          6695 => x"60",
          6696 => x"04",
          6697 => x"00",
          6698 => x"00",
          6699 => x"60",
          6700 => x"05",
          6701 => x"00",
          6702 => x"00",
          6703 => x"60",
          6704 => x"05",
          6705 => x"00",
          6706 => x"00",
          6707 => x"60",
          6708 => x"05",
          6709 => x"00",
          6710 => x"00",
          6711 => x"60",
          6712 => x"05",
          6713 => x"00",
          6714 => x"00",
          6715 => x"60",
          6716 => x"05",
          6717 => x"00",
          6718 => x"00",
          6719 => x"60",
          6720 => x"05",
          6721 => x"00",
          6722 => x"00",
          6723 => x"60",
          6724 => x"06",
          6725 => x"00",
          6726 => x"00",
          6727 => x"60",
          6728 => x"06",
          6729 => x"00",
          6730 => x"00",
          6731 => x"60",
          6732 => x"07",
          6733 => x"00",
          6734 => x"00",
          6735 => x"60",
          6736 => x"07",
          6737 => x"00",
          6738 => x"00",
          6739 => x"60",
          6740 => x"08",
          6741 => x"00",
          6742 => x"00",
          6743 => x"60",
          6744 => x"08",
          6745 => x"00",
          6746 => x"00",
          6747 => x"60",
          6748 => x"08",
          6749 => x"00",
          6750 => x"00",
          6751 => x"60",
          6752 => x"08",
          6753 => x"00",
          6754 => x"00",
          6755 => x"60",
          6756 => x"08",
          6757 => x"00",
          6758 => x"00",
          6759 => x"60",
          6760 => x"08",
          6761 => x"00",
          6762 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"89",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"84",
            11 => x"0b",
            12 => x"04",
            13 => x"84",
            14 => x"0b",
            15 => x"04",
            16 => x"84",
            17 => x"0b",
            18 => x"04",
            19 => x"84",
            20 => x"0b",
            21 => x"04",
            22 => x"84",
            23 => x"0b",
            24 => x"04",
            25 => x"85",
            26 => x"0b",
            27 => x"04",
            28 => x"85",
            29 => x"0b",
            30 => x"04",
            31 => x"85",
            32 => x"0b",
            33 => x"04",
            34 => x"85",
            35 => x"0b",
            36 => x"04",
            37 => x"86",
            38 => x"0b",
            39 => x"04",
            40 => x"86",
            41 => x"0b",
            42 => x"04",
            43 => x"86",
            44 => x"0b",
            45 => x"04",
            46 => x"86",
            47 => x"0b",
            48 => x"04",
            49 => x"87",
            50 => x"0b",
            51 => x"04",
            52 => x"87",
            53 => x"0b",
            54 => x"04",
            55 => x"87",
            56 => x"0b",
            57 => x"04",
            58 => x"87",
            59 => x"0b",
            60 => x"04",
            61 => x"88",
            62 => x"0b",
            63 => x"04",
            64 => x"88",
            65 => x"0b",
            66 => x"04",
            67 => x"88",
            68 => x"0b",
            69 => x"04",
            70 => x"88",
            71 => x"0b",
            72 => x"04",
            73 => x"89",
            74 => x"0b",
            75 => x"04",
            76 => x"89",
            77 => x"0b",
            78 => x"04",
            79 => x"89",
            80 => x"0b",
            81 => x"04",
            82 => x"89",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"84",
           129 => x"d3",
           130 => x"e7",
           131 => x"b8",
           132 => x"90",
           133 => x"b8",
           134 => x"2d",
           135 => x"08",
           136 => x"04",
           137 => x"0c",
           138 => x"81",
           139 => x"83",
           140 => x"81",
           141 => x"a0",
           142 => x"d3",
           143 => x"80",
           144 => x"d3",
           145 => x"de",
           146 => x"b8",
           147 => x"90",
           148 => x"b8",
           149 => x"2d",
           150 => x"08",
           151 => x"04",
           152 => x"0c",
           153 => x"81",
           154 => x"83",
           155 => x"81",
           156 => x"a8",
           157 => x"d3",
           158 => x"80",
           159 => x"d3",
           160 => x"a5",
           161 => x"b8",
           162 => x"90",
           163 => x"b8",
           164 => x"2d",
           165 => x"08",
           166 => x"04",
           167 => x"0c",
           168 => x"81",
           169 => x"83",
           170 => x"81",
           171 => x"a6",
           172 => x"d3",
           173 => x"80",
           174 => x"d3",
           175 => x"e7",
           176 => x"b8",
           177 => x"90",
           178 => x"b8",
           179 => x"2d",
           180 => x"08",
           181 => x"04",
           182 => x"0c",
           183 => x"81",
           184 => x"83",
           185 => x"81",
           186 => x"90",
           187 => x"d3",
           188 => x"80",
           189 => x"d3",
           190 => x"d1",
           191 => x"b8",
           192 => x"90",
           193 => x"b8",
           194 => x"d9",
           195 => x"b8",
           196 => x"90",
           197 => x"b8",
           198 => x"d0",
           199 => x"b8",
           200 => x"90",
           201 => x"b8",
           202 => x"df",
           203 => x"b8",
           204 => x"90",
           205 => x"b8",
           206 => x"c6",
           207 => x"b8",
           208 => x"90",
           209 => x"b8",
           210 => x"f9",
           211 => x"b8",
           212 => x"90",
           213 => x"b8",
           214 => x"ed",
           215 => x"b8",
           216 => x"90",
           217 => x"b8",
           218 => x"81",
           219 => x"b8",
           220 => x"90",
           221 => x"b8",
           222 => x"a4",
           223 => x"b8",
           224 => x"90",
           225 => x"b8",
           226 => x"c8",
           227 => x"b8",
           228 => x"90",
           229 => x"b8",
           230 => x"f1",
           231 => x"b8",
           232 => x"90",
           233 => x"b8",
           234 => x"81",
           235 => x"b8",
           236 => x"90",
           237 => x"b8",
           238 => x"f9",
           239 => x"b8",
           240 => x"90",
           241 => x"b8",
           242 => x"da",
           243 => x"b8",
           244 => x"90",
           245 => x"b8",
           246 => x"e7",
           247 => x"b8",
           248 => x"90",
           249 => x"b8",
           250 => x"de",
           251 => x"b8",
           252 => x"90",
           253 => x"b8",
           254 => x"e4",
           255 => x"b8",
           256 => x"90",
           257 => x"b8",
           258 => x"b0",
           259 => x"b8",
           260 => x"90",
           261 => x"b8",
           262 => x"89",
           263 => x"b8",
           264 => x"90",
           265 => x"b8",
           266 => x"b3",
           267 => x"b8",
           268 => x"90",
           269 => x"b8",
           270 => x"c1",
           271 => x"b8",
           272 => x"90",
           273 => x"b8",
           274 => x"dd",
           275 => x"b8",
           276 => x"90",
           277 => x"b8",
           278 => x"e8",
           279 => x"b8",
           280 => x"90",
           281 => x"b8",
           282 => x"d5",
           283 => x"b8",
           284 => x"90",
           285 => x"b8",
           286 => x"ea",
           287 => x"b8",
           288 => x"90",
           289 => x"b8",
           290 => x"c6",
           291 => x"b8",
           292 => x"90",
           293 => x"b8",
           294 => x"2d",
           295 => x"08",
           296 => x"04",
           297 => x"0c",
           298 => x"81",
           299 => x"83",
           300 => x"81",
           301 => x"b1",
           302 => x"d3",
           303 => x"80",
           304 => x"d3",
           305 => x"e8",
           306 => x"b8",
           307 => x"90",
           308 => x"b8",
           309 => x"2d",
           310 => x"08",
           311 => x"04",
           312 => x"0c",
           313 => x"81",
           314 => x"83",
           315 => x"81",
           316 => x"81",
           317 => x"81",
           318 => x"83",
           319 => x"81",
           320 => x"81",
           321 => x"8e",
           322 => x"70",
           323 => x"0c",
           324 => x"8a",
           325 => x"80",
           326 => x"c1",
           327 => x"81",
           328 => x"02",
           329 => x"0c",
           330 => x"80",
           331 => x"b8",
           332 => x"08",
           333 => x"b8",
           334 => x"08",
           335 => x"3f",
           336 => x"08",
           337 => x"ac",
           338 => x"3d",
           339 => x"b8",
           340 => x"d3",
           341 => x"81",
           342 => x"fd",
           343 => x"53",
           344 => x"08",
           345 => x"52",
           346 => x"08",
           347 => x"51",
           348 => x"d3",
           349 => x"81",
           350 => x"54",
           351 => x"81",
           352 => x"04",
           353 => x"08",
           354 => x"b8",
           355 => x"0d",
           356 => x"d3",
           357 => x"05",
           358 => x"81",
           359 => x"f8",
           360 => x"d3",
           361 => x"05",
           362 => x"b8",
           363 => x"08",
           364 => x"81",
           365 => x"fc",
           366 => x"2e",
           367 => x"0b",
           368 => x"08",
           369 => x"24",
           370 => x"d3",
           371 => x"05",
           372 => x"d3",
           373 => x"05",
           374 => x"b8",
           375 => x"08",
           376 => x"b8",
           377 => x"0c",
           378 => x"81",
           379 => x"fc",
           380 => x"2e",
           381 => x"81",
           382 => x"8c",
           383 => x"d3",
           384 => x"05",
           385 => x"38",
           386 => x"08",
           387 => x"81",
           388 => x"8c",
           389 => x"81",
           390 => x"88",
           391 => x"d3",
           392 => x"05",
           393 => x"b8",
           394 => x"08",
           395 => x"b8",
           396 => x"0c",
           397 => x"08",
           398 => x"81",
           399 => x"b8",
           400 => x"0c",
           401 => x"08",
           402 => x"81",
           403 => x"b8",
           404 => x"0c",
           405 => x"81",
           406 => x"90",
           407 => x"2e",
           408 => x"d3",
           409 => x"05",
           410 => x"d3",
           411 => x"05",
           412 => x"39",
           413 => x"08",
           414 => x"70",
           415 => x"08",
           416 => x"51",
           417 => x"08",
           418 => x"81",
           419 => x"85",
           420 => x"d3",
           421 => x"fc",
           422 => x"79",
           423 => x"05",
           424 => x"57",
           425 => x"83",
           426 => x"38",
           427 => x"51",
           428 => x"a4",
           429 => x"52",
           430 => x"93",
           431 => x"70",
           432 => x"34",
           433 => x"71",
           434 => x"81",
           435 => x"74",
           436 => x"0c",
           437 => x"04",
           438 => x"2b",
           439 => x"71",
           440 => x"51",
           441 => x"72",
           442 => x"72",
           443 => x"05",
           444 => x"71",
           445 => x"53",
           446 => x"70",
           447 => x"0c",
           448 => x"84",
           449 => x"f0",
           450 => x"8f",
           451 => x"83",
           452 => x"38",
           453 => x"84",
           454 => x"fc",
           455 => x"83",
           456 => x"70",
           457 => x"39",
           458 => x"77",
           459 => x"07",
           460 => x"54",
           461 => x"38",
           462 => x"08",
           463 => x"71",
           464 => x"80",
           465 => x"75",
           466 => x"33",
           467 => x"06",
           468 => x"80",
           469 => x"72",
           470 => x"75",
           471 => x"06",
           472 => x"12",
           473 => x"33",
           474 => x"06",
           475 => x"52",
           476 => x"72",
           477 => x"81",
           478 => x"81",
           479 => x"71",
           480 => x"ac",
           481 => x"87",
           482 => x"71",
           483 => x"fb",
           484 => x"06",
           485 => x"82",
           486 => x"51",
           487 => x"97",
           488 => x"84",
           489 => x"54",
           490 => x"75",
           491 => x"38",
           492 => x"52",
           493 => x"80",
           494 => x"ac",
           495 => x"0d",
           496 => x"0d",
           497 => x"52",
           498 => x"52",
           499 => x"81",
           500 => x"81",
           501 => x"07",
           502 => x"52",
           503 => x"e8",
           504 => x"d3",
           505 => x"3d",
           506 => x"3d",
           507 => x"08",
           508 => x"55",
           509 => x"80",
           510 => x"33",
           511 => x"2e",
           512 => x"8c",
           513 => x"70",
           514 => x"70",
           515 => x"38",
           516 => x"39",
           517 => x"80",
           518 => x"53",
           519 => x"83",
           520 => x"70",
           521 => x"2a",
           522 => x"51",
           523 => x"71",
           524 => x"a0",
           525 => x"06",
           526 => x"72",
           527 => x"54",
           528 => x"0c",
           529 => x"81",
           530 => x"86",
           531 => x"fc",
           532 => x"53",
           533 => x"2e",
           534 => x"3d",
           535 => x"72",
           536 => x"3f",
           537 => x"08",
           538 => x"53",
           539 => x"53",
           540 => x"ac",
           541 => x"0d",
           542 => x"0d",
           543 => x"33",
           544 => x"5c",
           545 => x"8b",
           546 => x"38",
           547 => x"ff",
           548 => x"5b",
           549 => x"81",
           550 => x"1c",
           551 => x"5b",
           552 => x"81",
           553 => x"1c",
           554 => x"5b",
           555 => x"81",
           556 => x"1c",
           557 => x"5b",
           558 => x"81",
           559 => x"1c",
           560 => x"5b",
           561 => x"26",
           562 => x"8a",
           563 => x"87",
           564 => x"e7",
           565 => x"38",
           566 => x"59",
           567 => x"58",
           568 => x"57",
           569 => x"56",
           570 => x"55",
           571 => x"54",
           572 => x"53",
           573 => x"81",
           574 => x"94",
           575 => x"c0",
           576 => x"81",
           577 => x"22",
           578 => x"bc",
           579 => x"33",
           580 => x"b8",
           581 => x"33",
           582 => x"b4",
           583 => x"33",
           584 => x"b0",
           585 => x"33",
           586 => x"ac",
           587 => x"33",
           588 => x"a8",
           589 => x"22",
           590 => x"a4",
           591 => x"22",
           592 => x"a0",
           593 => x"0c",
           594 => x"81",
           595 => x"8d",
           596 => x"f5",
           597 => x"5a",
           598 => x"9c",
           599 => x"0c",
           600 => x"bc",
           601 => x"7a",
           602 => x"98",
           603 => x"7a",
           604 => x"87",
           605 => x"08",
           606 => x"1b",
           607 => x"98",
           608 => x"7a",
           609 => x"87",
           610 => x"08",
           611 => x"1b",
           612 => x"98",
           613 => x"7a",
           614 => x"87",
           615 => x"08",
           616 => x"1b",
           617 => x"98",
           618 => x"7a",
           619 => x"80",
           620 => x"1a",
           621 => x"1a",
           622 => x"1a",
           623 => x"1a",
           624 => x"1a",
           625 => x"1a",
           626 => x"1a",
           627 => x"22",
           628 => x"8c",
           629 => x"3f",
           630 => x"04",
           631 => x"02",
           632 => x"70",
           633 => x"2a",
           634 => x"70",
           635 => x"cb",
           636 => x"3d",
           637 => x"3d",
           638 => x"0b",
           639 => x"33",
           640 => x"c0",
           641 => x"72",
           642 => x"38",
           643 => x"94",
           644 => x"70",
           645 => x"81",
           646 => x"52",
           647 => x"8c",
           648 => x"2a",
           649 => x"51",
           650 => x"38",
           651 => x"81",
           652 => x"06",
           653 => x"80",
           654 => x"71",
           655 => x"81",
           656 => x"70",
           657 => x"0b",
           658 => x"a4",
           659 => x"c0",
           660 => x"70",
           661 => x"38",
           662 => x"90",
           663 => x"0c",
           664 => x"ac",
           665 => x"0d",
           666 => x"0d",
           667 => x"33",
           668 => x"cb",
           669 => x"54",
           670 => x"84",
           671 => x"2e",
           672 => x"c0",
           673 => x"70",
           674 => x"2a",
           675 => x"51",
           676 => x"80",
           677 => x"71",
           678 => x"81",
           679 => x"70",
           680 => x"96",
           681 => x"70",
           682 => x"51",
           683 => x"8d",
           684 => x"2a",
           685 => x"51",
           686 => x"bc",
           687 => x"81",
           688 => x"51",
           689 => x"80",
           690 => x"2e",
           691 => x"c0",
           692 => x"73",
           693 => x"3d",
           694 => x"3d",
           695 => x"80",
           696 => x"56",
           697 => x"80",
           698 => x"70",
           699 => x"33",
           700 => x"cb",
           701 => x"55",
           702 => x"84",
           703 => x"2e",
           704 => x"c0",
           705 => x"70",
           706 => x"2a",
           707 => x"51",
           708 => x"80",
           709 => x"71",
           710 => x"81",
           711 => x"70",
           712 => x"96",
           713 => x"70",
           714 => x"51",
           715 => x"8d",
           716 => x"2a",
           717 => x"51",
           718 => x"bc",
           719 => x"81",
           720 => x"51",
           721 => x"80",
           722 => x"2e",
           723 => x"c0",
           724 => x"74",
           725 => x"16",
           726 => x"56",
           727 => x"38",
           728 => x"ac",
           729 => x"0d",
           730 => x"0d",
           731 => x"cb",
           732 => x"87",
           733 => x"51",
           734 => x"86",
           735 => x"94",
           736 => x"08",
           737 => x"70",
           738 => x"51",
           739 => x"2e",
           740 => x"0b",
           741 => x"33",
           742 => x"94",
           743 => x"80",
           744 => x"87",
           745 => x"52",
           746 => x"81",
           747 => x"d3",
           748 => x"83",
           749 => x"ff",
           750 => x"0b",
           751 => x"33",
           752 => x"94",
           753 => x"80",
           754 => x"87",
           755 => x"52",
           756 => x"82",
           757 => x"06",
           758 => x"ff",
           759 => x"2e",
           760 => x"0b",
           761 => x"33",
           762 => x"94",
           763 => x"80",
           764 => x"87",
           765 => x"52",
           766 => x"98",
           767 => x"2c",
           768 => x"71",
           769 => x"0c",
           770 => x"04",
           771 => x"87",
           772 => x"70",
           773 => x"2a",
           774 => x"52",
           775 => x"2e",
           776 => x"81",
           777 => x"87",
           778 => x"08",
           779 => x"11",
           780 => x"a0",
           781 => x"52",
           782 => x"c0",
           783 => x"71",
           784 => x"11",
           785 => x"90",
           786 => x"52",
           787 => x"c0",
           788 => x"71",
           789 => x"11",
           790 => x"98",
           791 => x"52",
           792 => x"c0",
           793 => x"71",
           794 => x"11",
           795 => x"a8",
           796 => x"52",
           797 => x"c0",
           798 => x"71",
           799 => x"08",
           800 => x"a4",
           801 => x"12",
           802 => x"84",
           803 => x"51",
           804 => x"13",
           805 => x"52",
           806 => x"c0",
           807 => x"70",
           808 => x"51",
           809 => x"80",
           810 => x"81",
           811 => x"34",
           812 => x"c0",
           813 => x"70",
           814 => x"06",
           815 => x"70",
           816 => x"38",
           817 => x"81",
           818 => x"80",
           819 => x"9e",
           820 => x"80",
           821 => x"51",
           822 => x"80",
           823 => x"81",
           824 => x"cb",
           825 => x"0b",
           826 => x"88",
           827 => x"80",
           828 => x"52",
           829 => x"83",
           830 => x"71",
           831 => x"34",
           832 => x"c0",
           833 => x"70",
           834 => x"51",
           835 => x"80",
           836 => x"81",
           837 => x"cb",
           838 => x"0b",
           839 => x"88",
           840 => x"80",
           841 => x"52",
           842 => x"83",
           843 => x"71",
           844 => x"34",
           845 => x"c0",
           846 => x"70",
           847 => x"51",
           848 => x"80",
           849 => x"81",
           850 => x"cb",
           851 => x"0b",
           852 => x"88",
           853 => x"80",
           854 => x"52",
           855 => x"83",
           856 => x"71",
           857 => x"34",
           858 => x"52",
           859 => x"88",
           860 => x"80",
           861 => x"86",
           862 => x"52",
           863 => x"70",
           864 => x"34",
           865 => x"73",
           866 => x"06",
           867 => x"70",
           868 => x"38",
           869 => x"74",
           870 => x"87",
           871 => x"08",
           872 => x"51",
           873 => x"80",
           874 => x"81",
           875 => x"cb",
           876 => x"c0",
           877 => x"70",
           878 => x"51",
           879 => x"e0",
           880 => x"0d",
           881 => x"0d",
           882 => x"51",
           883 => x"81",
           884 => x"54",
           885 => x"88",
           886 => x"b8",
           887 => x"3f",
           888 => x"51",
           889 => x"81",
           890 => x"33",
           891 => x"80",
           892 => x"d7",
           893 => x"81",
           894 => x"52",
           895 => x"51",
           896 => x"81",
           897 => x"33",
           898 => x"80",
           899 => x"de",
           900 => x"da",
           901 => x"81",
           902 => x"89",
           903 => x"cb",
           904 => x"55",
           905 => x"38",
           906 => x"54",
           907 => x"93",
           908 => x"bc",
           909 => x"fc",
           910 => x"54",
           911 => x"51",
           912 => x"81",
           913 => x"54",
           914 => x"88",
           915 => x"d4",
           916 => x"3f",
           917 => x"33",
           918 => x"2e",
           919 => x"b7",
           920 => x"a8",
           921 => x"db",
           922 => x"80",
           923 => x"81",
           924 => x"83",
           925 => x"cb",
           926 => x"55",
           927 => x"2e",
           928 => x"15",
           929 => x"b7",
           930 => x"fa",
           931 => x"de",
           932 => x"80",
           933 => x"81",
           934 => x"82",
           935 => x"cb",
           936 => x"55",
           937 => x"2e",
           938 => x"15",
           939 => x"b8",
           940 => x"d2",
           941 => x"d0",
           942 => x"3f",
           943 => x"70",
           944 => x"05",
           945 => x"81",
           946 => x"55",
           947 => x"3f",
           948 => x"81",
           949 => x"88",
           950 => x"15",
           951 => x"b9",
           952 => x"a2",
           953 => x"22",
           954 => x"d4",
           955 => x"3f",
           956 => x"52",
           957 => x"51",
           958 => x"86",
           959 => x"ff",
           960 => x"8e",
           961 => x"71",
           962 => x"38",
           963 => x"0b",
           964 => x"a8",
           965 => x"08",
           966 => x"a4",
           967 => x"3f",
           968 => x"ba",
           969 => x"b2",
           970 => x"81",
           971 => x"f7",
           972 => x"39",
           973 => x"51",
           974 => x"91",
           975 => x"c0",
           976 => x"3f",
           977 => x"ba",
           978 => x"8e",
           979 => x"0d",
           980 => x"80",
           981 => x"0b",
           982 => x"84",
           983 => x"3d",
           984 => x"96",
           985 => x"52",
           986 => x"0c",
           987 => x"70",
           988 => x"0c",
           989 => x"3d",
           990 => x"3d",
           991 => x"96",
           992 => x"81",
           993 => x"52",
           994 => x"73",
           995 => x"cb",
           996 => x"70",
           997 => x"0c",
           998 => x"83",
           999 => x"81",
          1000 => x"87",
          1001 => x"0c",
          1002 => x"0d",
          1003 => x"33",
          1004 => x"2e",
          1005 => x"85",
          1006 => x"ed",
          1007 => x"c4",
          1008 => x"95",
          1009 => x"c4",
          1010 => x"72",
          1011 => x"c4",
          1012 => x"81",
          1013 => x"92",
          1014 => x"bc",
          1015 => x"8a",
          1016 => x"81",
          1017 => x"52",
          1018 => x"3d",
          1019 => x"3d",
          1020 => x"05",
          1021 => x"bc",
          1022 => x"d3",
          1023 => x"51",
          1024 => x"72",
          1025 => x"0c",
          1026 => x"04",
          1027 => x"74",
          1028 => x"53",
          1029 => x"91",
          1030 => x"81",
          1031 => x"51",
          1032 => x"72",
          1033 => x"f1",
          1034 => x"0d",
          1035 => x"0d",
          1036 => x"bc",
          1037 => x"d3",
          1038 => x"33",
          1039 => x"71",
          1040 => x"38",
          1041 => x"05",
          1042 => x"fe",
          1043 => x"33",
          1044 => x"38",
          1045 => x"bc",
          1046 => x"0d",
          1047 => x"0d",
          1048 => x"59",
          1049 => x"05",
          1050 => x"75",
          1051 => x"92",
          1052 => x"2e",
          1053 => x"51",
          1054 => x"e8",
          1055 => x"7a",
          1056 => x"5c",
          1057 => x"5a",
          1058 => x"09",
          1059 => x"38",
          1060 => x"81",
          1061 => x"57",
          1062 => x"75",
          1063 => x"81",
          1064 => x"82",
          1065 => x"05",
          1066 => x"5d",
          1067 => x"09",
          1068 => x"38",
          1069 => x"71",
          1070 => x"81",
          1071 => x"59",
          1072 => x"9f",
          1073 => x"53",
          1074 => x"97",
          1075 => x"29",
          1076 => x"79",
          1077 => x"5b",
          1078 => x"55",
          1079 => x"73",
          1080 => x"75",
          1081 => x"70",
          1082 => x"07",
          1083 => x"80",
          1084 => x"30",
          1085 => x"80",
          1086 => x"53",
          1087 => x"54",
          1088 => x"2e",
          1089 => x"84",
          1090 => x"81",
          1091 => x"57",
          1092 => x"2e",
          1093 => x"75",
          1094 => x"76",
          1095 => x"e0",
          1096 => x"ff",
          1097 => x"ff",
          1098 => x"72",
          1099 => x"98",
          1100 => x"10",
          1101 => x"05",
          1102 => x"04",
          1103 => x"71",
          1104 => x"53",
          1105 => x"54",
          1106 => x"2e",
          1107 => x"14",
          1108 => x"33",
          1109 => x"72",
          1110 => x"81",
          1111 => x"06",
          1112 => x"a3",
          1113 => x"15",
          1114 => x"7a",
          1115 => x"7c",
          1116 => x"06",
          1117 => x"fc",
          1118 => x"8b",
          1119 => x"15",
          1120 => x"73",
          1121 => x"74",
          1122 => x"3f",
          1123 => x"55",
          1124 => x"27",
          1125 => x"a0",
          1126 => x"3f",
          1127 => x"55",
          1128 => x"26",
          1129 => x"bc",
          1130 => x"1d",
          1131 => x"53",
          1132 => x"f5",
          1133 => x"39",
          1134 => x"39",
          1135 => x"39",
          1136 => x"39",
          1137 => x"39",
          1138 => x"dd",
          1139 => x"39",
          1140 => x"70",
          1141 => x"53",
          1142 => x"8b",
          1143 => x"1d",
          1144 => x"5d",
          1145 => x"74",
          1146 => x"09",
          1147 => x"38",
          1148 => x"71",
          1149 => x"53",
          1150 => x"84",
          1151 => x"59",
          1152 => x"80",
          1153 => x"30",
          1154 => x"80",
          1155 => x"7b",
          1156 => x"52",
          1157 => x"80",
          1158 => x"76",
          1159 => x"07",
          1160 => x"58",
          1161 => x"51",
          1162 => x"81",
          1163 => x"81",
          1164 => x"53",
          1165 => x"e5",
          1166 => x"d3",
          1167 => x"89",
          1168 => x"38",
          1169 => x"70",
          1170 => x"57",
          1171 => x"80",
          1172 => x"38",
          1173 => x"81",
          1174 => x"53",
          1175 => x"05",
          1176 => x"16",
          1177 => x"74",
          1178 => x"77",
          1179 => x"07",
          1180 => x"9f",
          1181 => x"51",
          1182 => x"72",
          1183 => x"7c",
          1184 => x"81",
          1185 => x"72",
          1186 => x"38",
          1187 => x"05",
          1188 => x"ad",
          1189 => x"18",
          1190 => x"81",
          1191 => x"b0",
          1192 => x"38",
          1193 => x"81",
          1194 => x"06",
          1195 => x"a3",
          1196 => x"15",
          1197 => x"7a",
          1198 => x"7c",
          1199 => x"06",
          1200 => x"f9",
          1201 => x"8b",
          1202 => x"15",
          1203 => x"73",
          1204 => x"ff",
          1205 => x"e0",
          1206 => x"33",
          1207 => x"f9",
          1208 => x"ef",
          1209 => x"15",
          1210 => x"7a",
          1211 => x"38",
          1212 => x"b5",
          1213 => x"15",
          1214 => x"73",
          1215 => x"fa",
          1216 => x"3d",
          1217 => x"3d",
          1218 => x"70",
          1219 => x"52",
          1220 => x"73",
          1221 => x"3f",
          1222 => x"04",
          1223 => x"74",
          1224 => x"0c",
          1225 => x"05",
          1226 => x"fa",
          1227 => x"d3",
          1228 => x"80",
          1229 => x"0b",
          1230 => x"0c",
          1231 => x"04",
          1232 => x"81",
          1233 => x"76",
          1234 => x"0c",
          1235 => x"05",
          1236 => x"53",
          1237 => x"72",
          1238 => x"0c",
          1239 => x"04",
          1240 => x"78",
          1241 => x"80",
          1242 => x"c0",
          1243 => x"80",
          1244 => x"39",
          1245 => x"f3",
          1246 => x"81",
          1247 => x"52",
          1248 => x"d3",
          1249 => x"ff",
          1250 => x"80",
          1251 => x"73",
          1252 => x"ca",
          1253 => x"32",
          1254 => x"30",
          1255 => x"9f",
          1256 => x"25",
          1257 => x"51",
          1258 => x"2e",
          1259 => x"15",
          1260 => x"06",
          1261 => x"f1",
          1262 => x"9f",
          1263 => x"bb",
          1264 => x"52",
          1265 => x"ff",
          1266 => x"15",
          1267 => x"34",
          1268 => x"81",
          1269 => x"55",
          1270 => x"ff",
          1271 => x"17",
          1272 => x"34",
          1273 => x"c1",
          1274 => x"72",
          1275 => x"0c",
          1276 => x"04",
          1277 => x"81",
          1278 => x"75",
          1279 => x"0c",
          1280 => x"52",
          1281 => x"3f",
          1282 => x"c0",
          1283 => x"0d",
          1284 => x"0d",
          1285 => x"55",
          1286 => x"0c",
          1287 => x"33",
          1288 => x"73",
          1289 => x"81",
          1290 => x"74",
          1291 => x"75",
          1292 => x"70",
          1293 => x"73",
          1294 => x"38",
          1295 => x"09",
          1296 => x"38",
          1297 => x"11",
          1298 => x"08",
          1299 => x"54",
          1300 => x"2e",
          1301 => x"80",
          1302 => x"08",
          1303 => x"0c",
          1304 => x"33",
          1305 => x"80",
          1306 => x"38",
          1307 => x"2e",
          1308 => x"a1",
          1309 => x"81",
          1310 => x"75",
          1311 => x"56",
          1312 => x"c1",
          1313 => x"08",
          1314 => x"0c",
          1315 => x"33",
          1316 => x"b1",
          1317 => x"a0",
          1318 => x"82",
          1319 => x"53",
          1320 => x"57",
          1321 => x"9d",
          1322 => x"39",
          1323 => x"80",
          1324 => x"26",
          1325 => x"8b",
          1326 => x"80",
          1327 => x"56",
          1328 => x"8a",
          1329 => x"a0",
          1330 => x"c5",
          1331 => x"74",
          1332 => x"e0",
          1333 => x"ff",
          1334 => x"d0",
          1335 => x"ff",
          1336 => x"90",
          1337 => x"38",
          1338 => x"81",
          1339 => x"53",
          1340 => x"c5",
          1341 => x"27",
          1342 => x"76",
          1343 => x"08",
          1344 => x"0c",
          1345 => x"33",
          1346 => x"73",
          1347 => x"bd",
          1348 => x"2e",
          1349 => x"30",
          1350 => x"0c",
          1351 => x"81",
          1352 => x"8a",
          1353 => x"f8",
          1354 => x"7c",
          1355 => x"70",
          1356 => x"08",
          1357 => x"54",
          1358 => x"2e",
          1359 => x"92",
          1360 => x"81",
          1361 => x"74",
          1362 => x"55",
          1363 => x"2e",
          1364 => x"ad",
          1365 => x"06",
          1366 => x"75",
          1367 => x"0c",
          1368 => x"33",
          1369 => x"73",
          1370 => x"81",
          1371 => x"38",
          1372 => x"05",
          1373 => x"08",
          1374 => x"53",
          1375 => x"2e",
          1376 => x"80",
          1377 => x"81",
          1378 => x"90",
          1379 => x"76",
          1380 => x"70",
          1381 => x"57",
          1382 => x"82",
          1383 => x"05",
          1384 => x"08",
          1385 => x"54",
          1386 => x"81",
          1387 => x"27",
          1388 => x"d0",
          1389 => x"56",
          1390 => x"73",
          1391 => x"80",
          1392 => x"14",
          1393 => x"72",
          1394 => x"e8",
          1395 => x"80",
          1396 => x"39",
          1397 => x"dc",
          1398 => x"80",
          1399 => x"27",
          1400 => x"80",
          1401 => x"89",
          1402 => x"70",
          1403 => x"55",
          1404 => x"70",
          1405 => x"55",
          1406 => x"27",
          1407 => x"14",
          1408 => x"06",
          1409 => x"74",
          1410 => x"73",
          1411 => x"38",
          1412 => x"14",
          1413 => x"05",
          1414 => x"08",
          1415 => x"54",
          1416 => x"26",
          1417 => x"77",
          1418 => x"38",
          1419 => x"75",
          1420 => x"56",
          1421 => x"ac",
          1422 => x"0d",
          1423 => x"0d",
          1424 => x"33",
          1425 => x"70",
          1426 => x"38",
          1427 => x"11",
          1428 => x"81",
          1429 => x"83",
          1430 => x"fd",
          1431 => x"97",
          1432 => x"84",
          1433 => x"33",
          1434 => x"51",
          1435 => x"80",
          1436 => x"90",
          1437 => x"92",
          1438 => x"88",
          1439 => x"2e",
          1440 => x"88",
          1441 => x"0c",
          1442 => x"87",
          1443 => x"05",
          1444 => x"0c",
          1445 => x"c0",
          1446 => x"70",
          1447 => x"98",
          1448 => x"08",
          1449 => x"51",
          1450 => x"2e",
          1451 => x"08",
          1452 => x"38",
          1453 => x"87",
          1454 => x"05",
          1455 => x"80",
          1456 => x"51",
          1457 => x"87",
          1458 => x"08",
          1459 => x"2e",
          1460 => x"81",
          1461 => x"34",
          1462 => x"13",
          1463 => x"81",
          1464 => x"85",
          1465 => x"f2",
          1466 => x"63",
          1467 => x"05",
          1468 => x"33",
          1469 => x"58",
          1470 => x"5b",
          1471 => x"81",
          1472 => x"81",
          1473 => x"52",
          1474 => x"38",
          1475 => x"5d",
          1476 => x"8c",
          1477 => x"87",
          1478 => x"11",
          1479 => x"84",
          1480 => x"5c",
          1481 => x"85",
          1482 => x"c0",
          1483 => x"7c",
          1484 => x"84",
          1485 => x"08",
          1486 => x"70",
          1487 => x"53",
          1488 => x"2e",
          1489 => x"08",
          1490 => x"70",
          1491 => x"34",
          1492 => x"73",
          1493 => x"71",
          1494 => x"38",
          1495 => x"71",
          1496 => x"08",
          1497 => x"2e",
          1498 => x"84",
          1499 => x"38",
          1500 => x"87",
          1501 => x"1e",
          1502 => x"70",
          1503 => x"52",
          1504 => x"ff",
          1505 => x"39",
          1506 => x"81",
          1507 => x"ff",
          1508 => x"5c",
          1509 => x"90",
          1510 => x"80",
          1511 => x"71",
          1512 => x"7d",
          1513 => x"38",
          1514 => x"80",
          1515 => x"80",
          1516 => x"81",
          1517 => x"73",
          1518 => x"0c",
          1519 => x"04",
          1520 => x"60",
          1521 => x"8c",
          1522 => x"33",
          1523 => x"57",
          1524 => x"5a",
          1525 => x"81",
          1526 => x"81",
          1527 => x"52",
          1528 => x"38",
          1529 => x"c0",
          1530 => x"84",
          1531 => x"92",
          1532 => x"c0",
          1533 => x"72",
          1534 => x"5a",
          1535 => x"0c",
          1536 => x"80",
          1537 => x"0c",
          1538 => x"0c",
          1539 => x"08",
          1540 => x"70",
          1541 => x"53",
          1542 => x"2e",
          1543 => x"70",
          1544 => x"33",
          1545 => x"13",
          1546 => x"2a",
          1547 => x"51",
          1548 => x"2e",
          1549 => x"08",
          1550 => x"38",
          1551 => x"71",
          1552 => x"38",
          1553 => x"2e",
          1554 => x"75",
          1555 => x"92",
          1556 => x"72",
          1557 => x"06",
          1558 => x"f7",
          1559 => x"5a",
          1560 => x"1c",
          1561 => x"06",
          1562 => x"5d",
          1563 => x"80",
          1564 => x"73",
          1565 => x"06",
          1566 => x"38",
          1567 => x"fe",
          1568 => x"fc",
          1569 => x"52",
          1570 => x"83",
          1571 => x"71",
          1572 => x"d3",
          1573 => x"3d",
          1574 => x"3d",
          1575 => x"84",
          1576 => x"33",
          1577 => x"b3",
          1578 => x"54",
          1579 => x"fb",
          1580 => x"d3",
          1581 => x"06",
          1582 => x"71",
          1583 => x"54",
          1584 => x"a2",
          1585 => x"24",
          1586 => x"80",
          1587 => x"a7",
          1588 => x"2e",
          1589 => x"39",
          1590 => x"87",
          1591 => x"05",
          1592 => x"52",
          1593 => x"80",
          1594 => x"80",
          1595 => x"81",
          1596 => x"80",
          1597 => x"84",
          1598 => x"d3",
          1599 => x"3d",
          1600 => x"3d",
          1601 => x"33",
          1602 => x"70",
          1603 => x"07",
          1604 => x"0c",
          1605 => x"83",
          1606 => x"fd",
          1607 => x"83",
          1608 => x"12",
          1609 => x"2b",
          1610 => x"07",
          1611 => x"71",
          1612 => x"71",
          1613 => x"81",
          1614 => x"51",
          1615 => x"52",
          1616 => x"04",
          1617 => x"73",
          1618 => x"92",
          1619 => x"52",
          1620 => x"81",
          1621 => x"70",
          1622 => x"70",
          1623 => x"3d",
          1624 => x"3d",
          1625 => x"52",
          1626 => x"70",
          1627 => x"34",
          1628 => x"51",
          1629 => x"81",
          1630 => x"70",
          1631 => x"70",
          1632 => x"05",
          1633 => x"88",
          1634 => x"72",
          1635 => x"0d",
          1636 => x"0d",
          1637 => x"54",
          1638 => x"80",
          1639 => x"71",
          1640 => x"53",
          1641 => x"81",
          1642 => x"ff",
          1643 => x"ef",
          1644 => x"0d",
          1645 => x"0d",
          1646 => x"54",
          1647 => x"72",
          1648 => x"54",
          1649 => x"51",
          1650 => x"84",
          1651 => x"fc",
          1652 => x"77",
          1653 => x"53",
          1654 => x"05",
          1655 => x"70",
          1656 => x"33",
          1657 => x"ff",
          1658 => x"52",
          1659 => x"2e",
          1660 => x"80",
          1661 => x"71",
          1662 => x"0c",
          1663 => x"04",
          1664 => x"74",
          1665 => x"53",
          1666 => x"80",
          1667 => x"70",
          1668 => x"38",
          1669 => x"33",
          1670 => x"80",
          1671 => x"70",
          1672 => x"81",
          1673 => x"71",
          1674 => x"ac",
          1675 => x"0d",
          1676 => x"81",
          1677 => x"04",
          1678 => x"d3",
          1679 => x"f9",
          1680 => x"56",
          1681 => x"17",
          1682 => x"74",
          1683 => x"d7",
          1684 => x"b0",
          1685 => x"b4",
          1686 => x"81",
          1687 => x"57",
          1688 => x"81",
          1689 => x"78",
          1690 => x"06",
          1691 => x"d3",
          1692 => x"17",
          1693 => x"08",
          1694 => x"31",
          1695 => x"17",
          1696 => x"38",
          1697 => x"55",
          1698 => x"09",
          1699 => x"38",
          1700 => x"16",
          1701 => x"08",
          1702 => x"52",
          1703 => x"51",
          1704 => x"83",
          1705 => x"77",
          1706 => x"0c",
          1707 => x"04",
          1708 => x"78",
          1709 => x"80",
          1710 => x"08",
          1711 => x"38",
          1712 => x"fb",
          1713 => x"ac",
          1714 => x"d3",
          1715 => x"38",
          1716 => x"53",
          1717 => x"81",
          1718 => x"f8",
          1719 => x"d3",
          1720 => x"2e",
          1721 => x"55",
          1722 => x"b0",
          1723 => x"81",
          1724 => x"88",
          1725 => x"f8",
          1726 => x"70",
          1727 => x"bf",
          1728 => x"ac",
          1729 => x"d3",
          1730 => x"91",
          1731 => x"55",
          1732 => x"09",
          1733 => x"f0",
          1734 => x"33",
          1735 => x"2e",
          1736 => x"80",
          1737 => x"80",
          1738 => x"ac",
          1739 => x"17",
          1740 => x"fd",
          1741 => x"d4",
          1742 => x"b2",
          1743 => x"84",
          1744 => x"85",
          1745 => x"75",
          1746 => x"3f",
          1747 => x"e4",
          1748 => x"98",
          1749 => x"8a",
          1750 => x"08",
          1751 => x"17",
          1752 => x"3f",
          1753 => x"52",
          1754 => x"51",
          1755 => x"a0",
          1756 => x"05",
          1757 => x"0c",
          1758 => x"75",
          1759 => x"33",
          1760 => x"3f",
          1761 => x"34",
          1762 => x"52",
          1763 => x"51",
          1764 => x"81",
          1765 => x"80",
          1766 => x"81",
          1767 => x"d3",
          1768 => x"3d",
          1769 => x"3d",
          1770 => x"1a",
          1771 => x"fe",
          1772 => x"54",
          1773 => x"73",
          1774 => x"8a",
          1775 => x"76",
          1776 => x"08",
          1777 => x"75",
          1778 => x"0c",
          1779 => x"04",
          1780 => x"7a",
          1781 => x"56",
          1782 => x"75",
          1783 => x"98",
          1784 => x"26",
          1785 => x"56",
          1786 => x"ff",
          1787 => x"56",
          1788 => x"80",
          1789 => x"82",
          1790 => x"72",
          1791 => x"38",
          1792 => x"72",
          1793 => x"8e",
          1794 => x"39",
          1795 => x"15",
          1796 => x"a4",
          1797 => x"53",
          1798 => x"fd",
          1799 => x"d3",
          1800 => x"9f",
          1801 => x"ff",
          1802 => x"11",
          1803 => x"70",
          1804 => x"18",
          1805 => x"76",
          1806 => x"53",
          1807 => x"81",
          1808 => x"80",
          1809 => x"83",
          1810 => x"b4",
          1811 => x"88",
          1812 => x"77",
          1813 => x"84",
          1814 => x"5a",
          1815 => x"80",
          1816 => x"9f",
          1817 => x"80",
          1818 => x"88",
          1819 => x"08",
          1820 => x"51",
          1821 => x"81",
          1822 => x"80",
          1823 => x"15",
          1824 => x"74",
          1825 => x"51",
          1826 => x"81",
          1827 => x"83",
          1828 => x"56",
          1829 => x"87",
          1830 => x"08",
          1831 => x"51",
          1832 => x"81",
          1833 => x"9b",
          1834 => x"2b",
          1835 => x"74",
          1836 => x"51",
          1837 => x"81",
          1838 => x"f0",
          1839 => x"83",
          1840 => x"75",
          1841 => x"0c",
          1842 => x"04",
          1843 => x"7b",
          1844 => x"55",
          1845 => x"81",
          1846 => x"af",
          1847 => x"16",
          1848 => x"a7",
          1849 => x"53",
          1850 => x"81",
          1851 => x"77",
          1852 => x"72",
          1853 => x"38",
          1854 => x"72",
          1855 => x"c9",
          1856 => x"39",
          1857 => x"14",
          1858 => x"a4",
          1859 => x"53",
          1860 => x"fb",
          1861 => x"d3",
          1862 => x"81",
          1863 => x"81",
          1864 => x"83",
          1865 => x"b4",
          1866 => x"76",
          1867 => x"5b",
          1868 => x"57",
          1869 => x"8f",
          1870 => x"2b",
          1871 => x"78",
          1872 => x"71",
          1873 => x"76",
          1874 => x"0b",
          1875 => x"78",
          1876 => x"16",
          1877 => x"74",
          1878 => x"3f",
          1879 => x"08",
          1880 => x"ac",
          1881 => x"38",
          1882 => x"06",
          1883 => x"75",
          1884 => x"84",
          1885 => x"51",
          1886 => x"38",
          1887 => x"78",
          1888 => x"06",
          1889 => x"06",
          1890 => x"78",
          1891 => x"83",
          1892 => x"f7",
          1893 => x"2a",
          1894 => x"05",
          1895 => x"fa",
          1896 => x"d3",
          1897 => x"81",
          1898 => x"80",
          1899 => x"83",
          1900 => x"52",
          1901 => x"ff",
          1902 => x"b4",
          1903 => x"84",
          1904 => x"83",
          1905 => x"c3",
          1906 => x"2a",
          1907 => x"05",
          1908 => x"f9",
          1909 => x"d3",
          1910 => x"81",
          1911 => x"ab",
          1912 => x"0a",
          1913 => x"2b",
          1914 => x"76",
          1915 => x"70",
          1916 => x"56",
          1917 => x"81",
          1918 => x"8f",
          1919 => x"07",
          1920 => x"f6",
          1921 => x"0b",
          1922 => x"76",
          1923 => x"0c",
          1924 => x"04",
          1925 => x"79",
          1926 => x"08",
          1927 => x"57",
          1928 => x"88",
          1929 => x"08",
          1930 => x"38",
          1931 => x"8e",
          1932 => x"2e",
          1933 => x"53",
          1934 => x"51",
          1935 => x"81",
          1936 => x"56",
          1937 => x"08",
          1938 => x"93",
          1939 => x"80",
          1940 => x"56",
          1941 => x"81",
          1942 => x"56",
          1943 => x"73",
          1944 => x"fa",
          1945 => x"d3",
          1946 => x"81",
          1947 => x"80",
          1948 => x"38",
          1949 => x"08",
          1950 => x"38",
          1951 => x"08",
          1952 => x"38",
          1953 => x"52",
          1954 => x"c0",
          1955 => x"ac",
          1956 => x"98",
          1957 => x"05",
          1958 => x"08",
          1959 => x"38",
          1960 => x"81",
          1961 => x"0c",
          1962 => x"81",
          1963 => x"84",
          1964 => x"54",
          1965 => x"76",
          1966 => x"38",
          1967 => x"81",
          1968 => x"89",
          1969 => x"f5",
          1970 => x"7f",
          1971 => x"5c",
          1972 => x"38",
          1973 => x"58",
          1974 => x"88",
          1975 => x"08",
          1976 => x"38",
          1977 => x"39",
          1978 => x"51",
          1979 => x"81",
          1980 => x"d3",
          1981 => x"82",
          1982 => x"d3",
          1983 => x"81",
          1984 => x"ff",
          1985 => x"38",
          1986 => x"08",
          1987 => x"08",
          1988 => x"08",
          1989 => x"38",
          1990 => x"55",
          1991 => x"75",
          1992 => x"38",
          1993 => x"7b",
          1994 => x"06",
          1995 => x"81",
          1996 => x"19",
          1997 => x"83",
          1998 => x"76",
          1999 => x"f9",
          2000 => x"d3",
          2001 => x"80",
          2002 => x"ac",
          2003 => x"09",
          2004 => x"38",
          2005 => x"08",
          2006 => x"32",
          2007 => x"72",
          2008 => x"70",
          2009 => x"53",
          2010 => x"54",
          2011 => x"38",
          2012 => x"95",
          2013 => x"08",
          2014 => x"27",
          2015 => x"98",
          2016 => x"83",
          2017 => x"80",
          2018 => x"de",
          2019 => x"81",
          2020 => x"19",
          2021 => x"89",
          2022 => x"76",
          2023 => x"b6",
          2024 => x"7b",
          2025 => x"3f",
          2026 => x"08",
          2027 => x"ac",
          2028 => x"b6",
          2029 => x"81",
          2030 => x"81",
          2031 => x"06",
          2032 => x"d3",
          2033 => x"75",
          2034 => x"30",
          2035 => x"80",
          2036 => x"07",
          2037 => x"54",
          2038 => x"38",
          2039 => x"09",
          2040 => x"ab",
          2041 => x"80",
          2042 => x"53",
          2043 => x"51",
          2044 => x"81",
          2045 => x"81",
          2046 => x"30",
          2047 => x"ac",
          2048 => x"25",
          2049 => x"7f",
          2050 => x"72",
          2051 => x"51",
          2052 => x"80",
          2053 => x"76",
          2054 => x"78",
          2055 => x"3f",
          2056 => x"08",
          2057 => x"38",
          2058 => x"0c",
          2059 => x"fe",
          2060 => x"19",
          2061 => x"89",
          2062 => x"08",
          2063 => x"1a",
          2064 => x"33",
          2065 => x"73",
          2066 => x"94",
          2067 => x"75",
          2068 => x"38",
          2069 => x"55",
          2070 => x"55",
          2071 => x"57",
          2072 => x"81",
          2073 => x"8d",
          2074 => x"f7",
          2075 => x"70",
          2076 => x"cb",
          2077 => x"81",
          2078 => x"80",
          2079 => x"52",
          2080 => x"a2",
          2081 => x"ac",
          2082 => x"ac",
          2083 => x"0c",
          2084 => x"53",
          2085 => x"17",
          2086 => x"f2",
          2087 => x"59",
          2088 => x"56",
          2089 => x"16",
          2090 => x"22",
          2091 => x"27",
          2092 => x"54",
          2093 => x"78",
          2094 => x"33",
          2095 => x"3f",
          2096 => x"08",
          2097 => x"38",
          2098 => x"18",
          2099 => x"74",
          2100 => x"38",
          2101 => x"55",
          2102 => x"ac",
          2103 => x"0d",
          2104 => x"0d",
          2105 => x"08",
          2106 => x"74",
          2107 => x"26",
          2108 => x"9f",
          2109 => x"80",
          2110 => x"82",
          2111 => x"39",
          2112 => x"0c",
          2113 => x"54",
          2114 => x"75",
          2115 => x"73",
          2116 => x"a8",
          2117 => x"73",
          2118 => x"85",
          2119 => x"0b",
          2120 => x"5a",
          2121 => x"27",
          2122 => x"a8",
          2123 => x"18",
          2124 => x"39",
          2125 => x"70",
          2126 => x"58",
          2127 => x"b6",
          2128 => x"76",
          2129 => x"3f",
          2130 => x"08",
          2131 => x"ac",
          2132 => x"bf",
          2133 => x"81",
          2134 => x"27",
          2135 => x"16",
          2136 => x"ac",
          2137 => x"38",
          2138 => x"c1",
          2139 => x"31",
          2140 => x"27",
          2141 => x"52",
          2142 => x"aa",
          2143 => x"ac",
          2144 => x"0c",
          2145 => x"0c",
          2146 => x"17",
          2147 => x"9d",
          2148 => x"81",
          2149 => x"74",
          2150 => x"18",
          2151 => x"18",
          2152 => x"ff",
          2153 => x"05",
          2154 => x"80",
          2155 => x"d3",
          2156 => x"3d",
          2157 => x"3d",
          2158 => x"71",
          2159 => x"08",
          2160 => x"59",
          2161 => x"80",
          2162 => x"86",
          2163 => x"98",
          2164 => x"53",
          2165 => x"80",
          2166 => x"38",
          2167 => x"06",
          2168 => x"c1",
          2169 => x"08",
          2170 => x"16",
          2171 => x"08",
          2172 => x"85",
          2173 => x"22",
          2174 => x"73",
          2175 => x"38",
          2176 => x"0c",
          2177 => x"ad",
          2178 => x"22",
          2179 => x"89",
          2180 => x"53",
          2181 => x"38",
          2182 => x"52",
          2183 => x"b0",
          2184 => x"ac",
          2185 => x"53",
          2186 => x"d3",
          2187 => x"81",
          2188 => x"53",
          2189 => x"08",
          2190 => x"f9",
          2191 => x"08",
          2192 => x"08",
          2193 => x"38",
          2194 => x"77",
          2195 => x"84",
          2196 => x"39",
          2197 => x"52",
          2198 => x"eb",
          2199 => x"ac",
          2200 => x"53",
          2201 => x"08",
          2202 => x"c9",
          2203 => x"81",
          2204 => x"81",
          2205 => x"81",
          2206 => x"ac",
          2207 => x"b5",
          2208 => x"ac",
          2209 => x"51",
          2210 => x"81",
          2211 => x"ac",
          2212 => x"73",
          2213 => x"73",
          2214 => x"f2",
          2215 => x"d3",
          2216 => x"16",
          2217 => x"16",
          2218 => x"ff",
          2219 => x"05",
          2220 => x"80",
          2221 => x"d3",
          2222 => x"3d",
          2223 => x"3d",
          2224 => x"71",
          2225 => x"56",
          2226 => x"51",
          2227 => x"81",
          2228 => x"54",
          2229 => x"08",
          2230 => x"81",
          2231 => x"57",
          2232 => x"52",
          2233 => x"c8",
          2234 => x"ac",
          2235 => x"d3",
          2236 => x"c7",
          2237 => x"ac",
          2238 => x"08",
          2239 => x"54",
          2240 => x"e5",
          2241 => x"06",
          2242 => x"55",
          2243 => x"80",
          2244 => x"51",
          2245 => x"2e",
          2246 => x"17",
          2247 => x"2e",
          2248 => x"39",
          2249 => x"52",
          2250 => x"8a",
          2251 => x"ac",
          2252 => x"d3",
          2253 => x"2e",
          2254 => x"73",
          2255 => x"81",
          2256 => x"87",
          2257 => x"d3",
          2258 => x"3d",
          2259 => x"3d",
          2260 => x"11",
          2261 => x"aa",
          2262 => x"ac",
          2263 => x"ff",
          2264 => x"33",
          2265 => x"71",
          2266 => x"81",
          2267 => x"94",
          2268 => x"8e",
          2269 => x"ac",
          2270 => x"73",
          2271 => x"81",
          2272 => x"85",
          2273 => x"fc",
          2274 => x"79",
          2275 => x"ff",
          2276 => x"12",
          2277 => x"eb",
          2278 => x"70",
          2279 => x"72",
          2280 => x"81",
          2281 => x"73",
          2282 => x"94",
          2283 => x"94",
          2284 => x"0d",
          2285 => x"0d",
          2286 => x"56",
          2287 => x"5a",
          2288 => x"08",
          2289 => x"86",
          2290 => x"08",
          2291 => x"ed",
          2292 => x"d3",
          2293 => x"81",
          2294 => x"80",
          2295 => x"16",
          2296 => x"56",
          2297 => x"38",
          2298 => x"e2",
          2299 => x"08",
          2300 => x"70",
          2301 => x"81",
          2302 => x"51",
          2303 => x"86",
          2304 => x"81",
          2305 => x"30",
          2306 => x"70",
          2307 => x"06",
          2308 => x"51",
          2309 => x"73",
          2310 => x"38",
          2311 => x"96",
          2312 => x"df",
          2313 => x"72",
          2314 => x"81",
          2315 => x"81",
          2316 => x"2e",
          2317 => x"52",
          2318 => x"fa",
          2319 => x"ac",
          2320 => x"d3",
          2321 => x"38",
          2322 => x"fe",
          2323 => x"80",
          2324 => x"80",
          2325 => x"0c",
          2326 => x"ac",
          2327 => x"0d",
          2328 => x"0d",
          2329 => x"59",
          2330 => x"75",
          2331 => x"3f",
          2332 => x"08",
          2333 => x"ac",
          2334 => x"38",
          2335 => x"57",
          2336 => x"98",
          2337 => x"77",
          2338 => x"3f",
          2339 => x"08",
          2340 => x"ac",
          2341 => x"38",
          2342 => x"70",
          2343 => x"73",
          2344 => x"38",
          2345 => x"8b",
          2346 => x"06",
          2347 => x"86",
          2348 => x"15",
          2349 => x"2a",
          2350 => x"51",
          2351 => x"93",
          2352 => x"a0",
          2353 => x"51",
          2354 => x"81",
          2355 => x"80",
          2356 => x"80",
          2357 => x"f9",
          2358 => x"d3",
          2359 => x"81",
          2360 => x"80",
          2361 => x"38",
          2362 => x"81",
          2363 => x"8a",
          2364 => x"fb",
          2365 => x"70",
          2366 => x"81",
          2367 => x"fb",
          2368 => x"d3",
          2369 => x"81",
          2370 => x"b4",
          2371 => x"08",
          2372 => x"eb",
          2373 => x"d3",
          2374 => x"81",
          2375 => x"a0",
          2376 => x"81",
          2377 => x"52",
          2378 => x"51",
          2379 => x"8b",
          2380 => x"52",
          2381 => x"51",
          2382 => x"81",
          2383 => x"34",
          2384 => x"ac",
          2385 => x"0d",
          2386 => x"0d",
          2387 => x"98",
          2388 => x"70",
          2389 => x"ea",
          2390 => x"d3",
          2391 => x"81",
          2392 => x"8d",
          2393 => x"08",
          2394 => x"34",
          2395 => x"16",
          2396 => x"d3",
          2397 => x"3d",
          2398 => x"3d",
          2399 => x"57",
          2400 => x"89",
          2401 => x"17",
          2402 => x"81",
          2403 => x"70",
          2404 => x"17",
          2405 => x"33",
          2406 => x"54",
          2407 => x"2e",
          2408 => x"85",
          2409 => x"06",
          2410 => x"e5",
          2411 => x"2e",
          2412 => x"8e",
          2413 => x"88",
          2414 => x"0b",
          2415 => x"81",
          2416 => x"15",
          2417 => x"72",
          2418 => x"81",
          2419 => x"74",
          2420 => x"75",
          2421 => x"52",
          2422 => x"13",
          2423 => x"08",
          2424 => x"33",
          2425 => x"9c",
          2426 => x"05",
          2427 => x"3f",
          2428 => x"08",
          2429 => x"17",
          2430 => x"51",
          2431 => x"81",
          2432 => x"86",
          2433 => x"17",
          2434 => x"51",
          2435 => x"81",
          2436 => x"84",
          2437 => x"3d",
          2438 => x"3d",
          2439 => x"08",
          2440 => x"5d",
          2441 => x"53",
          2442 => x"51",
          2443 => x"80",
          2444 => x"88",
          2445 => x"5a",
          2446 => x"09",
          2447 => x"df",
          2448 => x"70",
          2449 => x"71",
          2450 => x"30",
          2451 => x"73",
          2452 => x"51",
          2453 => x"57",
          2454 => x"38",
          2455 => x"75",
          2456 => x"18",
          2457 => x"75",
          2458 => x"30",
          2459 => x"32",
          2460 => x"73",
          2461 => x"53",
          2462 => x"55",
          2463 => x"89",
          2464 => x"75",
          2465 => x"e4",
          2466 => x"7c",
          2467 => x"a0",
          2468 => x"38",
          2469 => x"8b",
          2470 => x"54",
          2471 => x"78",
          2472 => x"81",
          2473 => x"54",
          2474 => x"82",
          2475 => x"af",
          2476 => x"77",
          2477 => x"70",
          2478 => x"25",
          2479 => x"07",
          2480 => x"51",
          2481 => x"2e",
          2482 => x"39",
          2483 => x"80",
          2484 => x"33",
          2485 => x"73",
          2486 => x"81",
          2487 => x"81",
          2488 => x"1a",
          2489 => x"55",
          2490 => x"dc",
          2491 => x"06",
          2492 => x"55",
          2493 => x"54",
          2494 => x"81",
          2495 => x"ae",
          2496 => x"70",
          2497 => x"7d",
          2498 => x"51",
          2499 => x"2e",
          2500 => x"8b",
          2501 => x"77",
          2502 => x"30",
          2503 => x"71",
          2504 => x"53",
          2505 => x"55",
          2506 => x"38",
          2507 => x"5a",
          2508 => x"75",
          2509 => x"73",
          2510 => x"38",
          2511 => x"06",
          2512 => x"11",
          2513 => x"75",
          2514 => x"3f",
          2515 => x"08",
          2516 => x"38",
          2517 => x"33",
          2518 => x"54",
          2519 => x"e5",
          2520 => x"d3",
          2521 => x"2e",
          2522 => x"1a",
          2523 => x"26",
          2524 => x"54",
          2525 => x"7a",
          2526 => x"74",
          2527 => x"7b",
          2528 => x"74",
          2529 => x"18",
          2530 => x"39",
          2531 => x"ba",
          2532 => x"ec",
          2533 => x"ac",
          2534 => x"38",
          2535 => x"54",
          2536 => x"89",
          2537 => x"70",
          2538 => x"57",
          2539 => x"54",
          2540 => x"81",
          2541 => x"e7",
          2542 => x"7c",
          2543 => x"77",
          2544 => x"38",
          2545 => x"73",
          2546 => x"09",
          2547 => x"38",
          2548 => x"84",
          2549 => x"27",
          2550 => x"39",
          2551 => x"39",
          2552 => x"39",
          2553 => x"8b",
          2554 => x"54",
          2555 => x"ac",
          2556 => x"0d",
          2557 => x"0d",
          2558 => x"58",
          2559 => x"70",
          2560 => x"55",
          2561 => x"83",
          2562 => x"80",
          2563 => x"51",
          2564 => x"80",
          2565 => x"38",
          2566 => x"74",
          2567 => x"80",
          2568 => x"94",
          2569 => x"17",
          2570 => x"81",
          2571 => x"7a",
          2572 => x"54",
          2573 => x"2e",
          2574 => x"83",
          2575 => x"80",
          2576 => x"51",
          2577 => x"80",
          2578 => x"81",
          2579 => x"81",
          2580 => x"07",
          2581 => x"38",
          2582 => x"17",
          2583 => x"33",
          2584 => x"9f",
          2585 => x"ff",
          2586 => x"17",
          2587 => x"75",
          2588 => x"3f",
          2589 => x"08",
          2590 => x"39",
          2591 => x"a5",
          2592 => x"84",
          2593 => x"51",
          2594 => x"81",
          2595 => x"55",
          2596 => x"08",
          2597 => x"75",
          2598 => x"3f",
          2599 => x"08",
          2600 => x"55",
          2601 => x"ac",
          2602 => x"80",
          2603 => x"d3",
          2604 => x"2e",
          2605 => x"80",
          2606 => x"85",
          2607 => x"06",
          2608 => x"80",
          2609 => x"73",
          2610 => x"81",
          2611 => x"72",
          2612 => x"ad",
          2613 => x"0b",
          2614 => x"80",
          2615 => x"39",
          2616 => x"70",
          2617 => x"53",
          2618 => x"85",
          2619 => x"73",
          2620 => x"81",
          2621 => x"72",
          2622 => x"16",
          2623 => x"2a",
          2624 => x"51",
          2625 => x"80",
          2626 => x"38",
          2627 => x"83",
          2628 => x"b4",
          2629 => x"51",
          2630 => x"81",
          2631 => x"88",
          2632 => x"dd",
          2633 => x"d3",
          2634 => x"3d",
          2635 => x"3d",
          2636 => x"ff",
          2637 => x"72",
          2638 => x"5a",
          2639 => x"81",
          2640 => x"70",
          2641 => x"33",
          2642 => x"70",
          2643 => x"26",
          2644 => x"06",
          2645 => x"53",
          2646 => x"72",
          2647 => x"81",
          2648 => x"38",
          2649 => x"11",
          2650 => x"89",
          2651 => x"82",
          2652 => x"ff",
          2653 => x"51",
          2654 => x"77",
          2655 => x"38",
          2656 => x"bb",
          2657 => x"77",
          2658 => x"70",
          2659 => x"57",
          2660 => x"70",
          2661 => x"33",
          2662 => x"05",
          2663 => x"9f",
          2664 => x"54",
          2665 => x"89",
          2666 => x"70",
          2667 => x"55",
          2668 => x"13",
          2669 => x"26",
          2670 => x"13",
          2671 => x"06",
          2672 => x"30",
          2673 => x"70",
          2674 => x"07",
          2675 => x"9f",
          2676 => x"55",
          2677 => x"ff",
          2678 => x"30",
          2679 => x"70",
          2680 => x"07",
          2681 => x"9f",
          2682 => x"55",
          2683 => x"80",
          2684 => x"81",
          2685 => x"78",
          2686 => x"38",
          2687 => x"83",
          2688 => x"77",
          2689 => x"5a",
          2690 => x"39",
          2691 => x"33",
          2692 => x"d3",
          2693 => x"3d",
          2694 => x"3d",
          2695 => x"80",
          2696 => x"34",
          2697 => x"17",
          2698 => x"75",
          2699 => x"3f",
          2700 => x"d3",
          2701 => x"84",
          2702 => x"16",
          2703 => x"3f",
          2704 => x"08",
          2705 => x"06",
          2706 => x"73",
          2707 => x"2e",
          2708 => x"80",
          2709 => x"0b",
          2710 => x"55",
          2711 => x"e9",
          2712 => x"06",
          2713 => x"55",
          2714 => x"32",
          2715 => x"80",
          2716 => x"51",
          2717 => x"8e",
          2718 => x"33",
          2719 => x"e8",
          2720 => x"06",
          2721 => x"53",
          2722 => x"52",
          2723 => x"51",
          2724 => x"81",
          2725 => x"55",
          2726 => x"08",
          2727 => x"38",
          2728 => x"ba",
          2729 => x"86",
          2730 => x"a3",
          2731 => x"ac",
          2732 => x"d3",
          2733 => x"2e",
          2734 => x"55",
          2735 => x"ac",
          2736 => x"0d",
          2737 => x"0d",
          2738 => x"05",
          2739 => x"33",
          2740 => x"74",
          2741 => x"fc",
          2742 => x"d3",
          2743 => x"8b",
          2744 => x"81",
          2745 => x"24",
          2746 => x"81",
          2747 => x"10",
          2748 => x"c8",
          2749 => x"56",
          2750 => x"74",
          2751 => x"88",
          2752 => x"0c",
          2753 => x"06",
          2754 => x"57",
          2755 => x"af",
          2756 => x"33",
          2757 => x"3f",
          2758 => x"08",
          2759 => x"70",
          2760 => x"54",
          2761 => x"76",
          2762 => x"38",
          2763 => x"70",
          2764 => x"53",
          2765 => x"86",
          2766 => x"56",
          2767 => x"80",
          2768 => x"81",
          2769 => x"52",
          2770 => x"51",
          2771 => x"81",
          2772 => x"81",
          2773 => x"81",
          2774 => x"83",
          2775 => x"a8",
          2776 => x"2e",
          2777 => x"82",
          2778 => x"06",
          2779 => x"56",
          2780 => x"38",
          2781 => x"75",
          2782 => x"9e",
          2783 => x"ac",
          2784 => x"06",
          2785 => x"2e",
          2786 => x"80",
          2787 => x"54",
          2788 => x"15",
          2789 => x"10",
          2790 => x"05",
          2791 => x"33",
          2792 => x"80",
          2793 => x"2e",
          2794 => x"fa",
          2795 => x"eb",
          2796 => x"ac",
          2797 => x"78",
          2798 => x"54",
          2799 => x"d0",
          2800 => x"8f",
          2801 => x"10",
          2802 => x"08",
          2803 => x"57",
          2804 => x"90",
          2805 => x"74",
          2806 => x"3f",
          2807 => x"08",
          2808 => x"57",
          2809 => x"89",
          2810 => x"54",
          2811 => x"d3",
          2812 => x"76",
          2813 => x"90",
          2814 => x"76",
          2815 => x"88",
          2816 => x"51",
          2817 => x"81",
          2818 => x"83",
          2819 => x"53",
          2820 => x"84",
          2821 => x"81",
          2822 => x"38",
          2823 => x"51",
          2824 => x"81",
          2825 => x"83",
          2826 => x"54",
          2827 => x"80",
          2828 => x"d9",
          2829 => x"d3",
          2830 => x"73",
          2831 => x"80",
          2832 => x"82",
          2833 => x"c4",
          2834 => x"05",
          2835 => x"72",
          2836 => x"b4",
          2837 => x"33",
          2838 => x"80",
          2839 => x"52",
          2840 => x"8a",
          2841 => x"83",
          2842 => x"53",
          2843 => x"8b",
          2844 => x"73",
          2845 => x"80",
          2846 => x"8d",
          2847 => x"39",
          2848 => x"51",
          2849 => x"81",
          2850 => x"88",
          2851 => x"d3",
          2852 => x"ff",
          2853 => x"06",
          2854 => x"72",
          2855 => x"80",
          2856 => x"d8",
          2857 => x"d3",
          2858 => x"ff",
          2859 => x"72",
          2860 => x"d4",
          2861 => x"e3",
          2862 => x"ac",
          2863 => x"c2",
          2864 => x"be",
          2865 => x"ac",
          2866 => x"ff",
          2867 => x"56",
          2868 => x"83",
          2869 => x"15",
          2870 => x"71",
          2871 => x"59",
          2872 => x"77",
          2873 => x"a0",
          2874 => x"22",
          2875 => x"31",
          2876 => x"ab",
          2877 => x"ac",
          2878 => x"56",
          2879 => x"08",
          2880 => x"84",
          2881 => x"81",
          2882 => x"80",
          2883 => x"f5",
          2884 => x"83",
          2885 => x"ff",
          2886 => x"38",
          2887 => x"9f",
          2888 => x"38",
          2889 => x"56",
          2890 => x"82",
          2891 => x"13",
          2892 => x"79",
          2893 => x"79",
          2894 => x"0c",
          2895 => x"16",
          2896 => x"2e",
          2897 => x"b7",
          2898 => x"15",
          2899 => x"3f",
          2900 => x"08",
          2901 => x"06",
          2902 => x"72",
          2903 => x"88",
          2904 => x"8d",
          2905 => x"a0",
          2906 => x"15",
          2907 => x"3f",
          2908 => x"08",
          2909 => x"98",
          2910 => x"2b",
          2911 => x"88",
          2912 => x"8d",
          2913 => x"2e",
          2914 => x"a4",
          2915 => x"a8",
          2916 => x"82",
          2917 => x"06",
          2918 => x"15",
          2919 => x"94",
          2920 => x"08",
          2921 => x"08",
          2922 => x"2a",
          2923 => x"81",
          2924 => x"53",
          2925 => x"89",
          2926 => x"56",
          2927 => x"08",
          2928 => x"38",
          2929 => x"16",
          2930 => x"8c",
          2931 => x"80",
          2932 => x"34",
          2933 => x"09",
          2934 => x"92",
          2935 => x"15",
          2936 => x"3f",
          2937 => x"08",
          2938 => x"06",
          2939 => x"2e",
          2940 => x"80",
          2941 => x"1a",
          2942 => x"d9",
          2943 => x"d3",
          2944 => x"ea",
          2945 => x"ac",
          2946 => x"34",
          2947 => x"51",
          2948 => x"81",
          2949 => x"83",
          2950 => x"53",
          2951 => x"d5",
          2952 => x"06",
          2953 => x"b4",
          2954 => x"ef",
          2955 => x"ac",
          2956 => x"85",
          2957 => x"09",
          2958 => x"38",
          2959 => x"51",
          2960 => x"81",
          2961 => x"86",
          2962 => x"f2",
          2963 => x"06",
          2964 => x"9c",
          2965 => x"c3",
          2966 => x"ac",
          2967 => x"0c",
          2968 => x"51",
          2969 => x"81",
          2970 => x"8c",
          2971 => x"75",
          2972 => x"d8",
          2973 => x"53",
          2974 => x"d8",
          2975 => x"16",
          2976 => x"94",
          2977 => x"56",
          2978 => x"ac",
          2979 => x"0d",
          2980 => x"0d",
          2981 => x"55",
          2982 => x"b5",
          2983 => x"80",
          2984 => x"73",
          2985 => x"53",
          2986 => x"2e",
          2987 => x"14",
          2988 => x"22",
          2989 => x"76",
          2990 => x"06",
          2991 => x"13",
          2992 => x"f9",
          2993 => x"ac",
          2994 => x"52",
          2995 => x"71",
          2996 => x"74",
          2997 => x"81",
          2998 => x"73",
          2999 => x"73",
          3000 => x"74",
          3001 => x"0c",
          3002 => x"04",
          3003 => x"02",
          3004 => x"7a",
          3005 => x"fc",
          3006 => x"f4",
          3007 => x"d3",
          3008 => x"8b",
          3009 => x"81",
          3010 => x"24",
          3011 => x"81",
          3012 => x"10",
          3013 => x"c8",
          3014 => x"51",
          3015 => x"2e",
          3016 => x"74",
          3017 => x"2e",
          3018 => x"54",
          3019 => x"74",
          3020 => x"d3",
          3021 => x"71",
          3022 => x"54",
          3023 => x"92",
          3024 => x"89",
          3025 => x"84",
          3026 => x"f9",
          3027 => x"ac",
          3028 => x"81",
          3029 => x"88",
          3030 => x"eb",
          3031 => x"02",
          3032 => x"e7",
          3033 => x"58",
          3034 => x"80",
          3035 => x"38",
          3036 => x"70",
          3037 => x"d0",
          3038 => x"3d",
          3039 => x"57",
          3040 => x"81",
          3041 => x"56",
          3042 => x"08",
          3043 => x"7a",
          3044 => x"97",
          3045 => x"51",
          3046 => x"81",
          3047 => x"56",
          3048 => x"08",
          3049 => x"80",
          3050 => x"70",
          3051 => x"59",
          3052 => x"83",
          3053 => x"76",
          3054 => x"74",
          3055 => x"c3",
          3056 => x"2e",
          3057 => x"84",
          3058 => x"06",
          3059 => x"3d",
          3060 => x"ea",
          3061 => x"d3",
          3062 => x"76",
          3063 => x"a0",
          3064 => x"05",
          3065 => x"55",
          3066 => x"85",
          3067 => x"90",
          3068 => x"2a",
          3069 => x"51",
          3070 => x"2e",
          3071 => x"56",
          3072 => x"38",
          3073 => x"70",
          3074 => x"55",
          3075 => x"81",
          3076 => x"52",
          3077 => x"b6",
          3078 => x"ac",
          3079 => x"88",
          3080 => x"62",
          3081 => x"d2",
          3082 => x"55",
          3083 => x"16",
          3084 => x"62",
          3085 => x"e6",
          3086 => x"52",
          3087 => x"51",
          3088 => x"7a",
          3089 => x"83",
          3090 => x"80",
          3091 => x"38",
          3092 => x"08",
          3093 => x"54",
          3094 => x"05",
          3095 => x"db",
          3096 => x"d3",
          3097 => x"81",
          3098 => x"82",
          3099 => x"52",
          3100 => x"bc",
          3101 => x"ac",
          3102 => x"1b",
          3103 => x"56",
          3104 => x"75",
          3105 => x"02",
          3106 => x"70",
          3107 => x"81",
          3108 => x"59",
          3109 => x"85",
          3110 => x"9c",
          3111 => x"2a",
          3112 => x"51",
          3113 => x"2e",
          3114 => x"b2",
          3115 => x"06",
          3116 => x"2e",
          3117 => x"56",
          3118 => x"38",
          3119 => x"70",
          3120 => x"55",
          3121 => x"86",
          3122 => x"c0",
          3123 => x"b0",
          3124 => x"1a",
          3125 => x"1a",
          3126 => x"81",
          3127 => x"52",
          3128 => x"ea",
          3129 => x"ac",
          3130 => x"0c",
          3131 => x"51",
          3132 => x"81",
          3133 => x"8c",
          3134 => x"78",
          3135 => x"22",
          3136 => x"76",
          3137 => x"75",
          3138 => x"75",
          3139 => x"75",
          3140 => x"84",
          3141 => x"52",
          3142 => x"d1",
          3143 => x"85",
          3144 => x"06",
          3145 => x"80",
          3146 => x"38",
          3147 => x"80",
          3148 => x"38",
          3149 => x"94",
          3150 => x"8a",
          3151 => x"89",
          3152 => x"08",
          3153 => x"5d",
          3154 => x"55",
          3155 => x"52",
          3156 => x"fc",
          3157 => x"ac",
          3158 => x"d3",
          3159 => x"26",
          3160 => x"56",
          3161 => x"09",
          3162 => x"38",
          3163 => x"7a",
          3164 => x"30",
          3165 => x"80",
          3166 => x"7d",
          3167 => x"51",
          3168 => x"38",
          3169 => x"0c",
          3170 => x"38",
          3171 => x"06",
          3172 => x"2e",
          3173 => x"52",
          3174 => x"8a",
          3175 => x"ac",
          3176 => x"82",
          3177 => x"78",
          3178 => x"d3",
          3179 => x"70",
          3180 => x"55",
          3181 => x"53",
          3182 => x"7a",
          3183 => x"52",
          3184 => x"3f",
          3185 => x"08",
          3186 => x"38",
          3187 => x"80",
          3188 => x"80",
          3189 => x"55",
          3190 => x"ac",
          3191 => x"0d",
          3192 => x"0d",
          3193 => x"63",
          3194 => x"57",
          3195 => x"8f",
          3196 => x"52",
          3197 => x"99",
          3198 => x"ac",
          3199 => x"d3",
          3200 => x"38",
          3201 => x"55",
          3202 => x"86",
          3203 => x"83",
          3204 => x"17",
          3205 => x"55",
          3206 => x"80",
          3207 => x"38",
          3208 => x"0b",
          3209 => x"82",
          3210 => x"39",
          3211 => x"18",
          3212 => x"83",
          3213 => x"0b",
          3214 => x"82",
          3215 => x"39",
          3216 => x"18",
          3217 => x"82",
          3218 => x"0b",
          3219 => x"81",
          3220 => x"39",
          3221 => x"18",
          3222 => x"82",
          3223 => x"17",
          3224 => x"08",
          3225 => x"79",
          3226 => x"74",
          3227 => x"2e",
          3228 => x"94",
          3229 => x"83",
          3230 => x"56",
          3231 => x"38",
          3232 => x"22",
          3233 => x"89",
          3234 => x"55",
          3235 => x"75",
          3236 => x"17",
          3237 => x"39",
          3238 => x"52",
          3239 => x"b0",
          3240 => x"ac",
          3241 => x"75",
          3242 => x"38",
          3243 => x"fe",
          3244 => x"98",
          3245 => x"17",
          3246 => x"51",
          3247 => x"81",
          3248 => x"80",
          3249 => x"38",
          3250 => x"08",
          3251 => x"2a",
          3252 => x"80",
          3253 => x"38",
          3254 => x"8a",
          3255 => x"56",
          3256 => x"27",
          3257 => x"7b",
          3258 => x"54",
          3259 => x"52",
          3260 => x"33",
          3261 => x"ef",
          3262 => x"ac",
          3263 => x"38",
          3264 => x"70",
          3265 => x"56",
          3266 => x"9b",
          3267 => x"08",
          3268 => x"74",
          3269 => x"38",
          3270 => x"a8",
          3271 => x"84",
          3272 => x"51",
          3273 => x"79",
          3274 => x"80",
          3275 => x"17",
          3276 => x"80",
          3277 => x"17",
          3278 => x"2b",
          3279 => x"80",
          3280 => x"81",
          3281 => x"08",
          3282 => x"52",
          3283 => x"33",
          3284 => x"ec",
          3285 => x"ac",
          3286 => x"38",
          3287 => x"80",
          3288 => x"74",
          3289 => x"81",
          3290 => x"a8",
          3291 => x"81",
          3292 => x"55",
          3293 => x"81",
          3294 => x"fd",
          3295 => x"9c",
          3296 => x"17",
          3297 => x"06",
          3298 => x"31",
          3299 => x"76",
          3300 => x"78",
          3301 => x"94",
          3302 => x"ff",
          3303 => x"05",
          3304 => x"cb",
          3305 => x"76",
          3306 => x"17",
          3307 => x"1d",
          3308 => x"18",
          3309 => x"5d",
          3310 => x"b7",
          3311 => x"75",
          3312 => x"0c",
          3313 => x"04",
          3314 => x"7f",
          3315 => x"5f",
          3316 => x"80",
          3317 => x"3d",
          3318 => x"76",
          3319 => x"3f",
          3320 => x"08",
          3321 => x"ac",
          3322 => x"91",
          3323 => x"74",
          3324 => x"38",
          3325 => x"82",
          3326 => x"33",
          3327 => x"70",
          3328 => x"56",
          3329 => x"74",
          3330 => x"ee",
          3331 => x"82",
          3332 => x"34",
          3333 => x"e2",
          3334 => x"91",
          3335 => x"56",
          3336 => x"81",
          3337 => x"34",
          3338 => x"ce",
          3339 => x"91",
          3340 => x"56",
          3341 => x"81",
          3342 => x"34",
          3343 => x"ba",
          3344 => x"91",
          3345 => x"56",
          3346 => x"94",
          3347 => x"55",
          3348 => x"08",
          3349 => x"94",
          3350 => x"59",
          3351 => x"83",
          3352 => x"17",
          3353 => x"ff",
          3354 => x"74",
          3355 => x"7d",
          3356 => x"ff",
          3357 => x"2a",
          3358 => x"7a",
          3359 => x"75",
          3360 => x"17",
          3361 => x"a3",
          3362 => x"76",
          3363 => x"3f",
          3364 => x"08",
          3365 => x"98",
          3366 => x"76",
          3367 => x"3f",
          3368 => x"08",
          3369 => x"2e",
          3370 => x"74",
          3371 => x"df",
          3372 => x"2e",
          3373 => x"74",
          3374 => x"88",
          3375 => x"38",
          3376 => x"0c",
          3377 => x"70",
          3378 => x"58",
          3379 => x"a5",
          3380 => x"9c",
          3381 => x"a8",
          3382 => x"81",
          3383 => x"55",
          3384 => x"81",
          3385 => x"fe",
          3386 => x"17",
          3387 => x"06",
          3388 => x"18",
          3389 => x"08",
          3390 => x"cd",
          3391 => x"d3",
          3392 => x"2e",
          3393 => x"81",
          3394 => x"1b",
          3395 => x"5b",
          3396 => x"2e",
          3397 => x"79",
          3398 => x"11",
          3399 => x"56",
          3400 => x"85",
          3401 => x"31",
          3402 => x"77",
          3403 => x"7d",
          3404 => x"52",
          3405 => x"3f",
          3406 => x"08",
          3407 => x"9c",
          3408 => x"31",
          3409 => x"27",
          3410 => x"80",
          3411 => x"80",
          3412 => x"a8",
          3413 => x"b9",
          3414 => x"33",
          3415 => x"55",
          3416 => x"34",
          3417 => x"56",
          3418 => x"9c",
          3419 => x"2e",
          3420 => x"17",
          3421 => x"08",
          3422 => x"81",
          3423 => x"a8",
          3424 => x"81",
          3425 => x"55",
          3426 => x"81",
          3427 => x"fd",
          3428 => x"9c",
          3429 => x"17",
          3430 => x"06",
          3431 => x"31",
          3432 => x"76",
          3433 => x"78",
          3434 => x"7b",
          3435 => x"08",
          3436 => x"17",
          3437 => x"c7",
          3438 => x"17",
          3439 => x"07",
          3440 => x"18",
          3441 => x"31",
          3442 => x"7e",
          3443 => x"94",
          3444 => x"70",
          3445 => x"8c",
          3446 => x"58",
          3447 => x"76",
          3448 => x"75",
          3449 => x"18",
          3450 => x"f6",
          3451 => x"33",
          3452 => x"55",
          3453 => x"34",
          3454 => x"81",
          3455 => x"8f",
          3456 => x"f7",
          3457 => x"8c",
          3458 => x"53",
          3459 => x"f1",
          3460 => x"d3",
          3461 => x"81",
          3462 => x"81",
          3463 => x"18",
          3464 => x"2a",
          3465 => x"51",
          3466 => x"80",
          3467 => x"38",
          3468 => x"55",
          3469 => x"a7",
          3470 => x"9c",
          3471 => x"a8",
          3472 => x"81",
          3473 => x"55",
          3474 => x"81",
          3475 => x"ac",
          3476 => x"38",
          3477 => x"80",
          3478 => x"74",
          3479 => x"a0",
          3480 => x"79",
          3481 => x"3f",
          3482 => x"08",
          3483 => x"ac",
          3484 => x"38",
          3485 => x"8b",
          3486 => x"07",
          3487 => x"8b",
          3488 => x"18",
          3489 => x"52",
          3490 => x"d9",
          3491 => x"18",
          3492 => x"16",
          3493 => x"3f",
          3494 => x"0a",
          3495 => x"51",
          3496 => x"76",
          3497 => x"51",
          3498 => x"79",
          3499 => x"83",
          3500 => x"51",
          3501 => x"81",
          3502 => x"90",
          3503 => x"bf",
          3504 => x"74",
          3505 => x"76",
          3506 => x"d3",
          3507 => x"3d",
          3508 => x"3d",
          3509 => x"52",
          3510 => x"3f",
          3511 => x"08",
          3512 => x"ac",
          3513 => x"86",
          3514 => x"52",
          3515 => x"a1",
          3516 => x"ac",
          3517 => x"d3",
          3518 => x"38",
          3519 => x"08",
          3520 => x"81",
          3521 => x"86",
          3522 => x"fe",
          3523 => x"3d",
          3524 => x"3f",
          3525 => x"0b",
          3526 => x"08",
          3527 => x"81",
          3528 => x"81",
          3529 => x"80",
          3530 => x"d3",
          3531 => x"3d",
          3532 => x"3d",
          3533 => x"93",
          3534 => x"52",
          3535 => x"e7",
          3536 => x"d3",
          3537 => x"81",
          3538 => x"80",
          3539 => x"58",
          3540 => x"3d",
          3541 => x"e1",
          3542 => x"d3",
          3543 => x"81",
          3544 => x"be",
          3545 => x"c7",
          3546 => x"98",
          3547 => x"73",
          3548 => x"38",
          3549 => x"12",
          3550 => x"39",
          3551 => x"33",
          3552 => x"70",
          3553 => x"55",
          3554 => x"2e",
          3555 => x"7f",
          3556 => x"54",
          3557 => x"81",
          3558 => x"94",
          3559 => x"39",
          3560 => x"84",
          3561 => x"06",
          3562 => x"55",
          3563 => x"ac",
          3564 => x"0d",
          3565 => x"0d",
          3566 => x"a3",
          3567 => x"5c",
          3568 => x"80",
          3569 => x"ff",
          3570 => x"a2",
          3571 => x"f5",
          3572 => x"ac",
          3573 => x"d3",
          3574 => x"93",
          3575 => x"7b",
          3576 => x"08",
          3577 => x"56",
          3578 => x"2e",
          3579 => x"96",
          3580 => x"3d",
          3581 => x"a0",
          3582 => x"d1",
          3583 => x"d3",
          3584 => x"81",
          3585 => x"81",
          3586 => x"52",
          3587 => x"a0",
          3588 => x"ac",
          3589 => x"d3",
          3590 => x"cb",
          3591 => x"7e",
          3592 => x"3f",
          3593 => x"08",
          3594 => x"7a",
          3595 => x"3f",
          3596 => x"08",
          3597 => x"ac",
          3598 => x"38",
          3599 => x"52",
          3600 => x"f1",
          3601 => x"ac",
          3602 => x"d3",
          3603 => x"38",
          3604 => x"51",
          3605 => x"81",
          3606 => x"75",
          3607 => x"76",
          3608 => x"d2",
          3609 => x"d3",
          3610 => x"81",
          3611 => x"80",
          3612 => x"76",
          3613 => x"81",
          3614 => x"82",
          3615 => x"ef",
          3616 => x"ff",
          3617 => x"d4",
          3618 => x"ee",
          3619 => x"3d",
          3620 => x"81",
          3621 => x"52",
          3622 => x"73",
          3623 => x"38",
          3624 => x"16",
          3625 => x"51",
          3626 => x"f4",
          3627 => x"54",
          3628 => x"85",
          3629 => x"af",
          3630 => x"2e",
          3631 => x"58",
          3632 => x"3d",
          3633 => x"18",
          3634 => x"58",
          3635 => x"14",
          3636 => x"75",
          3637 => x"19",
          3638 => x"11",
          3639 => x"74",
          3640 => x"74",
          3641 => x"76",
          3642 => x"78",
          3643 => x"81",
          3644 => x"ff",
          3645 => x"08",
          3646 => x"af",
          3647 => x"70",
          3648 => x"33",
          3649 => x"81",
          3650 => x"70",
          3651 => x"52",
          3652 => x"57",
          3653 => x"2e",
          3654 => x"16",
          3655 => x"33",
          3656 => x"73",
          3657 => x"16",
          3658 => x"26",
          3659 => x"58",
          3660 => x"94",
          3661 => x"54",
          3662 => x"70",
          3663 => x"34",
          3664 => x"75",
          3665 => x"38",
          3666 => x"81",
          3667 => x"81",
          3668 => x"83",
          3669 => x"76",
          3670 => x"3d",
          3671 => x"1a",
          3672 => x"33",
          3673 => x"05",
          3674 => x"79",
          3675 => x"80",
          3676 => x"81",
          3677 => x"a1",
          3678 => x"f4",
          3679 => x"60",
          3680 => x"05",
          3681 => x"59",
          3682 => x"3f",
          3683 => x"08",
          3684 => x"ac",
          3685 => x"91",
          3686 => x"79",
          3687 => x"38",
          3688 => x"f9",
          3689 => x"08",
          3690 => x"38",
          3691 => x"70",
          3692 => x"81",
          3693 => x"56",
          3694 => x"8c",
          3695 => x"94",
          3696 => x"80",
          3697 => x"0c",
          3698 => x"2e",
          3699 => x"7c",
          3700 => x"70",
          3701 => x"51",
          3702 => x"2e",
          3703 => x"52",
          3704 => x"ff",
          3705 => x"81",
          3706 => x"ff",
          3707 => x"70",
          3708 => x"ff",
          3709 => x"81",
          3710 => x"75",
          3711 => x"78",
          3712 => x"94",
          3713 => x"94",
          3714 => x"98",
          3715 => x"58",
          3716 => x"88",
          3717 => x"75",
          3718 => x"52",
          3719 => x"a7",
          3720 => x"ac",
          3721 => x"d3",
          3722 => x"2e",
          3723 => x"8b",
          3724 => x"91",
          3725 => x"55",
          3726 => x"81",
          3727 => x"ff",
          3728 => x"06",
          3729 => x"0b",
          3730 => x"81",
          3731 => x"39",
          3732 => x"08",
          3733 => x"75",
          3734 => x"75",
          3735 => x"a1",
          3736 => x"27",
          3737 => x"77",
          3738 => x"18",
          3739 => x"19",
          3740 => x"33",
          3741 => x"70",
          3742 => x"57",
          3743 => x"80",
          3744 => x"75",
          3745 => x"c8",
          3746 => x"d3",
          3747 => x"81",
          3748 => x"94",
          3749 => x"ac",
          3750 => x"39",
          3751 => x"51",
          3752 => x"81",
          3753 => x"56",
          3754 => x"81",
          3755 => x"76",
          3756 => x"7c",
          3757 => x"08",
          3758 => x"38",
          3759 => x"18",
          3760 => x"81",
          3761 => x"98",
          3762 => x"79",
          3763 => x"38",
          3764 => x"18",
          3765 => x"77",
          3766 => x"55",
          3767 => x"a1",
          3768 => x"7c",
          3769 => x"3f",
          3770 => x"08",
          3771 => x"0b",
          3772 => x"82",
          3773 => x"39",
          3774 => x"81",
          3775 => x"05",
          3776 => x"08",
          3777 => x"27",
          3778 => x"17",
          3779 => x"0c",
          3780 => x"80",
          3781 => x"74",
          3782 => x"94",
          3783 => x"ff",
          3784 => x"80",
          3785 => x"38",
          3786 => x"7b",
          3787 => x"38",
          3788 => x"70",
          3789 => x"5c",
          3790 => x"b0",
          3791 => x"9c",
          3792 => x"a8",
          3793 => x"81",
          3794 => x"55",
          3795 => x"3f",
          3796 => x"08",
          3797 => x"38",
          3798 => x"18",
          3799 => x"bd",
          3800 => x"33",
          3801 => x"55",
          3802 => x"34",
          3803 => x"53",
          3804 => x"7c",
          3805 => x"52",
          3806 => x"eb",
          3807 => x"ac",
          3808 => x"93",
          3809 => x"91",
          3810 => x"55",
          3811 => x"0b",
          3812 => x"81",
          3813 => x"7a",
          3814 => x"79",
          3815 => x"d3",
          3816 => x"3d",
          3817 => x"3d",
          3818 => x"89",
          3819 => x"2e",
          3820 => x"80",
          3821 => x"fc",
          3822 => x"3d",
          3823 => x"de",
          3824 => x"d3",
          3825 => x"81",
          3826 => x"80",
          3827 => x"76",
          3828 => x"75",
          3829 => x"3f",
          3830 => x"08",
          3831 => x"ac",
          3832 => x"38",
          3833 => x"70",
          3834 => x"57",
          3835 => x"a6",
          3836 => x"33",
          3837 => x"70",
          3838 => x"55",
          3839 => x"2e",
          3840 => x"16",
          3841 => x"51",
          3842 => x"81",
          3843 => x"88",
          3844 => x"39",
          3845 => x"95",
          3846 => x"86",
          3847 => x"17",
          3848 => x"75",
          3849 => x"3f",
          3850 => x"08",
          3851 => x"2e",
          3852 => x"83",
          3853 => x"74",
          3854 => x"38",
          3855 => x"74",
          3856 => x"d3",
          3857 => x"3d",
          3858 => x"3d",
          3859 => x"3d",
          3860 => x"70",
          3861 => x"b9",
          3862 => x"ac",
          3863 => x"d3",
          3864 => x"38",
          3865 => x"08",
          3866 => x"81",
          3867 => x"86",
          3868 => x"fb",
          3869 => x"79",
          3870 => x"05",
          3871 => x"56",
          3872 => x"3f",
          3873 => x"08",
          3874 => x"ac",
          3875 => x"38",
          3876 => x"81",
          3877 => x"52",
          3878 => x"c5",
          3879 => x"ac",
          3880 => x"39",
          3881 => x"51",
          3882 => x"81",
          3883 => x"53",
          3884 => x"08",
          3885 => x"81",
          3886 => x"80",
          3887 => x"38",
          3888 => x"51",
          3889 => x"72",
          3890 => x"c9",
          3891 => x"d3",
          3892 => x"81",
          3893 => x"84",
          3894 => x"06",
          3895 => x"53",
          3896 => x"ac",
          3897 => x"0d",
          3898 => x"0d",
          3899 => x"53",
          3900 => x"53",
          3901 => x"54",
          3902 => x"81",
          3903 => x"55",
          3904 => x"08",
          3905 => x"52",
          3906 => x"e9",
          3907 => x"ac",
          3908 => x"d3",
          3909 => x"38",
          3910 => x"05",
          3911 => x"2b",
          3912 => x"80",
          3913 => x"86",
          3914 => x"75",
          3915 => x"38",
          3916 => x"3d",
          3917 => x"d0",
          3918 => x"81",
          3919 => x"93",
          3920 => x"f2",
          3921 => x"63",
          3922 => x"53",
          3923 => x"05",
          3924 => x"51",
          3925 => x"81",
          3926 => x"59",
          3927 => x"08",
          3928 => x"7a",
          3929 => x"08",
          3930 => x"fe",
          3931 => x"90",
          3932 => x"26",
          3933 => x"15",
          3934 => x"81",
          3935 => x"59",
          3936 => x"82",
          3937 => x"39",
          3938 => x"33",
          3939 => x"73",
          3940 => x"81",
          3941 => x"38",
          3942 => x"56",
          3943 => x"3d",
          3944 => x"ff",
          3945 => x"81",
          3946 => x"ff",
          3947 => x"81",
          3948 => x"81",
          3949 => x"81",
          3950 => x"30",
          3951 => x"ac",
          3952 => x"25",
          3953 => x"18",
          3954 => x"58",
          3955 => x"08",
          3956 => x"38",
          3957 => x"7a",
          3958 => x"a4",
          3959 => x"57",
          3960 => x"74",
          3961 => x"52",
          3962 => x"52",
          3963 => x"c0",
          3964 => x"ac",
          3965 => x"d3",
          3966 => x"d5",
          3967 => x"33",
          3968 => x"82",
          3969 => x"06",
          3970 => x"15",
          3971 => x"ff",
          3972 => x"81",
          3973 => x"83",
          3974 => x"70",
          3975 => x"25",
          3976 => x"58",
          3977 => x"9d",
          3978 => x"b4",
          3979 => x"b5",
          3980 => x"d3",
          3981 => x"0a",
          3982 => x"70",
          3983 => x"84",
          3984 => x"51",
          3985 => x"ff",
          3986 => x"57",
          3987 => x"93",
          3988 => x"0c",
          3989 => x"12",
          3990 => x"84",
          3991 => x"07",
          3992 => x"84",
          3993 => x"81",
          3994 => x"90",
          3995 => x"f8",
          3996 => x"8b",
          3997 => x"53",
          3998 => x"e0",
          3999 => x"d3",
          4000 => x"81",
          4001 => x"8a",
          4002 => x"33",
          4003 => x"2e",
          4004 => x"56",
          4005 => x"90",
          4006 => x"81",
          4007 => x"06",
          4008 => x"87",
          4009 => x"2e",
          4010 => x"94",
          4011 => x"19",
          4012 => x"bc",
          4013 => x"08",
          4014 => x"53",
          4015 => x"52",
          4016 => x"be",
          4017 => x"d3",
          4018 => x"80",
          4019 => x"0c",
          4020 => x"98",
          4021 => x"77",
          4022 => x"f4",
          4023 => x"ac",
          4024 => x"ac",
          4025 => x"70",
          4026 => x"07",
          4027 => x"57",
          4028 => x"d3",
          4029 => x"2e",
          4030 => x"83",
          4031 => x"76",
          4032 => x"55",
          4033 => x"08",
          4034 => x"98",
          4035 => x"75",
          4036 => x"ff",
          4037 => x"81",
          4038 => x"57",
          4039 => x"8c",
          4040 => x"18",
          4041 => x"07",
          4042 => x"19",
          4043 => x"38",
          4044 => x"55",
          4045 => x"ab",
          4046 => x"9c",
          4047 => x"a8",
          4048 => x"81",
          4049 => x"55",
          4050 => x"3f",
          4051 => x"08",
          4052 => x"38",
          4053 => x"39",
          4054 => x"80",
          4055 => x"74",
          4056 => x"76",
          4057 => x"38",
          4058 => x"34",
          4059 => x"39",
          4060 => x"81",
          4061 => x"8a",
          4062 => x"e3",
          4063 => x"ba",
          4064 => x"96",
          4065 => x"53",
          4066 => x"a4",
          4067 => x"3d",
          4068 => x"3f",
          4069 => x"08",
          4070 => x"ac",
          4071 => x"38",
          4072 => x"51",
          4073 => x"3f",
          4074 => x"52",
          4075 => x"05",
          4076 => x"3f",
          4077 => x"08",
          4078 => x"52",
          4079 => x"9a",
          4080 => x"ae",
          4081 => x"f7",
          4082 => x"85",
          4083 => x"06",
          4084 => x"73",
          4085 => x"38",
          4086 => x"82",
          4087 => x"ba",
          4088 => x"95",
          4089 => x"80",
          4090 => x"70",
          4091 => x"55",
          4092 => x"85",
          4093 => x"90",
          4094 => x"d2",
          4095 => x"06",
          4096 => x"2e",
          4097 => x"56",
          4098 => x"38",
          4099 => x"51",
          4100 => x"81",
          4101 => x"02",
          4102 => x"d2",
          4103 => x"84",
          4104 => x"06",
          4105 => x"57",
          4106 => x"80",
          4107 => x"bb",
          4108 => x"95",
          4109 => x"78",
          4110 => x"14",
          4111 => x"80",
          4112 => x"bb",
          4113 => x"95",
          4114 => x"59",
          4115 => x"bb",
          4116 => x"95",
          4117 => x"52",
          4118 => x"52",
          4119 => x"3f",
          4120 => x"08",
          4121 => x"ac",
          4122 => x"38",
          4123 => x"08",
          4124 => x"c6",
          4125 => x"d3",
          4126 => x"81",
          4127 => x"83",
          4128 => x"75",
          4129 => x"30",
          4130 => x"9f",
          4131 => x"58",
          4132 => x"80",
          4133 => x"bb",
          4134 => x"94",
          4135 => x"3d",
          4136 => x"c9",
          4137 => x"d3",
          4138 => x"d3",
          4139 => x"70",
          4140 => x"08",
          4141 => x"79",
          4142 => x"07",
          4143 => x"06",
          4144 => x"56",
          4145 => x"2e",
          4146 => x"bb",
          4147 => x"94",
          4148 => x"53",
          4149 => x"3d",
          4150 => x"ff",
          4151 => x"81",
          4152 => x"56",
          4153 => x"77",
          4154 => x"8b",
          4155 => x"ac",
          4156 => x"bb",
          4157 => x"93",
          4158 => x"81",
          4159 => x"9f",
          4160 => x"ea",
          4161 => x"53",
          4162 => x"05",
          4163 => x"51",
          4164 => x"81",
          4165 => x"55",
          4166 => x"08",
          4167 => x"77",
          4168 => x"98",
          4169 => x"51",
          4170 => x"81",
          4171 => x"55",
          4172 => x"08",
          4173 => x"55",
          4174 => x"09",
          4175 => x"93",
          4176 => x"db",
          4177 => x"85",
          4178 => x"06",
          4179 => x"73",
          4180 => x"38",
          4181 => x"84",
          4182 => x"06",
          4183 => x"77",
          4184 => x"98",
          4185 => x"51",
          4186 => x"3f",
          4187 => x"08",
          4188 => x"81",
          4189 => x"75",
          4190 => x"06",
          4191 => x"55",
          4192 => x"09",
          4193 => x"38",
          4194 => x"ff",
          4195 => x"06",
          4196 => x"55",
          4197 => x"0a",
          4198 => x"aa",
          4199 => x"77",
          4200 => x"c7",
          4201 => x"ac",
          4202 => x"d3",
          4203 => x"96",
          4204 => x"a0",
          4205 => x"51",
          4206 => x"3f",
          4207 => x"0b",
          4208 => x"77",
          4209 => x"bf",
          4210 => x"52",
          4211 => x"51",
          4212 => x"3f",
          4213 => x"18",
          4214 => x"c3",
          4215 => x"53",
          4216 => x"80",
          4217 => x"ff",
          4218 => x"77",
          4219 => x"80",
          4220 => x"7e",
          4221 => x"18",
          4222 => x"c3",
          4223 => x"54",
          4224 => x"15",
          4225 => x"d4",
          4226 => x"e7",
          4227 => x"ac",
          4228 => x"d3",
          4229 => x"38",
          4230 => x"96",
          4231 => x"ae",
          4232 => x"53",
          4233 => x"51",
          4234 => x"63",
          4235 => x"8b",
          4236 => x"54",
          4237 => x"15",
          4238 => x"ff",
          4239 => x"81",
          4240 => x"55",
          4241 => x"53",
          4242 => x"3d",
          4243 => x"ff",
          4244 => x"74",
          4245 => x"0c",
          4246 => x"04",
          4247 => x"a8",
          4248 => x"51",
          4249 => x"82",
          4250 => x"ff",
          4251 => x"a8",
          4252 => x"d1",
          4253 => x"ac",
          4254 => x"d3",
          4255 => x"d7",
          4256 => x"a8",
          4257 => x"a7",
          4258 => x"51",
          4259 => x"81",
          4260 => x"55",
          4261 => x"08",
          4262 => x"02",
          4263 => x"33",
          4264 => x"54",
          4265 => x"83",
          4266 => x"74",
          4267 => x"a0",
          4268 => x"08",
          4269 => x"ff",
          4270 => x"ff",
          4271 => x"ac",
          4272 => x"d4",
          4273 => x"3d",
          4274 => x"ff",
          4275 => x"a9",
          4276 => x"73",
          4277 => x"3f",
          4278 => x"08",
          4279 => x"ac",
          4280 => x"62",
          4281 => x"81",
          4282 => x"84",
          4283 => x"3d",
          4284 => x"38",
          4285 => x"84",
          4286 => x"06",
          4287 => x"a7",
          4288 => x"05",
          4289 => x"3f",
          4290 => x"08",
          4291 => x"ac",
          4292 => x"38",
          4293 => x"53",
          4294 => x"95",
          4295 => x"16",
          4296 => x"ed",
          4297 => x"05",
          4298 => x"34",
          4299 => x"70",
          4300 => x"81",
          4301 => x"57",
          4302 => x"76",
          4303 => x"73",
          4304 => x"77",
          4305 => x"83",
          4306 => x"16",
          4307 => x"2a",
          4308 => x"51",
          4309 => x"80",
          4310 => x"38",
          4311 => x"80",
          4312 => x"52",
          4313 => x"bf",
          4314 => x"d3",
          4315 => x"77",
          4316 => x"b2",
          4317 => x"81",
          4318 => x"80",
          4319 => x"81",
          4320 => x"52",
          4321 => x"ae",
          4322 => x"d3",
          4323 => x"d4",
          4324 => x"81",
          4325 => x"bf",
          4326 => x"33",
          4327 => x"2e",
          4328 => x"92",
          4329 => x"75",
          4330 => x"ff",
          4331 => x"77",
          4332 => x"83",
          4333 => x"9f",
          4334 => x"d4",
          4335 => x"89",
          4336 => x"ac",
          4337 => x"d3",
          4338 => x"38",
          4339 => x"ae",
          4340 => x"d3",
          4341 => x"74",
          4342 => x"0c",
          4343 => x"04",
          4344 => x"02",
          4345 => x"33",
          4346 => x"80",
          4347 => x"57",
          4348 => x"95",
          4349 => x"52",
          4350 => x"cd",
          4351 => x"d3",
          4352 => x"81",
          4353 => x"80",
          4354 => x"5a",
          4355 => x"3d",
          4356 => x"c7",
          4357 => x"d3",
          4358 => x"81",
          4359 => x"bd",
          4360 => x"cf",
          4361 => x"a0",
          4362 => x"80",
          4363 => x"86",
          4364 => x"38",
          4365 => x"61",
          4366 => x"12",
          4367 => x"7a",
          4368 => x"51",
          4369 => x"74",
          4370 => x"78",
          4371 => x"83",
          4372 => x"51",
          4373 => x"3f",
          4374 => x"08",
          4375 => x"d3",
          4376 => x"3d",
          4377 => x"3d",
          4378 => x"82",
          4379 => x"d0",
          4380 => x"3d",
          4381 => x"3f",
          4382 => x"08",
          4383 => x"ac",
          4384 => x"38",
          4385 => x"52",
          4386 => x"05",
          4387 => x"3f",
          4388 => x"08",
          4389 => x"ac",
          4390 => x"02",
          4391 => x"33",
          4392 => x"54",
          4393 => x"83",
          4394 => x"74",
          4395 => x"16",
          4396 => x"22",
          4397 => x"72",
          4398 => x"54",
          4399 => x"51",
          4400 => x"3f",
          4401 => x"0b",
          4402 => x"77",
          4403 => x"a7",
          4404 => x"ac",
          4405 => x"81",
          4406 => x"94",
          4407 => x"ea",
          4408 => x"6b",
          4409 => x"53",
          4410 => x"05",
          4411 => x"51",
          4412 => x"81",
          4413 => x"81",
          4414 => x"30",
          4415 => x"ac",
          4416 => x"25",
          4417 => x"7d",
          4418 => x"72",
          4419 => x"51",
          4420 => x"80",
          4421 => x"38",
          4422 => x"5f",
          4423 => x"3d",
          4424 => x"ff",
          4425 => x"81",
          4426 => x"56",
          4427 => x"08",
          4428 => x"81",
          4429 => x"ff",
          4430 => x"81",
          4431 => x"56",
          4432 => x"08",
          4433 => x"d3",
          4434 => x"d3",
          4435 => x"5c",
          4436 => x"17",
          4437 => x"1a",
          4438 => x"74",
          4439 => x"81",
          4440 => x"77",
          4441 => x"77",
          4442 => x"74",
          4443 => x"2e",
          4444 => x"18",
          4445 => x"33",
          4446 => x"73",
          4447 => x"38",
          4448 => x"09",
          4449 => x"38",
          4450 => x"80",
          4451 => x"70",
          4452 => x"25",
          4453 => x"7e",
          4454 => x"72",
          4455 => x"51",
          4456 => x"2e",
          4457 => x"a0",
          4458 => x"51",
          4459 => x"3f",
          4460 => x"08",
          4461 => x"ac",
          4462 => x"7b",
          4463 => x"54",
          4464 => x"73",
          4465 => x"38",
          4466 => x"73",
          4467 => x"38",
          4468 => x"18",
          4469 => x"ff",
          4470 => x"81",
          4471 => x"7b",
          4472 => x"d3",
          4473 => x"3d",
          4474 => x"3d",
          4475 => x"9a",
          4476 => x"05",
          4477 => x"51",
          4478 => x"81",
          4479 => x"55",
          4480 => x"08",
          4481 => x"8b",
          4482 => x"9a",
          4483 => x"05",
          4484 => x"a1",
          4485 => x"70",
          4486 => x"57",
          4487 => x"74",
          4488 => x"38",
          4489 => x"81",
          4490 => x"81",
          4491 => x"56",
          4492 => x"3f",
          4493 => x"08",
          4494 => x"38",
          4495 => x"70",
          4496 => x"ff",
          4497 => x"81",
          4498 => x"80",
          4499 => x"75",
          4500 => x"07",
          4501 => x"4c",
          4502 => x"80",
          4503 => x"16",
          4504 => x"26",
          4505 => x"16",
          4506 => x"ff",
          4507 => x"80",
          4508 => x"87",
          4509 => x"dc",
          4510 => x"75",
          4511 => x"38",
          4512 => x"bc",
          4513 => x"a6",
          4514 => x"d3",
          4515 => x"38",
          4516 => x"27",
          4517 => x"89",
          4518 => x"8b",
          4519 => x"27",
          4520 => x"55",
          4521 => x"81",
          4522 => x"93",
          4523 => x"77",
          4524 => x"05",
          4525 => x"55",
          4526 => x"34",
          4527 => x"9a",
          4528 => x"ff",
          4529 => x"75",
          4530 => x"17",
          4531 => x"56",
          4532 => x"9f",
          4533 => x"38",
          4534 => x"54",
          4535 => x"81",
          4536 => x"ea",
          4537 => x"2e",
          4538 => x"9f",
          4539 => x"12",
          4540 => x"52",
          4541 => x"a0",
          4542 => x"06",
          4543 => x"17",
          4544 => x"2e",
          4545 => x"15",
          4546 => x"54",
          4547 => x"ee",
          4548 => x"80",
          4549 => x"8f",
          4550 => x"55",
          4551 => x"3f",
          4552 => x"08",
          4553 => x"ac",
          4554 => x"38",
          4555 => x"51",
          4556 => x"3f",
          4557 => x"08",
          4558 => x"ac",
          4559 => x"76",
          4560 => x"38",
          4561 => x"3d",
          4562 => x"52",
          4563 => x"a4",
          4564 => x"39",
          4565 => x"74",
          4566 => x"81",
          4567 => x"34",
          4568 => x"a7",
          4569 => x"d3",
          4570 => x"80",
          4571 => x"d3",
          4572 => x"2e",
          4573 => x"80",
          4574 => x"54",
          4575 => x"80",
          4576 => x"52",
          4577 => x"05",
          4578 => x"b2",
          4579 => x"ac",
          4580 => x"d3",
          4581 => x"38",
          4582 => x"d3",
          4583 => x"65",
          4584 => x"91",
          4585 => x"88",
          4586 => x"34",
          4587 => x"3d",
          4588 => x"52",
          4589 => x"a3",
          4590 => x"54",
          4591 => x"15",
          4592 => x"ff",
          4593 => x"81",
          4594 => x"54",
          4595 => x"81",
          4596 => x"9a",
          4597 => x"f1",
          4598 => x"63",
          4599 => x"80",
          4600 => x"94",
          4601 => x"55",
          4602 => x"5c",
          4603 => x"3f",
          4604 => x"08",
          4605 => x"ac",
          4606 => x"91",
          4607 => x"76",
          4608 => x"38",
          4609 => x"b7",
          4610 => x"2e",
          4611 => x"18",
          4612 => x"90",
          4613 => x"81",
          4614 => x"06",
          4615 => x"73",
          4616 => x"54",
          4617 => x"82",
          4618 => x"39",
          4619 => x"84",
          4620 => x"11",
          4621 => x"2b",
          4622 => x"54",
          4623 => x"fe",
          4624 => x"ff",
          4625 => x"70",
          4626 => x"07",
          4627 => x"d3",
          4628 => x"62",
          4629 => x"5d",
          4630 => x"55",
          4631 => x"79",
          4632 => x"98",
          4633 => x"26",
          4634 => x"59",
          4635 => x"5d",
          4636 => x"52",
          4637 => x"a6",
          4638 => x"d3",
          4639 => x"16",
          4640 => x"56",
          4641 => x"75",
          4642 => x"82",
          4643 => x"2e",
          4644 => x"75",
          4645 => x"94",
          4646 => x"38",
          4647 => x"79",
          4648 => x"38",
          4649 => x"5d",
          4650 => x"79",
          4651 => x"06",
          4652 => x"57",
          4653 => x"38",
          4654 => x"b9",
          4655 => x"57",
          4656 => x"2e",
          4657 => x"15",
          4658 => x"2e",
          4659 => x"83",
          4660 => x"73",
          4661 => x"7f",
          4662 => x"f0",
          4663 => x"ac",
          4664 => x"d3",
          4665 => x"38",
          4666 => x"ff",
          4667 => x"5f",
          4668 => x"84",
          4669 => x"5f",
          4670 => x"38",
          4671 => x"12",
          4672 => x"80",
          4673 => x"7c",
          4674 => x"7a",
          4675 => x"90",
          4676 => x"c0",
          4677 => x"90",
          4678 => x"98",
          4679 => x"05",
          4680 => x"15",
          4681 => x"95",
          4682 => x"08",
          4683 => x"16",
          4684 => x"11",
          4685 => x"55",
          4686 => x"16",
          4687 => x"73",
          4688 => x"0c",
          4689 => x"04",
          4690 => x"6a",
          4691 => x"80",
          4692 => x"9b",
          4693 => x"58",
          4694 => x"3f",
          4695 => x"08",
          4696 => x"80",
          4697 => x"ac",
          4698 => x"d1",
          4699 => x"ac",
          4700 => x"81",
          4701 => x"55",
          4702 => x"2e",
          4703 => x"08",
          4704 => x"34",
          4705 => x"06",
          4706 => x"79",
          4707 => x"cb",
          4708 => x"ac",
          4709 => x"06",
          4710 => x"56",
          4711 => x"74",
          4712 => x"75",
          4713 => x"81",
          4714 => x"8a",
          4715 => x"8d",
          4716 => x"fc",
          4717 => x"52",
          4718 => x"9d",
          4719 => x"d3",
          4720 => x"38",
          4721 => x"93",
          4722 => x"80",
          4723 => x"38",
          4724 => x"67",
          4725 => x"80",
          4726 => x"81",
          4727 => x"5e",
          4728 => x"86",
          4729 => x"26",
          4730 => x"81",
          4731 => x"8b",
          4732 => x"78",
          4733 => x"80",
          4734 => x"93",
          4735 => x"39",
          4736 => x"51",
          4737 => x"3f",
          4738 => x"08",
          4739 => x"6e",
          4740 => x"fe",
          4741 => x"81",
          4742 => x"7e",
          4743 => x"08",
          4744 => x"70",
          4745 => x"25",
          4746 => x"08",
          4747 => x"d3",
          4748 => x"80",
          4749 => x"52",
          4750 => x"46",
          4751 => x"75",
          4752 => x"98",
          4753 => x"53",
          4754 => x"51",
          4755 => x"3f",
          4756 => x"d3",
          4757 => x"e5",
          4758 => x"2a",
          4759 => x"51",
          4760 => x"74",
          4761 => x"81",
          4762 => x"bf",
          4763 => x"63",
          4764 => x"c9",
          4765 => x"31",
          4766 => x"80",
          4767 => x"8a",
          4768 => x"57",
          4769 => x"26",
          4770 => x"7c",
          4771 => x"81",
          4772 => x"74",
          4773 => x"38",
          4774 => x"55",
          4775 => x"88",
          4776 => x"06",
          4777 => x"38",
          4778 => x"39",
          4779 => x"55",
          4780 => x"42",
          4781 => x"8a",
          4782 => x"59",
          4783 => x"09",
          4784 => x"f1",
          4785 => x"38",
          4786 => x"78",
          4787 => x"0b",
          4788 => x"70",
          4789 => x"58",
          4790 => x"80",
          4791 => x"74",
          4792 => x"38",
          4793 => x"10",
          4794 => x"70",
          4795 => x"5a",
          4796 => x"2e",
          4797 => x"75",
          4798 => x"78",
          4799 => x"fe",
          4800 => x"81",
          4801 => x"81",
          4802 => x"10",
          4803 => x"54",
          4804 => x"56",
          4805 => x"3f",
          4806 => x"08",
          4807 => x"80",
          4808 => x"8a",
          4809 => x"fd",
          4810 => x"75",
          4811 => x"38",
          4812 => x"89",
          4813 => x"38",
          4814 => x"78",
          4815 => x"0b",
          4816 => x"70",
          4817 => x"58",
          4818 => x"80",
          4819 => x"74",
          4820 => x"38",
          4821 => x"10",
          4822 => x"70",
          4823 => x"5a",
          4824 => x"2e",
          4825 => x"75",
          4826 => x"78",
          4827 => x"fe",
          4828 => x"81",
          4829 => x"10",
          4830 => x"81",
          4831 => x"9f",
          4832 => x"38",
          4833 => x"d3",
          4834 => x"29",
          4835 => x"2a",
          4836 => x"58",
          4837 => x"76",
          4838 => x"51",
          4839 => x"3f",
          4840 => x"08",
          4841 => x"53",
          4842 => x"80",
          4843 => x"ef",
          4844 => x"ac",
          4845 => x"ff",
          4846 => x"1b",
          4847 => x"05",
          4848 => x"05",
          4849 => x"72",
          4850 => x"52",
          4851 => x"40",
          4852 => x"09",
          4853 => x"38",
          4854 => x"18",
          4855 => x"39",
          4856 => x"78",
          4857 => x"70",
          4858 => x"55",
          4859 => x"87",
          4860 => x"7b",
          4861 => x"79",
          4862 => x"31",
          4863 => x"f2",
          4864 => x"d3",
          4865 => x"61",
          4866 => x"81",
          4867 => x"81",
          4868 => x"83",
          4869 => x"91",
          4870 => x"38",
          4871 => x"58",
          4872 => x"38",
          4873 => x"95",
          4874 => x"2e",
          4875 => x"80",
          4876 => x"ff",
          4877 => x"b4",
          4878 => x"38",
          4879 => x"74",
          4880 => x"86",
          4881 => x"fc",
          4882 => x"81",
          4883 => x"55",
          4884 => x"86",
          4885 => x"fc",
          4886 => x"8b",
          4887 => x"58",
          4888 => x"27",
          4889 => x"8e",
          4890 => x"39",
          4891 => x"26",
          4892 => x"8b",
          4893 => x"58",
          4894 => x"27",
          4895 => x"8e",
          4896 => x"39",
          4897 => x"81",
          4898 => x"06",
          4899 => x"55",
          4900 => x"26",
          4901 => x"8e",
          4902 => x"a1",
          4903 => x"80",
          4904 => x"ff",
          4905 => x"8b",
          4906 => x"98",
          4907 => x"ff",
          4908 => x"7d",
          4909 => x"51",
          4910 => x"3f",
          4911 => x"05",
          4912 => x"ff",
          4913 => x"8e",
          4914 => x"98",
          4915 => x"7f",
          4916 => x"61",
          4917 => x"30",
          4918 => x"84",
          4919 => x"51",
          4920 => x"51",
          4921 => x"3f",
          4922 => x"ff",
          4923 => x"02",
          4924 => x"22",
          4925 => x"51",
          4926 => x"3f",
          4927 => x"52",
          4928 => x"ff",
          4929 => x"f8",
          4930 => x"34",
          4931 => x"1f",
          4932 => x"b0",
          4933 => x"52",
          4934 => x"ff",
          4935 => x"63",
          4936 => x"51",
          4937 => x"3f",
          4938 => x"09",
          4939 => x"cf",
          4940 => x"b2",
          4941 => x"c3",
          4942 => x"98",
          4943 => x"52",
          4944 => x"ff",
          4945 => x"82",
          4946 => x"51",
          4947 => x"3f",
          4948 => x"1f",
          4949 => x"ec",
          4950 => x"b2",
          4951 => x"97",
          4952 => x"80",
          4953 => x"05",
          4954 => x"80",
          4955 => x"93",
          4956 => x"a4",
          4957 => x"1f",
          4958 => x"95",
          4959 => x"82",
          4960 => x"52",
          4961 => x"ff",
          4962 => x"7b",
          4963 => x"06",
          4964 => x"51",
          4965 => x"3f",
          4966 => x"a4",
          4967 => x"7f",
          4968 => x"93",
          4969 => x"b8",
          4970 => x"51",
          4971 => x"3f",
          4972 => x"52",
          4973 => x"51",
          4974 => x"3f",
          4975 => x"53",
          4976 => x"51",
          4977 => x"3f",
          4978 => x"d3",
          4979 => x"ed",
          4980 => x"2e",
          4981 => x"80",
          4982 => x"54",
          4983 => x"53",
          4984 => x"51",
          4985 => x"3f",
          4986 => x"52",
          4987 => x"97",
          4988 => x"8b",
          4989 => x"52",
          4990 => x"96",
          4991 => x"8a",
          4992 => x"52",
          4993 => x"51",
          4994 => x"3f",
          4995 => x"83",
          4996 => x"ff",
          4997 => x"82",
          4998 => x"1f",
          4999 => x"c2",
          5000 => x"d5",
          5001 => x"1f",
          5002 => x"98",
          5003 => x"63",
          5004 => x"7e",
          5005 => x"ff",
          5006 => x"81",
          5007 => x"05",
          5008 => x"79",
          5009 => x"f8",
          5010 => x"80",
          5011 => x"ff",
          5012 => x"7f",
          5013 => x"61",
          5014 => x"81",
          5015 => x"f8",
          5016 => x"ff",
          5017 => x"ff",
          5018 => x"51",
          5019 => x"3f",
          5020 => x"88",
          5021 => x"95",
          5022 => x"39",
          5023 => x"f8",
          5024 => x"2e",
          5025 => x"55",
          5026 => x"51",
          5027 => x"3f",
          5028 => x"57",
          5029 => x"83",
          5030 => x"76",
          5031 => x"7e",
          5032 => x"ff",
          5033 => x"81",
          5034 => x"82",
          5035 => x"53",
          5036 => x"51",
          5037 => x"3f",
          5038 => x"78",
          5039 => x"74",
          5040 => x"1b",
          5041 => x"2e",
          5042 => x"78",
          5043 => x"2e",
          5044 => x"55",
          5045 => x"61",
          5046 => x"74",
          5047 => x"75",
          5048 => x"79",
          5049 => x"d8",
          5050 => x"ac",
          5051 => x"38",
          5052 => x"78",
          5053 => x"74",
          5054 => x"57",
          5055 => x"93",
          5056 => x"65",
          5057 => x"26",
          5058 => x"57",
          5059 => x"83",
          5060 => x"7c",
          5061 => x"06",
          5062 => x"ff",
          5063 => x"77",
          5064 => x"ff",
          5065 => x"82",
          5066 => x"83",
          5067 => x"ff",
          5068 => x"83",
          5069 => x"77",
          5070 => x"0b",
          5071 => x"81",
          5072 => x"34",
          5073 => x"34",
          5074 => x"34",
          5075 => x"57",
          5076 => x"52",
          5077 => x"eb",
          5078 => x"0b",
          5079 => x"81",
          5080 => x"82",
          5081 => x"55",
          5082 => x"34",
          5083 => x"08",
          5084 => x"63",
          5085 => x"1f",
          5086 => x"e6",
          5087 => x"83",
          5088 => x"ff",
          5089 => x"81",
          5090 => x"7e",
          5091 => x"ff",
          5092 => x"81",
          5093 => x"ac",
          5094 => x"80",
          5095 => x"79",
          5096 => x"f6",
          5097 => x"81",
          5098 => x"91",
          5099 => x"8e",
          5100 => x"81",
          5101 => x"81",
          5102 => x"80",
          5103 => x"d3",
          5104 => x"3d",
          5105 => x"3d",
          5106 => x"71",
          5107 => x"e2",
          5108 => x"10",
          5109 => x"05",
          5110 => x"04",
          5111 => x"51",
          5112 => x"3f",
          5113 => x"81",
          5114 => x"ff",
          5115 => x"81",
          5116 => x"c1",
          5117 => x"80",
          5118 => x"be",
          5119 => x"90",
          5120 => x"88",
          5121 => x"39",
          5122 => x"51",
          5123 => x"3f",
          5124 => x"81",
          5125 => x"fe",
          5126 => x"81",
          5127 => x"c2",
          5128 => x"ff",
          5129 => x"92",
          5130 => x"d4",
          5131 => x"dc",
          5132 => x"39",
          5133 => x"51",
          5134 => x"3f",
          5135 => x"81",
          5136 => x"fe",
          5137 => x"80",
          5138 => x"c3",
          5139 => x"ff",
          5140 => x"e6",
          5141 => x"b8",
          5142 => x"b0",
          5143 => x"39",
          5144 => x"51",
          5145 => x"3f",
          5146 => x"81",
          5147 => x"fe",
          5148 => x"80",
          5149 => x"c4",
          5150 => x"ff",
          5151 => x"39",
          5152 => x"51",
          5153 => x"3f",
          5154 => x"c4",
          5155 => x"fe",
          5156 => x"39",
          5157 => x"51",
          5158 => x"3f",
          5159 => x"c4",
          5160 => x"fe",
          5161 => x"39",
          5162 => x"51",
          5163 => x"3f",
          5164 => x"c5",
          5165 => x"fe",
          5166 => x"3d",
          5167 => x"3d",
          5168 => x"56",
          5169 => x"e7",
          5170 => x"74",
          5171 => x"e8",
          5172 => x"e8",
          5173 => x"d3",
          5174 => x"9a",
          5175 => x"52",
          5176 => x"e8",
          5177 => x"d3",
          5178 => x"75",
          5179 => x"af",
          5180 => x"ac",
          5181 => x"54",
          5182 => x"52",
          5183 => x"51",
          5184 => x"3f",
          5185 => x"04",
          5186 => x"0d",
          5187 => x"08",
          5188 => x"08",
          5189 => x"84",
          5190 => x"71",
          5191 => x"75",
          5192 => x"87",
          5193 => x"07",
          5194 => x"5c",
          5195 => x"55",
          5196 => x"38",
          5197 => x"52",
          5198 => x"fb",
          5199 => x"ff",
          5200 => x"81",
          5201 => x"58",
          5202 => x"08",
          5203 => x"d3",
          5204 => x"c0",
          5205 => x"81",
          5206 => x"59",
          5207 => x"fb",
          5208 => x"55",
          5209 => x"76",
          5210 => x"15",
          5211 => x"3f",
          5212 => x"08",
          5213 => x"ac",
          5214 => x"7a",
          5215 => x"38",
          5216 => x"18",
          5217 => x"39",
          5218 => x"fb",
          5219 => x"ca",
          5220 => x"30",
          5221 => x"80",
          5222 => x"70",
          5223 => x"06",
          5224 => x"56",
          5225 => x"90",
          5226 => x"c8",
          5227 => x"98",
          5228 => x"78",
          5229 => x"3f",
          5230 => x"81",
          5231 => x"81",
          5232 => x"04",
          5233 => x"02",
          5234 => x"57",
          5235 => x"59",
          5236 => x"52",
          5237 => x"b0",
          5238 => x"ac",
          5239 => x"76",
          5240 => x"38",
          5241 => x"98",
          5242 => x"61",
          5243 => x"81",
          5244 => x"7f",
          5245 => x"75",
          5246 => x"ac",
          5247 => x"39",
          5248 => x"81",
          5249 => x"8a",
          5250 => x"fb",
          5251 => x"9f",
          5252 => x"c5",
          5253 => x"c5",
          5254 => x"ff",
          5255 => x"81",
          5256 => x"22",
          5257 => x"f9",
          5258 => x"c5",
          5259 => x"c5",
          5260 => x"15",
          5261 => x"c5",
          5262 => x"81",
          5263 => x"80",
          5264 => x"fe",
          5265 => x"87",
          5266 => x"fe",
          5267 => x"c0",
          5268 => x"53",
          5269 => x"3f",
          5270 => x"ee",
          5271 => x"c6",
          5272 => x"f0",
          5273 => x"51",
          5274 => x"3f",
          5275 => x"70",
          5276 => x"52",
          5277 => x"95",
          5278 => x"fe",
          5279 => x"81",
          5280 => x"fe",
          5281 => x"80",
          5282 => x"d0",
          5283 => x"2a",
          5284 => x"51",
          5285 => x"2e",
          5286 => x"51",
          5287 => x"3f",
          5288 => x"51",
          5289 => x"3f",
          5290 => x"ee",
          5291 => x"83",
          5292 => x"06",
          5293 => x"80",
          5294 => x"81",
          5295 => x"9c",
          5296 => x"d4",
          5297 => x"92",
          5298 => x"fe",
          5299 => x"72",
          5300 => x"81",
          5301 => x"71",
          5302 => x"38",
          5303 => x"ed",
          5304 => x"c6",
          5305 => x"ef",
          5306 => x"51",
          5307 => x"3f",
          5308 => x"70",
          5309 => x"52",
          5310 => x"95",
          5311 => x"fe",
          5312 => x"81",
          5313 => x"fe",
          5314 => x"80",
          5315 => x"cc",
          5316 => x"2a",
          5317 => x"51",
          5318 => x"2e",
          5319 => x"51",
          5320 => x"3f",
          5321 => x"51",
          5322 => x"3f",
          5323 => x"ed",
          5324 => x"87",
          5325 => x"06",
          5326 => x"80",
          5327 => x"81",
          5328 => x"98",
          5329 => x"a4",
          5330 => x"8e",
          5331 => x"fe",
          5332 => x"72",
          5333 => x"81",
          5334 => x"71",
          5335 => x"38",
          5336 => x"ec",
          5337 => x"c7",
          5338 => x"ee",
          5339 => x"51",
          5340 => x"3f",
          5341 => x"3f",
          5342 => x"04",
          5343 => x"78",
          5344 => x"55",
          5345 => x"80",
          5346 => x"38",
          5347 => x"77",
          5348 => x"33",
          5349 => x"39",
          5350 => x"80",
          5351 => x"54",
          5352 => x"83",
          5353 => x"72",
          5354 => x"2a",
          5355 => x"53",
          5356 => x"74",
          5357 => x"a0",
          5358 => x"06",
          5359 => x"75",
          5360 => x"57",
          5361 => x"75",
          5362 => x"cb",
          5363 => x"08",
          5364 => x"52",
          5365 => x"d0",
          5366 => x"ac",
          5367 => x"84",
          5368 => x"72",
          5369 => x"a6",
          5370 => x"70",
          5371 => x"57",
          5372 => x"27",
          5373 => x"53",
          5374 => x"ac",
          5375 => x"0d",
          5376 => x"0d",
          5377 => x"f6",
          5378 => x"0c",
          5379 => x"8c",
          5380 => x"7b",
          5381 => x"c3",
          5382 => x"ac",
          5383 => x"06",
          5384 => x"2e",
          5385 => x"9f",
          5386 => x"f8",
          5387 => x"70",
          5388 => x"fd",
          5389 => x"53",
          5390 => x"b0",
          5391 => x"b5",
          5392 => x"d3",
          5393 => x"79",
          5394 => x"38",
          5395 => x"51",
          5396 => x"3f",
          5397 => x"70",
          5398 => x"c8",
          5399 => x"f7",
          5400 => x"3d",
          5401 => x"80",
          5402 => x"5a",
          5403 => x"51",
          5404 => x"3f",
          5405 => x"51",
          5406 => x"3f",
          5407 => x"f8",
          5408 => x"f8",
          5409 => x"ac",
          5410 => x"70",
          5411 => x"59",
          5412 => x"26",
          5413 => x"78",
          5414 => x"b1",
          5415 => x"78",
          5416 => x"3d",
          5417 => x"53",
          5418 => x"51",
          5419 => x"3f",
          5420 => x"08",
          5421 => x"c8",
          5422 => x"fc",
          5423 => x"9a",
          5424 => x"fe",
          5425 => x"fe",
          5426 => x"fe",
          5427 => x"81",
          5428 => x"80",
          5429 => x"81",
          5430 => x"38",
          5431 => x"bf",
          5432 => x"02",
          5433 => x"33",
          5434 => x"ef",
          5435 => x"ac",
          5436 => x"06",
          5437 => x"38",
          5438 => x"51",
          5439 => x"3f",
          5440 => x"d6",
          5441 => x"d8",
          5442 => x"80",
          5443 => x"39",
          5444 => x"f4",
          5445 => x"f8",
          5446 => x"fd",
          5447 => x"d3",
          5448 => x"2e",
          5449 => x"80",
          5450 => x"02",
          5451 => x"33",
          5452 => x"e6",
          5453 => x"ac",
          5454 => x"c8",
          5455 => x"fb",
          5456 => x"96",
          5457 => x"fe",
          5458 => x"fe",
          5459 => x"fe",
          5460 => x"81",
          5461 => x"80",
          5462 => x"60",
          5463 => x"fa",
          5464 => x"fe",
          5465 => x"fe",
          5466 => x"fe",
          5467 => x"81",
          5468 => x"86",
          5469 => x"ac",
          5470 => x"53",
          5471 => x"52",
          5472 => x"52",
          5473 => x"94",
          5474 => x"05",
          5475 => x"52",
          5476 => x"29",
          5477 => x"05",
          5478 => x"d0",
          5479 => x"ac",
          5480 => x"8c",
          5481 => x"ac",
          5482 => x"9a",
          5483 => x"39",
          5484 => x"51",
          5485 => x"3f",
          5486 => x"9e",
          5487 => x"fe",
          5488 => x"fe",
          5489 => x"81",
          5490 => x"b5",
          5491 => x"05",
          5492 => x"e4",
          5493 => x"53",
          5494 => x"08",
          5495 => x"f6",
          5496 => x"d3",
          5497 => x"2e",
          5498 => x"81",
          5499 => x"51",
          5500 => x"fc",
          5501 => x"3d",
          5502 => x"51",
          5503 => x"3f",
          5504 => x"08",
          5505 => x"f8",
          5506 => x"fe",
          5507 => x"81",
          5508 => x"b5",
          5509 => x"05",
          5510 => x"e4",
          5511 => x"d3",
          5512 => x"3d",
          5513 => x"52",
          5514 => x"a3",
          5515 => x"a8",
          5516 => x"e0",
          5517 => x"80",
          5518 => x"ac",
          5519 => x"06",
          5520 => x"79",
          5521 => x"f6",
          5522 => x"d3",
          5523 => x"2e",
          5524 => x"81",
          5525 => x"51",
          5526 => x"fb",
          5527 => x"c8",
          5528 => x"f3",
          5529 => x"51",
          5530 => x"3f",
          5531 => x"81",
          5532 => x"fe",
          5533 => x"a2",
          5534 => x"e2",
          5535 => x"39",
          5536 => x"0b",
          5537 => x"84",
          5538 => x"81",
          5539 => x"94",
          5540 => x"c9",
          5541 => x"f2",
          5542 => x"be",
          5543 => x"c0",
          5544 => x"e8",
          5545 => x"83",
          5546 => x"94",
          5547 => x"80",
          5548 => x"c0",
          5549 => x"fb",
          5550 => x"3d",
          5551 => x"53",
          5552 => x"51",
          5553 => x"3f",
          5554 => x"08",
          5555 => x"8a",
          5556 => x"81",
          5557 => x"fe",
          5558 => x"60",
          5559 => x"b4",
          5560 => x"11",
          5561 => x"05",
          5562 => x"a5",
          5563 => x"ac",
          5564 => x"fa",
          5565 => x"52",
          5566 => x"51",
          5567 => x"3f",
          5568 => x"2d",
          5569 => x"08",
          5570 => x"ac",
          5571 => x"fa",
          5572 => x"d3",
          5573 => x"81",
          5574 => x"fe",
          5575 => x"fa",
          5576 => x"ca",
          5577 => x"f1",
          5578 => x"d1",
          5579 => x"aa",
          5580 => x"c4",
          5581 => x"d4",
          5582 => x"ff",
          5583 => x"ed",
          5584 => x"96",
          5585 => x"33",
          5586 => x"80",
          5587 => x"38",
          5588 => x"59",
          5589 => x"80",
          5590 => x"3d",
          5591 => x"51",
          5592 => x"3f",
          5593 => x"56",
          5594 => x"08",
          5595 => x"dc",
          5596 => x"81",
          5597 => x"a0",
          5598 => x"59",
          5599 => x"3f",
          5600 => x"58",
          5601 => x"57",
          5602 => x"81",
          5603 => x"55",
          5604 => x"80",
          5605 => x"80",
          5606 => x"51",
          5607 => x"81",
          5608 => x"5e",
          5609 => x"7c",
          5610 => x"59",
          5611 => x"7d",
          5612 => x"81",
          5613 => x"38",
          5614 => x"51",
          5615 => x"3f",
          5616 => x"80",
          5617 => x"0b",
          5618 => x"34",
          5619 => x"e4",
          5620 => x"94",
          5621 => x"90",
          5622 => x"87",
          5623 => x"0c",
          5624 => x"0b",
          5625 => x"84",
          5626 => x"83",
          5627 => x"94",
          5628 => x"f4",
          5629 => x"bc",
          5630 => x"0b",
          5631 => x"0c",
          5632 => x"3f",
          5633 => x"3f",
          5634 => x"51",
          5635 => x"3f",
          5636 => x"51",
          5637 => x"3f",
          5638 => x"51",
          5639 => x"3f",
          5640 => x"e7",
          5641 => x"3f",
          5642 => x"00",
          5643 => x"00",
          5644 => x"00",
          5645 => x"00",
          5646 => x"00",
          5647 => x"00",
          5648 => x"00",
          5649 => x"00",
          5650 => x"00",
          5651 => x"00",
          5652 => x"00",
          5653 => x"00",
          5654 => x"00",
          5655 => x"00",
          5656 => x"00",
          5657 => x"00",
          5658 => x"00",
          5659 => x"00",
          5660 => x"00",
          5661 => x"00",
          5662 => x"00",
          5663 => x"00",
          5664 => x"00",
          5665 => x"00",
          5666 => x"00",
          5667 => x"00",
          5668 => x"00",
          5669 => x"00",
          5670 => x"00",
          5671 => x"00",
          5672 => x"00",
          5673 => x"00",
          5674 => x"00",
          5675 => x"00",
          5676 => x"00",
          5677 => x"00",
          5678 => x"00",
          5679 => x"00",
          5680 => x"00",
          5681 => x"00",
          5682 => x"00",
          5683 => x"00",
          5684 => x"00",
          5685 => x"00",
          5686 => x"00",
          5687 => x"00",
          5688 => x"00",
          5689 => x"00",
          5690 => x"00",
          5691 => x"00",
          5692 => x"00",
          5693 => x"00",
          5694 => x"00",
          5695 => x"00",
          5696 => x"00",
          5697 => x"00",
          5698 => x"00",
          5699 => x"00",
          5700 => x"00",
          5701 => x"00",
          5702 => x"00",
          5703 => x"00",
          5704 => x"00",
          5705 => x"00",
          5706 => x"00",
          5707 => x"00",
          5708 => x"00",
          5709 => x"00",
          5710 => x"00",
          5711 => x"00",
          5712 => x"00",
          5713 => x"00",
          5714 => x"00",
          5715 => x"00",
          5716 => x"00",
          5717 => x"00",
          5718 => x"00",
          5719 => x"00",
          5720 => x"00",
          5721 => x"00",
          5722 => x"00",
          5723 => x"00",
          5724 => x"00",
          5725 => x"00",
          5726 => x"00",
          5727 => x"00",
          5728 => x"00",
          5729 => x"00",
          5730 => x"00",
          5731 => x"00",
          5732 => x"00",
          5733 => x"00",
          5734 => x"00",
          5735 => x"00",
          5736 => x"00",
          5737 => x"00",
          5738 => x"00",
          5739 => x"00",
          5740 => x"00",
          5741 => x"00",
          5742 => x"00",
          5743 => x"00",
          5744 => x"00",
          5745 => x"00",
          5746 => x"00",
          5747 => x"00",
          5748 => x"00",
          5749 => x"00",
          5750 => x"00",
          5751 => x"00",
          5752 => x"00",
          5753 => x"00",
          5754 => x"00",
          5755 => x"00",
          5756 => x"00",
          5757 => x"00",
          5758 => x"00",
          5759 => x"00",
          5760 => x"00",
          5761 => x"00",
          5762 => x"00",
          5763 => x"00",
          5764 => x"00",
          5765 => x"00",
          5766 => x"00",
          5767 => x"00",
          5768 => x"00",
          5769 => x"00",
          5770 => x"00",
          5771 => x"00",
          5772 => x"00",
          5773 => x"00",
          5774 => x"00",
          5775 => x"00",
          5776 => x"00",
          5777 => x"00",
          5778 => x"00",
          5779 => x"00",
          5780 => x"00",
          5781 => x"00",
          5782 => x"00",
          5783 => x"00",
          5784 => x"00",
          5785 => x"00",
          5786 => x"00",
          5787 => x"00",
          5788 => x"00",
          5789 => x"00",
          5790 => x"00",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"00",
          5815 => x"00",
          5816 => x"00",
          5817 => x"00",
          5818 => x"00",
          5819 => x"00",
          5820 => x"00",
          5821 => x"00",
          5822 => x"00",
          5823 => x"00",
          5824 => x"00",
          5825 => x"00",
          5826 => x"00",
          5827 => x"64",
          5828 => x"2f",
          5829 => x"25",
          5830 => x"64",
          5831 => x"2e",
          5832 => x"64",
          5833 => x"6f",
          5834 => x"6f",
          5835 => x"67",
          5836 => x"74",
          5837 => x"00",
          5838 => x"28",
          5839 => x"6d",
          5840 => x"43",
          5841 => x"6e",
          5842 => x"29",
          5843 => x"0a",
          5844 => x"69",
          5845 => x"20",
          5846 => x"6c",
          5847 => x"6e",
          5848 => x"3a",
          5849 => x"20",
          5850 => x"4e",
          5851 => x"42",
          5852 => x"20",
          5853 => x"61",
          5854 => x"25",
          5855 => x"2c",
          5856 => x"7a",
          5857 => x"30",
          5858 => x"2e",
          5859 => x"20",
          5860 => x"52",
          5861 => x"28",
          5862 => x"72",
          5863 => x"30",
          5864 => x"20",
          5865 => x"65",
          5866 => x"38",
          5867 => x"0a",
          5868 => x"20",
          5869 => x"41",
          5870 => x"53",
          5871 => x"74",
          5872 => x"38",
          5873 => x"53",
          5874 => x"3d",
          5875 => x"58",
          5876 => x"00",
          5877 => x"20",
          5878 => x"4f",
          5879 => x"0a",
          5880 => x"20",
          5881 => x"53",
          5882 => x"00",
          5883 => x"20",
          5884 => x"50",
          5885 => x"00",
          5886 => x"20",
          5887 => x"44",
          5888 => x"72",
          5889 => x"44",
          5890 => x"63",
          5891 => x"25",
          5892 => x"29",
          5893 => x"00",
          5894 => x"20",
          5895 => x"4e",
          5896 => x"52",
          5897 => x"20",
          5898 => x"54",
          5899 => x"4c",
          5900 => x"00",
          5901 => x"20",
          5902 => x"49",
          5903 => x"31",
          5904 => x"69",
          5905 => x"73",
          5906 => x"31",
          5907 => x"0a",
          5908 => x"64",
          5909 => x"73",
          5910 => x"3a",
          5911 => x"20",
          5912 => x"50",
          5913 => x"65",
          5914 => x"20",
          5915 => x"74",
          5916 => x"41",
          5917 => x"65",
          5918 => x"3d",
          5919 => x"38",
          5920 => x"00",
          5921 => x"20",
          5922 => x"50",
          5923 => x"65",
          5924 => x"79",
          5925 => x"61",
          5926 => x"41",
          5927 => x"65",
          5928 => x"3d",
          5929 => x"38",
          5930 => x"00",
          5931 => x"20",
          5932 => x"74",
          5933 => x"20",
          5934 => x"72",
          5935 => x"64",
          5936 => x"73",
          5937 => x"20",
          5938 => x"3d",
          5939 => x"38",
          5940 => x"00",
          5941 => x"20",
          5942 => x"50",
          5943 => x"64",
          5944 => x"20",
          5945 => x"20",
          5946 => x"20",
          5947 => x"20",
          5948 => x"3d",
          5949 => x"38",
          5950 => x"00",
          5951 => x"20",
          5952 => x"79",
          5953 => x"6d",
          5954 => x"6f",
          5955 => x"46",
          5956 => x"20",
          5957 => x"20",
          5958 => x"3d",
          5959 => x"38",
          5960 => x"00",
          5961 => x"6d",
          5962 => x"00",
          5963 => x"65",
          5964 => x"6d",
          5965 => x"6c",
          5966 => x"00",
          5967 => x"56",
          5968 => x"56",
          5969 => x"6e",
          5970 => x"6e",
          5971 => x"77",
          5972 => x"44",
          5973 => x"2a",
          5974 => x"3b",
          5975 => x"3f",
          5976 => x"7f",
          5977 => x"41",
          5978 => x"41",
          5979 => x"00",
          5980 => x"0a",
          5981 => x"0a",
          5982 => x"0a",
          5983 => x"0a",
          5984 => x"0a",
          5985 => x"0a",
          5986 => x"0a",
          5987 => x"0a",
          5988 => x"0a",
          5989 => x"30",
          5990 => x"fe",
          5991 => x"44",
          5992 => x"2e",
          5993 => x"4f",
          5994 => x"4d",
          5995 => x"20",
          5996 => x"54",
          5997 => x"20",
          5998 => x"4f",
          5999 => x"4d",
          6000 => x"20",
          6001 => x"54",
          6002 => x"20",
          6003 => x"00",
          6004 => x"00",
          6005 => x"00",
          6006 => x"00",
          6007 => x"9a",
          6008 => x"41",
          6009 => x"45",
          6010 => x"49",
          6011 => x"92",
          6012 => x"4f",
          6013 => x"99",
          6014 => x"9d",
          6015 => x"49",
          6016 => x"a5",
          6017 => x"a9",
          6018 => x"ad",
          6019 => x"b1",
          6020 => x"b5",
          6021 => x"b9",
          6022 => x"bd",
          6023 => x"c1",
          6024 => x"c5",
          6025 => x"c9",
          6026 => x"cd",
          6027 => x"d1",
          6028 => x"d5",
          6029 => x"d9",
          6030 => x"dd",
          6031 => x"e1",
          6032 => x"e5",
          6033 => x"e9",
          6034 => x"ed",
          6035 => x"f1",
          6036 => x"f5",
          6037 => x"f9",
          6038 => x"fd",
          6039 => x"2e",
          6040 => x"5b",
          6041 => x"22",
          6042 => x"3e",
          6043 => x"00",
          6044 => x"01",
          6045 => x"10",
          6046 => x"00",
          6047 => x"00",
          6048 => x"01",
          6049 => x"04",
          6050 => x"10",
          6051 => x"00",
          6052 => x"41",
          6053 => x"00",
          6054 => x"41",
          6055 => x"00",
          6056 => x"78",
          6057 => x"00",
          6058 => x"49",
          6059 => x"49",
          6060 => x"4f",
          6061 => x"4f",
          6062 => x"00",
          6063 => x"49",
          6064 => x"42",
          6065 => x"45",
          6066 => x"4f",
          6067 => x"4f",
          6068 => x"00",
          6069 => x"49",
          6070 => x"59",
          6071 => x"4d",
          6072 => x"4e",
          6073 => x"4c",
          6074 => x"45",
          6075 => x"59",
          6076 => x"41",
          6077 => x"41",
          6078 => x"00",
          6079 => x"45",
          6080 => x"4e",
          6081 => x"58",
          6082 => x"54",
          6083 => x"00",
          6084 => x"49",
          6085 => x"43",
          6086 => x"41",
          6087 => x"00",
          6088 => x"64",
          6089 => x"00",
          6090 => x"69",
          6091 => x"00",
          6092 => x"73",
          6093 => x"00",
          6094 => x"69",
          6095 => x"6c",
          6096 => x"64",
          6097 => x"00",
          6098 => x"65",
          6099 => x"00",
          6100 => x"72",
          6101 => x"00",
          6102 => x"77",
          6103 => x"65",
          6104 => x"66",
          6105 => x"00",
          6106 => x"6c",
          6107 => x"00",
          6108 => x"69",
          6109 => x"00",
          6110 => x"6f",
          6111 => x"00",
          6112 => x"63",
          6113 => x"65",
          6114 => x"73",
          6115 => x"00",
          6116 => x"72",
          6117 => x"00",
          6118 => x"69",
          6119 => x"65",
          6120 => x"00",
          6121 => x"77",
          6122 => x"65",
          6123 => x"74",
          6124 => x"63",
          6125 => x"61",
          6126 => x"63",
          6127 => x"61",
          6128 => x"00",
          6129 => x"74",
          6130 => x"00",
          6131 => x"72",
          6132 => x"6d",
          6133 => x"64",
          6134 => x"00",
          6135 => x"6d",
          6136 => x"72",
          6137 => x"73",
          6138 => x"00",
          6139 => x"64",
          6140 => x"00",
          6141 => x"63",
          6142 => x"00",
          6143 => x"63",
          6144 => x"63",
          6145 => x"61",
          6146 => x"78",
          6147 => x"63",
          6148 => x"6c",
          6149 => x"00",
          6150 => x"65",
          6151 => x"00",
          6152 => x"73",
          6153 => x"00",
          6154 => x"64",
          6155 => x"00",
          6156 => x"63",
          6157 => x"64",
          6158 => x"65",
          6159 => x"73",
          6160 => x"64",
          6161 => x"00",
          6162 => x"6c",
          6163 => x"6c",
          6164 => x"6d",
          6165 => x"00",
          6166 => x"63",
          6167 => x"00",
          6168 => x"64",
          6169 => x"00",
          6170 => x"65",
          6171 => x"65",
          6172 => x"65",
          6173 => x"69",
          6174 => x"69",
          6175 => x"72",
          6176 => x"74",
          6177 => x"66",
          6178 => x"66",
          6179 => x"68",
          6180 => x"00",
          6181 => x"6f",
          6182 => x"61",
          6183 => x"00",
          6184 => x"61",
          6185 => x"00",
          6186 => x"6d",
          6187 => x"65",
          6188 => x"72",
          6189 => x"65",
          6190 => x"00",
          6191 => x"65",
          6192 => x"00",
          6193 => x"6e",
          6194 => x"00",
          6195 => x"69",
          6196 => x"00",
          6197 => x"65",
          6198 => x"00",
          6199 => x"69",
          6200 => x"45",
          6201 => x"72",
          6202 => x"6e",
          6203 => x"6e",
          6204 => x"65",
          6205 => x"72",
          6206 => x"00",
          6207 => x"69",
          6208 => x"6e",
          6209 => x"72",
          6210 => x"79",
          6211 => x"00",
          6212 => x"6f",
          6213 => x"6c",
          6214 => x"6f",
          6215 => x"2e",
          6216 => x"6f",
          6217 => x"74",
          6218 => x"6f",
          6219 => x"2e",
          6220 => x"6e",
          6221 => x"69",
          6222 => x"69",
          6223 => x"61",
          6224 => x"0a",
          6225 => x"63",
          6226 => x"73",
          6227 => x"6e",
          6228 => x"2e",
          6229 => x"69",
          6230 => x"61",
          6231 => x"61",
          6232 => x"65",
          6233 => x"74",
          6234 => x"00",
          6235 => x"69",
          6236 => x"68",
          6237 => x"6c",
          6238 => x"6e",
          6239 => x"69",
          6240 => x"00",
          6241 => x"44",
          6242 => x"20",
          6243 => x"74",
          6244 => x"72",
          6245 => x"63",
          6246 => x"2e",
          6247 => x"72",
          6248 => x"20",
          6249 => x"62",
          6250 => x"69",
          6251 => x"6e",
          6252 => x"69",
          6253 => x"00",
          6254 => x"69",
          6255 => x"6e",
          6256 => x"65",
          6257 => x"6c",
          6258 => x"0a",
          6259 => x"6f",
          6260 => x"6d",
          6261 => x"69",
          6262 => x"20",
          6263 => x"65",
          6264 => x"74",
          6265 => x"66",
          6266 => x"64",
          6267 => x"20",
          6268 => x"6b",
          6269 => x"00",
          6270 => x"6f",
          6271 => x"74",
          6272 => x"6f",
          6273 => x"64",
          6274 => x"00",
          6275 => x"69",
          6276 => x"75",
          6277 => x"6f",
          6278 => x"61",
          6279 => x"6e",
          6280 => x"6e",
          6281 => x"6c",
          6282 => x"0a",
          6283 => x"69",
          6284 => x"69",
          6285 => x"6f",
          6286 => x"64",
          6287 => x"00",
          6288 => x"6e",
          6289 => x"66",
          6290 => x"65",
          6291 => x"6d",
          6292 => x"72",
          6293 => x"00",
          6294 => x"6f",
          6295 => x"61",
          6296 => x"6f",
          6297 => x"20",
          6298 => x"65",
          6299 => x"00",
          6300 => x"61",
          6301 => x"65",
          6302 => x"73",
          6303 => x"63",
          6304 => x"65",
          6305 => x"0a",
          6306 => x"75",
          6307 => x"73",
          6308 => x"00",
          6309 => x"6e",
          6310 => x"77",
          6311 => x"72",
          6312 => x"2e",
          6313 => x"25",
          6314 => x"62",
          6315 => x"73",
          6316 => x"20",
          6317 => x"25",
          6318 => x"62",
          6319 => x"73",
          6320 => x"63",
          6321 => x"00",
          6322 => x"65",
          6323 => x"00",
          6324 => x"50",
          6325 => x"00",
          6326 => x"2a",
          6327 => x"73",
          6328 => x"00",
          6329 => x"38",
          6330 => x"2f",
          6331 => x"39",
          6332 => x"31",
          6333 => x"00",
          6334 => x"5a",
          6335 => x"20",
          6336 => x"20",
          6337 => x"78",
          6338 => x"73",
          6339 => x"20",
          6340 => x"0a",
          6341 => x"50",
          6342 => x"20",
          6343 => x"65",
          6344 => x"70",
          6345 => x"61",
          6346 => x"65",
          6347 => x"00",
          6348 => x"69",
          6349 => x"20",
          6350 => x"65",
          6351 => x"70",
          6352 => x"00",
          6353 => x"53",
          6354 => x"6e",
          6355 => x"72",
          6356 => x"0a",
          6357 => x"4f",
          6358 => x"20",
          6359 => x"69",
          6360 => x"72",
          6361 => x"74",
          6362 => x"4f",
          6363 => x"20",
          6364 => x"69",
          6365 => x"72",
          6366 => x"74",
          6367 => x"41",
          6368 => x"20",
          6369 => x"69",
          6370 => x"72",
          6371 => x"74",
          6372 => x"41",
          6373 => x"20",
          6374 => x"69",
          6375 => x"72",
          6376 => x"74",
          6377 => x"41",
          6378 => x"20",
          6379 => x"69",
          6380 => x"72",
          6381 => x"74",
          6382 => x"41",
          6383 => x"20",
          6384 => x"69",
          6385 => x"72",
          6386 => x"74",
          6387 => x"65",
          6388 => x"6e",
          6389 => x"70",
          6390 => x"6d",
          6391 => x"2e",
          6392 => x"00",
          6393 => x"6e",
          6394 => x"69",
          6395 => x"74",
          6396 => x"72",
          6397 => x"0a",
          6398 => x"3a",
          6399 => x"61",
          6400 => x"64",
          6401 => x"20",
          6402 => x"74",
          6403 => x"69",
          6404 => x"73",
          6405 => x"61",
          6406 => x"30",
          6407 => x"6c",
          6408 => x"65",
          6409 => x"69",
          6410 => x"61",
          6411 => x"6c",
          6412 => x"0a",
          6413 => x"20",
          6414 => x"61",
          6415 => x"69",
          6416 => x"69",
          6417 => x"00",
          6418 => x"6e",
          6419 => x"61",
          6420 => x"65",
          6421 => x"00",
          6422 => x"61",
          6423 => x"64",
          6424 => x"20",
          6425 => x"74",
          6426 => x"69",
          6427 => x"0a",
          6428 => x"63",
          6429 => x"0a",
          6430 => x"75",
          6431 => x"69",
          6432 => x"6c",
          6433 => x"20",
          6434 => x"65",
          6435 => x"70",
          6436 => x"00",
          6437 => x"6e",
          6438 => x"69",
          6439 => x"69",
          6440 => x"72",
          6441 => x"74",
          6442 => x"00",
          6443 => x"69",
          6444 => x"6c",
          6445 => x"75",
          6446 => x"20",
          6447 => x"6f",
          6448 => x"6e",
          6449 => x"69",
          6450 => x"75",
          6451 => x"20",
          6452 => x"6f",
          6453 => x"78",
          6454 => x"74",
          6455 => x"20",
          6456 => x"65",
          6457 => x"25",
          6458 => x"20",
          6459 => x"0a",
          6460 => x"61",
          6461 => x"6e",
          6462 => x"6f",
          6463 => x"40",
          6464 => x"38",
          6465 => x"2e",
          6466 => x"00",
          6467 => x"61",
          6468 => x"72",
          6469 => x"72",
          6470 => x"20",
          6471 => x"65",
          6472 => x"64",
          6473 => x"00",
          6474 => x"65",
          6475 => x"72",
          6476 => x"67",
          6477 => x"70",
          6478 => x"61",
          6479 => x"6e",
          6480 => x"0a",
          6481 => x"6f",
          6482 => x"72",
          6483 => x"6f",
          6484 => x"67",
          6485 => x"0a",
          6486 => x"50",
          6487 => x"69",
          6488 => x"64",
          6489 => x"73",
          6490 => x"2e",
          6491 => x"00",
          6492 => x"61",
          6493 => x"6f",
          6494 => x"6e",
          6495 => x"00",
          6496 => x"75",
          6497 => x"6e",
          6498 => x"2e",
          6499 => x"6e",
          6500 => x"69",
          6501 => x"69",
          6502 => x"72",
          6503 => x"74",
          6504 => x"2e",
          6505 => x"00",
          6506 => x"00",
          6507 => x"00",
          6508 => x"00",
          6509 => x"00",
          6510 => x"01",
          6511 => x"00",
          6512 => x"00",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"f5",
          6517 => x"01",
          6518 => x"01",
          6519 => x"01",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"00",
          6524 => x"01",
          6525 => x"00",
          6526 => x"00",
          6527 => x"00",
          6528 => x"02",
          6529 => x"00",
          6530 => x"00",
          6531 => x"00",
          6532 => x"03",
          6533 => x"00",
          6534 => x"00",
          6535 => x"00",
          6536 => x"04",
          6537 => x"00",
          6538 => x"00",
          6539 => x"00",
          6540 => x"0a",
          6541 => x"00",
          6542 => x"00",
          6543 => x"00",
          6544 => x"0b",
          6545 => x"00",
          6546 => x"00",
          6547 => x"00",
          6548 => x"0c",
          6549 => x"00",
          6550 => x"00",
          6551 => x"00",
          6552 => x"0d",
          6553 => x"00",
          6554 => x"00",
          6555 => x"00",
          6556 => x"0e",
          6557 => x"00",
          6558 => x"00",
          6559 => x"00",
          6560 => x"0f",
          6561 => x"00",
          6562 => x"00",
          6563 => x"00",
          6564 => x"14",
          6565 => x"00",
          6566 => x"00",
          6567 => x"00",
          6568 => x"17",
          6569 => x"00",
          6570 => x"00",
          6571 => x"00",
          6572 => x"18",
          6573 => x"00",
          6574 => x"00",
          6575 => x"00",
          6576 => x"19",
          6577 => x"00",
          6578 => x"00",
          6579 => x"00",
          6580 => x"1a",
          6581 => x"00",
          6582 => x"00",
          6583 => x"00",
          6584 => x"1c",
          6585 => x"00",
          6586 => x"00",
          6587 => x"00",
          6588 => x"1d",
          6589 => x"00",
          6590 => x"00",
          6591 => x"00",
          6592 => x"1e",
          6593 => x"00",
          6594 => x"00",
          6595 => x"00",
          6596 => x"22",
          6597 => x"00",
          6598 => x"00",
          6599 => x"00",
          6600 => x"23",
          6601 => x"00",
          6602 => x"00",
          6603 => x"00",
          6604 => x"24",
          6605 => x"00",
          6606 => x"00",
          6607 => x"00",
          6608 => x"1f",
          6609 => x"00",
          6610 => x"00",
          6611 => x"00",
          6612 => x"20",
          6613 => x"00",
          6614 => x"00",
          6615 => x"00",
          6616 => x"21",
          6617 => x"00",
          6618 => x"00",
          6619 => x"00",
          6620 => x"15",
          6621 => x"00",
          6622 => x"00",
          6623 => x"00",
          6624 => x"16",
          6625 => x"00",
          6626 => x"00",
          6627 => x"00",
          6628 => x"1b",
          6629 => x"00",
          6630 => x"00",
          6631 => x"00",
          6632 => x"25",
          6633 => x"00",
          6634 => x"00",
          6635 => x"00",
          6636 => x"2d",
          6637 => x"00",
          6638 => x"00",
          6639 => x"00",
          6640 => x"2e",
          6641 => x"00",
          6642 => x"00",
          6643 => x"00",
          6644 => x"2b",
          6645 => x"00",
          6646 => x"00",
          6647 => x"00",
          6648 => x"30",
          6649 => x"00",
          6650 => x"00",
          6651 => x"00",
          6652 => x"2f",
          6653 => x"00",
          6654 => x"00",
          6655 => x"00",
          6656 => x"2c",
          6657 => x"00",
          6658 => x"00",
          6659 => x"00",
          6660 => x"26",
          6661 => x"00",
          6662 => x"00",
          6663 => x"00",
          6664 => x"27",
          6665 => x"00",
          6666 => x"00",
          6667 => x"00",
          6668 => x"28",
          6669 => x"00",
          6670 => x"00",
          6671 => x"00",
          6672 => x"29",
          6673 => x"00",
          6674 => x"00",
          6675 => x"00",
          6676 => x"2a",
          6677 => x"00",
          6678 => x"00",
          6679 => x"00",
          6680 => x"3c",
          6681 => x"00",
          6682 => x"00",
          6683 => x"00",
          6684 => x"3d",
          6685 => x"00",
          6686 => x"00",
          6687 => x"00",
          6688 => x"3e",
          6689 => x"00",
          6690 => x"00",
          6691 => x"00",
          6692 => x"3f",
          6693 => x"00",
          6694 => x"00",
          6695 => x"00",
          6696 => x"40",
          6697 => x"00",
          6698 => x"00",
          6699 => x"00",
          6700 => x"50",
          6701 => x"00",
          6702 => x"00",
          6703 => x"00",
          6704 => x"51",
          6705 => x"00",
          6706 => x"00",
          6707 => x"00",
          6708 => x"52",
          6709 => x"00",
          6710 => x"00",
          6711 => x"00",
          6712 => x"53",
          6713 => x"00",
          6714 => x"00",
          6715 => x"00",
          6716 => x"54",
          6717 => x"00",
          6718 => x"00",
          6719 => x"00",
          6720 => x"55",
          6721 => x"00",
          6722 => x"00",
          6723 => x"00",
          6724 => x"64",
          6725 => x"00",
          6726 => x"00",
          6727 => x"00",
          6728 => x"65",
          6729 => x"00",
          6730 => x"00",
          6731 => x"00",
          6732 => x"79",
          6733 => x"00",
          6734 => x"00",
          6735 => x"00",
          6736 => x"78",
          6737 => x"00",
          6738 => x"00",
          6739 => x"00",
          6740 => x"82",
          6741 => x"00",
          6742 => x"00",
          6743 => x"00",
          6744 => x"83",
          6745 => x"00",
          6746 => x"00",
          6747 => x"00",
          6748 => x"84",
          6749 => x"00",
          6750 => x"00",
          6751 => x"00",
          6752 => x"85",
          6753 => x"00",
          6754 => x"00",
          6755 => x"00",
          6756 => x"86",
          6757 => x"00",
          6758 => x"00",
          6759 => x"00",
          6760 => x"87",
          6761 => x"00",
          6762 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"0b",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"0b",
            11 => x"0b",
            12 => x"93",
            13 => x"0b",
            14 => x"0b",
            15 => x"b1",
            16 => x"0b",
            17 => x"0b",
            18 => x"cf",
            19 => x"0b",
            20 => x"0b",
            21 => x"ed",
            22 => x"0b",
            23 => x"0b",
            24 => x"8b",
            25 => x"0b",
            26 => x"0b",
            27 => x"a9",
            28 => x"0b",
            29 => x"0b",
            30 => x"c7",
            31 => x"0b",
            32 => x"0b",
            33 => x"e5",
            34 => x"0b",
            35 => x"0b",
            36 => x"83",
            37 => x"0b",
            38 => x"0b",
            39 => x"a3",
            40 => x"0b",
            41 => x"0b",
            42 => x"c3",
            43 => x"0b",
            44 => x"0b",
            45 => x"e3",
            46 => x"0b",
            47 => x"0b",
            48 => x"83",
            49 => x"0b",
            50 => x"0b",
            51 => x"a3",
            52 => x"0b",
            53 => x"0b",
            54 => x"c3",
            55 => x"0b",
            56 => x"0b",
            57 => x"e3",
            58 => x"0b",
            59 => x"0b",
            60 => x"83",
            61 => x"0b",
            62 => x"0b",
            63 => x"a3",
            64 => x"0b",
            65 => x"0b",
            66 => x"c3",
            67 => x"0b",
            68 => x"0b",
            69 => x"e3",
            70 => x"0b",
            71 => x"0b",
            72 => x"83",
            73 => x"0b",
            74 => x"0b",
            75 => x"a2",
            76 => x"0b",
            77 => x"0b",
            78 => x"c0",
            79 => x"0b",
            80 => x"0b",
            81 => x"de",
            82 => x"0b",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"81",
           130 => x"94",
           131 => x"d3",
           132 => x"80",
           133 => x"d3",
           134 => x"a7",
           135 => x"b8",
           136 => x"90",
           137 => x"b8",
           138 => x"2d",
           139 => x"08",
           140 => x"04",
           141 => x"0c",
           142 => x"81",
           143 => x"83",
           144 => x"81",
           145 => x"a6",
           146 => x"d3",
           147 => x"80",
           148 => x"d3",
           149 => x"f2",
           150 => x"b8",
           151 => x"90",
           152 => x"b8",
           153 => x"2d",
           154 => x"08",
           155 => x"04",
           156 => x"0c",
           157 => x"81",
           158 => x"83",
           159 => x"81",
           160 => x"aa",
           161 => x"d3",
           162 => x"80",
           163 => x"d3",
           164 => x"84",
           165 => x"b8",
           166 => x"90",
           167 => x"b8",
           168 => x"2d",
           169 => x"08",
           170 => x"04",
           171 => x"0c",
           172 => x"81",
           173 => x"83",
           174 => x"81",
           175 => x"96",
           176 => x"d3",
           177 => x"80",
           178 => x"d3",
           179 => x"b5",
           180 => x"b8",
           181 => x"90",
           182 => x"b8",
           183 => x"2d",
           184 => x"08",
           185 => x"04",
           186 => x"0c",
           187 => x"81",
           188 => x"83",
           189 => x"81",
           190 => x"92",
           191 => x"d3",
           192 => x"80",
           193 => x"d3",
           194 => x"de",
           195 => x"d3",
           196 => x"80",
           197 => x"d3",
           198 => x"ed",
           199 => x"d3",
           200 => x"80",
           201 => x"d3",
           202 => x"e3",
           203 => x"d3",
           204 => x"80",
           205 => x"d3",
           206 => x"e7",
           207 => x"d3",
           208 => x"80",
           209 => x"d3",
           210 => x"f2",
           211 => x"d3",
           212 => x"80",
           213 => x"d3",
           214 => x"fc",
           215 => x"d3",
           216 => x"80",
           217 => x"d3",
           218 => x"ec",
           219 => x"d3",
           220 => x"80",
           221 => x"d3",
           222 => x"f7",
           223 => x"d3",
           224 => x"80",
           225 => x"d3",
           226 => x"f8",
           227 => x"d3",
           228 => x"80",
           229 => x"d3",
           230 => x"f8",
           231 => x"d3",
           232 => x"80",
           233 => x"d3",
           234 => x"82",
           235 => x"d3",
           236 => x"80",
           237 => x"d3",
           238 => x"fe",
           239 => x"d3",
           240 => x"80",
           241 => x"d3",
           242 => x"84",
           243 => x"d3",
           244 => x"80",
           245 => x"d3",
           246 => x"f9",
           247 => x"d3",
           248 => x"80",
           249 => x"d3",
           250 => x"87",
           251 => x"d3",
           252 => x"80",
           253 => x"d3",
           254 => x"88",
           255 => x"d3",
           256 => x"80",
           257 => x"d3",
           258 => x"ee",
           259 => x"d3",
           260 => x"80",
           261 => x"d3",
           262 => x"ee",
           263 => x"d3",
           264 => x"80",
           265 => x"d3",
           266 => x"ef",
           267 => x"d3",
           268 => x"80",
           269 => x"d3",
           270 => x"fa",
           271 => x"d3",
           272 => x"80",
           273 => x"d3",
           274 => x"89",
           275 => x"d3",
           276 => x"80",
           277 => x"d3",
           278 => x"8b",
           279 => x"d3",
           280 => x"80",
           281 => x"d3",
           282 => x"8f",
           283 => x"d3",
           284 => x"80",
           285 => x"d3",
           286 => x"dd",
           287 => x"d3",
           288 => x"80",
           289 => x"d3",
           290 => x"92",
           291 => x"d3",
           292 => x"80",
           293 => x"d3",
           294 => x"e5",
           295 => x"b8",
           296 => x"90",
           297 => x"b8",
           298 => x"2d",
           299 => x"08",
           300 => x"04",
           301 => x"0c",
           302 => x"81",
           303 => x"83",
           304 => x"81",
           305 => x"8f",
           306 => x"d3",
           307 => x"80",
           308 => x"d3",
           309 => x"cd",
           310 => x"b8",
           311 => x"90",
           312 => x"b8",
           313 => x"2d",
           314 => x"08",
           315 => x"04",
           316 => x"0c",
           317 => x"2d",
           318 => x"08",
           319 => x"04",
           320 => x"70",
           321 => x"27",
           322 => x"71",
           323 => x"53",
           324 => x"0b",
           325 => x"84",
           326 => x"af",
           327 => x"04",
           328 => x"08",
           329 => x"b8",
           330 => x"0d",
           331 => x"d3",
           332 => x"05",
           333 => x"d3",
           334 => x"05",
           335 => x"c5",
           336 => x"ac",
           337 => x"d3",
           338 => x"85",
           339 => x"d3",
           340 => x"81",
           341 => x"02",
           342 => x"0c",
           343 => x"81",
           344 => x"b8",
           345 => x"08",
           346 => x"b8",
           347 => x"08",
           348 => x"81",
           349 => x"70",
           350 => x"0c",
           351 => x"0d",
           352 => x"0c",
           353 => x"b8",
           354 => x"d3",
           355 => x"3d",
           356 => x"81",
           357 => x"fc",
           358 => x"0b",
           359 => x"08",
           360 => x"81",
           361 => x"8c",
           362 => x"d3",
           363 => x"05",
           364 => x"38",
           365 => x"08",
           366 => x"80",
           367 => x"80",
           368 => x"b8",
           369 => x"08",
           370 => x"81",
           371 => x"8c",
           372 => x"81",
           373 => x"8c",
           374 => x"d3",
           375 => x"05",
           376 => x"d3",
           377 => x"05",
           378 => x"39",
           379 => x"08",
           380 => x"80",
           381 => x"38",
           382 => x"08",
           383 => x"81",
           384 => x"88",
           385 => x"ad",
           386 => x"b8",
           387 => x"08",
           388 => x"08",
           389 => x"31",
           390 => x"08",
           391 => x"81",
           392 => x"f8",
           393 => x"d3",
           394 => x"05",
           395 => x"d3",
           396 => x"05",
           397 => x"b8",
           398 => x"08",
           399 => x"d3",
           400 => x"05",
           401 => x"b8",
           402 => x"08",
           403 => x"d3",
           404 => x"05",
           405 => x"39",
           406 => x"08",
           407 => x"80",
           408 => x"81",
           409 => x"88",
           410 => x"81",
           411 => x"f4",
           412 => x"91",
           413 => x"b8",
           414 => x"08",
           415 => x"b8",
           416 => x"0c",
           417 => x"b8",
           418 => x"08",
           419 => x"0c",
           420 => x"81",
           421 => x"04",
           422 => x"76",
           423 => x"8c",
           424 => x"33",
           425 => x"55",
           426 => x"8a",
           427 => x"06",
           428 => x"2e",
           429 => x"12",
           430 => x"2e",
           431 => x"73",
           432 => x"55",
           433 => x"52",
           434 => x"09",
           435 => x"38",
           436 => x"ac",
           437 => x"0d",
           438 => x"88",
           439 => x"70",
           440 => x"07",
           441 => x"8f",
           442 => x"38",
           443 => x"84",
           444 => x"72",
           445 => x"05",
           446 => x"71",
           447 => x"53",
           448 => x"70",
           449 => x"0c",
           450 => x"71",
           451 => x"38",
           452 => x"90",
           453 => x"70",
           454 => x"0c",
           455 => x"71",
           456 => x"38",
           457 => x"8e",
           458 => x"0d",
           459 => x"72",
           460 => x"53",
           461 => x"93",
           462 => x"73",
           463 => x"54",
           464 => x"2e",
           465 => x"73",
           466 => x"71",
           467 => x"ff",
           468 => x"70",
           469 => x"38",
           470 => x"70",
           471 => x"81",
           472 => x"81",
           473 => x"71",
           474 => x"ff",
           475 => x"54",
           476 => x"38",
           477 => x"73",
           478 => x"75",
           479 => x"71",
           480 => x"d3",
           481 => x"52",
           482 => x"04",
           483 => x"f7",
           484 => x"14",
           485 => x"84",
           486 => x"06",
           487 => x"70",
           488 => x"14",
           489 => x"08",
           490 => x"71",
           491 => x"dc",
           492 => x"54",
           493 => x"39",
           494 => x"d3",
           495 => x"3d",
           496 => x"3d",
           497 => x"54",
           498 => x"2b",
           499 => x"3f",
           500 => x"08",
           501 => x"72",
           502 => x"54",
           503 => x"25",
           504 => x"81",
           505 => x"84",
           506 => x"fc",
           507 => x"70",
           508 => x"55",
           509 => x"2e",
           510 => x"73",
           511 => x"a0",
           512 => x"06",
           513 => x"14",
           514 => x"54",
           515 => x"f6",
           516 => x"84",
           517 => x"52",
           518 => x"52",
           519 => x"2e",
           520 => x"53",
           521 => x"9f",
           522 => x"51",
           523 => x"38",
           524 => x"70",
           525 => x"81",
           526 => x"80",
           527 => x"05",
           528 => x"75",
           529 => x"70",
           530 => x"0c",
           531 => x"04",
           532 => x"76",
           533 => x"80",
           534 => x"86",
           535 => x"52",
           536 => x"c4",
           537 => x"ac",
           538 => x"80",
           539 => x"74",
           540 => x"d3",
           541 => x"3d",
           542 => x"3d",
           543 => x"11",
           544 => x"5b",
           545 => x"79",
           546 => x"bf",
           547 => x"33",
           548 => x"82",
           549 => x"26",
           550 => x"84",
           551 => x"83",
           552 => x"26",
           553 => x"85",
           554 => x"84",
           555 => x"26",
           556 => x"86",
           557 => x"85",
           558 => x"26",
           559 => x"88",
           560 => x"86",
           561 => x"e7",
           562 => x"38",
           563 => x"5a",
           564 => x"87",
           565 => x"f3",
           566 => x"22",
           567 => x"22",
           568 => x"33",
           569 => x"33",
           570 => x"33",
           571 => x"33",
           572 => x"33",
           573 => x"52",
           574 => x"51",
           575 => x"87",
           576 => x"5b",
           577 => x"7b",
           578 => x"98",
           579 => x"1c",
           580 => x"98",
           581 => x"1c",
           582 => x"98",
           583 => x"1c",
           584 => x"98",
           585 => x"1c",
           586 => x"98",
           587 => x"1c",
           588 => x"98",
           589 => x"1c",
           590 => x"98",
           591 => x"1c",
           592 => x"98",
           593 => x"7b",
           594 => x"7a",
           595 => x"0c",
           596 => x"04",
           597 => x"7d",
           598 => x"98",
           599 => x"7c",
           600 => x"98",
           601 => x"7a",
           602 => x"c0",
           603 => x"5b",
           604 => x"34",
           605 => x"b4",
           606 => x"83",
           607 => x"c0",
           608 => x"5b",
           609 => x"34",
           610 => x"ac",
           611 => x"85",
           612 => x"c0",
           613 => x"5b",
           614 => x"34",
           615 => x"a4",
           616 => x"88",
           617 => x"c0",
           618 => x"5b",
           619 => x"23",
           620 => x"8a",
           621 => x"88",
           622 => x"86",
           623 => x"85",
           624 => x"84",
           625 => x"83",
           626 => x"82",
           627 => x"79",
           628 => x"b6",
           629 => x"af",
           630 => x"0d",
           631 => x"0d",
           632 => x"33",
           633 => x"9f",
           634 => x"51",
           635 => x"81",
           636 => x"82",
           637 => x"fd",
           638 => x"0b",
           639 => x"a4",
           640 => x"87",
           641 => x"51",
           642 => x"86",
           643 => x"94",
           644 => x"08",
           645 => x"70",
           646 => x"52",
           647 => x"2e",
           648 => x"91",
           649 => x"06",
           650 => x"d7",
           651 => x"2a",
           652 => x"81",
           653 => x"70",
           654 => x"38",
           655 => x"70",
           656 => x"51",
           657 => x"38",
           658 => x"cb",
           659 => x"87",
           660 => x"52",
           661 => x"86",
           662 => x"94",
           663 => x"72",
           664 => x"d3",
           665 => x"3d",
           666 => x"3d",
           667 => x"05",
           668 => x"81",
           669 => x"54",
           670 => x"94",
           671 => x"80",
           672 => x"87",
           673 => x"51",
           674 => x"96",
           675 => x"06",
           676 => x"70",
           677 => x"38",
           678 => x"70",
           679 => x"51",
           680 => x"71",
           681 => x"32",
           682 => x"51",
           683 => x"2e",
           684 => x"93",
           685 => x"06",
           686 => x"ff",
           687 => x"0b",
           688 => x"33",
           689 => x"94",
           690 => x"80",
           691 => x"87",
           692 => x"52",
           693 => x"85",
           694 => x"fb",
           695 => x"54",
           696 => x"52",
           697 => x"2e",
           698 => x"73",
           699 => x"55",
           700 => x"81",
           701 => x"54",
           702 => x"94",
           703 => x"80",
           704 => x"87",
           705 => x"51",
           706 => x"96",
           707 => x"06",
           708 => x"70",
           709 => x"38",
           710 => x"70",
           711 => x"51",
           712 => x"71",
           713 => x"32",
           714 => x"51",
           715 => x"2e",
           716 => x"93",
           717 => x"06",
           718 => x"ff",
           719 => x"0b",
           720 => x"33",
           721 => x"94",
           722 => x"80",
           723 => x"87",
           724 => x"52",
           725 => x"81",
           726 => x"52",
           727 => x"8b",
           728 => x"d3",
           729 => x"3d",
           730 => x"3d",
           731 => x"81",
           732 => x"52",
           733 => x"84",
           734 => x"2e",
           735 => x"c0",
           736 => x"70",
           737 => x"2a",
           738 => x"51",
           739 => x"80",
           740 => x"0b",
           741 => x"a4",
           742 => x"c0",
           743 => x"70",
           744 => x"38",
           745 => x"90",
           746 => x"70",
           747 => x"81",
           748 => x"51",
           749 => x"04",
           750 => x"0b",
           751 => x"a4",
           752 => x"c0",
           753 => x"70",
           754 => x"38",
           755 => x"94",
           756 => x"70",
           757 => x"81",
           758 => x"51",
           759 => x"80",
           760 => x"0b",
           761 => x"a4",
           762 => x"c0",
           763 => x"70",
           764 => x"38",
           765 => x"90",
           766 => x"70",
           767 => x"98",
           768 => x"51",
           769 => x"ac",
           770 => x"0d",
           771 => x"0d",
           772 => x"80",
           773 => x"9c",
           774 => x"51",
           775 => x"80",
           776 => x"38",
           777 => x"0b",
           778 => x"9c",
           779 => x"84",
           780 => x"9e",
           781 => x"0c",
           782 => x"87",
           783 => x"08",
           784 => x"8c",
           785 => x"9e",
           786 => x"0c",
           787 => x"87",
           788 => x"08",
           789 => x"94",
           790 => x"9e",
           791 => x"0c",
           792 => x"87",
           793 => x"08",
           794 => x"9c",
           795 => x"9e",
           796 => x"0c",
           797 => x"87",
           798 => x"08",
           799 => x"73",
           800 => x"70",
           801 => x"a8",
           802 => x"9e",
           803 => x"0c",
           804 => x"ac",
           805 => x"12",
           806 => x"87",
           807 => x"08",
           808 => x"06",
           809 => x"70",
           810 => x"38",
           811 => x"72",
           812 => x"87",
           813 => x"08",
           814 => x"80",
           815 => x"52",
           816 => x"83",
           817 => x"71",
           818 => x"34",
           819 => x"c0",
           820 => x"70",
           821 => x"06",
           822 => x"70",
           823 => x"38",
           824 => x"81",
           825 => x"80",
           826 => x"9e",
           827 => x"90",
           828 => x"52",
           829 => x"2e",
           830 => x"52",
           831 => x"d8",
           832 => x"87",
           833 => x"08",
           834 => x"06",
           835 => x"70",
           836 => x"38",
           837 => x"81",
           838 => x"80",
           839 => x"9e",
           840 => x"84",
           841 => x"52",
           842 => x"2e",
           843 => x"52",
           844 => x"da",
           845 => x"87",
           846 => x"08",
           847 => x"06",
           848 => x"70",
           849 => x"38",
           850 => x"81",
           851 => x"80",
           852 => x"9e",
           853 => x"81",
           854 => x"52",
           855 => x"2e",
           856 => x"52",
           857 => x"dc",
           858 => x"dd",
           859 => x"9e",
           860 => x"70",
           861 => x"70",
           862 => x"51",
           863 => x"72",
           864 => x"54",
           865 => x"80",
           866 => x"90",
           867 => x"52",
           868 => x"83",
           869 => x"71",
           870 => x"0b",
           871 => x"88",
           872 => x"06",
           873 => x"70",
           874 => x"38",
           875 => x"81",
           876 => x"87",
           877 => x"08",
           878 => x"51",
           879 => x"cb",
           880 => x"3d",
           881 => x"3d",
           882 => x"a4",
           883 => x"3f",
           884 => x"33",
           885 => x"2e",
           886 => x"b6",
           887 => x"ad",
           888 => x"cc",
           889 => x"3f",
           890 => x"70",
           891 => x"73",
           892 => x"38",
           893 => x"53",
           894 => x"08",
           895 => x"e4",
           896 => x"3f",
           897 => x"70",
           898 => x"73",
           899 => x"38",
           900 => x"53",
           901 => x"52",
           902 => x"51",
           903 => x"81",
           904 => x"33",
           905 => x"8a",
           906 => x"33",
           907 => x"2e",
           908 => x"cb",
           909 => x"54",
           910 => x"53",
           911 => x"b0",
           912 => x"3f",
           913 => x"33",
           914 => x"2e",
           915 => x"b7",
           916 => x"b9",
           917 => x"da",
           918 => x"80",
           919 => x"81",
           920 => x"83",
           921 => x"cb",
           922 => x"73",
           923 => x"38",
           924 => x"51",
           925 => x"81",
           926 => x"33",
           927 => x"80",
           928 => x"81",
           929 => x"81",
           930 => x"88",
           931 => x"cb",
           932 => x"73",
           933 => x"38",
           934 => x"51",
           935 => x"81",
           936 => x"33",
           937 => x"80",
           938 => x"81",
           939 => x"81",
           940 => x"88",
           941 => x"b8",
           942 => x"d1",
           943 => x"c0",
           944 => x"84",
           945 => x"54",
           946 => x"53",
           947 => x"b7",
           948 => x"52",
           949 => x"51",
           950 => x"88",
           951 => x"81",
           952 => x"88",
           953 => x"15",
           954 => x"b9",
           955 => x"97",
           956 => x"08",
           957 => x"fc",
           958 => x"3f",
           959 => x"04",
           960 => x"02",
           961 => x"52",
           962 => x"bb",
           963 => x"10",
           964 => x"b0",
           965 => x"71",
           966 => x"ba",
           967 => x"bb",
           968 => x"81",
           969 => x"f7",
           970 => x"39",
           971 => x"51",
           972 => x"9a",
           973 => x"bc",
           974 => x"3f",
           975 => x"ba",
           976 => x"97",
           977 => x"81",
           978 => x"f7",
           979 => x"3d",
           980 => x"88",
           981 => x"80",
           982 => x"96",
           983 => x"ff",
           984 => x"c0",
           985 => x"08",
           986 => x"72",
           987 => x"07",
           988 => x"e4",
           989 => x"83",
           990 => x"ff",
           991 => x"c0",
           992 => x"08",
           993 => x"0c",
           994 => x"0c",
           995 => x"81",
           996 => x"06",
           997 => x"e4",
           998 => x"51",
           999 => x"04",
          1000 => x"08",
          1001 => x"84",
          1002 => x"3d",
          1003 => x"05",
          1004 => x"8a",
          1005 => x"06",
          1006 => x"51",
          1007 => x"d3",
          1008 => x"2e",
          1009 => x"d3",
          1010 => x"72",
          1011 => x"d3",
          1012 => x"05",
          1013 => x"0c",
          1014 => x"d3",
          1015 => x"2e",
          1016 => x"51",
          1017 => x"08",
          1018 => x"84",
          1019 => x"fe",
          1020 => x"97",
          1021 => x"d3",
          1022 => x"81",
          1023 => x"54",
          1024 => x"3f",
          1025 => x"bc",
          1026 => x"0d",
          1027 => x"0d",
          1028 => x"53",
          1029 => x"2e",
          1030 => x"70",
          1031 => x"33",
          1032 => x"3f",
          1033 => x"71",
          1034 => x"3d",
          1035 => x"3d",
          1036 => x"d3",
          1037 => x"81",
          1038 => x"71",
          1039 => x"53",
          1040 => x"91",
          1041 => x"81",
          1042 => x"51",
          1043 => x"72",
          1044 => x"f1",
          1045 => x"d3",
          1046 => x"3d",
          1047 => x"3d",
          1048 => x"5d",
          1049 => x"81",
          1050 => x"56",
          1051 => x"85",
          1052 => x"a5",
          1053 => x"75",
          1054 => x"3f",
          1055 => x"70",
          1056 => x"05",
          1057 => x"5e",
          1058 => x"2e",
          1059 => x"8c",
          1060 => x"70",
          1061 => x"33",
          1062 => x"39",
          1063 => x"09",
          1064 => x"38",
          1065 => x"81",
          1066 => x"57",
          1067 => x"2e",
          1068 => x"92",
          1069 => x"1d",
          1070 => x"70",
          1071 => x"33",
          1072 => x"53",
          1073 => x"16",
          1074 => x"26",
          1075 => x"8a",
          1076 => x"05",
          1077 => x"05",
          1078 => x"11",
          1079 => x"89",
          1080 => x"38",
          1081 => x"32",
          1082 => x"72",
          1083 => x"78",
          1084 => x"70",
          1085 => x"07",
          1086 => x"07",
          1087 => x"52",
          1088 => x"80",
          1089 => x"7c",
          1090 => x"70",
          1091 => x"33",
          1092 => x"80",
          1093 => x"38",
          1094 => x"e0",
          1095 => x"38",
          1096 => x"81",
          1097 => x"53",
          1098 => x"53",
          1099 => x"81",
          1100 => x"10",
          1101 => x"c0",
          1102 => x"08",
          1103 => x"1d",
          1104 => x"5d",
          1105 => x"33",
          1106 => x"74",
          1107 => x"81",
          1108 => x"70",
          1109 => x"54",
          1110 => x"7c",
          1111 => x"81",
          1112 => x"72",
          1113 => x"81",
          1114 => x"72",
          1115 => x"38",
          1116 => x"81",
          1117 => x"51",
          1118 => x"75",
          1119 => x"81",
          1120 => x"79",
          1121 => x"38",
          1122 => x"81",
          1123 => x"15",
          1124 => x"7a",
          1125 => x"38",
          1126 => x"8e",
          1127 => x"15",
          1128 => x"73",
          1129 => x"fd",
          1130 => x"84",
          1131 => x"33",
          1132 => x"fb",
          1133 => x"ad",
          1134 => x"95",
          1135 => x"91",
          1136 => x"8d",
          1137 => x"89",
          1138 => x"fb",
          1139 => x"95",
          1140 => x"2a",
          1141 => x"51",
          1142 => x"2e",
          1143 => x"84",
          1144 => x"59",
          1145 => x"39",
          1146 => x"2e",
          1147 => x"8b",
          1148 => x"1d",
          1149 => x"5d",
          1150 => x"7b",
          1151 => x"08",
          1152 => x"74",
          1153 => x"70",
          1154 => x"07",
          1155 => x"80",
          1156 => x"51",
          1157 => x"72",
          1158 => x"38",
          1159 => x"90",
          1160 => x"80",
          1161 => x"76",
          1162 => x"3f",
          1163 => x"08",
          1164 => x"7b",
          1165 => x"55",
          1166 => x"81",
          1167 => x"57",
          1168 => x"99",
          1169 => x"16",
          1170 => x"06",
          1171 => x"75",
          1172 => x"89",
          1173 => x"70",
          1174 => x"56",
          1175 => x"78",
          1176 => x"b0",
          1177 => x"72",
          1178 => x"18",
          1179 => x"79",
          1180 => x"70",
          1181 => x"06",
          1182 => x"58",
          1183 => x"38",
          1184 => x"70",
          1185 => x"53",
          1186 => x"8e",
          1187 => x"78",
          1188 => x"53",
          1189 => x"81",
          1190 => x"7d",
          1191 => x"54",
          1192 => x"83",
          1193 => x"7c",
          1194 => x"81",
          1195 => x"72",
          1196 => x"81",
          1197 => x"72",
          1198 => x"38",
          1199 => x"81",
          1200 => x"51",
          1201 => x"75",
          1202 => x"81",
          1203 => x"79",
          1204 => x"38",
          1205 => x"3d",
          1206 => x"70",
          1207 => x"58",
          1208 => x"77",
          1209 => x"81",
          1210 => x"72",
          1211 => x"f5",
          1212 => x"f9",
          1213 => x"81",
          1214 => x"79",
          1215 => x"38",
          1216 => x"96",
          1217 => x"fd",
          1218 => x"3d",
          1219 => x"05",
          1220 => x"52",
          1221 => x"c6",
          1222 => x"0d",
          1223 => x"0d",
          1224 => x"c4",
          1225 => x"88",
          1226 => x"51",
          1227 => x"81",
          1228 => x"53",
          1229 => x"80",
          1230 => x"c4",
          1231 => x"0d",
          1232 => x"0d",
          1233 => x"08",
          1234 => x"bc",
          1235 => x"88",
          1236 => x"52",
          1237 => x"3f",
          1238 => x"bc",
          1239 => x"0d",
          1240 => x"0d",
          1241 => x"57",
          1242 => x"d3",
          1243 => x"2e",
          1244 => x"86",
          1245 => x"80",
          1246 => x"55",
          1247 => x"08",
          1248 => x"81",
          1249 => x"81",
          1250 => x"73",
          1251 => x"38",
          1252 => x"80",
          1253 => x"88",
          1254 => x"76",
          1255 => x"07",
          1256 => x"80",
          1257 => x"54",
          1258 => x"80",
          1259 => x"ff",
          1260 => x"ff",
          1261 => x"f7",
          1262 => x"39",
          1263 => x"ff",
          1264 => x"16",
          1265 => x"25",
          1266 => x"76",
          1267 => x"72",
          1268 => x"74",
          1269 => x"52",
          1270 => x"3f",
          1271 => x"74",
          1272 => x"72",
          1273 => x"f7",
          1274 => x"53",
          1275 => x"ac",
          1276 => x"0d",
          1277 => x"0d",
          1278 => x"08",
          1279 => x"c0",
          1280 => x"76",
          1281 => x"d9",
          1282 => x"d3",
          1283 => x"3d",
          1284 => x"3d",
          1285 => x"5a",
          1286 => x"7a",
          1287 => x"70",
          1288 => x"58",
          1289 => x"09",
          1290 => x"38",
          1291 => x"05",
          1292 => x"08",
          1293 => x"53",
          1294 => x"f0",
          1295 => x"2e",
          1296 => x"8e",
          1297 => x"08",
          1298 => x"75",
          1299 => x"56",
          1300 => x"b0",
          1301 => x"06",
          1302 => x"74",
          1303 => x"75",
          1304 => x"70",
          1305 => x"73",
          1306 => x"9a",
          1307 => x"f8",
          1308 => x"06",
          1309 => x"0b",
          1310 => x"0c",
          1311 => x"33",
          1312 => x"80",
          1313 => x"75",
          1314 => x"76",
          1315 => x"70",
          1316 => x"57",
          1317 => x"56",
          1318 => x"81",
          1319 => x"14",
          1320 => x"88",
          1321 => x"27",
          1322 => x"f3",
          1323 => x"53",
          1324 => x"89",
          1325 => x"38",
          1326 => x"56",
          1327 => x"80",
          1328 => x"39",
          1329 => x"56",
          1330 => x"80",
          1331 => x"e0",
          1332 => x"38",
          1333 => x"81",
          1334 => x"53",
          1335 => x"81",
          1336 => x"53",
          1337 => x"8e",
          1338 => x"70",
          1339 => x"55",
          1340 => x"27",
          1341 => x"77",
          1342 => x"76",
          1343 => x"75",
          1344 => x"76",
          1345 => x"70",
          1346 => x"56",
          1347 => x"ff",
          1348 => x"80",
          1349 => x"75",
          1350 => x"79",
          1351 => x"75",
          1352 => x"0c",
          1353 => x"04",
          1354 => x"7a",
          1355 => x"80",
          1356 => x"75",
          1357 => x"56",
          1358 => x"a0",
          1359 => x"06",
          1360 => x"08",
          1361 => x"0c",
          1362 => x"33",
          1363 => x"a0",
          1364 => x"73",
          1365 => x"81",
          1366 => x"81",
          1367 => x"76",
          1368 => x"70",
          1369 => x"58",
          1370 => x"09",
          1371 => x"d3",
          1372 => x"81",
          1373 => x"74",
          1374 => x"55",
          1375 => x"e2",
          1376 => x"73",
          1377 => x"09",
          1378 => x"38",
          1379 => x"14",
          1380 => x"08",
          1381 => x"54",
          1382 => x"39",
          1383 => x"81",
          1384 => x"75",
          1385 => x"56",
          1386 => x"39",
          1387 => x"74",
          1388 => x"38",
          1389 => x"80",
          1390 => x"89",
          1391 => x"38",
          1392 => x"d0",
          1393 => x"56",
          1394 => x"80",
          1395 => x"39",
          1396 => x"e1",
          1397 => x"80",
          1398 => x"57",
          1399 => x"74",
          1400 => x"38",
          1401 => x"27",
          1402 => x"14",
          1403 => x"06",
          1404 => x"14",
          1405 => x"06",
          1406 => x"74",
          1407 => x"f9",
          1408 => x"ff",
          1409 => x"89",
          1410 => x"38",
          1411 => x"c5",
          1412 => x"29",
          1413 => x"81",
          1414 => x"75",
          1415 => x"56",
          1416 => x"a0",
          1417 => x"38",
          1418 => x"84",
          1419 => x"56",
          1420 => x"81",
          1421 => x"d3",
          1422 => x"3d",
          1423 => x"3d",
          1424 => x"05",
          1425 => x"52",
          1426 => x"87",
          1427 => x"e8",
          1428 => x"71",
          1429 => x"0c",
          1430 => x"04",
          1431 => x"02",
          1432 => x"02",
          1433 => x"05",
          1434 => x"83",
          1435 => x"26",
          1436 => x"72",
          1437 => x"c0",
          1438 => x"51",
          1439 => x"80",
          1440 => x"81",
          1441 => x"71",
          1442 => x"29",
          1443 => x"8c",
          1444 => x"71",
          1445 => x"87",
          1446 => x"0c",
          1447 => x"c0",
          1448 => x"71",
          1449 => x"06",
          1450 => x"80",
          1451 => x"73",
          1452 => x"ef",
          1453 => x"29",
          1454 => x"8c",
          1455 => x"fc",
          1456 => x"53",
          1457 => x"38",
          1458 => x"8c",
          1459 => x"80",
          1460 => x"71",
          1461 => x"14",
          1462 => x"e8",
          1463 => x"70",
          1464 => x"0c",
          1465 => x"04",
          1466 => x"61",
          1467 => x"8c",
          1468 => x"05",
          1469 => x"5d",
          1470 => x"52",
          1471 => x"3f",
          1472 => x"08",
          1473 => x"55",
          1474 => x"ac",
          1475 => x"58",
          1476 => x"98",
          1477 => x"2b",
          1478 => x"8c",
          1479 => x"92",
          1480 => x"42",
          1481 => x"56",
          1482 => x"87",
          1483 => x"1a",
          1484 => x"52",
          1485 => x"74",
          1486 => x"2a",
          1487 => x"51",
          1488 => x"80",
          1489 => x"78",
          1490 => x"78",
          1491 => x"5a",
          1492 => x"57",
          1493 => x"52",
          1494 => x"87",
          1495 => x"52",
          1496 => x"75",
          1497 => x"80",
          1498 => x"76",
          1499 => x"99",
          1500 => x"0c",
          1501 => x"8c",
          1502 => x"08",
          1503 => x"51",
          1504 => x"38",
          1505 => x"8d",
          1506 => x"1c",
          1507 => x"81",
          1508 => x"53",
          1509 => x"2e",
          1510 => x"fc",
          1511 => x"52",
          1512 => x"7e",
          1513 => x"80",
          1514 => x"80",
          1515 => x"71",
          1516 => x"38",
          1517 => x"54",
          1518 => x"ac",
          1519 => x"0d",
          1520 => x"0d",
          1521 => x"02",
          1522 => x"05",
          1523 => x"5c",
          1524 => x"52",
          1525 => x"3f",
          1526 => x"08",
          1527 => x"55",
          1528 => x"ae",
          1529 => x"87",
          1530 => x"73",
          1531 => x"c0",
          1532 => x"87",
          1533 => x"12",
          1534 => x"57",
          1535 => x"76",
          1536 => x"92",
          1537 => x"71",
          1538 => x"75",
          1539 => x"74",
          1540 => x"2a",
          1541 => x"51",
          1542 => x"80",
          1543 => x"76",
          1544 => x"58",
          1545 => x"81",
          1546 => x"81",
          1547 => x"06",
          1548 => x"80",
          1549 => x"75",
          1550 => x"d3",
          1551 => x"52",
          1552 => x"87",
          1553 => x"80",
          1554 => x"81",
          1555 => x"c0",
          1556 => x"53",
          1557 => x"82",
          1558 => x"71",
          1559 => x"1a",
          1560 => x"81",
          1561 => x"ff",
          1562 => x"1d",
          1563 => x"79",
          1564 => x"38",
          1565 => x"80",
          1566 => x"87",
          1567 => x"26",
          1568 => x"73",
          1569 => x"06",
          1570 => x"2e",
          1571 => x"52",
          1572 => x"81",
          1573 => x"8f",
          1574 => x"f7",
          1575 => x"02",
          1576 => x"05",
          1577 => x"05",
          1578 => x"71",
          1579 => x"56",
          1580 => x"81",
          1581 => x"81",
          1582 => x"54",
          1583 => x"81",
          1584 => x"2e",
          1585 => x"74",
          1586 => x"72",
          1587 => x"38",
          1588 => x"83",
          1589 => x"a0",
          1590 => x"29",
          1591 => x"8c",
          1592 => x"51",
          1593 => x"88",
          1594 => x"0c",
          1595 => x"39",
          1596 => x"0c",
          1597 => x"39",
          1598 => x"81",
          1599 => x"8b",
          1600 => x"ff",
          1601 => x"70",
          1602 => x"33",
          1603 => x"72",
          1604 => x"ac",
          1605 => x"52",
          1606 => x"04",
          1607 => x"75",
          1608 => x"82",
          1609 => x"90",
          1610 => x"2b",
          1611 => x"33",
          1612 => x"33",
          1613 => x"07",
          1614 => x"0c",
          1615 => x"54",
          1616 => x"0d",
          1617 => x"0d",
          1618 => x"05",
          1619 => x"52",
          1620 => x"70",
          1621 => x"34",
          1622 => x"51",
          1623 => x"83",
          1624 => x"ff",
          1625 => x"75",
          1626 => x"72",
          1627 => x"54",
          1628 => x"2a",
          1629 => x"70",
          1630 => x"34",
          1631 => x"51",
          1632 => x"81",
          1633 => x"70",
          1634 => x"70",
          1635 => x"3d",
          1636 => x"3d",
          1637 => x"77",
          1638 => x"70",
          1639 => x"38",
          1640 => x"05",
          1641 => x"70",
          1642 => x"34",
          1643 => x"70",
          1644 => x"3d",
          1645 => x"3d",
          1646 => x"76",
          1647 => x"72",
          1648 => x"05",
          1649 => x"11",
          1650 => x"38",
          1651 => x"04",
          1652 => x"78",
          1653 => x"56",
          1654 => x"81",
          1655 => x"74",
          1656 => x"56",
          1657 => x"31",
          1658 => x"52",
          1659 => x"80",
          1660 => x"71",
          1661 => x"38",
          1662 => x"ac",
          1663 => x"0d",
          1664 => x"0d",
          1665 => x"33",
          1666 => x"70",
          1667 => x"38",
          1668 => x"94",
          1669 => x"70",
          1670 => x"70",
          1671 => x"38",
          1672 => x"09",
          1673 => x"38",
          1674 => x"d3",
          1675 => x"3d",
          1676 => x"0b",
          1677 => x"0c",
          1678 => x"81",
          1679 => x"04",
          1680 => x"79",
          1681 => x"83",
          1682 => x"58",
          1683 => x"80",
          1684 => x"54",
          1685 => x"53",
          1686 => x"53",
          1687 => x"52",
          1688 => x"3f",
          1689 => x"08",
          1690 => x"81",
          1691 => x"81",
          1692 => x"83",
          1693 => x"16",
          1694 => x"08",
          1695 => x"9c",
          1696 => x"a4",
          1697 => x"33",
          1698 => x"2e",
          1699 => x"98",
          1700 => x"b0",
          1701 => x"17",
          1702 => x"76",
          1703 => x"33",
          1704 => x"3f",
          1705 => x"58",
          1706 => x"ac",
          1707 => x"0d",
          1708 => x"0d",
          1709 => x"57",
          1710 => x"17",
          1711 => x"af",
          1712 => x"fe",
          1713 => x"d3",
          1714 => x"81",
          1715 => x"9f",
          1716 => x"74",
          1717 => x"52",
          1718 => x"51",
          1719 => x"81",
          1720 => x"80",
          1721 => x"ff",
          1722 => x"74",
          1723 => x"75",
          1724 => x"0c",
          1725 => x"04",
          1726 => x"7a",
          1727 => x"fe",
          1728 => x"d3",
          1729 => x"81",
          1730 => x"81",
          1731 => x"33",
          1732 => x"2e",
          1733 => x"80",
          1734 => x"17",
          1735 => x"81",
          1736 => x"06",
          1737 => x"84",
          1738 => x"d3",
          1739 => x"b4",
          1740 => x"56",
          1741 => x"82",
          1742 => x"84",
          1743 => x"fc",
          1744 => x"8b",
          1745 => x"52",
          1746 => x"97",
          1747 => x"85",
          1748 => x"84",
          1749 => x"fc",
          1750 => x"17",
          1751 => x"9c",
          1752 => x"ff",
          1753 => x"08",
          1754 => x"17",
          1755 => x"3f",
          1756 => x"81",
          1757 => x"19",
          1758 => x"53",
          1759 => x"17",
          1760 => x"bd",
          1761 => x"18",
          1762 => x"80",
          1763 => x"33",
          1764 => x"3f",
          1765 => x"08",
          1766 => x"38",
          1767 => x"81",
          1768 => x"8a",
          1769 => x"fb",
          1770 => x"fe",
          1771 => x"08",
          1772 => x"56",
          1773 => x"74",
          1774 => x"38",
          1775 => x"70",
          1776 => x"16",
          1777 => x"53",
          1778 => x"ac",
          1779 => x"0d",
          1780 => x"0d",
          1781 => x"08",
          1782 => x"81",
          1783 => x"38",
          1784 => x"75",
          1785 => x"81",
          1786 => x"39",
          1787 => x"54",
          1788 => x"2e",
          1789 => x"72",
          1790 => x"38",
          1791 => x"8d",
          1792 => x"39",
          1793 => x"81",
          1794 => x"b6",
          1795 => x"2a",
          1796 => x"2a",
          1797 => x"05",
          1798 => x"57",
          1799 => x"81",
          1800 => x"81",
          1801 => x"83",
          1802 => x"b4",
          1803 => x"19",
          1804 => x"a4",
          1805 => x"55",
          1806 => x"59",
          1807 => x"3f",
          1808 => x"08",
          1809 => x"76",
          1810 => x"14",
          1811 => x"70",
          1812 => x"07",
          1813 => x"71",
          1814 => x"52",
          1815 => x"72",
          1816 => x"77",
          1817 => x"56",
          1818 => x"74",
          1819 => x"15",
          1820 => x"73",
          1821 => x"3f",
          1822 => x"08",
          1823 => x"74",
          1824 => x"06",
          1825 => x"05",
          1826 => x"3f",
          1827 => x"08",
          1828 => x"06",
          1829 => x"74",
          1830 => x"15",
          1831 => x"73",
          1832 => x"3f",
          1833 => x"08",
          1834 => x"82",
          1835 => x"06",
          1836 => x"05",
          1837 => x"3f",
          1838 => x"08",
          1839 => x"56",
          1840 => x"56",
          1841 => x"ac",
          1842 => x"0d",
          1843 => x"0d",
          1844 => x"58",
          1845 => x"57",
          1846 => x"82",
          1847 => x"98",
          1848 => x"82",
          1849 => x"33",
          1850 => x"2e",
          1851 => x"72",
          1852 => x"38",
          1853 => x"8d",
          1854 => x"39",
          1855 => x"81",
          1856 => x"88",
          1857 => x"2a",
          1858 => x"2a",
          1859 => x"05",
          1860 => x"59",
          1861 => x"81",
          1862 => x"57",
          1863 => x"08",
          1864 => x"78",
          1865 => x"15",
          1866 => x"1b",
          1867 => x"56",
          1868 => x"75",
          1869 => x"2e",
          1870 => x"84",
          1871 => x"06",
          1872 => x"06",
          1873 => x"53",
          1874 => x"81",
          1875 => x"34",
          1876 => x"a4",
          1877 => x"52",
          1878 => x"d5",
          1879 => x"ac",
          1880 => x"d3",
          1881 => x"a4",
          1882 => x"ff",
          1883 => x"11",
          1884 => x"78",
          1885 => x"55",
          1886 => x"8f",
          1887 => x"2a",
          1888 => x"8f",
          1889 => x"f0",
          1890 => x"73",
          1891 => x"0b",
          1892 => x"80",
          1893 => x"88",
          1894 => x"08",
          1895 => x"51",
          1896 => x"81",
          1897 => x"57",
          1898 => x"08",
          1899 => x"75",
          1900 => x"06",
          1901 => x"83",
          1902 => x"05",
          1903 => x"f7",
          1904 => x"0b",
          1905 => x"80",
          1906 => x"87",
          1907 => x"08",
          1908 => x"51",
          1909 => x"81",
          1910 => x"57",
          1911 => x"08",
          1912 => x"f0",
          1913 => x"82",
          1914 => x"06",
          1915 => x"05",
          1916 => x"54",
          1917 => x"3f",
          1918 => x"08",
          1919 => x"76",
          1920 => x"51",
          1921 => x"81",
          1922 => x"34",
          1923 => x"ac",
          1924 => x"0d",
          1925 => x"0d",
          1926 => x"72",
          1927 => x"55",
          1928 => x"27",
          1929 => x"15",
          1930 => x"86",
          1931 => x"81",
          1932 => x"80",
          1933 => x"ff",
          1934 => x"74",
          1935 => x"3f",
          1936 => x"08",
          1937 => x"ac",
          1938 => x"38",
          1939 => x"56",
          1940 => x"81",
          1941 => x"39",
          1942 => x"08",
          1943 => x"39",
          1944 => x"51",
          1945 => x"81",
          1946 => x"56",
          1947 => x"08",
          1948 => x"c9",
          1949 => x"ac",
          1950 => x"d2",
          1951 => x"ac",
          1952 => x"cf",
          1953 => x"73",
          1954 => x"fc",
          1955 => x"d3",
          1956 => x"38",
          1957 => x"fe",
          1958 => x"15",
          1959 => x"93",
          1960 => x"08",
          1961 => x"16",
          1962 => x"33",
          1963 => x"73",
          1964 => x"75",
          1965 => x"08",
          1966 => x"a4",
          1967 => x"75",
          1968 => x"0c",
          1969 => x"04",
          1970 => x"7d",
          1971 => x"5b",
          1972 => x"95",
          1973 => x"08",
          1974 => x"2e",
          1975 => x"19",
          1976 => x"b7",
          1977 => x"b3",
          1978 => x"7b",
          1979 => x"3f",
          1980 => x"81",
          1981 => x"27",
          1982 => x"81",
          1983 => x"55",
          1984 => x"08",
          1985 => x"db",
          1986 => x"ac",
          1987 => x"19",
          1988 => x"ac",
          1989 => x"cb",
          1990 => x"80",
          1991 => x"08",
          1992 => x"bf",
          1993 => x"77",
          1994 => x"81",
          1995 => x"38",
          1996 => x"98",
          1997 => x"26",
          1998 => x"57",
          1999 => x"51",
          2000 => x"81",
          2001 => x"56",
          2002 => x"d3",
          2003 => x"2e",
          2004 => x"86",
          2005 => x"ac",
          2006 => x"ff",
          2007 => x"70",
          2008 => x"25",
          2009 => x"79",
          2010 => x"56",
          2011 => x"f3",
          2012 => x"2e",
          2013 => x"19",
          2014 => x"76",
          2015 => x"75",
          2016 => x"27",
          2017 => x"58",
          2018 => x"80",
          2019 => x"57",
          2020 => x"98",
          2021 => x"26",
          2022 => x"57",
          2023 => x"81",
          2024 => x"52",
          2025 => x"a9",
          2026 => x"ac",
          2027 => x"d3",
          2028 => x"2e",
          2029 => x"5a",
          2030 => x"08",
          2031 => x"81",
          2032 => x"81",
          2033 => x"5a",
          2034 => x"70",
          2035 => x"07",
          2036 => x"7d",
          2037 => x"56",
          2038 => x"ff",
          2039 => x"2e",
          2040 => x"ff",
          2041 => x"55",
          2042 => x"ff",
          2043 => x"78",
          2044 => x"3f",
          2045 => x"08",
          2046 => x"08",
          2047 => x"d3",
          2048 => x"80",
          2049 => x"70",
          2050 => x"2a",
          2051 => x"57",
          2052 => x"74",
          2053 => x"38",
          2054 => x"52",
          2055 => x"ad",
          2056 => x"ac",
          2057 => x"a6",
          2058 => x"1a",
          2059 => x"08",
          2060 => x"90",
          2061 => x"26",
          2062 => x"19",
          2063 => x"90",
          2064 => x"19",
          2065 => x"54",
          2066 => x"34",
          2067 => x"57",
          2068 => x"8d",
          2069 => x"80",
          2070 => x"75",
          2071 => x"81",
          2072 => x"74",
          2073 => x"0c",
          2074 => x"04",
          2075 => x"7b",
          2076 => x"f3",
          2077 => x"55",
          2078 => x"08",
          2079 => x"7c",
          2080 => x"f6",
          2081 => x"d3",
          2082 => x"d3",
          2083 => x"19",
          2084 => x"80",
          2085 => x"b4",
          2086 => x"55",
          2087 => x"74",
          2088 => x"80",
          2089 => x"77",
          2090 => x"17",
          2091 => x"75",
          2092 => x"77",
          2093 => x"53",
          2094 => x"17",
          2095 => x"81",
          2096 => x"ac",
          2097 => x"df",
          2098 => x"8a",
          2099 => x"58",
          2100 => x"83",
          2101 => x"77",
          2102 => x"d3",
          2103 => x"3d",
          2104 => x"3d",
          2105 => x"71",
          2106 => x"57",
          2107 => x"0a",
          2108 => x"74",
          2109 => x"72",
          2110 => x"38",
          2111 => x"ae",
          2112 => x"18",
          2113 => x"08",
          2114 => x"38",
          2115 => x"82",
          2116 => x"38",
          2117 => x"54",
          2118 => x"74",
          2119 => x"82",
          2120 => x"22",
          2121 => x"79",
          2122 => x"38",
          2123 => x"98",
          2124 => x"d1",
          2125 => x"22",
          2126 => x"54",
          2127 => x"26",
          2128 => x"52",
          2129 => x"89",
          2130 => x"ac",
          2131 => x"d3",
          2132 => x"2e",
          2133 => x"0b",
          2134 => x"08",
          2135 => x"98",
          2136 => x"d3",
          2137 => x"86",
          2138 => x"80",
          2139 => x"73",
          2140 => x"73",
          2141 => x"73",
          2142 => x"f4",
          2143 => x"d3",
          2144 => x"18",
          2145 => x"18",
          2146 => x"98",
          2147 => x"2e",
          2148 => x"39",
          2149 => x"39",
          2150 => x"98",
          2151 => x"98",
          2152 => x"83",
          2153 => x"b4",
          2154 => x"0c",
          2155 => x"81",
          2156 => x"8a",
          2157 => x"f9",
          2158 => x"7b",
          2159 => x"13",
          2160 => x"59",
          2161 => x"f0",
          2162 => x"27",
          2163 => x"0b",
          2164 => x"84",
          2165 => x"08",
          2166 => x"da",
          2167 => x"ff",
          2168 => x"81",
          2169 => x"15",
          2170 => x"98",
          2171 => x"15",
          2172 => x"75",
          2173 => x"18",
          2174 => x"77",
          2175 => x"a6",
          2176 => x"16",
          2177 => x"81",
          2178 => x"17",
          2179 => x"77",
          2180 => x"51",
          2181 => x"8e",
          2182 => x"08",
          2183 => x"f3",
          2184 => x"d3",
          2185 => x"82",
          2186 => x"81",
          2187 => x"27",
          2188 => x"81",
          2189 => x"ac",
          2190 => x"80",
          2191 => x"17",
          2192 => x"ac",
          2193 => x"cc",
          2194 => x"38",
          2195 => x"0c",
          2196 => x"e2",
          2197 => x"08",
          2198 => x"f8",
          2199 => x"d3",
          2200 => x"87",
          2201 => x"ac",
          2202 => x"80",
          2203 => x"53",
          2204 => x"08",
          2205 => x"38",
          2206 => x"d3",
          2207 => x"2e",
          2208 => x"d3",
          2209 => x"76",
          2210 => x"3f",
          2211 => x"d3",
          2212 => x"38",
          2213 => x"0c",
          2214 => x"51",
          2215 => x"81",
          2216 => x"98",
          2217 => x"90",
          2218 => x"83",
          2219 => x"b4",
          2220 => x"0c",
          2221 => x"81",
          2222 => x"89",
          2223 => x"f8",
          2224 => x"7c",
          2225 => x"5a",
          2226 => x"75",
          2227 => x"3f",
          2228 => x"08",
          2229 => x"ac",
          2230 => x"38",
          2231 => x"08",
          2232 => x"08",
          2233 => x"ef",
          2234 => x"d3",
          2235 => x"81",
          2236 => x"80",
          2237 => x"d3",
          2238 => x"17",
          2239 => x"51",
          2240 => x"81",
          2241 => x"81",
          2242 => x"81",
          2243 => x"70",
          2244 => x"07",
          2245 => x"80",
          2246 => x"81",
          2247 => x"79",
          2248 => x"83",
          2249 => x"81",
          2250 => x"fd",
          2251 => x"d3",
          2252 => x"81",
          2253 => x"80",
          2254 => x"38",
          2255 => x"09",
          2256 => x"38",
          2257 => x"81",
          2258 => x"8a",
          2259 => x"fd",
          2260 => x"9a",
          2261 => x"eb",
          2262 => x"d3",
          2263 => x"ff",
          2264 => x"70",
          2265 => x"53",
          2266 => x"09",
          2267 => x"38",
          2268 => x"eb",
          2269 => x"d3",
          2270 => x"2b",
          2271 => x"72",
          2272 => x"0c",
          2273 => x"04",
          2274 => x"77",
          2275 => x"ff",
          2276 => x"9a",
          2277 => x"55",
          2278 => x"76",
          2279 => x"53",
          2280 => x"09",
          2281 => x"38",
          2282 => x"52",
          2283 => x"eb",
          2284 => x"3d",
          2285 => x"3d",
          2286 => x"5b",
          2287 => x"08",
          2288 => x"16",
          2289 => x"81",
          2290 => x"16",
          2291 => x"51",
          2292 => x"81",
          2293 => x"58",
          2294 => x"08",
          2295 => x"9c",
          2296 => x"33",
          2297 => x"86",
          2298 => x"80",
          2299 => x"16",
          2300 => x"33",
          2301 => x"70",
          2302 => x"5a",
          2303 => x"72",
          2304 => x"74",
          2305 => x"70",
          2306 => x"32",
          2307 => x"73",
          2308 => x"53",
          2309 => x"54",
          2310 => x"9b",
          2311 => x"2e",
          2312 => x"77",
          2313 => x"54",
          2314 => x"09",
          2315 => x"38",
          2316 => x"7a",
          2317 => x"80",
          2318 => x"fa",
          2319 => x"d3",
          2320 => x"81",
          2321 => x"87",
          2322 => x"08",
          2323 => x"77",
          2324 => x"38",
          2325 => x"17",
          2326 => x"d3",
          2327 => x"3d",
          2328 => x"3d",
          2329 => x"08",
          2330 => x"52",
          2331 => x"f2",
          2332 => x"ac",
          2333 => x"d3",
          2334 => x"ef",
          2335 => x"84",
          2336 => x"39",
          2337 => x"52",
          2338 => x"a5",
          2339 => x"ac",
          2340 => x"d3",
          2341 => x"d1",
          2342 => x"08",
          2343 => x"54",
          2344 => x"db",
          2345 => x"08",
          2346 => x"bf",
          2347 => x"73",
          2348 => x"8b",
          2349 => x"83",
          2350 => x"06",
          2351 => x"73",
          2352 => x"53",
          2353 => x"74",
          2354 => x"3f",
          2355 => x"08",
          2356 => x"38",
          2357 => x"51",
          2358 => x"81",
          2359 => x"57",
          2360 => x"08",
          2361 => x"9c",
          2362 => x"73",
          2363 => x"0c",
          2364 => x"04",
          2365 => x"77",
          2366 => x"54",
          2367 => x"51",
          2368 => x"81",
          2369 => x"55",
          2370 => x"08",
          2371 => x"14",
          2372 => x"51",
          2373 => x"81",
          2374 => x"55",
          2375 => x"08",
          2376 => x"53",
          2377 => x"08",
          2378 => x"08",
          2379 => x"3f",
          2380 => x"14",
          2381 => x"08",
          2382 => x"3f",
          2383 => x"17",
          2384 => x"d3",
          2385 => x"3d",
          2386 => x"3d",
          2387 => x"08",
          2388 => x"54",
          2389 => x"53",
          2390 => x"81",
          2391 => x"54",
          2392 => x"08",
          2393 => x"13",
          2394 => x"73",
          2395 => x"83",
          2396 => x"81",
          2397 => x"86",
          2398 => x"fa",
          2399 => x"7a",
          2400 => x"0b",
          2401 => x"98",
          2402 => x"2e",
          2403 => x"80",
          2404 => x"9c",
          2405 => x"70",
          2406 => x"56",
          2407 => x"a0",
          2408 => x"72",
          2409 => x"81",
          2410 => x"81",
          2411 => x"89",
          2412 => x"06",
          2413 => x"15",
          2414 => x"ae",
          2415 => x"34",
          2416 => x"75",
          2417 => x"52",
          2418 => x"34",
          2419 => x"8a",
          2420 => x"38",
          2421 => x"05",
          2422 => x"81",
          2423 => x"17",
          2424 => x"12",
          2425 => x"34",
          2426 => x"9c",
          2427 => x"ac",
          2428 => x"ac",
          2429 => x"9c",
          2430 => x"05",
          2431 => x"3f",
          2432 => x"08",
          2433 => x"9c",
          2434 => x"05",
          2435 => x"3f",
          2436 => x"08",
          2437 => x"88",
          2438 => x"f5",
          2439 => x"70",
          2440 => x"05",
          2441 => x"8b",
          2442 => x"7a",
          2443 => x"3f",
          2444 => x"58",
          2445 => x"55",
          2446 => x"2e",
          2447 => x"80",
          2448 => x"17",
          2449 => x"19",
          2450 => x"70",
          2451 => x"2a",
          2452 => x"07",
          2453 => x"59",
          2454 => x"8c",
          2455 => x"54",
          2456 => x"81",
          2457 => x"39",
          2458 => x"70",
          2459 => x"dc",
          2460 => x"70",
          2461 => x"2a",
          2462 => x"51",
          2463 => x"2e",
          2464 => x"54",
          2465 => x"82",
          2466 => x"19",
          2467 => x"54",
          2468 => x"83",
          2469 => x"73",
          2470 => x"80",
          2471 => x"39",
          2472 => x"33",
          2473 => x"57",
          2474 => x"27",
          2475 => x"75",
          2476 => x"30",
          2477 => x"32",
          2478 => x"80",
          2479 => x"25",
          2480 => x"56",
          2481 => x"80",
          2482 => x"84",
          2483 => x"57",
          2484 => x"70",
          2485 => x"5a",
          2486 => x"09",
          2487 => x"38",
          2488 => x"77",
          2489 => x"51",
          2490 => x"80",
          2491 => x"81",
          2492 => x"81",
          2493 => x"07",
          2494 => x"38",
          2495 => x"75",
          2496 => x"30",
          2497 => x"7a",
          2498 => x"51",
          2499 => x"80",
          2500 => x"79",
          2501 => x"30",
          2502 => x"70",
          2503 => x"25",
          2504 => x"07",
          2505 => x"51",
          2506 => x"b1",
          2507 => x"8b",
          2508 => x"39",
          2509 => x"54",
          2510 => x"8c",
          2511 => x"ff",
          2512 => x"dc",
          2513 => x"54",
          2514 => x"e6",
          2515 => x"ac",
          2516 => x"b9",
          2517 => x"70",
          2518 => x"71",
          2519 => x"54",
          2520 => x"81",
          2521 => x"80",
          2522 => x"ff",
          2523 => x"78",
          2524 => x"86",
          2525 => x"39",
          2526 => x"75",
          2527 => x"18",
          2528 => x"58",
          2529 => x"81",
          2530 => x"94",
          2531 => x"81",
          2532 => x"e4",
          2533 => x"d3",
          2534 => x"c5",
          2535 => x"16",
          2536 => x"26",
          2537 => x"16",
          2538 => x"06",
          2539 => x"18",
          2540 => x"34",
          2541 => x"fd",
          2542 => x"19",
          2543 => x"54",
          2544 => x"a9",
          2545 => x"54",
          2546 => x"2e",
          2547 => x"84",
          2548 => x"34",
          2549 => x"76",
          2550 => x"89",
          2551 => x"8d",
          2552 => x"89",
          2553 => x"73",
          2554 => x"80",
          2555 => x"d3",
          2556 => x"3d",
          2557 => x"3d",
          2558 => x"08",
          2559 => x"7a",
          2560 => x"54",
          2561 => x"2e",
          2562 => x"55",
          2563 => x"33",
          2564 => x"72",
          2565 => x"83",
          2566 => x"74",
          2567 => x"72",
          2568 => x"38",
          2569 => x"88",
          2570 => x"39",
          2571 => x"80",
          2572 => x"51",
          2573 => x"af",
          2574 => x"06",
          2575 => x"55",
          2576 => x"33",
          2577 => x"72",
          2578 => x"09",
          2579 => x"38",
          2580 => x"74",
          2581 => x"d4",
          2582 => x"88",
          2583 => x"70",
          2584 => x"72",
          2585 => x"38",
          2586 => x"ab",
          2587 => x"52",
          2588 => x"ee",
          2589 => x"ac",
          2590 => x"aa",
          2591 => x"81",
          2592 => x"3d",
          2593 => x"75",
          2594 => x"3f",
          2595 => x"08",
          2596 => x"ac",
          2597 => x"38",
          2598 => x"c6",
          2599 => x"ac",
          2600 => x"33",
          2601 => x"d3",
          2602 => x"2e",
          2603 => x"81",
          2604 => x"84",
          2605 => x"06",
          2606 => x"73",
          2607 => x"81",
          2608 => x"72",
          2609 => x"38",
          2610 => x"70",
          2611 => x"53",
          2612 => x"ff",
          2613 => x"80",
          2614 => x"34",
          2615 => x"c6",
          2616 => x"2a",
          2617 => x"51",
          2618 => x"38",
          2619 => x"39",
          2620 => x"70",
          2621 => x"53",
          2622 => x"86",
          2623 => x"84",
          2624 => x"06",
          2625 => x"72",
          2626 => x"f1",
          2627 => x"08",
          2628 => x"17",
          2629 => x"76",
          2630 => x"3f",
          2631 => x"08",
          2632 => x"fe",
          2633 => x"81",
          2634 => x"88",
          2635 => x"f6",
          2636 => x"59",
          2637 => x"70",
          2638 => x"56",
          2639 => x"2e",
          2640 => x"76",
          2641 => x"58",
          2642 => x"32",
          2643 => x"a0",
          2644 => x"2a",
          2645 => x"52",
          2646 => x"38",
          2647 => x"09",
          2648 => x"a9",
          2649 => x"d0",
          2650 => x"70",
          2651 => x"38",
          2652 => x"81",
          2653 => x"11",
          2654 => x"70",
          2655 => x"ff",
          2656 => x"81",
          2657 => x"58",
          2658 => x"1b",
          2659 => x"08",
          2660 => x"75",
          2661 => x"57",
          2662 => x"81",
          2663 => x"ff",
          2664 => x"54",
          2665 => x"26",
          2666 => x"14",
          2667 => x"06",
          2668 => x"9f",
          2669 => x"99",
          2670 => x"e0",
          2671 => x"ff",
          2672 => x"73",
          2673 => x"32",
          2674 => x"72",
          2675 => x"73",
          2676 => x"53",
          2677 => x"70",
          2678 => x"73",
          2679 => x"32",
          2680 => x"72",
          2681 => x"73",
          2682 => x"53",
          2683 => x"70",
          2684 => x"38",
          2685 => x"83",
          2686 => x"8c",
          2687 => x"77",
          2688 => x"38",
          2689 => x"0c",
          2690 => x"86",
          2691 => x"dc",
          2692 => x"81",
          2693 => x"8c",
          2694 => x"fb",
          2695 => x"56",
          2696 => x"17",
          2697 => x"b0",
          2698 => x"52",
          2699 => x"81",
          2700 => x"81",
          2701 => x"81",
          2702 => x"b2",
          2703 => x"c3",
          2704 => x"ac",
          2705 => x"ff",
          2706 => x"55",
          2707 => x"d5",
          2708 => x"06",
          2709 => x"80",
          2710 => x"33",
          2711 => x"81",
          2712 => x"81",
          2713 => x"81",
          2714 => x"eb",
          2715 => x"70",
          2716 => x"07",
          2717 => x"73",
          2718 => x"16",
          2719 => x"81",
          2720 => x"81",
          2721 => x"83",
          2722 => x"e4",
          2723 => x"16",
          2724 => x"3f",
          2725 => x"08",
          2726 => x"ac",
          2727 => x"9d",
          2728 => x"81",
          2729 => x"81",
          2730 => x"de",
          2731 => x"d3",
          2732 => x"81",
          2733 => x"80",
          2734 => x"82",
          2735 => x"d3",
          2736 => x"3d",
          2737 => x"3d",
          2738 => x"84",
          2739 => x"05",
          2740 => x"80",
          2741 => x"51",
          2742 => x"81",
          2743 => x"58",
          2744 => x"0b",
          2745 => x"08",
          2746 => x"38",
          2747 => x"08",
          2748 => x"d3",
          2749 => x"08",
          2750 => x"56",
          2751 => x"87",
          2752 => x"74",
          2753 => x"fe",
          2754 => x"54",
          2755 => x"2e",
          2756 => x"15",
          2757 => x"a6",
          2758 => x"ac",
          2759 => x"06",
          2760 => x"54",
          2761 => x"38",
          2762 => x"8f",
          2763 => x"2a",
          2764 => x"51",
          2765 => x"72",
          2766 => x"80",
          2767 => x"39",
          2768 => x"77",
          2769 => x"81",
          2770 => x"33",
          2771 => x"3f",
          2772 => x"08",
          2773 => x"70",
          2774 => x"54",
          2775 => x"86",
          2776 => x"80",
          2777 => x"73",
          2778 => x"81",
          2779 => x"8a",
          2780 => x"95",
          2781 => x"53",
          2782 => x"fd",
          2783 => x"d3",
          2784 => x"ff",
          2785 => x"82",
          2786 => x"06",
          2787 => x"79",
          2788 => x"29",
          2789 => x"75",
          2790 => x"f0",
          2791 => x"12",
          2792 => x"56",
          2793 => x"77",
          2794 => x"83",
          2795 => x"da",
          2796 => x"d3",
          2797 => x"76",
          2798 => x"14",
          2799 => x"27",
          2800 => x"54",
          2801 => x"10",
          2802 => x"11",
          2803 => x"83",
          2804 => x"2e",
          2805 => x"52",
          2806 => x"bf",
          2807 => x"ac",
          2808 => x"06",
          2809 => x"27",
          2810 => x"14",
          2811 => x"27",
          2812 => x"56",
          2813 => x"85",
          2814 => x"56",
          2815 => x"85",
          2816 => x"15",
          2817 => x"3f",
          2818 => x"08",
          2819 => x"06",
          2820 => x"72",
          2821 => x"09",
          2822 => x"ed",
          2823 => x"15",
          2824 => x"3f",
          2825 => x"08",
          2826 => x"06",
          2827 => x"38",
          2828 => x"51",
          2829 => x"81",
          2830 => x"54",
          2831 => x"0c",
          2832 => x"33",
          2833 => x"80",
          2834 => x"ff",
          2835 => x"56",
          2836 => x"84",
          2837 => x"15",
          2838 => x"29",
          2839 => x"33",
          2840 => x"72",
          2841 => x"72",
          2842 => x"06",
          2843 => x"2e",
          2844 => x"13",
          2845 => x"72",
          2846 => x"38",
          2847 => x"89",
          2848 => x"15",
          2849 => x"3f",
          2850 => x"08",
          2851 => x"81",
          2852 => x"83",
          2853 => x"8f",
          2854 => x"56",
          2855 => x"38",
          2856 => x"51",
          2857 => x"81",
          2858 => x"83",
          2859 => x"53",
          2860 => x"80",
          2861 => x"d8",
          2862 => x"d3",
          2863 => x"80",
          2864 => x"d8",
          2865 => x"d3",
          2866 => x"ff",
          2867 => x"8d",
          2868 => x"2e",
          2869 => x"88",
          2870 => x"1a",
          2871 => x"05",
          2872 => x"56",
          2873 => x"83",
          2874 => x"15",
          2875 => x"78",
          2876 => x"b0",
          2877 => x"d3",
          2878 => x"8d",
          2879 => x"ac",
          2880 => x"83",
          2881 => x"57",
          2882 => x"08",
          2883 => x"ff",
          2884 => x"38",
          2885 => x"83",
          2886 => x"83",
          2887 => x"72",
          2888 => x"83",
          2889 => x"8d",
          2890 => x"2e",
          2891 => x"82",
          2892 => x"0c",
          2893 => x"0c",
          2894 => x"16",
          2895 => x"ac",
          2896 => x"83",
          2897 => x"06",
          2898 => x"de",
          2899 => x"b3",
          2900 => x"ac",
          2901 => x"ff",
          2902 => x"56",
          2903 => x"38",
          2904 => x"53",
          2905 => x"82",
          2906 => x"e0",
          2907 => x"ac",
          2908 => x"ac",
          2909 => x"0c",
          2910 => x"82",
          2911 => x"39",
          2912 => x"53",
          2913 => x"80",
          2914 => x"38",
          2915 => x"14",
          2916 => x"76",
          2917 => x"81",
          2918 => x"98",
          2919 => x"53",
          2920 => x"15",
          2921 => x"16",
          2922 => x"81",
          2923 => x"08",
          2924 => x"51",
          2925 => x"13",
          2926 => x"8d",
          2927 => x"16",
          2928 => x"c5",
          2929 => x"90",
          2930 => x"0b",
          2931 => x"ff",
          2932 => x"16",
          2933 => x"2e",
          2934 => x"81",
          2935 => x"e4",
          2936 => x"9f",
          2937 => x"ac",
          2938 => x"ff",
          2939 => x"81",
          2940 => x"06",
          2941 => x"81",
          2942 => x"51",
          2943 => x"81",
          2944 => x"80",
          2945 => x"d3",
          2946 => x"16",
          2947 => x"15",
          2948 => x"3f",
          2949 => x"08",
          2950 => x"06",
          2951 => x"d4",
          2952 => x"81",
          2953 => x"38",
          2954 => x"d5",
          2955 => x"d3",
          2956 => x"8b",
          2957 => x"2e",
          2958 => x"b3",
          2959 => x"15",
          2960 => x"3f",
          2961 => x"08",
          2962 => x"e4",
          2963 => x"81",
          2964 => x"84",
          2965 => x"d5",
          2966 => x"d3",
          2967 => x"16",
          2968 => x"15",
          2969 => x"3f",
          2970 => x"08",
          2971 => x"76",
          2972 => x"d3",
          2973 => x"05",
          2974 => x"d3",
          2975 => x"86",
          2976 => x"0b",
          2977 => x"80",
          2978 => x"d3",
          2979 => x"3d",
          2980 => x"3d",
          2981 => x"89",
          2982 => x"2e",
          2983 => x"08",
          2984 => x"38",
          2985 => x"33",
          2986 => x"80",
          2987 => x"84",
          2988 => x"14",
          2989 => x"71",
          2990 => x"81",
          2991 => x"81",
          2992 => x"ce",
          2993 => x"d3",
          2994 => x"06",
          2995 => x"38",
          2996 => x"53",
          2997 => x"09",
          2998 => x"38",
          2999 => x"78",
          3000 => x"52",
          3001 => x"ac",
          3002 => x"0d",
          3003 => x"0d",
          3004 => x"33",
          3005 => x"3d",
          3006 => x"56",
          3007 => x"81",
          3008 => x"55",
          3009 => x"0b",
          3010 => x"08",
          3011 => x"38",
          3012 => x"08",
          3013 => x"d3",
          3014 => x"08",
          3015 => x"80",
          3016 => x"80",
          3017 => x"80",
          3018 => x"78",
          3019 => x"34",
          3020 => x"81",
          3021 => x"79",
          3022 => x"75",
          3023 => x"2e",
          3024 => x"53",
          3025 => x"53",
          3026 => x"f6",
          3027 => x"d3",
          3028 => x"73",
          3029 => x"0c",
          3030 => x"04",
          3031 => x"67",
          3032 => x"80",
          3033 => x"58",
          3034 => x"77",
          3035 => x"e9",
          3036 => x"06",
          3037 => x"3d",
          3038 => x"99",
          3039 => x"52",
          3040 => x"3f",
          3041 => x"08",
          3042 => x"ac",
          3043 => x"38",
          3044 => x"52",
          3045 => x"05",
          3046 => x"3f",
          3047 => x"08",
          3048 => x"ac",
          3049 => x"02",
          3050 => x"33",
          3051 => x"56",
          3052 => x"25",
          3053 => x"56",
          3054 => x"55",
          3055 => x"81",
          3056 => x"80",
          3057 => x"75",
          3058 => x"81",
          3059 => x"97",
          3060 => x"51",
          3061 => x"81",
          3062 => x"56",
          3063 => x"57",
          3064 => x"b2",
          3065 => x"06",
          3066 => x"2e",
          3067 => x"56",
          3068 => x"82",
          3069 => x"06",
          3070 => x"80",
          3071 => x"88",
          3072 => x"d0",
          3073 => x"2a",
          3074 => x"51",
          3075 => x"2e",
          3076 => x"62",
          3077 => x"e6",
          3078 => x"d3",
          3079 => x"82",
          3080 => x"52",
          3081 => x"51",
          3082 => x"62",
          3083 => x"8b",
          3084 => x"53",
          3085 => x"51",
          3086 => x"75",
          3087 => x"05",
          3088 => x"3f",
          3089 => x"0b",
          3090 => x"78",
          3091 => x"e9",
          3092 => x"11",
          3093 => x"7a",
          3094 => x"d4",
          3095 => x"55",
          3096 => x"81",
          3097 => x"56",
          3098 => x"08",
          3099 => x"74",
          3100 => x"d4",
          3101 => x"d3",
          3102 => x"ff",
          3103 => x"0c",
          3104 => x"39",
          3105 => x"38",
          3106 => x"33",
          3107 => x"70",
          3108 => x"56",
          3109 => x"2e",
          3110 => x"56",
          3111 => x"81",
          3112 => x"06",
          3113 => x"80",
          3114 => x"02",
          3115 => x"81",
          3116 => x"80",
          3117 => x"87",
          3118 => x"98",
          3119 => x"2a",
          3120 => x"51",
          3121 => x"2e",
          3122 => x"80",
          3123 => x"7a",
          3124 => x"a0",
          3125 => x"a4",
          3126 => x"75",
          3127 => x"62",
          3128 => x"e4",
          3129 => x"d3",
          3130 => x"19",
          3131 => x"05",
          3132 => x"3f",
          3133 => x"08",
          3134 => x"74",
          3135 => x"15",
          3136 => x"23",
          3137 => x"34",
          3138 => x"34",
          3139 => x"0c",
          3140 => x"0c",
          3141 => x"75",
          3142 => x"51",
          3143 => x"76",
          3144 => x"81",
          3145 => x"74",
          3146 => x"a3",
          3147 => x"08",
          3148 => x"9b",
          3149 => x"08",
          3150 => x"7a",
          3151 => x"70",
          3152 => x"1b",
          3153 => x"08",
          3154 => x"51",
          3155 => x"76",
          3156 => x"d4",
          3157 => x"d3",
          3158 => x"81",
          3159 => x"81",
          3160 => x"82",
          3161 => x"2e",
          3162 => x"83",
          3163 => x"78",
          3164 => x"75",
          3165 => x"07",
          3166 => x"7b",
          3167 => x"51",
          3168 => x"cb",
          3169 => x"19",
          3170 => x"c8",
          3171 => x"ff",
          3172 => x"80",
          3173 => x"76",
          3174 => x"d4",
          3175 => x"d3",
          3176 => x"38",
          3177 => x"39",
          3178 => x"81",
          3179 => x"05",
          3180 => x"0c",
          3181 => x"74",
          3182 => x"52",
          3183 => x"33",
          3184 => x"a4",
          3185 => x"ac",
          3186 => x"83",
          3187 => x"75",
          3188 => x"38",
          3189 => x"75",
          3190 => x"d3",
          3191 => x"3d",
          3192 => x"3d",
          3193 => x"64",
          3194 => x"5a",
          3195 => x"0c",
          3196 => x"05",
          3197 => x"f9",
          3198 => x"d3",
          3199 => x"81",
          3200 => x"8a",
          3201 => x"33",
          3202 => x"2e",
          3203 => x"56",
          3204 => x"90",
          3205 => x"06",
          3206 => x"74",
          3207 => x"a0",
          3208 => x"82",
          3209 => x"34",
          3210 => x"94",
          3211 => x"91",
          3212 => x"56",
          3213 => x"82",
          3214 => x"34",
          3215 => x"80",
          3216 => x"91",
          3217 => x"56",
          3218 => x"81",
          3219 => x"34",
          3220 => x"ec",
          3221 => x"91",
          3222 => x"56",
          3223 => x"8c",
          3224 => x"18",
          3225 => x"74",
          3226 => x"38",
          3227 => x"80",
          3228 => x"38",
          3229 => x"70",
          3230 => x"56",
          3231 => x"83",
          3232 => x"11",
          3233 => x"77",
          3234 => x"5c",
          3235 => x"38",
          3236 => x"88",
          3237 => x"8f",
          3238 => x"08",
          3239 => x"d2",
          3240 => x"d3",
          3241 => x"81",
          3242 => x"f7",
          3243 => x"2e",
          3244 => x"74",
          3245 => x"98",
          3246 => x"7d",
          3247 => x"3f",
          3248 => x"08",
          3249 => x"ef",
          3250 => x"ac",
          3251 => x"89",
          3252 => x"79",
          3253 => x"d7",
          3254 => x"7e",
          3255 => x"51",
          3256 => x"76",
          3257 => x"74",
          3258 => x"79",
          3259 => x"7b",
          3260 => x"11",
          3261 => x"c7",
          3262 => x"d3",
          3263 => x"c1",
          3264 => x"33",
          3265 => x"56",
          3266 => x"25",
          3267 => x"17",
          3268 => x"55",
          3269 => x"90",
          3270 => x"53",
          3271 => x"74",
          3272 => x"1c",
          3273 => x"3f",
          3274 => x"56",
          3275 => x"9c",
          3276 => x"2e",
          3277 => x"90",
          3278 => x"98",
          3279 => x"74",
          3280 => x"38",
          3281 => x"17",
          3282 => x"17",
          3283 => x"11",
          3284 => x"c8",
          3285 => x"d3",
          3286 => x"ef",
          3287 => x"33",
          3288 => x"55",
          3289 => x"34",
          3290 => x"53",
          3291 => x"7d",
          3292 => x"52",
          3293 => x"3f",
          3294 => x"08",
          3295 => x"77",
          3296 => x"94",
          3297 => x"ff",
          3298 => x"71",
          3299 => x"78",
          3300 => x"38",
          3301 => x"53",
          3302 => x"83",
          3303 => x"a8",
          3304 => x"51",
          3305 => x"78",
          3306 => x"08",
          3307 => x"76",
          3308 => x"08",
          3309 => x"0c",
          3310 => x"fd",
          3311 => x"56",
          3312 => x"ac",
          3313 => x"0d",
          3314 => x"0d",
          3315 => x"63",
          3316 => x"57",
          3317 => x"8f",
          3318 => x"52",
          3319 => x"b2",
          3320 => x"ac",
          3321 => x"d3",
          3322 => x"38",
          3323 => x"55",
          3324 => x"86",
          3325 => x"84",
          3326 => x"17",
          3327 => x"2a",
          3328 => x"51",
          3329 => x"56",
          3330 => x"83",
          3331 => x"39",
          3332 => x"18",
          3333 => x"83",
          3334 => x"0b",
          3335 => x"81",
          3336 => x"39",
          3337 => x"18",
          3338 => x"83",
          3339 => x"0b",
          3340 => x"82",
          3341 => x"39",
          3342 => x"18",
          3343 => x"83",
          3344 => x"0b",
          3345 => x"81",
          3346 => x"39",
          3347 => x"19",
          3348 => x"18",
          3349 => x"38",
          3350 => x"09",
          3351 => x"2e",
          3352 => x"94",
          3353 => x"83",
          3354 => x"56",
          3355 => x"38",
          3356 => x"22",
          3357 => x"89",
          3358 => x"55",
          3359 => x"38",
          3360 => x"88",
          3361 => x"74",
          3362 => x"52",
          3363 => x"b8",
          3364 => x"ac",
          3365 => x"39",
          3366 => x"52",
          3367 => x"a8",
          3368 => x"ac",
          3369 => x"80",
          3370 => x"38",
          3371 => x"fe",
          3372 => x"ff",
          3373 => x"38",
          3374 => x"0c",
          3375 => x"85",
          3376 => x"18",
          3377 => x"33",
          3378 => x"56",
          3379 => x"25",
          3380 => x"54",
          3381 => x"53",
          3382 => x"7d",
          3383 => x"52",
          3384 => x"3f",
          3385 => x"08",
          3386 => x"90",
          3387 => x"ff",
          3388 => x"90",
          3389 => x"17",
          3390 => x"51",
          3391 => x"81",
          3392 => x"80",
          3393 => x"38",
          3394 => x"08",
          3395 => x"2a",
          3396 => x"80",
          3397 => x"38",
          3398 => x"8a",
          3399 => x"56",
          3400 => x"27",
          3401 => x"7b",
          3402 => x"54",
          3403 => x"52",
          3404 => x"33",
          3405 => x"89",
          3406 => x"ac",
          3407 => x"38",
          3408 => x"78",
          3409 => x"7a",
          3410 => x"84",
          3411 => x"84",
          3412 => x"52",
          3413 => x"c8",
          3414 => x"17",
          3415 => x"06",
          3416 => x"18",
          3417 => x"2b",
          3418 => x"39",
          3419 => x"78",
          3420 => x"94",
          3421 => x"18",
          3422 => x"38",
          3423 => x"53",
          3424 => x"7d",
          3425 => x"52",
          3426 => x"3f",
          3427 => x"08",
          3428 => x"77",
          3429 => x"94",
          3430 => x"ff",
          3431 => x"71",
          3432 => x"78",
          3433 => x"38",
          3434 => x"53",
          3435 => x"17",
          3436 => x"06",
          3437 => x"51",
          3438 => x"90",
          3439 => x"80",
          3440 => x"90",
          3441 => x"76",
          3442 => x"17",
          3443 => x"1d",
          3444 => x"18",
          3445 => x"0c",
          3446 => x"58",
          3447 => x"74",
          3448 => x"38",
          3449 => x"8c",
          3450 => x"fc",
          3451 => x"17",
          3452 => x"07",
          3453 => x"18",
          3454 => x"75",
          3455 => x"0c",
          3456 => x"04",
          3457 => x"7b",
          3458 => x"05",
          3459 => x"58",
          3460 => x"81",
          3461 => x"57",
          3462 => x"08",
          3463 => x"90",
          3464 => x"86",
          3465 => x"06",
          3466 => x"74",
          3467 => x"98",
          3468 => x"2b",
          3469 => x"25",
          3470 => x"54",
          3471 => x"53",
          3472 => x"79",
          3473 => x"52",
          3474 => x"3f",
          3475 => x"d3",
          3476 => x"f6",
          3477 => x"33",
          3478 => x"55",
          3479 => x"34",
          3480 => x"52",
          3481 => x"c9",
          3482 => x"ac",
          3483 => x"d3",
          3484 => x"d4",
          3485 => x"08",
          3486 => x"a0",
          3487 => x"74",
          3488 => x"88",
          3489 => x"75",
          3490 => x"51",
          3491 => x"8c",
          3492 => x"9c",
          3493 => x"cb",
          3494 => x"b2",
          3495 => x"16",
          3496 => x"3f",
          3497 => x"16",
          3498 => x"3f",
          3499 => x"0b",
          3500 => x"79",
          3501 => x"3f",
          3502 => x"08",
          3503 => x"81",
          3504 => x"57",
          3505 => x"34",
          3506 => x"81",
          3507 => x"8b",
          3508 => x"fc",
          3509 => x"70",
          3510 => x"a8",
          3511 => x"ac",
          3512 => x"d3",
          3513 => x"38",
          3514 => x"05",
          3515 => x"ef",
          3516 => x"d3",
          3517 => x"81",
          3518 => x"87",
          3519 => x"ac",
          3520 => x"72",
          3521 => x"0c",
          3522 => x"04",
          3523 => x"85",
          3524 => x"9b",
          3525 => x"80",
          3526 => x"ac",
          3527 => x"38",
          3528 => x"08",
          3529 => x"34",
          3530 => x"81",
          3531 => x"84",
          3532 => x"ef",
          3533 => x"53",
          3534 => x"05",
          3535 => x"51",
          3536 => x"81",
          3537 => x"55",
          3538 => x"08",
          3539 => x"76",
          3540 => x"93",
          3541 => x"51",
          3542 => x"81",
          3543 => x"55",
          3544 => x"08",
          3545 => x"80",
          3546 => x"70",
          3547 => x"56",
          3548 => x"89",
          3549 => x"94",
          3550 => x"a7",
          3551 => x"05",
          3552 => x"2a",
          3553 => x"51",
          3554 => x"80",
          3555 => x"76",
          3556 => x"52",
          3557 => x"3f",
          3558 => x"08",
          3559 => x"83",
          3560 => x"74",
          3561 => x"81",
          3562 => x"85",
          3563 => x"d3",
          3564 => x"3d",
          3565 => x"3d",
          3566 => x"08",
          3567 => x"5b",
          3568 => x"34",
          3569 => x"3d",
          3570 => x"52",
          3571 => x"e5",
          3572 => x"d3",
          3573 => x"81",
          3574 => x"83",
          3575 => x"46",
          3576 => x"11",
          3577 => x"68",
          3578 => x"80",
          3579 => x"38",
          3580 => x"94",
          3581 => x"5b",
          3582 => x"51",
          3583 => x"81",
          3584 => x"57",
          3585 => x"08",
          3586 => x"6b",
          3587 => x"c5",
          3588 => x"d3",
          3589 => x"81",
          3590 => x"81",
          3591 => x"52",
          3592 => x"ab",
          3593 => x"ac",
          3594 => x"52",
          3595 => x"b2",
          3596 => x"ac",
          3597 => x"d3",
          3598 => x"ac",
          3599 => x"80",
          3600 => x"d6",
          3601 => x"d3",
          3602 => x"81",
          3603 => x"a4",
          3604 => x"7e",
          3605 => x"3f",
          3606 => x"08",
          3607 => x"38",
          3608 => x"51",
          3609 => x"81",
          3610 => x"57",
          3611 => x"08",
          3612 => x"38",
          3613 => x"09",
          3614 => x"38",
          3615 => x"81",
          3616 => x"3d",
          3617 => x"53",
          3618 => x"d9",
          3619 => x"93",
          3620 => x"12",
          3621 => x"51",
          3622 => x"56",
          3623 => x"8e",
          3624 => x"70",
          3625 => x"33",
          3626 => x"73",
          3627 => x"16",
          3628 => x"27",
          3629 => x"57",
          3630 => x"80",
          3631 => x"7d",
          3632 => x"a3",
          3633 => x"ff",
          3634 => x"57",
          3635 => x"81",
          3636 => x"34",
          3637 => x"ff",
          3638 => x"08",
          3639 => x"af",
          3640 => x"55",
          3641 => x"38",
          3642 => x"38",
          3643 => x"09",
          3644 => x"38",
          3645 => x"3d",
          3646 => x"59",
          3647 => x"80",
          3648 => x"dc",
          3649 => x"10",
          3650 => x"05",
          3651 => x"33",
          3652 => x"57",
          3653 => x"78",
          3654 => x"81",
          3655 => x"70",
          3656 => x"56",
          3657 => x"82",
          3658 => x"79",
          3659 => x"80",
          3660 => x"27",
          3661 => x"15",
          3662 => x"7a",
          3663 => x"5c",
          3664 => x"58",
          3665 => x"ee",
          3666 => x"70",
          3667 => x"34",
          3668 => x"77",
          3669 => x"57",
          3670 => x"a2",
          3671 => x"81",
          3672 => x"73",
          3673 => x"81",
          3674 => x"7b",
          3675 => x"38",
          3676 => x"76",
          3677 => x"0c",
          3678 => x"04",
          3679 => x"7e",
          3680 => x"fc",
          3681 => x"53",
          3682 => x"86",
          3683 => x"ac",
          3684 => x"d3",
          3685 => x"38",
          3686 => x"5a",
          3687 => x"86",
          3688 => x"83",
          3689 => x"17",
          3690 => x"94",
          3691 => x"33",
          3692 => x"70",
          3693 => x"56",
          3694 => x"38",
          3695 => x"58",
          3696 => x"56",
          3697 => x"19",
          3698 => x"7b",
          3699 => x"38",
          3700 => x"22",
          3701 => x"5b",
          3702 => x"7b",
          3703 => x"78",
          3704 => x"51",
          3705 => x"3f",
          3706 => x"08",
          3707 => x"54",
          3708 => x"55",
          3709 => x"3f",
          3710 => x"08",
          3711 => x"38",
          3712 => x"06",
          3713 => x"77",
          3714 => x"31",
          3715 => x"57",
          3716 => x"39",
          3717 => x"56",
          3718 => x"75",
          3719 => x"c9",
          3720 => x"d3",
          3721 => x"81",
          3722 => x"81",
          3723 => x"06",
          3724 => x"0b",
          3725 => x"82",
          3726 => x"39",
          3727 => x"08",
          3728 => x"81",
          3729 => x"81",
          3730 => x"34",
          3731 => x"ce",
          3732 => x"ac",
          3733 => x"0c",
          3734 => x"0c",
          3735 => x"81",
          3736 => x"78",
          3737 => x"38",
          3738 => x"94",
          3739 => x"94",
          3740 => x"18",
          3741 => x"2a",
          3742 => x"51",
          3743 => x"74",
          3744 => x"38",
          3745 => x"51",
          3746 => x"81",
          3747 => x"56",
          3748 => x"08",
          3749 => x"d3",
          3750 => x"b5",
          3751 => x"76",
          3752 => x"3f",
          3753 => x"08",
          3754 => x"2e",
          3755 => x"81",
          3756 => x"38",
          3757 => x"15",
          3758 => x"8b",
          3759 => x"91",
          3760 => x"55",
          3761 => x"75",
          3762 => x"77",
          3763 => x"98",
          3764 => x"08",
          3765 => x"0c",
          3766 => x"06",
          3767 => x"2e",
          3768 => x"52",
          3769 => x"bf",
          3770 => x"ac",
          3771 => x"82",
          3772 => x"34",
          3773 => x"a6",
          3774 => x"2a",
          3775 => x"08",
          3776 => x"17",
          3777 => x"08",
          3778 => x"94",
          3779 => x"18",
          3780 => x"33",
          3781 => x"55",
          3782 => x"34",
          3783 => x"83",
          3784 => x"74",
          3785 => x"f4",
          3786 => x"08",
          3787 => x"ec",
          3788 => x"33",
          3789 => x"56",
          3790 => x"25",
          3791 => x"54",
          3792 => x"53",
          3793 => x"7c",
          3794 => x"52",
          3795 => x"f1",
          3796 => x"ac",
          3797 => x"8a",
          3798 => x"91",
          3799 => x"55",
          3800 => x"17",
          3801 => x"06",
          3802 => x"18",
          3803 => x"7a",
          3804 => x"52",
          3805 => x"33",
          3806 => x"b6",
          3807 => x"d3",
          3808 => x"2e",
          3809 => x"0b",
          3810 => x"81",
          3811 => x"81",
          3812 => x"34",
          3813 => x"39",
          3814 => x"0c",
          3815 => x"81",
          3816 => x"8e",
          3817 => x"f9",
          3818 => x"56",
          3819 => x"80",
          3820 => x"38",
          3821 => x"3d",
          3822 => x"8a",
          3823 => x"51",
          3824 => x"81",
          3825 => x"55",
          3826 => x"08",
          3827 => x"77",
          3828 => x"52",
          3829 => x"9e",
          3830 => x"ac",
          3831 => x"d3",
          3832 => x"ca",
          3833 => x"33",
          3834 => x"55",
          3835 => x"24",
          3836 => x"16",
          3837 => x"2a",
          3838 => x"51",
          3839 => x"80",
          3840 => x"9c",
          3841 => x"77",
          3842 => x"3f",
          3843 => x"08",
          3844 => x"83",
          3845 => x"74",
          3846 => x"54",
          3847 => x"84",
          3848 => x"52",
          3849 => x"ba",
          3850 => x"ac",
          3851 => x"84",
          3852 => x"06",
          3853 => x"55",
          3854 => x"84",
          3855 => x"0c",
          3856 => x"81",
          3857 => x"89",
          3858 => x"fc",
          3859 => x"87",
          3860 => x"53",
          3861 => x"e4",
          3862 => x"d3",
          3863 => x"81",
          3864 => x"87",
          3865 => x"ac",
          3866 => x"72",
          3867 => x"0c",
          3868 => x"04",
          3869 => x"77",
          3870 => x"fc",
          3871 => x"53",
          3872 => x"8e",
          3873 => x"ac",
          3874 => x"d3",
          3875 => x"d1",
          3876 => x"38",
          3877 => x"08",
          3878 => x"c8",
          3879 => x"d3",
          3880 => x"bd",
          3881 => x"73",
          3882 => x"3f",
          3883 => x"08",
          3884 => x"ac",
          3885 => x"09",
          3886 => x"38",
          3887 => x"a1",
          3888 => x"73",
          3889 => x"3f",
          3890 => x"51",
          3891 => x"81",
          3892 => x"53",
          3893 => x"08",
          3894 => x"81",
          3895 => x"80",
          3896 => x"d3",
          3897 => x"3d",
          3898 => x"3d",
          3899 => x"80",
          3900 => x"70",
          3901 => x"52",
          3902 => x"3f",
          3903 => x"08",
          3904 => x"ac",
          3905 => x"63",
          3906 => x"d5",
          3907 => x"d3",
          3908 => x"81",
          3909 => x"a3",
          3910 => x"c7",
          3911 => x"98",
          3912 => x"73",
          3913 => x"38",
          3914 => x"39",
          3915 => x"8b",
          3916 => x"93",
          3917 => x"51",
          3918 => x"74",
          3919 => x"0c",
          3920 => x"04",
          3921 => x"61",
          3922 => x"80",
          3923 => x"ec",
          3924 => x"3d",
          3925 => x"3f",
          3926 => x"08",
          3927 => x"ac",
          3928 => x"38",
          3929 => x"73",
          3930 => x"08",
          3931 => x"55",
          3932 => x"74",
          3933 => x"90",
          3934 => x"0c",
          3935 => x"81",
          3936 => x"39",
          3937 => x"ca",
          3938 => x"70",
          3939 => x"57",
          3940 => x"09",
          3941 => x"c0",
          3942 => x"5d",
          3943 => x"90",
          3944 => x"51",
          3945 => x"3f",
          3946 => x"08",
          3947 => x"38",
          3948 => x"08",
          3949 => x"38",
          3950 => x"08",
          3951 => x"d3",
          3952 => x"80",
          3953 => x"81",
          3954 => x"58",
          3955 => x"14",
          3956 => x"c9",
          3957 => x"39",
          3958 => x"08",
          3959 => x"5a",
          3960 => x"55",
          3961 => x"77",
          3962 => x"7b",
          3963 => x"b9",
          3964 => x"d3",
          3965 => x"81",
          3966 => x"80",
          3967 => x"70",
          3968 => x"73",
          3969 => x"81",
          3970 => x"7a",
          3971 => x"51",
          3972 => x"3f",
          3973 => x"08",
          3974 => x"06",
          3975 => x"80",
          3976 => x"18",
          3977 => x"54",
          3978 => x"15",
          3979 => x"ff",
          3980 => x"81",
          3981 => x"f0",
          3982 => x"30",
          3983 => x"19",
          3984 => x"59",
          3985 => x"83",
          3986 => x"17",
          3987 => x"ff",
          3988 => x"7a",
          3989 => x"90",
          3990 => x"7a",
          3991 => x"81",
          3992 => x"73",
          3993 => x"78",
          3994 => x"0c",
          3995 => x"04",
          3996 => x"7a",
          3997 => x"05",
          3998 => x"58",
          3999 => x"81",
          4000 => x"57",
          4001 => x"08",
          4002 => x"18",
          4003 => x"80",
          4004 => x"76",
          4005 => x"39",
          4006 => x"70",
          4007 => x"81",
          4008 => x"56",
          4009 => x"80",
          4010 => x"38",
          4011 => x"8c",
          4012 => x"81",
          4013 => x"18",
          4014 => x"80",
          4015 => x"08",
          4016 => x"ff",
          4017 => x"81",
          4018 => x"57",
          4019 => x"19",
          4020 => x"39",
          4021 => x"52",
          4022 => x"b9",
          4023 => x"d3",
          4024 => x"d3",
          4025 => x"32",
          4026 => x"72",
          4027 => x"52",
          4028 => x"81",
          4029 => x"81",
          4030 => x"06",
          4031 => x"57",
          4032 => x"78",
          4033 => x"16",
          4034 => x"38",
          4035 => x"53",
          4036 => x"51",
          4037 => x"3f",
          4038 => x"08",
          4039 => x"08",
          4040 => x"90",
          4041 => x"c0",
          4042 => x"90",
          4043 => x"b9",
          4044 => x"2b",
          4045 => x"25",
          4046 => x"54",
          4047 => x"53",
          4048 => x"78",
          4049 => x"52",
          4050 => x"f5",
          4051 => x"ac",
          4052 => x"85",
          4053 => x"8c",
          4054 => x"33",
          4055 => x"55",
          4056 => x"34",
          4057 => x"89",
          4058 => x"19",
          4059 => x"83",
          4060 => x"75",
          4061 => x"0c",
          4062 => x"04",
          4063 => x"81",
          4064 => x"ff",
          4065 => x"82",
          4066 => x"ff",
          4067 => x"a0",
          4068 => x"b2",
          4069 => x"ac",
          4070 => x"d3",
          4071 => x"d3",
          4072 => x"f4",
          4073 => x"b3",
          4074 => x"6f",
          4075 => x"d4",
          4076 => x"c2",
          4077 => x"ac",
          4078 => x"f8",
          4079 => x"96",
          4080 => x"82",
          4081 => x"80",
          4082 => x"70",
          4083 => x"81",
          4084 => x"55",
          4085 => x"83",
          4086 => x"75",
          4087 => x"81",
          4088 => x"ff",
          4089 => x"02",
          4090 => x"33",
          4091 => x"55",
          4092 => x"25",
          4093 => x"56",
          4094 => x"80",
          4095 => x"81",
          4096 => x"80",
          4097 => x"87",
          4098 => x"e7",
          4099 => x"77",
          4100 => x"3f",
          4101 => x"08",
          4102 => x"80",
          4103 => x"70",
          4104 => x"81",
          4105 => x"56",
          4106 => x"2e",
          4107 => x"81",
          4108 => x"ff",
          4109 => x"87",
          4110 => x"94",
          4111 => x"2e",
          4112 => x"81",
          4113 => x"ff",
          4114 => x"77",
          4115 => x"81",
          4116 => x"ff",
          4117 => x"80",
          4118 => x"70",
          4119 => x"82",
          4120 => x"ac",
          4121 => x"d3",
          4122 => x"87",
          4123 => x"ac",
          4124 => x"51",
          4125 => x"81",
          4126 => x"56",
          4127 => x"08",
          4128 => x"56",
          4129 => x"70",
          4130 => x"07",
          4131 => x"06",
          4132 => x"75",
          4133 => x"81",
          4134 => x"ff",
          4135 => x"9f",
          4136 => x"51",
          4137 => x"81",
          4138 => x"81",
          4139 => x"30",
          4140 => x"ac",
          4141 => x"25",
          4142 => x"7b",
          4143 => x"72",
          4144 => x"51",
          4145 => x"80",
          4146 => x"81",
          4147 => x"ff",
          4148 => x"80",
          4149 => x"9f",
          4150 => x"51",
          4151 => x"3f",
          4152 => x"08",
          4153 => x"38",
          4154 => x"b4",
          4155 => x"d3",
          4156 => x"81",
          4157 => x"ff",
          4158 => x"75",
          4159 => x"0c",
          4160 => x"04",
          4161 => x"82",
          4162 => x"c0",
          4163 => x"3d",
          4164 => x"3f",
          4165 => x"08",
          4166 => x"ac",
          4167 => x"38",
          4168 => x"52",
          4169 => x"05",
          4170 => x"3f",
          4171 => x"08",
          4172 => x"ac",
          4173 => x"88",
          4174 => x"2e",
          4175 => x"82",
          4176 => x"80",
          4177 => x"70",
          4178 => x"81",
          4179 => x"56",
          4180 => x"83",
          4181 => x"74",
          4182 => x"81",
          4183 => x"38",
          4184 => x"52",
          4185 => x"05",
          4186 => x"dc",
          4187 => x"ac",
          4188 => x"55",
          4189 => x"08",
          4190 => x"81",
          4191 => x"87",
          4192 => x"2e",
          4193 => x"83",
          4194 => x"75",
          4195 => x"81",
          4196 => x"81",
          4197 => x"b2",
          4198 => x"81",
          4199 => x"52",
          4200 => x"bd",
          4201 => x"d3",
          4202 => x"81",
          4203 => x"81",
          4204 => x"53",
          4205 => x"18",
          4206 => x"fa",
          4207 => x"ae",
          4208 => x"34",
          4209 => x"0b",
          4210 => x"76",
          4211 => x"18",
          4212 => x"8f",
          4213 => x"b4",
          4214 => x"51",
          4215 => x"a0",
          4216 => x"52",
          4217 => x"51",
          4218 => x"3f",
          4219 => x"0b",
          4220 => x"34",
          4221 => x"d4",
          4222 => x"51",
          4223 => x"77",
          4224 => x"83",
          4225 => x"3d",
          4226 => x"c5",
          4227 => x"d3",
          4228 => x"81",
          4229 => x"af",
          4230 => x"63",
          4231 => x"ff",
          4232 => x"75",
          4233 => x"77",
          4234 => x"3f",
          4235 => x"0b",
          4236 => x"77",
          4237 => x"83",
          4238 => x"51",
          4239 => x"3f",
          4240 => x"08",
          4241 => x"80",
          4242 => x"98",
          4243 => x"51",
          4244 => x"3f",
          4245 => x"ac",
          4246 => x"0d",
          4247 => x"0d",
          4248 => x"05",
          4249 => x"3f",
          4250 => x"3d",
          4251 => x"52",
          4252 => x"d0",
          4253 => x"d3",
          4254 => x"81",
          4255 => x"82",
          4256 => x"4c",
          4257 => x"52",
          4258 => x"05",
          4259 => x"3f",
          4260 => x"08",
          4261 => x"ac",
          4262 => x"38",
          4263 => x"05",
          4264 => x"06",
          4265 => x"2e",
          4266 => x"55",
          4267 => x"38",
          4268 => x"3d",
          4269 => x"3d",
          4270 => x"51",
          4271 => x"3f",
          4272 => x"3d",
          4273 => x"91",
          4274 => x"54",
          4275 => x"3f",
          4276 => x"52",
          4277 => x"9e",
          4278 => x"ac",
          4279 => x"d3",
          4280 => x"38",
          4281 => x"09",
          4282 => x"38",
          4283 => x"a1",
          4284 => x"83",
          4285 => x"74",
          4286 => x"81",
          4287 => x"38",
          4288 => x"a8",
          4289 => x"ec",
          4290 => x"ac",
          4291 => x"d3",
          4292 => x"c4",
          4293 => x"93",
          4294 => x"ff",
          4295 => x"8d",
          4296 => x"ac",
          4297 => x"ab",
          4298 => x"17",
          4299 => x"33",
          4300 => x"70",
          4301 => x"55",
          4302 => x"38",
          4303 => x"54",
          4304 => x"34",
          4305 => x"0b",
          4306 => x"8b",
          4307 => x"84",
          4308 => x"06",
          4309 => x"73",
          4310 => x"db",
          4311 => x"2e",
          4312 => x"75",
          4313 => x"ff",
          4314 => x"81",
          4315 => x"52",
          4316 => x"b0",
          4317 => x"55",
          4318 => x"08",
          4319 => x"38",
          4320 => x"08",
          4321 => x"ff",
          4322 => x"81",
          4323 => x"80",
          4324 => x"55",
          4325 => x"08",
          4326 => x"16",
          4327 => x"ae",
          4328 => x"06",
          4329 => x"53",
          4330 => x"51",
          4331 => x"3f",
          4332 => x"0b",
          4333 => x"74",
          4334 => x"3d",
          4335 => x"c3",
          4336 => x"d3",
          4337 => x"81",
          4338 => x"8c",
          4339 => x"ff",
          4340 => x"81",
          4341 => x"55",
          4342 => x"ac",
          4343 => x"0d",
          4344 => x"0d",
          4345 => x"05",
          4346 => x"05",
          4347 => x"33",
          4348 => x"53",
          4349 => x"05",
          4350 => x"51",
          4351 => x"81",
          4352 => x"55",
          4353 => x"08",
          4354 => x"78",
          4355 => x"95",
          4356 => x"51",
          4357 => x"81",
          4358 => x"55",
          4359 => x"08",
          4360 => x"80",
          4361 => x"81",
          4362 => x"73",
          4363 => x"38",
          4364 => x"aa",
          4365 => x"06",
          4366 => x"8b",
          4367 => x"06",
          4368 => x"07",
          4369 => x"56",
          4370 => x"34",
          4371 => x"0b",
          4372 => x"78",
          4373 => x"a0",
          4374 => x"ac",
          4375 => x"81",
          4376 => x"95",
          4377 => x"ee",
          4378 => x"56",
          4379 => x"3d",
          4380 => x"95",
          4381 => x"ce",
          4382 => x"ac",
          4383 => x"d3",
          4384 => x"d3",
          4385 => x"64",
          4386 => x"d4",
          4387 => x"e6",
          4388 => x"ac",
          4389 => x"d3",
          4390 => x"38",
          4391 => x"05",
          4392 => x"06",
          4393 => x"2e",
          4394 => x"55",
          4395 => x"86",
          4396 => x"17",
          4397 => x"2b",
          4398 => x"57",
          4399 => x"05",
          4400 => x"9f",
          4401 => x"81",
          4402 => x"34",
          4403 => x"ac",
          4404 => x"d3",
          4405 => x"74",
          4406 => x"0c",
          4407 => x"04",
          4408 => x"69",
          4409 => x"80",
          4410 => x"d0",
          4411 => x"3d",
          4412 => x"3f",
          4413 => x"08",
          4414 => x"08",
          4415 => x"d3",
          4416 => x"80",
          4417 => x"70",
          4418 => x"2a",
          4419 => x"57",
          4420 => x"74",
          4421 => x"f6",
          4422 => x"80",
          4423 => x"8d",
          4424 => x"54",
          4425 => x"3f",
          4426 => x"08",
          4427 => x"ac",
          4428 => x"38",
          4429 => x"51",
          4430 => x"3f",
          4431 => x"08",
          4432 => x"ac",
          4433 => x"81",
          4434 => x"81",
          4435 => x"65",
          4436 => x"79",
          4437 => x"7a",
          4438 => x"55",
          4439 => x"34",
          4440 => x"8a",
          4441 => x"38",
          4442 => x"80",
          4443 => x"80",
          4444 => x"ff",
          4445 => x"70",
          4446 => x"58",
          4447 => x"e8",
          4448 => x"2e",
          4449 => x"86",
          4450 => x"34",
          4451 => x"30",
          4452 => x"80",
          4453 => x"70",
          4454 => x"2a",
          4455 => x"56",
          4456 => x"80",
          4457 => x"7b",
          4458 => x"53",
          4459 => x"81",
          4460 => x"ac",
          4461 => x"d3",
          4462 => x"38",
          4463 => x"51",
          4464 => x"58",
          4465 => x"8b",
          4466 => x"58",
          4467 => x"83",
          4468 => x"7b",
          4469 => x"51",
          4470 => x"3f",
          4471 => x"08",
          4472 => x"81",
          4473 => x"98",
          4474 => x"e8",
          4475 => x"53",
          4476 => x"b8",
          4477 => x"3d",
          4478 => x"3f",
          4479 => x"08",
          4480 => x"ac",
          4481 => x"38",
          4482 => x"52",
          4483 => x"bc",
          4484 => x"a7",
          4485 => x"6b",
          4486 => x"52",
          4487 => x"9f",
          4488 => x"b5",
          4489 => x"6b",
          4490 => x"70",
          4491 => x"52",
          4492 => x"fe",
          4493 => x"ac",
          4494 => x"a2",
          4495 => x"33",
          4496 => x"54",
          4497 => x"3f",
          4498 => x"08",
          4499 => x"38",
          4500 => x"74",
          4501 => x"05",
          4502 => x"39",
          4503 => x"9f",
          4504 => x"99",
          4505 => x"e0",
          4506 => x"ff",
          4507 => x"54",
          4508 => x"27",
          4509 => x"ba",
          4510 => x"56",
          4511 => x"a3",
          4512 => x"81",
          4513 => x"ff",
          4514 => x"81",
          4515 => x"93",
          4516 => x"76",
          4517 => x"76",
          4518 => x"38",
          4519 => x"77",
          4520 => x"86",
          4521 => x"39",
          4522 => x"27",
          4523 => x"3d",
          4524 => x"bc",
          4525 => x"2a",
          4526 => x"75",
          4527 => x"57",
          4528 => x"05",
          4529 => x"54",
          4530 => x"81",
          4531 => x"33",
          4532 => x"73",
          4533 => x"cd",
          4534 => x"33",
          4535 => x"73",
          4536 => x"81",
          4537 => x"80",
          4538 => x"02",
          4539 => x"78",
          4540 => x"51",
          4541 => x"73",
          4542 => x"81",
          4543 => x"ff",
          4544 => x"80",
          4545 => x"76",
          4546 => x"51",
          4547 => x"2e",
          4548 => x"5f",
          4549 => x"52",
          4550 => x"52",
          4551 => x"c2",
          4552 => x"ac",
          4553 => x"d3",
          4554 => x"a1",
          4555 => x"74",
          4556 => x"82",
          4557 => x"ac",
          4558 => x"d3",
          4559 => x"38",
          4560 => x"91",
          4561 => x"9a",
          4562 => x"05",
          4563 => x"ff",
          4564 => x"86",
          4565 => x"e5",
          4566 => x"54",
          4567 => x"15",
          4568 => x"ff",
          4569 => x"81",
          4570 => x"54",
          4571 => x"81",
          4572 => x"84",
          4573 => x"06",
          4574 => x"80",
          4575 => x"2e",
          4576 => x"81",
          4577 => x"d4",
          4578 => x"b6",
          4579 => x"d3",
          4580 => x"81",
          4581 => x"b5",
          4582 => x"81",
          4583 => x"52",
          4584 => x"a4",
          4585 => x"54",
          4586 => x"15",
          4587 => x"9a",
          4588 => x"05",
          4589 => x"ff",
          4590 => x"77",
          4591 => x"83",
          4592 => x"51",
          4593 => x"3f",
          4594 => x"08",
          4595 => x"74",
          4596 => x"0c",
          4597 => x"04",
          4598 => x"61",
          4599 => x"05",
          4600 => x"33",
          4601 => x"05",
          4602 => x"5e",
          4603 => x"a2",
          4604 => x"ac",
          4605 => x"d3",
          4606 => x"38",
          4607 => x"57",
          4608 => x"86",
          4609 => x"82",
          4610 => x"80",
          4611 => x"8c",
          4612 => x"38",
          4613 => x"70",
          4614 => x"81",
          4615 => x"55",
          4616 => x"87",
          4617 => x"39",
          4618 => x"89",
          4619 => x"81",
          4620 => x"8a",
          4621 => x"89",
          4622 => x"7d",
          4623 => x"54",
          4624 => x"3f",
          4625 => x"06",
          4626 => x"72",
          4627 => x"81",
          4628 => x"05",
          4629 => x"08",
          4630 => x"55",
          4631 => x"81",
          4632 => x"38",
          4633 => x"79",
          4634 => x"82",
          4635 => x"56",
          4636 => x"74",
          4637 => x"ff",
          4638 => x"81",
          4639 => x"81",
          4640 => x"56",
          4641 => x"08",
          4642 => x"38",
          4643 => x"81",
          4644 => x"38",
          4645 => x"ff",
          4646 => x"8b",
          4647 => x"5a",
          4648 => x"91",
          4649 => x"74",
          4650 => x"74",
          4651 => x"81",
          4652 => x"87",
          4653 => x"86",
          4654 => x"2e",
          4655 => x"7e",
          4656 => x"80",
          4657 => x"81",
          4658 => x"81",
          4659 => x"06",
          4660 => x"54",
          4661 => x"52",
          4662 => x"a7",
          4663 => x"d3",
          4664 => x"81",
          4665 => x"91",
          4666 => x"16",
          4667 => x"56",
          4668 => x"38",
          4669 => x"1d",
          4670 => x"c2",
          4671 => x"8c",
          4672 => x"7b",
          4673 => x"38",
          4674 => x"0c",
          4675 => x"0c",
          4676 => x"80",
          4677 => x"73",
          4678 => x"7f",
          4679 => x"fe",
          4680 => x"90",
          4681 => x"26",
          4682 => x"15",
          4683 => x"90",
          4684 => x"84",
          4685 => x"07",
          4686 => x"84",
          4687 => x"54",
          4688 => x"ac",
          4689 => x"0d",
          4690 => x"0d",
          4691 => x"05",
          4692 => x"33",
          4693 => x"5e",
          4694 => x"d3",
          4695 => x"ac",
          4696 => x"57",
          4697 => x"d3",
          4698 => x"8c",
          4699 => x"d3",
          4700 => x"10",
          4701 => x"05",
          4702 => x"80",
          4703 => x"74",
          4704 => x"75",
          4705 => x"ff",
          4706 => x"52",
          4707 => x"99",
          4708 => x"d3",
          4709 => x"ff",
          4710 => x"06",
          4711 => x"57",
          4712 => x"38",
          4713 => x"70",
          4714 => x"55",
          4715 => x"8c",
          4716 => x"3d",
          4717 => x"83",
          4718 => x"ff",
          4719 => x"81",
          4720 => x"98",
          4721 => x"2e",
          4722 => x"82",
          4723 => x"8c",
          4724 => x"05",
          4725 => x"74",
          4726 => x"38",
          4727 => x"80",
          4728 => x"2e",
          4729 => x"78",
          4730 => x"77",
          4731 => x"26",
          4732 => x"18",
          4733 => x"74",
          4734 => x"38",
          4735 => x"be",
          4736 => x"77",
          4737 => x"98",
          4738 => x"ac",
          4739 => x"54",
          4740 => x"58",
          4741 => x"3f",
          4742 => x"08",
          4743 => x"ac",
          4744 => x"30",
          4745 => x"80",
          4746 => x"ac",
          4747 => x"81",
          4748 => x"07",
          4749 => x"07",
          4750 => x"58",
          4751 => x"57",
          4752 => x"38",
          4753 => x"05",
          4754 => x"79",
          4755 => x"cb",
          4756 => x"81",
          4757 => x"8a",
          4758 => x"83",
          4759 => x"06",
          4760 => x"44",
          4761 => x"09",
          4762 => x"38",
          4763 => x"57",
          4764 => x"8a",
          4765 => x"64",
          4766 => x"57",
          4767 => x"27",
          4768 => x"93",
          4769 => x"80",
          4770 => x"38",
          4771 => x"70",
          4772 => x"55",
          4773 => x"95",
          4774 => x"06",
          4775 => x"2e",
          4776 => x"81",
          4777 => x"85",
          4778 => x"8f",
          4779 => x"06",
          4780 => x"82",
          4781 => x"2e",
          4782 => x"77",
          4783 => x"2e",
          4784 => x"80",
          4785 => x"b4",
          4786 => x"2a",
          4787 => x"81",
          4788 => x"80",
          4789 => x"52",
          4790 => x"74",
          4791 => x"38",
          4792 => x"98",
          4793 => x"79",
          4794 => x"18",
          4795 => x"57",
          4796 => x"80",
          4797 => x"76",
          4798 => x"38",
          4799 => x"51",
          4800 => x"3f",
          4801 => x"08",
          4802 => x"08",
          4803 => x"7f",
          4804 => x"52",
          4805 => x"88",
          4806 => x"ac",
          4807 => x"5b",
          4808 => x"80",
          4809 => x"43",
          4810 => x"0a",
          4811 => x"8b",
          4812 => x"89",
          4813 => x"b4",
          4814 => x"2a",
          4815 => x"81",
          4816 => x"f0",
          4817 => x"52",
          4818 => x"74",
          4819 => x"38",
          4820 => x"98",
          4821 => x"79",
          4822 => x"18",
          4823 => x"57",
          4824 => x"80",
          4825 => x"76",
          4826 => x"38",
          4827 => x"51",
          4828 => x"3f",
          4829 => x"08",
          4830 => x"57",
          4831 => x"08",
          4832 => x"92",
          4833 => x"81",
          4834 => x"83",
          4835 => x"72",
          4836 => x"51",
          4837 => x"52",
          4838 => x"05",
          4839 => x"80",
          4840 => x"ac",
          4841 => x"7e",
          4842 => x"80",
          4843 => x"f2",
          4844 => x"d3",
          4845 => x"ff",
          4846 => x"63",
          4847 => x"64",
          4848 => x"ff",
          4849 => x"70",
          4850 => x"31",
          4851 => x"57",
          4852 => x"2e",
          4853 => x"89",
          4854 => x"60",
          4855 => x"84",
          4856 => x"5c",
          4857 => x"16",
          4858 => x"51",
          4859 => x"26",
          4860 => x"65",
          4861 => x"31",
          4862 => x"64",
          4863 => x"fe",
          4864 => x"81",
          4865 => x"56",
          4866 => x"09",
          4867 => x"38",
          4868 => x"08",
          4869 => x"26",
          4870 => x"89",
          4871 => x"2a",
          4872 => x"97",
          4873 => x"87",
          4874 => x"82",
          4875 => x"06",
          4876 => x"83",
          4877 => x"27",
          4878 => x"8f",
          4879 => x"55",
          4880 => x"26",
          4881 => x"58",
          4882 => x"7c",
          4883 => x"06",
          4884 => x"2e",
          4885 => x"42",
          4886 => x"77",
          4887 => x"19",
          4888 => x"78",
          4889 => x"38",
          4890 => x"d2",
          4891 => x"f5",
          4892 => x"77",
          4893 => x"19",
          4894 => x"78",
          4895 => x"38",
          4896 => x"ba",
          4897 => x"61",
          4898 => x"81",
          4899 => x"61",
          4900 => x"f5",
          4901 => x"55",
          4902 => x"86",
          4903 => x"53",
          4904 => x"51",
          4905 => x"3f",
          4906 => x"bb",
          4907 => x"51",
          4908 => x"3f",
          4909 => x"1f",
          4910 => x"89",
          4911 => x"8d",
          4912 => x"83",
          4913 => x"52",
          4914 => x"ff",
          4915 => x"81",
          4916 => x"34",
          4917 => x"70",
          4918 => x"2a",
          4919 => x"54",
          4920 => x"1f",
          4921 => x"dd",
          4922 => x"ff",
          4923 => x"38",
          4924 => x"05",
          4925 => x"1f",
          4926 => x"c9",
          4927 => x"65",
          4928 => x"51",
          4929 => x"3f",
          4930 => x"05",
          4931 => x"98",
          4932 => x"98",
          4933 => x"ff",
          4934 => x"51",
          4935 => x"3f",
          4936 => x"1f",
          4937 => x"bb",
          4938 => x"2e",
          4939 => x"80",
          4940 => x"88",
          4941 => x"80",
          4942 => x"ff",
          4943 => x"7b",
          4944 => x"51",
          4945 => x"3f",
          4946 => x"1f",
          4947 => x"93",
          4948 => x"b0",
          4949 => x"97",
          4950 => x"52",
          4951 => x"ff",
          4952 => x"ff",
          4953 => x"c0",
          4954 => x"7f",
          4955 => x"34",
          4956 => x"bb",
          4957 => x"c7",
          4958 => x"98",
          4959 => x"39",
          4960 => x"0a",
          4961 => x"51",
          4962 => x"3f",
          4963 => x"ff",
          4964 => x"1f",
          4965 => x"ad",
          4966 => x"7f",
          4967 => x"a9",
          4968 => x"34",
          4969 => x"bb",
          4970 => x"1f",
          4971 => x"e2",
          4972 => x"d5",
          4973 => x"1f",
          4974 => x"89",
          4975 => x"63",
          4976 => x"79",
          4977 => x"f9",
          4978 => x"81",
          4979 => x"83",
          4980 => x"83",
          4981 => x"06",
          4982 => x"81",
          4983 => x"05",
          4984 => x"79",
          4985 => x"d9",
          4986 => x"80",
          4987 => x"ff",
          4988 => x"84",
          4989 => x"d2",
          4990 => x"ff",
          4991 => x"86",
          4992 => x"f2",
          4993 => x"1f",
          4994 => x"d7",
          4995 => x"52",
          4996 => x"51",
          4997 => x"3f",
          4998 => x"ec",
          4999 => x"96",
          5000 => x"d4",
          5001 => x"fe",
          5002 => x"96",
          5003 => x"54",
          5004 => x"53",
          5005 => x"51",
          5006 => x"3f",
          5007 => x"81",
          5008 => x"52",
          5009 => x"92",
          5010 => x"53",
          5011 => x"51",
          5012 => x"3f",
          5013 => x"5b",
          5014 => x"09",
          5015 => x"38",
          5016 => x"51",
          5017 => x"3f",
          5018 => x"1f",
          5019 => x"f3",
          5020 => x"52",
          5021 => x"ff",
          5022 => x"95",
          5023 => x"ff",
          5024 => x"81",
          5025 => x"f8",
          5026 => x"7e",
          5027 => x"d3",
          5028 => x"60",
          5029 => x"26",
          5030 => x"57",
          5031 => x"53",
          5032 => x"51",
          5033 => x"3f",
          5034 => x"08",
          5035 => x"7d",
          5036 => x"7e",
          5037 => x"fe",
          5038 => x"75",
          5039 => x"56",
          5040 => x"81",
          5041 => x"80",
          5042 => x"38",
          5043 => x"83",
          5044 => x"62",
          5045 => x"74",
          5046 => x"38",
          5047 => x"54",
          5048 => x"52",
          5049 => x"91",
          5050 => x"d3",
          5051 => x"c8",
          5052 => x"75",
          5053 => x"56",
          5054 => x"8c",
          5055 => x"2e",
          5056 => x"57",
          5057 => x"ff",
          5058 => x"84",
          5059 => x"2e",
          5060 => x"57",
          5061 => x"81",
          5062 => x"80",
          5063 => x"53",
          5064 => x"51",
          5065 => x"3f",
          5066 => x"52",
          5067 => x"51",
          5068 => x"3f",
          5069 => x"56",
          5070 => x"81",
          5071 => x"34",
          5072 => x"17",
          5073 => x"17",
          5074 => x"17",
          5075 => x"05",
          5076 => x"c1",
          5077 => x"fe",
          5078 => x"fe",
          5079 => x"34",
          5080 => x"08",
          5081 => x"07",
          5082 => x"17",
          5083 => x"ac",
          5084 => x"34",
          5085 => x"c6",
          5086 => x"93",
          5087 => x"52",
          5088 => x"51",
          5089 => x"3f",
          5090 => x"53",
          5091 => x"51",
          5092 => x"3f",
          5093 => x"d3",
          5094 => x"38",
          5095 => x"52",
          5096 => x"91",
          5097 => x"57",
          5098 => x"08",
          5099 => x"39",
          5100 => x"39",
          5101 => x"39",
          5102 => x"39",
          5103 => x"81",
          5104 => x"98",
          5105 => x"ff",
          5106 => x"52",
          5107 => x"81",
          5108 => x"10",
          5109 => x"9c",
          5110 => x"08",
          5111 => x"dc",
          5112 => x"a9",
          5113 => x"39",
          5114 => x"51",
          5115 => x"3f",
          5116 => x"81",
          5117 => x"ff",
          5118 => x"81",
          5119 => x"c2",
          5120 => x"80",
          5121 => x"b3",
          5122 => x"a0",
          5123 => x"fd",
          5124 => x"39",
          5125 => x"51",
          5126 => x"3f",
          5127 => x"81",
          5128 => x"fe",
          5129 => x"81",
          5130 => x"c2",
          5131 => x"ff",
          5132 => x"87",
          5133 => x"ec",
          5134 => x"d1",
          5135 => x"39",
          5136 => x"51",
          5137 => x"3f",
          5138 => x"81",
          5139 => x"fe",
          5140 => x"80",
          5141 => x"c3",
          5142 => x"ff",
          5143 => x"db",
          5144 => x"cc",
          5145 => x"a5",
          5146 => x"39",
          5147 => x"51",
          5148 => x"3f",
          5149 => x"81",
          5150 => x"fe",
          5151 => x"bb",
          5152 => x"ac",
          5153 => x"85",
          5154 => x"81",
          5155 => x"fe",
          5156 => x"a7",
          5157 => x"d8",
          5158 => x"f1",
          5159 => x"81",
          5160 => x"fe",
          5161 => x"93",
          5162 => x"88",
          5163 => x"dd",
          5164 => x"81",
          5165 => x"fe",
          5166 => x"83",
          5167 => x"fb",
          5168 => x"79",
          5169 => x"87",
          5170 => x"38",
          5171 => x"87",
          5172 => x"fe",
          5173 => x"81",
          5174 => x"55",
          5175 => x"e8",
          5176 => x"fe",
          5177 => x"81",
          5178 => x"52",
          5179 => x"e8",
          5180 => x"d3",
          5181 => x"74",
          5182 => x"75",
          5183 => x"a4",
          5184 => x"83",
          5185 => x"0d",
          5186 => x"3d",
          5187 => x"3d",
          5188 => x"3d",
          5189 => x"05",
          5190 => x"33",
          5191 => x"70",
          5192 => x"25",
          5193 => x"27",
          5194 => x"5a",
          5195 => x"93",
          5196 => x"87",
          5197 => x"77",
          5198 => x"3d",
          5199 => x"51",
          5200 => x"3f",
          5201 => x"08",
          5202 => x"ac",
          5203 => x"81",
          5204 => x"87",
          5205 => x"0c",
          5206 => x"08",
          5207 => x"3d",
          5208 => x"55",
          5209 => x"53",
          5210 => x"d8",
          5211 => x"f2",
          5212 => x"ac",
          5213 => x"d3",
          5214 => x"38",
          5215 => x"89",
          5216 => x"7b",
          5217 => x"d5",
          5218 => x"3d",
          5219 => x"51",
          5220 => x"77",
          5221 => x"07",
          5222 => x"30",
          5223 => x"72",
          5224 => x"51",
          5225 => x"2e",
          5226 => x"c5",
          5227 => x"c0",
          5228 => x"52",
          5229 => x"87",
          5230 => x"74",
          5231 => x"0c",
          5232 => x"0d",
          5233 => x"0d",
          5234 => x"33",
          5235 => x"57",
          5236 => x"7b",
          5237 => x"fe",
          5238 => x"d3",
          5239 => x"38",
          5240 => x"88",
          5241 => x"2e",
          5242 => x"39",
          5243 => x"54",
          5244 => x"53",
          5245 => x"51",
          5246 => x"d3",
          5247 => x"83",
          5248 => x"78",
          5249 => x"0c",
          5250 => x"04",
          5251 => x"02",
          5252 => x"81",
          5253 => x"81",
          5254 => x"56",
          5255 => x"3f",
          5256 => x"70",
          5257 => x"fe",
          5258 => x"81",
          5259 => x"81",
          5260 => x"81",
          5261 => x"81",
          5262 => x"ff",
          5263 => x"75",
          5264 => x"38",
          5265 => x"3f",
          5266 => x"04",
          5267 => x"87",
          5268 => x"08",
          5269 => x"ff",
          5270 => x"fe",
          5271 => x"81",
          5272 => x"fe",
          5273 => x"80",
          5274 => x"f1",
          5275 => x"2a",
          5276 => x"51",
          5277 => x"2e",
          5278 => x"51",
          5279 => x"3f",
          5280 => x"51",
          5281 => x"3f",
          5282 => x"ee",
          5283 => x"82",
          5284 => x"06",
          5285 => x"80",
          5286 => x"81",
          5287 => x"bd",
          5288 => x"c4",
          5289 => x"b3",
          5290 => x"fe",
          5291 => x"72",
          5292 => x"81",
          5293 => x"71",
          5294 => x"38",
          5295 => x"ee",
          5296 => x"c6",
          5297 => x"f0",
          5298 => x"51",
          5299 => x"3f",
          5300 => x"70",
          5301 => x"52",
          5302 => x"95",
          5303 => x"fe",
          5304 => x"81",
          5305 => x"fe",
          5306 => x"80",
          5307 => x"ed",
          5308 => x"2a",
          5309 => x"51",
          5310 => x"2e",
          5311 => x"51",
          5312 => x"3f",
          5313 => x"51",
          5314 => x"3f",
          5315 => x"ed",
          5316 => x"86",
          5317 => x"06",
          5318 => x"80",
          5319 => x"81",
          5320 => x"b9",
          5321 => x"90",
          5322 => x"af",
          5323 => x"fe",
          5324 => x"72",
          5325 => x"81",
          5326 => x"71",
          5327 => x"38",
          5328 => x"ed",
          5329 => x"c7",
          5330 => x"ef",
          5331 => x"51",
          5332 => x"3f",
          5333 => x"70",
          5334 => x"52",
          5335 => x"95",
          5336 => x"fe",
          5337 => x"81",
          5338 => x"fe",
          5339 => x"80",
          5340 => x"e9",
          5341 => x"a8",
          5342 => x"0d",
          5343 => x"0d",
          5344 => x"70",
          5345 => x"74",
          5346 => x"ed",
          5347 => x"74",
          5348 => x"14",
          5349 => x"e1",
          5350 => x"55",
          5351 => x"54",
          5352 => x"2e",
          5353 => x"54",
          5354 => x"9f",
          5355 => x"51",
          5356 => x"38",
          5357 => x"72",
          5358 => x"81",
          5359 => x"80",
          5360 => x"05",
          5361 => x"56",
          5362 => x"81",
          5363 => x"77",
          5364 => x"08",
          5365 => x"e6",
          5366 => x"d3",
          5367 => x"38",
          5368 => x"53",
          5369 => x"ff",
          5370 => x"16",
          5371 => x"06",
          5372 => x"76",
          5373 => x"ff",
          5374 => x"d3",
          5375 => x"3d",
          5376 => x"3d",
          5377 => x"81",
          5378 => x"71",
          5379 => x"5c",
          5380 => x"52",
          5381 => x"84",
          5382 => x"d3",
          5383 => x"ff",
          5384 => x"7c",
          5385 => x"06",
          5386 => x"c7",
          5387 => x"3d",
          5388 => x"fe",
          5389 => x"7b",
          5390 => x"ea",
          5391 => x"ff",
          5392 => x"81",
          5393 => x"5a",
          5394 => x"8b",
          5395 => x"fc",
          5396 => x"b3",
          5397 => x"81",
          5398 => x"81",
          5399 => x"fe",
          5400 => x"96",
          5401 => x"59",
          5402 => x"54",
          5403 => x"78",
          5404 => x"a4",
          5405 => x"61",
          5406 => x"e5",
          5407 => x"fe",
          5408 => x"fd",
          5409 => x"d3",
          5410 => x"2b",
          5411 => x"51",
          5412 => x"87",
          5413 => x"38",
          5414 => x"81",
          5415 => x"59",
          5416 => x"b4",
          5417 => x"11",
          5418 => x"05",
          5419 => x"e2",
          5420 => x"ac",
          5421 => x"81",
          5422 => x"fe",
          5423 => x"ff",
          5424 => x"3d",
          5425 => x"53",
          5426 => x"51",
          5427 => x"3f",
          5428 => x"08",
          5429 => x"38",
          5430 => x"83",
          5431 => x"02",
          5432 => x"52",
          5433 => x"05",
          5434 => x"82",
          5435 => x"d3",
          5436 => x"ff",
          5437 => x"8e",
          5438 => x"c8",
          5439 => x"8d",
          5440 => x"fe",
          5441 => x"c8",
          5442 => x"f6",
          5443 => x"cb",
          5444 => x"fe",
          5445 => x"fe",
          5446 => x"fe",
          5447 => x"81",
          5448 => x"80",
          5449 => x"38",
          5450 => x"52",
          5451 => x"05",
          5452 => x"86",
          5453 => x"d3",
          5454 => x"81",
          5455 => x"fe",
          5456 => x"fe",
          5457 => x"3d",
          5458 => x"53",
          5459 => x"51",
          5460 => x"3f",
          5461 => x"08",
          5462 => x"38",
          5463 => x"fd",
          5464 => x"3d",
          5465 => x"53",
          5466 => x"51",
          5467 => x"3f",
          5468 => x"08",
          5469 => x"d3",
          5470 => x"60",
          5471 => x"f8",
          5472 => x"70",
          5473 => x"fb",
          5474 => x"bf",
          5475 => x"78",
          5476 => x"b4",
          5477 => x"dc",
          5478 => x"b2",
          5479 => x"d3",
          5480 => x"2e",
          5481 => x"d3",
          5482 => x"f4",
          5483 => x"ab",
          5484 => x"c8",
          5485 => x"d5",
          5486 => x"fd",
          5487 => x"3d",
          5488 => x"51",
          5489 => x"3f",
          5490 => x"08",
          5491 => x"f8",
          5492 => x"fe",
          5493 => x"81",
          5494 => x"ac",
          5495 => x"51",
          5496 => x"81",
          5497 => x"80",
          5498 => x"38",
          5499 => x"08",
          5500 => x"3f",
          5501 => x"b4",
          5502 => x"05",
          5503 => x"eb",
          5504 => x"ac",
          5505 => x"fe",
          5506 => x"5b",
          5507 => x"3f",
          5508 => x"08",
          5509 => x"f8",
          5510 => x"fe",
          5511 => x"81",
          5512 => x"b5",
          5513 => x"05",
          5514 => x"e4",
          5515 => x"cb",
          5516 => x"d3",
          5517 => x"56",
          5518 => x"d3",
          5519 => x"ff",
          5520 => x"53",
          5521 => x"51",
          5522 => x"81",
          5523 => x"80",
          5524 => x"38",
          5525 => x"08",
          5526 => x"3f",
          5527 => x"81",
          5528 => x"fe",
          5529 => x"82",
          5530 => x"8f",
          5531 => x"39",
          5532 => x"51",
          5533 => x"3f",
          5534 => x"f1",
          5535 => x"db",
          5536 => x"81",
          5537 => x"94",
          5538 => x"80",
          5539 => x"c0",
          5540 => x"81",
          5541 => x"fe",
          5542 => x"fb",
          5543 => x"c9",
          5544 => x"f2",
          5545 => x"80",
          5546 => x"c0",
          5547 => x"8c",
          5548 => x"87",
          5549 => x"0c",
          5550 => x"b4",
          5551 => x"11",
          5552 => x"05",
          5553 => x"ca",
          5554 => x"ac",
          5555 => x"fb",
          5556 => x"52",
          5557 => x"51",
          5558 => x"3f",
          5559 => x"04",
          5560 => x"f4",
          5561 => x"f8",
          5562 => x"fa",
          5563 => x"d3",
          5564 => x"2e",
          5565 => x"60",
          5566 => x"f0",
          5567 => x"87",
          5568 => x"78",
          5569 => x"ac",
          5570 => x"d3",
          5571 => x"2e",
          5572 => x"81",
          5573 => x"52",
          5574 => x"51",
          5575 => x"3f",
          5576 => x"81",
          5577 => x"fe",
          5578 => x"fe",
          5579 => x"fa",
          5580 => x"ca",
          5581 => x"f1",
          5582 => x"59",
          5583 => x"fe",
          5584 => x"fa",
          5585 => x"70",
          5586 => x"78",
          5587 => x"8b",
          5588 => x"06",
          5589 => x"2e",
          5590 => x"b4",
          5591 => x"05",
          5592 => x"87",
          5593 => x"d8",
          5594 => x"ac",
          5595 => x"ca",
          5596 => x"53",
          5597 => x"52",
          5598 => x"52",
          5599 => x"9d",
          5600 => x"a8",
          5601 => x"e0",
          5602 => x"61",
          5603 => x"61",
          5604 => x"83",
          5605 => x"83",
          5606 => x"78",
          5607 => x"3f",
          5608 => x"08",
          5609 => x"32",
          5610 => x"07",
          5611 => x"38",
          5612 => x"09",
          5613 => x"a3",
          5614 => x"f0",
          5615 => x"c7",
          5616 => x"39",
          5617 => x"80",
          5618 => x"e0",
          5619 => x"86",
          5620 => x"c0",
          5621 => x"9b",
          5622 => x"0b",
          5623 => x"9c",
          5624 => x"83",
          5625 => x"94",
          5626 => x"80",
          5627 => x"c0",
          5628 => x"93",
          5629 => x"d3",
          5630 => x"e7",
          5631 => x"c0",
          5632 => x"89",
          5633 => x"cf",
          5634 => x"80",
          5635 => x"cb",
          5636 => x"8c",
          5637 => x"f5",
          5638 => x"c9",
          5639 => x"b2",
          5640 => x"f3",
          5641 => x"da",
          5642 => x"00",
          5643 => x"00",
          5644 => x"00",
          5645 => x"00",
          5646 => x"00",
          5647 => x"00",
          5648 => x"00",
          5649 => x"00",
          5650 => x"00",
          5651 => x"00",
          5652 => x"00",
          5653 => x"00",
          5654 => x"00",
          5655 => x"00",
          5656 => x"00",
          5657 => x"00",
          5658 => x"00",
          5659 => x"00",
          5660 => x"00",
          5661 => x"00",
          5662 => x"00",
          5663 => x"00",
          5664 => x"00",
          5665 => x"00",
          5666 => x"00",
          5667 => x"00",
          5668 => x"00",
          5669 => x"00",
          5670 => x"00",
          5671 => x"00",
          5672 => x"00",
          5673 => x"00",
          5674 => x"00",
          5675 => x"00",
          5676 => x"00",
          5677 => x"00",
          5678 => x"00",
          5679 => x"00",
          5680 => x"00",
          5681 => x"00",
          5682 => x"00",
          5683 => x"00",
          5684 => x"00",
          5685 => x"00",
          5686 => x"00",
          5687 => x"00",
          5688 => x"00",
          5689 => x"00",
          5690 => x"00",
          5691 => x"00",
          5692 => x"00",
          5693 => x"00",
          5694 => x"00",
          5695 => x"00",
          5696 => x"00",
          5697 => x"00",
          5698 => x"00",
          5699 => x"00",
          5700 => x"00",
          5701 => x"00",
          5702 => x"00",
          5703 => x"00",
          5704 => x"00",
          5705 => x"00",
          5706 => x"00",
          5707 => x"00",
          5708 => x"00",
          5709 => x"00",
          5710 => x"00",
          5711 => x"00",
          5712 => x"00",
          5713 => x"00",
          5714 => x"00",
          5715 => x"00",
          5716 => x"00",
          5717 => x"00",
          5718 => x"00",
          5719 => x"00",
          5720 => x"00",
          5721 => x"00",
          5722 => x"00",
          5723 => x"00",
          5724 => x"00",
          5725 => x"00",
          5726 => x"00",
          5727 => x"00",
          5728 => x"00",
          5729 => x"00",
          5730 => x"00",
          5731 => x"00",
          5732 => x"00",
          5733 => x"00",
          5734 => x"00",
          5735 => x"00",
          5736 => x"00",
          5737 => x"00",
          5738 => x"00",
          5739 => x"00",
          5740 => x"00",
          5741 => x"00",
          5742 => x"00",
          5743 => x"00",
          5744 => x"00",
          5745 => x"00",
          5746 => x"00",
          5747 => x"00",
          5748 => x"00",
          5749 => x"00",
          5750 => x"00",
          5751 => x"00",
          5752 => x"00",
          5753 => x"00",
          5754 => x"00",
          5755 => x"00",
          5756 => x"00",
          5757 => x"00",
          5758 => x"00",
          5759 => x"00",
          5760 => x"00",
          5761 => x"00",
          5762 => x"00",
          5763 => x"00",
          5764 => x"00",
          5765 => x"00",
          5766 => x"00",
          5767 => x"00",
          5768 => x"00",
          5769 => x"00",
          5770 => x"00",
          5771 => x"00",
          5772 => x"00",
          5773 => x"00",
          5774 => x"00",
          5775 => x"00",
          5776 => x"00",
          5777 => x"00",
          5778 => x"00",
          5779 => x"00",
          5780 => x"00",
          5781 => x"00",
          5782 => x"00",
          5783 => x"00",
          5784 => x"00",
          5785 => x"00",
          5786 => x"00",
          5787 => x"00",
          5788 => x"00",
          5789 => x"00",
          5790 => x"00",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"00",
          5815 => x"00",
          5816 => x"00",
          5817 => x"00",
          5818 => x"00",
          5819 => x"00",
          5820 => x"00",
          5821 => x"00",
          5822 => x"00",
          5823 => x"00",
          5824 => x"00",
          5825 => x"00",
          5826 => x"00",
          5827 => x"25",
          5828 => x"64",
          5829 => x"20",
          5830 => x"25",
          5831 => x"64",
          5832 => x"25",
          5833 => x"53",
          5834 => x"43",
          5835 => x"69",
          5836 => x"61",
          5837 => x"6e",
          5838 => x"20",
          5839 => x"6f",
          5840 => x"6f",
          5841 => x"6f",
          5842 => x"67",
          5843 => x"3a",
          5844 => x"76",
          5845 => x"73",
          5846 => x"70",
          5847 => x"65",
          5848 => x"64",
          5849 => x"20",
          5850 => x"49",
          5851 => x"20",
          5852 => x"4d",
          5853 => x"74",
          5854 => x"3d",
          5855 => x"58",
          5856 => x"69",
          5857 => x"25",
          5858 => x"29",
          5859 => x"20",
          5860 => x"42",
          5861 => x"20",
          5862 => x"61",
          5863 => x"25",
          5864 => x"2c",
          5865 => x"7a",
          5866 => x"30",
          5867 => x"2e",
          5868 => x"20",
          5869 => x"52",
          5870 => x"28",
          5871 => x"72",
          5872 => x"30",
          5873 => x"20",
          5874 => x"65",
          5875 => x"38",
          5876 => x"0a",
          5877 => x"20",
          5878 => x"49",
          5879 => x"4c",
          5880 => x"20",
          5881 => x"50",
          5882 => x"00",
          5883 => x"20",
          5884 => x"53",
          5885 => x"00",
          5886 => x"20",
          5887 => x"53",
          5888 => x"61",
          5889 => x"28",
          5890 => x"69",
          5891 => x"3d",
          5892 => x"58",
          5893 => x"00",
          5894 => x"20",
          5895 => x"49",
          5896 => x"52",
          5897 => x"54",
          5898 => x"4e",
          5899 => x"4c",
          5900 => x"0a",
          5901 => x"20",
          5902 => x"54",
          5903 => x"52",
          5904 => x"54",
          5905 => x"72",
          5906 => x"30",
          5907 => x"2e",
          5908 => x"41",
          5909 => x"65",
          5910 => x"73",
          5911 => x"20",
          5912 => x"43",
          5913 => x"52",
          5914 => x"74",
          5915 => x"63",
          5916 => x"20",
          5917 => x"72",
          5918 => x"20",
          5919 => x"30",
          5920 => x"00",
          5921 => x"20",
          5922 => x"43",
          5923 => x"4d",
          5924 => x"72",
          5925 => x"74",
          5926 => x"20",
          5927 => x"72",
          5928 => x"20",
          5929 => x"30",
          5930 => x"00",
          5931 => x"20",
          5932 => x"53",
          5933 => x"6b",
          5934 => x"61",
          5935 => x"41",
          5936 => x"65",
          5937 => x"20",
          5938 => x"20",
          5939 => x"30",
          5940 => x"00",
          5941 => x"20",
          5942 => x"5a",
          5943 => x"49",
          5944 => x"20",
          5945 => x"20",
          5946 => x"20",
          5947 => x"20",
          5948 => x"20",
          5949 => x"30",
          5950 => x"00",
          5951 => x"20",
          5952 => x"53",
          5953 => x"65",
          5954 => x"6c",
          5955 => x"20",
          5956 => x"71",
          5957 => x"20",
          5958 => x"20",
          5959 => x"30",
          5960 => x"00",
          5961 => x"53",
          5962 => x"6c",
          5963 => x"4d",
          5964 => x"75",
          5965 => x"46",
          5966 => x"00",
          5967 => x"45",
          5968 => x"45",
          5969 => x"69",
          5970 => x"55",
          5971 => x"6f",
          5972 => x"53",
          5973 => x"22",
          5974 => x"3a",
          5975 => x"3e",
          5976 => x"7c",
          5977 => x"46",
          5978 => x"46",
          5979 => x"32",
          5980 => x"30",
          5981 => x"31",
          5982 => x"32",
          5983 => x"33",
          5984 => x"35",
          5985 => x"36",
          5986 => x"37",
          5987 => x"38",
          5988 => x"39",
          5989 => x"31",
          5990 => x"eb",
          5991 => x"53",
          5992 => x"35",
          5993 => x"4e",
          5994 => x"41",
          5995 => x"20",
          5996 => x"41",
          5997 => x"20",
          5998 => x"4e",
          5999 => x"41",
          6000 => x"20",
          6001 => x"41",
          6002 => x"20",
          6003 => x"00",
          6004 => x"00",
          6005 => x"00",
          6006 => x"00",
          6007 => x"80",
          6008 => x"8e",
          6009 => x"45",
          6010 => x"49",
          6011 => x"90",
          6012 => x"99",
          6013 => x"59",
          6014 => x"9c",
          6015 => x"41",
          6016 => x"a5",
          6017 => x"a8",
          6018 => x"ac",
          6019 => x"b0",
          6020 => x"b4",
          6021 => x"b8",
          6022 => x"bc",
          6023 => x"c0",
          6024 => x"c4",
          6025 => x"c8",
          6026 => x"cc",
          6027 => x"d0",
          6028 => x"d4",
          6029 => x"d8",
          6030 => x"dc",
          6031 => x"e0",
          6032 => x"e4",
          6033 => x"e8",
          6034 => x"ec",
          6035 => x"f0",
          6036 => x"f4",
          6037 => x"f8",
          6038 => x"fc",
          6039 => x"2b",
          6040 => x"3d",
          6041 => x"5c",
          6042 => x"3c",
          6043 => x"7f",
          6044 => x"00",
          6045 => x"00",
          6046 => x"01",
          6047 => x"00",
          6048 => x"00",
          6049 => x"00",
          6050 => x"00",
          6051 => x"00",
          6052 => x"46",
          6053 => x"32",
          6054 => x"46",
          6055 => x"36",
          6056 => x"65",
          6057 => x"54",
          6058 => x"44",
          6059 => x"20",
          6060 => x"43",
          6061 => x"52",
          6062 => x"00",
          6063 => x"44",
          6064 => x"20",
          6065 => x"46",
          6066 => x"43",
          6067 => x"52",
          6068 => x"00",
          6069 => x"46",
          6070 => x"53",
          6071 => x"45",
          6072 => x"4f",
          6073 => x"4f",
          6074 => x"4d",
          6075 => x"52",
          6076 => x"48",
          6077 => x"57",
          6078 => x"00",
          6079 => x"54",
          6080 => x"49",
          6081 => x"45",
          6082 => x"55",
          6083 => x"4e",
          6084 => x"4d",
          6085 => x"20",
          6086 => x"4d",
          6087 => x"53",
          6088 => x"64",
          6089 => x"70",
          6090 => x"64",
          6091 => x"74",
          6092 => x"64",
          6093 => x"74",
          6094 => x"64",
          6095 => x"74",
          6096 => x"62",
          6097 => x"70",
          6098 => x"62",
          6099 => x"74",
          6100 => x"62",
          6101 => x"64",
          6102 => x"62",
          6103 => x"74",
          6104 => x"62",
          6105 => x"6c",
          6106 => x"62",
          6107 => x"00",
          6108 => x"66",
          6109 => x"74",
          6110 => x"66",
          6111 => x"6e",
          6112 => x"66",
          6113 => x"73",
          6114 => x"66",
          6115 => x"6b",
          6116 => x"66",
          6117 => x"64",
          6118 => x"66",
          6119 => x"70",
          6120 => x"00",
          6121 => x"66",
          6122 => x"74",
          6123 => x"66",
          6124 => x"6e",
          6125 => x"66",
          6126 => x"6f",
          6127 => x"66",
          6128 => x"72",
          6129 => x"66",
          6130 => x"65",
          6131 => x"66",
          6132 => x"61",
          6133 => x"66",
          6134 => x"00",
          6135 => x"66",
          6136 => x"69",
          6137 => x"66",
          6138 => x"74",
          6139 => x"66",
          6140 => x"00",
          6141 => x"66",
          6142 => x"00",
          6143 => x"66",
          6144 => x"66",
          6145 => x"63",
          6146 => x"66",
          6147 => x"61",
          6148 => x"66",
          6149 => x"64",
          6150 => x"66",
          6151 => x"63",
          6152 => x"66",
          6153 => x"65",
          6154 => x"66",
          6155 => x"70",
          6156 => x"66",
          6157 => x"66",
          6158 => x"76",
          6159 => x"66",
          6160 => x"77",
          6161 => x"00",
          6162 => x"66",
          6163 => x"65",
          6164 => x"66",
          6165 => x"73",
          6166 => x"6d",
          6167 => x"00",
          6168 => x"6d",
          6169 => x"70",
          6170 => x"6d",
          6171 => x"6d",
          6172 => x"6d",
          6173 => x"68",
          6174 => x"68",
          6175 => x"68",
          6176 => x"68",
          6177 => x"68",
          6178 => x"68",
          6179 => x"64",
          6180 => x"00",
          6181 => x"63",
          6182 => x"6d",
          6183 => x"00",
          6184 => x"63",
          6185 => x"00",
          6186 => x"6a",
          6187 => x"72",
          6188 => x"61",
          6189 => x"72",
          6190 => x"74",
          6191 => x"68",
          6192 => x"00",
          6193 => x"69",
          6194 => x"00",
          6195 => x"74",
          6196 => x"00",
          6197 => x"74",
          6198 => x"00",
          6199 => x"44",
          6200 => x"20",
          6201 => x"6f",
          6202 => x"49",
          6203 => x"72",
          6204 => x"20",
          6205 => x"6f",
          6206 => x"00",
          6207 => x"44",
          6208 => x"20",
          6209 => x"20",
          6210 => x"64",
          6211 => x"00",
          6212 => x"4e",
          6213 => x"69",
          6214 => x"66",
          6215 => x"64",
          6216 => x"4e",
          6217 => x"61",
          6218 => x"66",
          6219 => x"64",
          6220 => x"49",
          6221 => x"6c",
          6222 => x"66",
          6223 => x"6e",
          6224 => x"2e",
          6225 => x"41",
          6226 => x"73",
          6227 => x"65",
          6228 => x"64",
          6229 => x"46",
          6230 => x"20",
          6231 => x"65",
          6232 => x"20",
          6233 => x"73",
          6234 => x"0a",
          6235 => x"46",
          6236 => x"20",
          6237 => x"64",
          6238 => x"69",
          6239 => x"6c",
          6240 => x"0a",
          6241 => x"53",
          6242 => x"73",
          6243 => x"69",
          6244 => x"70",
          6245 => x"65",
          6246 => x"64",
          6247 => x"44",
          6248 => x"65",
          6249 => x"6d",
          6250 => x"20",
          6251 => x"69",
          6252 => x"6c",
          6253 => x"0a",
          6254 => x"44",
          6255 => x"20",
          6256 => x"20",
          6257 => x"62",
          6258 => x"2e",
          6259 => x"4e",
          6260 => x"6f",
          6261 => x"74",
          6262 => x"65",
          6263 => x"6c",
          6264 => x"73",
          6265 => x"20",
          6266 => x"6e",
          6267 => x"6e",
          6268 => x"73",
          6269 => x"00",
          6270 => x"46",
          6271 => x"61",
          6272 => x"62",
          6273 => x"65",
          6274 => x"00",
          6275 => x"54",
          6276 => x"6f",
          6277 => x"20",
          6278 => x"72",
          6279 => x"6f",
          6280 => x"61",
          6281 => x"6c",
          6282 => x"2e",
          6283 => x"46",
          6284 => x"20",
          6285 => x"6c",
          6286 => x"65",
          6287 => x"00",
          6288 => x"49",
          6289 => x"66",
          6290 => x"69",
          6291 => x"20",
          6292 => x"6f",
          6293 => x"0a",
          6294 => x"54",
          6295 => x"6d",
          6296 => x"20",
          6297 => x"6e",
          6298 => x"6c",
          6299 => x"0a",
          6300 => x"50",
          6301 => x"6d",
          6302 => x"72",
          6303 => x"6e",
          6304 => x"72",
          6305 => x"2e",
          6306 => x"53",
          6307 => x"65",
          6308 => x"0a",
          6309 => x"55",
          6310 => x"6f",
          6311 => x"65",
          6312 => x"72",
          6313 => x"0a",
          6314 => x"20",
          6315 => x"65",
          6316 => x"73",
          6317 => x"20",
          6318 => x"20",
          6319 => x"65",
          6320 => x"65",
          6321 => x"00",
          6322 => x"72",
          6323 => x"00",
          6324 => x"5a",
          6325 => x"41",
          6326 => x"0a",
          6327 => x"25",
          6328 => x"00",
          6329 => x"31",
          6330 => x"37",
          6331 => x"31",
          6332 => x"76",
          6333 => x"00",
          6334 => x"20",
          6335 => x"2c",
          6336 => x"76",
          6337 => x"32",
          6338 => x"25",
          6339 => x"73",
          6340 => x"0a",
          6341 => x"5a",
          6342 => x"41",
          6343 => x"74",
          6344 => x"75",
          6345 => x"48",
          6346 => x"6c",
          6347 => x"00",
          6348 => x"54",
          6349 => x"72",
          6350 => x"74",
          6351 => x"75",
          6352 => x"00",
          6353 => x"50",
          6354 => x"69",
          6355 => x"72",
          6356 => x"74",
          6357 => x"49",
          6358 => x"4c",
          6359 => x"20",
          6360 => x"65",
          6361 => x"70",
          6362 => x"49",
          6363 => x"4c",
          6364 => x"20",
          6365 => x"65",
          6366 => x"70",
          6367 => x"55",
          6368 => x"30",
          6369 => x"20",
          6370 => x"65",
          6371 => x"70",
          6372 => x"55",
          6373 => x"30",
          6374 => x"20",
          6375 => x"65",
          6376 => x"70",
          6377 => x"55",
          6378 => x"31",
          6379 => x"20",
          6380 => x"65",
          6381 => x"70",
          6382 => x"55",
          6383 => x"31",
          6384 => x"20",
          6385 => x"65",
          6386 => x"70",
          6387 => x"53",
          6388 => x"69",
          6389 => x"75",
          6390 => x"69",
          6391 => x"2e",
          6392 => x"00",
          6393 => x"45",
          6394 => x"6c",
          6395 => x"20",
          6396 => x"65",
          6397 => x"2e",
          6398 => x"30",
          6399 => x"46",
          6400 => x"65",
          6401 => x"6f",
          6402 => x"69",
          6403 => x"6c",
          6404 => x"20",
          6405 => x"63",
          6406 => x"20",
          6407 => x"70",
          6408 => x"73",
          6409 => x"6e",
          6410 => x"6d",
          6411 => x"61",
          6412 => x"2e",
          6413 => x"2a",
          6414 => x"42",
          6415 => x"64",
          6416 => x"20",
          6417 => x"0a",
          6418 => x"49",
          6419 => x"69",
          6420 => x"73",
          6421 => x"0a",
          6422 => x"46",
          6423 => x"65",
          6424 => x"6f",
          6425 => x"69",
          6426 => x"6c",
          6427 => x"2e",
          6428 => x"72",
          6429 => x"64",
          6430 => x"25",
          6431 => x"44",
          6432 => x"62",
          6433 => x"67",
          6434 => x"74",
          6435 => x"75",
          6436 => x"0a",
          6437 => x"45",
          6438 => x"6c",
          6439 => x"20",
          6440 => x"65",
          6441 => x"70",
          6442 => x"00",
          6443 => x"44",
          6444 => x"62",
          6445 => x"20",
          6446 => x"74",
          6447 => x"66",
          6448 => x"45",
          6449 => x"6c",
          6450 => x"20",
          6451 => x"74",
          6452 => x"66",
          6453 => x"45",
          6454 => x"75",
          6455 => x"67",
          6456 => x"64",
          6457 => x"20",
          6458 => x"78",
          6459 => x"2e",
          6460 => x"43",
          6461 => x"69",
          6462 => x"63",
          6463 => x"20",
          6464 => x"30",
          6465 => x"2e",
          6466 => x"00",
          6467 => x"43",
          6468 => x"20",
          6469 => x"75",
          6470 => x"64",
          6471 => x"64",
          6472 => x"25",
          6473 => x"0a",
          6474 => x"52",
          6475 => x"61",
          6476 => x"6e",
          6477 => x"70",
          6478 => x"63",
          6479 => x"6f",
          6480 => x"2e",
          6481 => x"43",
          6482 => x"20",
          6483 => x"6f",
          6484 => x"6e",
          6485 => x"2e",
          6486 => x"5a",
          6487 => x"62",
          6488 => x"25",
          6489 => x"25",
          6490 => x"73",
          6491 => x"00",
          6492 => x"42",
          6493 => x"63",
          6494 => x"61",
          6495 => x"0a",
          6496 => x"52",
          6497 => x"69",
          6498 => x"2e",
          6499 => x"45",
          6500 => x"6c",
          6501 => x"20",
          6502 => x"65",
          6503 => x"70",
          6504 => x"2e",
          6505 => x"00",
          6506 => x"00",
          6507 => x"00",
          6508 => x"00",
          6509 => x"00",
          6510 => x"00",
          6511 => x"00",
          6512 => x"00",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"05",
          6517 => x"00",
          6518 => x"01",
          6519 => x"80",
          6520 => x"01",
          6521 => x"00",
          6522 => x"01",
          6523 => x"00",
          6524 => x"00",
          6525 => x"00",
          6526 => x"00",
          6527 => x"00",
          6528 => x"01",
          6529 => x"00",
          6530 => x"00",
          6531 => x"00",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"00",
          6536 => x"01",
          6537 => x"00",
          6538 => x"00",
          6539 => x"00",
          6540 => x"00",
          6541 => x"00",
          6542 => x"00",
          6543 => x"00",
          6544 => x"00",
          6545 => x"00",
          6546 => x"00",
          6547 => x"00",
          6548 => x"00",
          6549 => x"00",
          6550 => x"00",
          6551 => x"00",
          6552 => x"00",
          6553 => x"00",
          6554 => x"00",
          6555 => x"00",
          6556 => x"00",
          6557 => x"00",
          6558 => x"00",
          6559 => x"00",
          6560 => x"00",
          6561 => x"00",
          6562 => x"00",
          6563 => x"00",
          6564 => x"01",
          6565 => x"00",
          6566 => x"00",
          6567 => x"00",
          6568 => x"00",
          6569 => x"00",
          6570 => x"00",
          6571 => x"00",
          6572 => x"00",
          6573 => x"00",
          6574 => x"00",
          6575 => x"00",
          6576 => x"00",
          6577 => x"00",
          6578 => x"00",
          6579 => x"00",
          6580 => x"00",
          6581 => x"00",
          6582 => x"00",
          6583 => x"00",
          6584 => x"00",
          6585 => x"00",
          6586 => x"00",
          6587 => x"00",
          6588 => x"00",
          6589 => x"00",
          6590 => x"00",
          6591 => x"00",
          6592 => x"00",
          6593 => x"00",
          6594 => x"00",
          6595 => x"00",
          6596 => x"00",
          6597 => x"00",
          6598 => x"00",
          6599 => x"00",
          6600 => x"00",
          6601 => x"00",
          6602 => x"00",
          6603 => x"00",
          6604 => x"00",
          6605 => x"00",
          6606 => x"00",
          6607 => x"00",
          6608 => x"00",
          6609 => x"00",
          6610 => x"00",
          6611 => x"00",
          6612 => x"00",
          6613 => x"00",
          6614 => x"00",
          6615 => x"00",
          6616 => x"00",
          6617 => x"00",
          6618 => x"00",
          6619 => x"00",
          6620 => x"00",
          6621 => x"00",
          6622 => x"00",
          6623 => x"00",
          6624 => x"00",
          6625 => x"00",
          6626 => x"00",
          6627 => x"00",
          6628 => x"00",
          6629 => x"00",
          6630 => x"00",
          6631 => x"00",
          6632 => x"00",
          6633 => x"00",
          6634 => x"00",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"00",
          6639 => x"00",
          6640 => x"00",
          6641 => x"00",
          6642 => x"00",
          6643 => x"00",
          6644 => x"01",
          6645 => x"00",
          6646 => x"00",
          6647 => x"00",
          6648 => x"01",
          6649 => x"00",
          6650 => x"00",
          6651 => x"00",
          6652 => x"00",
          6653 => x"00",
          6654 => x"00",
          6655 => x"00",
          6656 => x"00",
          6657 => x"00",
          6658 => x"00",
          6659 => x"00",
          6660 => x"00",
          6661 => x"00",
          6662 => x"00",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"00",
          6667 => x"00",
          6668 => x"00",
          6669 => x"00",
          6670 => x"00",
          6671 => x"00",
          6672 => x"00",
          6673 => x"00",
          6674 => x"00",
          6675 => x"00",
          6676 => x"00",
          6677 => x"00",
          6678 => x"00",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"00",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"00",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"00",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"00",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"00",
          6699 => x"00",
          6700 => x"01",
          6701 => x"00",
          6702 => x"00",
          6703 => x"00",
          6704 => x"01",
          6705 => x"00",
          6706 => x"00",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"00",
          6711 => x"00",
          6712 => x"00",
          6713 => x"00",
          6714 => x"00",
          6715 => x"00",
          6716 => x"01",
          6717 => x"00",
          6718 => x"00",
          6719 => x"00",
          6720 => x"01",
          6721 => x"00",
          6722 => x"00",
          6723 => x"00",
          6724 => x"00",
          6725 => x"00",
          6726 => x"00",
          6727 => x"00",
          6728 => x"00",
          6729 => x"00",
          6730 => x"00",
          6731 => x"00",
          6732 => x"01",
          6733 => x"00",
          6734 => x"00",
          6735 => x"00",
          6736 => x"01",
          6737 => x"00",
          6738 => x"00",
          6739 => x"00",
          6740 => x"01",
          6741 => x"00",
          6742 => x"00",
          6743 => x"00",
          6744 => x"01",
          6745 => x"00",
          6746 => x"00",
          6747 => x"00",
          6748 => x"00",
          6749 => x"00",
          6750 => x"00",
          6751 => x"00",
          6752 => x"01",
          6753 => x"00",
          6754 => x"00",
          6755 => x"00",
          6756 => x"00",
          6757 => x"00",
          6758 => x"00",
          6759 => x"00",
          6760 => x"01",
          6761 => x"00",
          6762 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
