-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8b",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"a0",
           281 => x"38",
           282 => x"84",
           283 => x"0b",
           284 => x"e2",
           285 => x"51",
           286 => x"00",
           287 => x"88",
           288 => x"00",
           289 => x"02",
           290 => x"3d",
           291 => x"94",
           292 => x"08",
           293 => x"88",
           294 => x"82",
           295 => x"08",
           296 => x"54",
           297 => x"94",
           298 => x"08",
           299 => x"fd",
           300 => x"53",
           301 => x"05",
           302 => x"08",
           303 => x"51",
           304 => x"88",
           305 => x"0c",
           306 => x"0d",
           307 => x"94",
           308 => x"0c",
           309 => x"80",
           310 => x"fc",
           311 => x"08",
           312 => x"80",
           313 => x"94",
           314 => x"08",
           315 => x"88",
           316 => x"0b",
           317 => x"05",
           318 => x"fc",
           319 => x"38",
           320 => x"08",
           321 => x"94",
           322 => x"08",
           323 => x"05",
           324 => x"8c",
           325 => x"25",
           326 => x"08",
           327 => x"30",
           328 => x"05",
           329 => x"94",
           330 => x"0c",
           331 => x"05",
           332 => x"81",
           333 => x"f0",
           334 => x"08",
           335 => x"94",
           336 => x"0c",
           337 => x"08",
           338 => x"52",
           339 => x"05",
           340 => x"a7",
           341 => x"70",
           342 => x"05",
           343 => x"08",
           344 => x"80",
           345 => x"94",
           346 => x"08",
           347 => x"f8",
           348 => x"08",
           349 => x"70",
           350 => x"89",
           351 => x"0c",
           352 => x"02",
           353 => x"3d",
           354 => x"94",
           355 => x"0c",
           356 => x"05",
           357 => x"93",
           358 => x"88",
           359 => x"94",
           360 => x"0c",
           361 => x"08",
           362 => x"94",
           363 => x"08",
           364 => x"38",
           365 => x"05",
           366 => x"08",
           367 => x"81",
           368 => x"8c",
           369 => x"94",
           370 => x"08",
           371 => x"88",
           372 => x"08",
           373 => x"54",
           374 => x"05",
           375 => x"8c",
           376 => x"f8",
           377 => x"94",
           378 => x"0c",
           379 => x"05",
           380 => x"0c",
           381 => x"0d",
           382 => x"94",
           383 => x"0c",
           384 => x"81",
           385 => x"fc",
           386 => x"0b",
           387 => x"05",
           388 => x"8c",
           389 => x"08",
           390 => x"27",
           391 => x"08",
           392 => x"80",
           393 => x"80",
           394 => x"8c",
           395 => x"99",
           396 => x"8c",
           397 => x"94",
           398 => x"0c",
           399 => x"05",
           400 => x"08",
           401 => x"c9",
           402 => x"fc",
           403 => x"2e",
           404 => x"94",
           405 => x"08",
           406 => x"05",
           407 => x"38",
           408 => x"05",
           409 => x"8c",
           410 => x"94",
           411 => x"0c",
           412 => x"05",
           413 => x"fc",
           414 => x"94",
           415 => x"0c",
           416 => x"05",
           417 => x"94",
           418 => x"0c",
           419 => x"05",
           420 => x"94",
           421 => x"0c",
           422 => x"94",
           423 => x"08",
           424 => x"38",
           425 => x"05",
           426 => x"08",
           427 => x"51",
           428 => x"08",
           429 => x"70",
           430 => x"05",
           431 => x"08",
           432 => x"88",
           433 => x"0d",
           434 => x"ff",
           435 => x"88",
           436 => x"92",
           437 => x"0b",
           438 => x"8c",
           439 => x"87",
           440 => x"0c",
           441 => x"8c",
           442 => x"06",
           443 => x"80",
           444 => x"87",
           445 => x"08",
           446 => x"38",
           447 => x"8c",
           448 => x"80",
           449 => x"93",
           450 => x"98",
           451 => x"70",
           452 => x"38",
           453 => x"0b",
           454 => x"0b",
           455 => x"f0",
           456 => x"83",
           457 => x"fa",
           458 => x"7b",
           459 => x"56",
           460 => x"0b",
           461 => x"33",
           462 => x"55",
           463 => x"75",
           464 => x"06",
           465 => x"85",
           466 => x"98",
           467 => x"87",
           468 => x"0c",
           469 => x"c0",
           470 => x"87",
           471 => x"08",
           472 => x"70",
           473 => x"52",
           474 => x"2e",
           475 => x"c0",
           476 => x"70",
           477 => x"76",
           478 => x"53",
           479 => x"2e",
           480 => x"80",
           481 => x"71",
           482 => x"05",
           483 => x"14",
           484 => x"55",
           485 => x"51",
           486 => x"8b",
           487 => x"98",
           488 => x"70",
           489 => x"87",
           490 => x"08",
           491 => x"38",
           492 => x"c0",
           493 => x"87",
           494 => x"08",
           495 => x"51",
           496 => x"38",
           497 => x"80",
           498 => x"52",
           499 => x"09",
           500 => x"38",
           501 => x"8c",
           502 => x"72",
           503 => x"06",
           504 => x"52",
           505 => x"88",
           506 => x"fe",
           507 => x"81",
           508 => x"33",
           509 => x"07",
           510 => x"51",
           511 => x"04",
           512 => x"75",
           513 => x"82",
           514 => x"90",
           515 => x"2b",
           516 => x"33",
           517 => x"88",
           518 => x"71",
           519 => x"52",
           520 => x"54",
           521 => x"0d",
           522 => x"0d",
           523 => x"0b",
           524 => x"57",
           525 => x"27",
           526 => x"76",
           527 => x"27",
           528 => x"75",
           529 => x"82",
           530 => x"74",
           531 => x"38",
           532 => x"74",
           533 => x"83",
           534 => x"76",
           535 => x"17",
           536 => x"88",
           537 => x"55",
           538 => x"88",
           539 => x"74",
           540 => x"3f",
           541 => x"ff",
           542 => x"ad",
           543 => x"76",
           544 => x"fc",
           545 => x"87",
           546 => x"08",
           547 => x"3d",
           548 => x"fd",
           549 => x"08",
           550 => x"51",
           551 => x"88",
           552 => x"06",
           553 => x"81",
           554 => x"0c",
           555 => x"04",
           556 => x"0b",
           557 => x"f4",
           558 => x"88",
           559 => x"05",
           560 => x"80",
           561 => x"27",
           562 => x"14",
           563 => x"29",
           564 => x"05",
           565 => x"88",
           566 => x"0d",
           567 => x"0d",
           568 => x"0b",
           569 => x"9f",
           570 => x"33",
           571 => x"71",
           572 => x"81",
           573 => x"94",
           574 => x"ef",
           575 => x"90",
           576 => x"14",
           577 => x"3f",
           578 => x"ff",
           579 => x"07",
           580 => x"3d",
           581 => x"3d",
           582 => x"0b",
           583 => x"08",
           584 => x"75",
           585 => x"08",
           586 => x"2e",
           587 => x"14",
           588 => x"85",
           589 => x"b0",
           590 => x"38",
           591 => x"71",
           592 => x"81",
           593 => x"90",
           594 => x"72",
           595 => x"72",
           596 => x"38",
           597 => x"d8",
           598 => x"52",
           599 => x"14",
           600 => x"90",
           601 => x"52",
           602 => x"86",
           603 => x"fa",
           604 => x"0b",
           605 => x"f4",
           606 => x"81",
           607 => x"ff",
           608 => x"54",
           609 => x"80",
           610 => x"90",
           611 => x"72",
           612 => x"52",
           613 => x"73",
           614 => x"71",
           615 => x"81",
           616 => x"0c",
           617 => x"53",
           618 => x"83",
           619 => x"22",
           620 => x"76",
           621 => x"b5",
           622 => x"33",
           623 => x"84",
           624 => x"71",
           625 => x"51",
           626 => x"81",
           627 => x"08",
           628 => x"83",
           629 => x"88",
           630 => x"96",
           631 => x"8c",
           632 => x"08",
           633 => x"3f",
           634 => x"16",
           635 => x"23",
           636 => x"88",
           637 => x"0d",
           638 => x"0d",
           639 => x"58",
           640 => x"33",
           641 => x"2e",
           642 => x"88",
           643 => x"70",
           644 => x"39",
           645 => x"56",
           646 => x"2e",
           647 => x"84",
           648 => x"43",
           649 => x"1d",
           650 => x"33",
           651 => x"9f",
           652 => x"7b",
           653 => x"3f",
           654 => x"80",
           655 => x"d3",
           656 => x"84",
           657 => x"58",
           658 => x"55",
           659 => x"81",
           660 => x"ff",
           661 => x"ff",
           662 => x"06",
           663 => x"70",
           664 => x"7f",
           665 => x"7a",
           666 => x"81",
           667 => x"13",
           668 => x"af",
           669 => x"a0",
           670 => x"80",
           671 => x"51",
           672 => x"5d",
           673 => x"80",
           674 => x"ae",
           675 => x"06",
           676 => x"55",
           677 => x"75",
           678 => x"80",
           679 => x"79",
           680 => x"30",
           681 => x"70",
           682 => x"07",
           683 => x"51",
           684 => x"75",
           685 => x"58",
           686 => x"ab",
           687 => x"19",
           688 => x"06",
           689 => x"5a",
           690 => x"75",
           691 => x"39",
           692 => x"0c",
           693 => x"a0",
           694 => x"81",
           695 => x"1a",
           696 => x"fc",
           697 => x"08",
           698 => x"a0",
           699 => x"70",
           700 => x"e0",
           701 => x"90",
           702 => x"7c",
           703 => x"3f",
           704 => x"88",
           705 => x"38",
           706 => x"74",
           707 => x"ee",
           708 => x"33",
           709 => x"70",
           710 => x"56",
           711 => x"38",
           712 => x"1e",
           713 => x"59",
           714 => x"ff",
           715 => x"ff",
           716 => x"79",
           717 => x"5b",
           718 => x"81",
           719 => x"71",
           720 => x"56",
           721 => x"2e",
           722 => x"39",
           723 => x"92",
           724 => x"fc",
           725 => x"8e",
           726 => x"56",
           727 => x"38",
           728 => x"56",
           729 => x"8b",
           730 => x"55",
           731 => x"8b",
           732 => x"84",
           733 => x"06",
           734 => x"74",
           735 => x"56",
           736 => x"56",
           737 => x"51",
           738 => x"88",
           739 => x"0c",
           740 => x"75",
           741 => x"3d",
           742 => x"3d",
           743 => x"59",
           744 => x"83",
           745 => x"52",
           746 => x"fb",
           747 => x"88",
           748 => x"38",
           749 => x"b3",
           750 => x"83",
           751 => x"55",
           752 => x"82",
           753 => x"09",
           754 => x"ce",
           755 => x"b6",
           756 => x"76",
           757 => x"3f",
           758 => x"88",
           759 => x"76",
           760 => x"3f",
           761 => x"ff",
           762 => x"74",
           763 => x"2e",
           764 => x"54",
           765 => x"77",
           766 => x"f6",
           767 => x"08",
           768 => x"94",
           769 => x"f7",
           770 => x"08",
           771 => x"06",
           772 => x"82",
           773 => x"38",
           774 => x"88",
           775 => x"0d",
           776 => x"0d",
           777 => x"0b",
           778 => x"9f",
           779 => x"9b",
           780 => x"81",
           781 => x"56",
           782 => x"38",
           783 => x"8d",
           784 => x"57",
           785 => x"3f",
           786 => x"ff",
           787 => x"81",
           788 => x"06",
           789 => x"54",
           790 => x"74",
           791 => x"f5",
           792 => x"08",
           793 => x"3d",
           794 => x"80",
           795 => x"95",
           796 => x"51",
           797 => x"88",
           798 => x"53",
           799 => x"fe",
           800 => x"08",
           801 => x"57",
           802 => x"09",
           803 => x"38",
           804 => x"99",
           805 => x"2e",
           806 => x"56",
           807 => x"a4",
           808 => x"79",
           809 => x"f4",
           810 => x"56",
           811 => x"fd",
           812 => x"e5",
           813 => x"b3",
           814 => x"83",
           815 => x"58",
           816 => x"95",
           817 => x"51",
           818 => x"88",
           819 => x"af",
           820 => x"71",
           821 => x"05",
           822 => x"54",
           823 => x"f6",
           824 => x"08",
           825 => x"06",
           826 => x"1a",
           827 => x"33",
           828 => x"95",
           829 => x"51",
           830 => x"88",
           831 => x"23",
           832 => x"05",
           833 => x"3f",
           834 => x"ff",
           835 => x"75",
           836 => x"3d",
           837 => x"f5",
           838 => x"08",
           839 => x"f5",
           840 => x"08",
           841 => x"06",
           842 => x"79",
           843 => x"22",
           844 => x"82",
           845 => x"72",
           846 => x"59",
           847 => x"ee",
           848 => x"08",
           849 => x"88",
           850 => x"08",
           851 => x"56",
           852 => x"df",
           853 => x"38",
           854 => x"ff",
           855 => x"85",
           856 => x"89",
           857 => x"76",
           858 => x"c1",
           859 => x"34",
           860 => x"09",
           861 => x"38",
           862 => x"05",
           863 => x"3f",
           864 => x"1a",
           865 => x"8c",
           866 => x"90",
           867 => x"83",
           868 => x"8c",
           869 => x"71",
           870 => x"94",
           871 => x"80",
           872 => x"34",
           873 => x"0b",
           874 => x"80",
           875 => x"0c",
           876 => x"04",
           877 => x"0b",
           878 => x"f4",
           879 => x"54",
           880 => x"80",
           881 => x"0b",
           882 => x"98",
           883 => x"45",
           884 => x"3d",
           885 => x"ec",
           886 => x"9d",
           887 => x"54",
           888 => x"c0",
           889 => x"33",
           890 => x"2e",
           891 => x"a7",
           892 => x"84",
           893 => x"06",
           894 => x"73",
           895 => x"38",
           896 => x"39",
           897 => x"d5",
           898 => x"a0",
           899 => x"3d",
           900 => x"f3",
           901 => x"08",
           902 => x"73",
           903 => x"81",
           904 => x"34",
           905 => x"98",
           906 => x"f6",
           907 => x"7f",
           908 => x"0b",
           909 => x"59",
           910 => x"80",
           911 => x"57",
           912 => x"81",
           913 => x"16",
           914 => x"55",
           915 => x"80",
           916 => x"38",
           917 => x"81",
           918 => x"39",
           919 => x"17",
           920 => x"81",
           921 => x"16",
           922 => x"08",
           923 => x"78",
           924 => x"74",
           925 => x"2e",
           926 => x"98",
           927 => x"83",
           928 => x"57",
           929 => x"38",
           930 => x"ff",
           931 => x"2a",
           932 => x"ff",
           933 => x"79",
           934 => x"87",
           935 => x"08",
           936 => x"a4",
           937 => x"f3",
           938 => x"08",
           939 => x"27",
           940 => x"74",
           941 => x"a4",
           942 => x"f3",
           943 => x"08",
           944 => x"80",
           945 => x"38",
           946 => x"a8",
           947 => x"16",
           948 => x"06",
           949 => x"31",
           950 => x"75",
           951 => x"77",
           952 => x"98",
           953 => x"ff",
           954 => x"16",
           955 => x"51",
           956 => x"88",
           957 => x"38",
           958 => x"15",
           959 => x"77",
           960 => x"08",
           961 => x"58",
           962 => x"fe",
           963 => x"19",
           964 => x"39",
           965 => x"88",
           966 => x"0d",
           967 => x"0d",
           968 => x"8c",
           969 => x"84",
           970 => x"51",
           971 => x"88",
           972 => x"87",
           973 => x"08",
           974 => x"84",
           975 => x"51",
           976 => x"73",
           977 => x"87",
           978 => x"0c",
           979 => x"9c",
           980 => x"84",
           981 => x"51",
           982 => x"88",
           983 => x"87",
           984 => x"08",
           985 => x"84",
           986 => x"51",
           987 => x"73",
           988 => x"87",
           989 => x"0c",
           990 => x"0b",
           991 => x"84",
           992 => x"83",
           993 => x"94",
           994 => x"f8",
           995 => x"3f",
           996 => x"38",
           997 => x"fc",
           998 => x"08",
           999 => x"80",
          1000 => x"87",
          1001 => x"0c",
          1002 => x"fc",
          1003 => x"80",
          1004 => x"fc",
          1005 => x"08",
          1006 => x"54",
          1007 => x"86",
          1008 => x"55",
          1009 => x"80",
          1010 => x"80",
          1011 => x"00",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"00",
          1016 => x"54",
          1017 => x"59",
          1018 => x"4d",
          1019 => x"00",
          1020 => x"00",
          2048 => x"a4",
          2049 => x"0b",
          2050 => x"04",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"a4",
          2057 => x"0b",
          2058 => x"04",
          2059 => x"a4",
          2060 => x"0b",
          2061 => x"04",
          2062 => x"a4",
          2063 => x"0b",
          2064 => x"04",
          2065 => x"a4",
          2066 => x"0b",
          2067 => x"04",
          2068 => x"a4",
          2069 => x"0b",
          2070 => x"04",
          2071 => x"a5",
          2072 => x"0b",
          2073 => x"04",
          2074 => x"a5",
          2075 => x"0b",
          2076 => x"04",
          2077 => x"a5",
          2078 => x"0b",
          2079 => x"04",
          2080 => x"a5",
          2081 => x"0b",
          2082 => x"04",
          2083 => x"a6",
          2084 => x"0b",
          2085 => x"04",
          2086 => x"a6",
          2087 => x"0b",
          2088 => x"04",
          2089 => x"a6",
          2090 => x"0b",
          2091 => x"04",
          2092 => x"a6",
          2093 => x"0b",
          2094 => x"04",
          2095 => x"a7",
          2096 => x"0b",
          2097 => x"04",
          2098 => x"a7",
          2099 => x"0b",
          2100 => x"04",
          2101 => x"a7",
          2102 => x"0b",
          2103 => x"04",
          2104 => x"a7",
          2105 => x"0b",
          2106 => x"04",
          2107 => x"a8",
          2108 => x"0b",
          2109 => x"04",
          2110 => x"a8",
          2111 => x"0b",
          2112 => x"04",
          2113 => x"a8",
          2114 => x"0b",
          2115 => x"04",
          2116 => x"a8",
          2117 => x"0b",
          2118 => x"04",
          2119 => x"a9",
          2120 => x"0b",
          2121 => x"04",
          2122 => x"a9",
          2123 => x"0b",
          2124 => x"04",
          2125 => x"a9",
          2126 => x"0b",
          2127 => x"04",
          2128 => x"a9",
          2129 => x"0b",
          2130 => x"04",
          2131 => x"aa",
          2132 => x"0b",
          2133 => x"04",
          2134 => x"aa",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"04",
          2177 => x"0c",
          2178 => x"82",
          2179 => x"83",
          2180 => x"82",
          2181 => x"80",
          2182 => x"82",
          2183 => x"83",
          2184 => x"82",
          2185 => x"80",
          2186 => x"82",
          2187 => x"83",
          2188 => x"82",
          2189 => x"80",
          2190 => x"82",
          2191 => x"83",
          2192 => x"82",
          2193 => x"80",
          2194 => x"82",
          2195 => x"83",
          2196 => x"82",
          2197 => x"80",
          2198 => x"82",
          2199 => x"83",
          2200 => x"82",
          2201 => x"80",
          2202 => x"82",
          2203 => x"83",
          2204 => x"82",
          2205 => x"80",
          2206 => x"82",
          2207 => x"83",
          2208 => x"82",
          2209 => x"80",
          2210 => x"82",
          2211 => x"83",
          2212 => x"82",
          2213 => x"80",
          2214 => x"82",
          2215 => x"83",
          2216 => x"82",
          2217 => x"80",
          2218 => x"82",
          2219 => x"83",
          2220 => x"82",
          2221 => x"80",
          2222 => x"82",
          2223 => x"83",
          2224 => x"82",
          2225 => x"80",
          2226 => x"82",
          2227 => x"83",
          2228 => x"82",
          2229 => x"ba",
          2230 => x"8c",
          2231 => x"80",
          2232 => x"8c",
          2233 => x"fe",
          2234 => x"e8",
          2235 => x"90",
          2236 => x"e8",
          2237 => x"2d",
          2238 => x"08",
          2239 => x"04",
          2240 => x"0c",
          2241 => x"82",
          2242 => x"83",
          2243 => x"82",
          2244 => x"b6",
          2245 => x"8c",
          2246 => x"80",
          2247 => x"8c",
          2248 => x"98",
          2249 => x"8c",
          2250 => x"80",
          2251 => x"8c",
          2252 => x"a5",
          2253 => x"8c",
          2254 => x"80",
          2255 => x"8c",
          2256 => x"9d",
          2257 => x"8c",
          2258 => x"80",
          2259 => x"8c",
          2260 => x"a0",
          2261 => x"8c",
          2262 => x"80",
          2263 => x"8c",
          2264 => x"aa",
          2265 => x"8c",
          2266 => x"80",
          2267 => x"8c",
          2268 => x"b3",
          2269 => x"8c",
          2270 => x"80",
          2271 => x"8c",
          2272 => x"a3",
          2273 => x"8c",
          2274 => x"80",
          2275 => x"8c",
          2276 => x"ad",
          2277 => x"8c",
          2278 => x"80",
          2279 => x"8c",
          2280 => x"ae",
          2281 => x"8c",
          2282 => x"80",
          2283 => x"8c",
          2284 => x"af",
          2285 => x"8c",
          2286 => x"80",
          2287 => x"8c",
          2288 => x"b6",
          2289 => x"8c",
          2290 => x"80",
          2291 => x"8c",
          2292 => x"b4",
          2293 => x"8c",
          2294 => x"80",
          2295 => x"8c",
          2296 => x"b9",
          2297 => x"8c",
          2298 => x"80",
          2299 => x"8c",
          2300 => x"b0",
          2301 => x"8c",
          2302 => x"80",
          2303 => x"8c",
          2304 => x"bc",
          2305 => x"8c",
          2306 => x"80",
          2307 => x"8c",
          2308 => x"bd",
          2309 => x"8c",
          2310 => x"80",
          2311 => x"8c",
          2312 => x"a5",
          2313 => x"8c",
          2314 => x"80",
          2315 => x"8c",
          2316 => x"a5",
          2317 => x"8c",
          2318 => x"80",
          2319 => x"8c",
          2320 => x"a6",
          2321 => x"8c",
          2322 => x"80",
          2323 => x"8c",
          2324 => x"b0",
          2325 => x"8c",
          2326 => x"80",
          2327 => x"8c",
          2328 => x"be",
          2329 => x"8c",
          2330 => x"80",
          2331 => x"8c",
          2332 => x"c0",
          2333 => x"8c",
          2334 => x"80",
          2335 => x"8c",
          2336 => x"c3",
          2337 => x"8c",
          2338 => x"80",
          2339 => x"8c",
          2340 => x"97",
          2341 => x"8c",
          2342 => x"80",
          2343 => x"8c",
          2344 => x"c6",
          2345 => x"8c",
          2346 => x"80",
          2347 => x"8c",
          2348 => x"d5",
          2349 => x"8c",
          2350 => x"80",
          2351 => x"8c",
          2352 => x"d3",
          2353 => x"8c",
          2354 => x"80",
          2355 => x"8c",
          2356 => x"e8",
          2357 => x"8c",
          2358 => x"80",
          2359 => x"8c",
          2360 => x"ea",
          2361 => x"8c",
          2362 => x"80",
          2363 => x"8c",
          2364 => x"ec",
          2365 => x"8c",
          2366 => x"80",
          2367 => x"8c",
          2368 => x"c3",
          2369 => x"e8",
          2370 => x"90",
          2371 => x"e8",
          2372 => x"2d",
          2373 => x"08",
          2374 => x"04",
          2375 => x"0c",
          2376 => x"82",
          2377 => x"83",
          2378 => x"82",
          2379 => x"81",
          2380 => x"82",
          2381 => x"83",
          2382 => x"82",
          2383 => x"82",
          2384 => x"8e",
          2385 => x"70",
          2386 => x"0c",
          2387 => x"aa",
          2388 => x"80",
          2389 => x"a0",
          2390 => x"82",
          2391 => x"02",
          2392 => x"0c",
          2393 => x"80",
          2394 => x"e8",
          2395 => x"08",
          2396 => x"e8",
          2397 => x"08",
          2398 => x"3f",
          2399 => x"08",
          2400 => x"dc",
          2401 => x"3d",
          2402 => x"e8",
          2403 => x"8c",
          2404 => x"82",
          2405 => x"fd",
          2406 => x"53",
          2407 => x"08",
          2408 => x"52",
          2409 => x"08",
          2410 => x"51",
          2411 => x"8c",
          2412 => x"82",
          2413 => x"54",
          2414 => x"82",
          2415 => x"04",
          2416 => x"08",
          2417 => x"e8",
          2418 => x"0d",
          2419 => x"8c",
          2420 => x"05",
          2421 => x"82",
          2422 => x"f8",
          2423 => x"8c",
          2424 => x"05",
          2425 => x"e8",
          2426 => x"08",
          2427 => x"82",
          2428 => x"fc",
          2429 => x"2e",
          2430 => x"0b",
          2431 => x"08",
          2432 => x"24",
          2433 => x"8c",
          2434 => x"05",
          2435 => x"8c",
          2436 => x"05",
          2437 => x"e8",
          2438 => x"08",
          2439 => x"e8",
          2440 => x"0c",
          2441 => x"82",
          2442 => x"fc",
          2443 => x"2e",
          2444 => x"82",
          2445 => x"8c",
          2446 => x"8c",
          2447 => x"05",
          2448 => x"38",
          2449 => x"08",
          2450 => x"82",
          2451 => x"8c",
          2452 => x"82",
          2453 => x"88",
          2454 => x"8c",
          2455 => x"05",
          2456 => x"e8",
          2457 => x"08",
          2458 => x"e8",
          2459 => x"0c",
          2460 => x"08",
          2461 => x"81",
          2462 => x"e8",
          2463 => x"0c",
          2464 => x"08",
          2465 => x"81",
          2466 => x"e8",
          2467 => x"0c",
          2468 => x"82",
          2469 => x"90",
          2470 => x"2e",
          2471 => x"8c",
          2472 => x"05",
          2473 => x"8c",
          2474 => x"05",
          2475 => x"39",
          2476 => x"08",
          2477 => x"70",
          2478 => x"08",
          2479 => x"51",
          2480 => x"08",
          2481 => x"82",
          2482 => x"85",
          2483 => x"8c",
          2484 => x"fc",
          2485 => x"70",
          2486 => x"55",
          2487 => x"72",
          2488 => x"72",
          2489 => x"06",
          2490 => x"2e",
          2491 => x"12",
          2492 => x"2e",
          2493 => x"70",
          2494 => x"33",
          2495 => x"05",
          2496 => x"12",
          2497 => x"2e",
          2498 => x"ea",
          2499 => x"8c",
          2500 => x"3d",
          2501 => x"51",
          2502 => x"05",
          2503 => x"70",
          2504 => x"0c",
          2505 => x"05",
          2506 => x"70",
          2507 => x"0c",
          2508 => x"05",
          2509 => x"70",
          2510 => x"0c",
          2511 => x"05",
          2512 => x"70",
          2513 => x"0c",
          2514 => x"71",
          2515 => x"38",
          2516 => x"95",
          2517 => x"84",
          2518 => x"71",
          2519 => x"53",
          2520 => x"52",
          2521 => x"ed",
          2522 => x"ff",
          2523 => x"3d",
          2524 => x"71",
          2525 => x"9f",
          2526 => x"55",
          2527 => x"72",
          2528 => x"74",
          2529 => x"70",
          2530 => x"38",
          2531 => x"71",
          2532 => x"38",
          2533 => x"81",
          2534 => x"ff",
          2535 => x"ff",
          2536 => x"06",
          2537 => x"82",
          2538 => x"86",
          2539 => x"74",
          2540 => x"75",
          2541 => x"90",
          2542 => x"54",
          2543 => x"27",
          2544 => x"71",
          2545 => x"53",
          2546 => x"70",
          2547 => x"0c",
          2548 => x"84",
          2549 => x"72",
          2550 => x"05",
          2551 => x"12",
          2552 => x"26",
          2553 => x"72",
          2554 => x"72",
          2555 => x"05",
          2556 => x"12",
          2557 => x"26",
          2558 => x"53",
          2559 => x"fc",
          2560 => x"70",
          2561 => x"07",
          2562 => x"54",
          2563 => x"80",
          2564 => x"70",
          2565 => x"70",
          2566 => x"ff",
          2567 => x"f8",
          2568 => x"80",
          2569 => x"53",
          2570 => x"a6",
          2571 => x"72",
          2572 => x"05",
          2573 => x"08",
          2574 => x"f7",
          2575 => x"13",
          2576 => x"84",
          2577 => x"06",
          2578 => x"53",
          2579 => x"2e",
          2580 => x"52",
          2581 => x"05",
          2582 => x"70",
          2583 => x"05",
          2584 => x"f0",
          2585 => x"8c",
          2586 => x"3d",
          2587 => x"3d",
          2588 => x"71",
          2589 => x"55",
          2590 => x"38",
          2591 => x"70",
          2592 => x"fd",
          2593 => x"70",
          2594 => x"81",
          2595 => x"51",
          2596 => x"9d",
          2597 => x"70",
          2598 => x"f7",
          2599 => x"12",
          2600 => x"84",
          2601 => x"06",
          2602 => x"53",
          2603 => x"e5",
          2604 => x"71",
          2605 => x"80",
          2606 => x"81",
          2607 => x"52",
          2608 => x"38",
          2609 => x"82",
          2610 => x"85",
          2611 => x"fa",
          2612 => x"7a",
          2613 => x"55",
          2614 => x"80",
          2615 => x"38",
          2616 => x"83",
          2617 => x"80",
          2618 => x"38",
          2619 => x"72",
          2620 => x"38",
          2621 => x"33",
          2622 => x"71",
          2623 => x"06",
          2624 => x"80",
          2625 => x"38",
          2626 => x"06",
          2627 => x"2e",
          2628 => x"81",
          2629 => x"ff",
          2630 => x"52",
          2631 => x"09",
          2632 => x"38",
          2633 => x"33",
          2634 => x"81",
          2635 => x"81",
          2636 => x"71",
          2637 => x"52",
          2638 => x"dc",
          2639 => x"0d",
          2640 => x"57",
          2641 => x"27",
          2642 => x"08",
          2643 => x"88",
          2644 => x"55",
          2645 => x"39",
          2646 => x"72",
          2647 => x"38",
          2648 => x"09",
          2649 => x"ff",
          2650 => x"f8",
          2651 => x"80",
          2652 => x"51",
          2653 => x"84",
          2654 => x"57",
          2655 => x"27",
          2656 => x"08",
          2657 => x"d0",
          2658 => x"55",
          2659 => x"39",
          2660 => x"8c",
          2661 => x"3d",
          2662 => x"3d",
          2663 => x"83",
          2664 => x"2b",
          2665 => x"3f",
          2666 => x"08",
          2667 => x"72",
          2668 => x"54",
          2669 => x"25",
          2670 => x"82",
          2671 => x"84",
          2672 => x"fb",
          2673 => x"70",
          2674 => x"53",
          2675 => x"2e",
          2676 => x"71",
          2677 => x"a0",
          2678 => x"06",
          2679 => x"12",
          2680 => x"71",
          2681 => x"81",
          2682 => x"73",
          2683 => x"ff",
          2684 => x"55",
          2685 => x"83",
          2686 => x"70",
          2687 => x"38",
          2688 => x"73",
          2689 => x"51",
          2690 => x"09",
          2691 => x"38",
          2692 => x"81",
          2693 => x"72",
          2694 => x"51",
          2695 => x"dc",
          2696 => x"0d",
          2697 => x"0d",
          2698 => x"08",
          2699 => x"38",
          2700 => x"05",
          2701 => x"9f",
          2702 => x"8c",
          2703 => x"38",
          2704 => x"39",
          2705 => x"82",
          2706 => x"86",
          2707 => x"fc",
          2708 => x"82",
          2709 => x"05",
          2710 => x"52",
          2711 => x"81",
          2712 => x"13",
          2713 => x"51",
          2714 => x"9e",
          2715 => x"38",
          2716 => x"51",
          2717 => x"97",
          2718 => x"38",
          2719 => x"51",
          2720 => x"bb",
          2721 => x"38",
          2722 => x"51",
          2723 => x"bb",
          2724 => x"38",
          2725 => x"55",
          2726 => x"87",
          2727 => x"d9",
          2728 => x"22",
          2729 => x"73",
          2730 => x"80",
          2731 => x"0b",
          2732 => x"9c",
          2733 => x"87",
          2734 => x"0c",
          2735 => x"87",
          2736 => x"0c",
          2737 => x"87",
          2738 => x"0c",
          2739 => x"87",
          2740 => x"0c",
          2741 => x"87",
          2742 => x"0c",
          2743 => x"87",
          2744 => x"0c",
          2745 => x"98",
          2746 => x"87",
          2747 => x"0c",
          2748 => x"c0",
          2749 => x"80",
          2750 => x"8c",
          2751 => x"3d",
          2752 => x"3d",
          2753 => x"87",
          2754 => x"5d",
          2755 => x"87",
          2756 => x"08",
          2757 => x"23",
          2758 => x"b8",
          2759 => x"82",
          2760 => x"c0",
          2761 => x"5a",
          2762 => x"34",
          2763 => x"b0",
          2764 => x"84",
          2765 => x"c0",
          2766 => x"5a",
          2767 => x"34",
          2768 => x"a8",
          2769 => x"86",
          2770 => x"c0",
          2771 => x"5c",
          2772 => x"23",
          2773 => x"a0",
          2774 => x"8a",
          2775 => x"7d",
          2776 => x"ff",
          2777 => x"7b",
          2778 => x"06",
          2779 => x"33",
          2780 => x"33",
          2781 => x"33",
          2782 => x"33",
          2783 => x"33",
          2784 => x"ff",
          2785 => x"81",
          2786 => x"98",
          2787 => x"3d",
          2788 => x"3d",
          2789 => x"05",
          2790 => x"70",
          2791 => x"52",
          2792 => x"0b",
          2793 => x"34",
          2794 => x"04",
          2795 => x"77",
          2796 => x"87",
          2797 => x"81",
          2798 => x"55",
          2799 => x"94",
          2800 => x"80",
          2801 => x"87",
          2802 => x"51",
          2803 => x"96",
          2804 => x"06",
          2805 => x"70",
          2806 => x"38",
          2807 => x"70",
          2808 => x"51",
          2809 => x"72",
          2810 => x"81",
          2811 => x"70",
          2812 => x"38",
          2813 => x"70",
          2814 => x"51",
          2815 => x"38",
          2816 => x"06",
          2817 => x"94",
          2818 => x"80",
          2819 => x"87",
          2820 => x"52",
          2821 => x"75",
          2822 => x"0c",
          2823 => x"04",
          2824 => x"02",
          2825 => x"0b",
          2826 => x"d4",
          2827 => x"ff",
          2828 => x"56",
          2829 => x"84",
          2830 => x"2e",
          2831 => x"c0",
          2832 => x"70",
          2833 => x"2a",
          2834 => x"53",
          2835 => x"80",
          2836 => x"71",
          2837 => x"81",
          2838 => x"70",
          2839 => x"81",
          2840 => x"06",
          2841 => x"80",
          2842 => x"71",
          2843 => x"81",
          2844 => x"70",
          2845 => x"73",
          2846 => x"51",
          2847 => x"80",
          2848 => x"2e",
          2849 => x"c0",
          2850 => x"75",
          2851 => x"3d",
          2852 => x"3d",
          2853 => x"80",
          2854 => x"81",
          2855 => x"53",
          2856 => x"2e",
          2857 => x"71",
          2858 => x"81",
          2859 => x"82",
          2860 => x"70",
          2861 => x"59",
          2862 => x"87",
          2863 => x"51",
          2864 => x"86",
          2865 => x"94",
          2866 => x"08",
          2867 => x"70",
          2868 => x"54",
          2869 => x"2e",
          2870 => x"91",
          2871 => x"06",
          2872 => x"d7",
          2873 => x"32",
          2874 => x"51",
          2875 => x"2e",
          2876 => x"93",
          2877 => x"06",
          2878 => x"ff",
          2879 => x"81",
          2880 => x"87",
          2881 => x"52",
          2882 => x"86",
          2883 => x"94",
          2884 => x"72",
          2885 => x"74",
          2886 => x"ff",
          2887 => x"57",
          2888 => x"38",
          2889 => x"dc",
          2890 => x"0d",
          2891 => x"0d",
          2892 => x"87",
          2893 => x"81",
          2894 => x"52",
          2895 => x"84",
          2896 => x"2e",
          2897 => x"c0",
          2898 => x"70",
          2899 => x"2a",
          2900 => x"51",
          2901 => x"80",
          2902 => x"71",
          2903 => x"51",
          2904 => x"80",
          2905 => x"2e",
          2906 => x"c0",
          2907 => x"71",
          2908 => x"ff",
          2909 => x"dc",
          2910 => x"3d",
          2911 => x"3d",
          2912 => x"82",
          2913 => x"70",
          2914 => x"52",
          2915 => x"94",
          2916 => x"80",
          2917 => x"87",
          2918 => x"52",
          2919 => x"82",
          2920 => x"06",
          2921 => x"ff",
          2922 => x"2e",
          2923 => x"81",
          2924 => x"87",
          2925 => x"52",
          2926 => x"86",
          2927 => x"94",
          2928 => x"08",
          2929 => x"70",
          2930 => x"53",
          2931 => x"8c",
          2932 => x"3d",
          2933 => x"3d",
          2934 => x"9e",
          2935 => x"9c",
          2936 => x"51",
          2937 => x"2e",
          2938 => x"87",
          2939 => x"08",
          2940 => x"0c",
          2941 => x"a8",
          2942 => x"dc",
          2943 => x"9e",
          2944 => x"87",
          2945 => x"c0",
          2946 => x"82",
          2947 => x"87",
          2948 => x"08",
          2949 => x"0c",
          2950 => x"a0",
          2951 => x"ec",
          2952 => x"9e",
          2953 => x"87",
          2954 => x"c0",
          2955 => x"82",
          2956 => x"87",
          2957 => x"08",
          2958 => x"0c",
          2959 => x"b8",
          2960 => x"fc",
          2961 => x"9e",
          2962 => x"88",
          2963 => x"c0",
          2964 => x"82",
          2965 => x"87",
          2966 => x"08",
          2967 => x"0c",
          2968 => x"80",
          2969 => x"82",
          2970 => x"87",
          2971 => x"08",
          2972 => x"0c",
          2973 => x"88",
          2974 => x"94",
          2975 => x"9e",
          2976 => x"88",
          2977 => x"0b",
          2978 => x"34",
          2979 => x"c0",
          2980 => x"70",
          2981 => x"06",
          2982 => x"70",
          2983 => x"38",
          2984 => x"82",
          2985 => x"80",
          2986 => x"9e",
          2987 => x"88",
          2988 => x"51",
          2989 => x"80",
          2990 => x"81",
          2991 => x"88",
          2992 => x"0b",
          2993 => x"90",
          2994 => x"80",
          2995 => x"52",
          2996 => x"2e",
          2997 => x"52",
          2998 => x"9f",
          2999 => x"87",
          3000 => x"08",
          3001 => x"80",
          3002 => x"52",
          3003 => x"83",
          3004 => x"71",
          3005 => x"34",
          3006 => x"c0",
          3007 => x"70",
          3008 => x"06",
          3009 => x"70",
          3010 => x"38",
          3011 => x"82",
          3012 => x"80",
          3013 => x"9e",
          3014 => x"90",
          3015 => x"51",
          3016 => x"80",
          3017 => x"81",
          3018 => x"88",
          3019 => x"0b",
          3020 => x"90",
          3021 => x"80",
          3022 => x"52",
          3023 => x"2e",
          3024 => x"52",
          3025 => x"a3",
          3026 => x"87",
          3027 => x"08",
          3028 => x"80",
          3029 => x"52",
          3030 => x"83",
          3031 => x"71",
          3032 => x"34",
          3033 => x"c0",
          3034 => x"70",
          3035 => x"06",
          3036 => x"70",
          3037 => x"38",
          3038 => x"82",
          3039 => x"80",
          3040 => x"9e",
          3041 => x"80",
          3042 => x"51",
          3043 => x"80",
          3044 => x"81",
          3045 => x"88",
          3046 => x"0b",
          3047 => x"90",
          3048 => x"80",
          3049 => x"52",
          3050 => x"83",
          3051 => x"71",
          3052 => x"34",
          3053 => x"90",
          3054 => x"80",
          3055 => x"2a",
          3056 => x"70",
          3057 => x"34",
          3058 => x"c0",
          3059 => x"70",
          3060 => x"51",
          3061 => x"80",
          3062 => x"81",
          3063 => x"88",
          3064 => x"c0",
          3065 => x"70",
          3066 => x"70",
          3067 => x"51",
          3068 => x"88",
          3069 => x"0b",
          3070 => x"90",
          3071 => x"06",
          3072 => x"70",
          3073 => x"38",
          3074 => x"82",
          3075 => x"87",
          3076 => x"08",
          3077 => x"51",
          3078 => x"88",
          3079 => x"3d",
          3080 => x"3d",
          3081 => x"fc",
          3082 => x"3f",
          3083 => x"33",
          3084 => x"2e",
          3085 => x"f2",
          3086 => x"cb",
          3087 => x"a4",
          3088 => x"3f",
          3089 => x"33",
          3090 => x"2e",
          3091 => x"87",
          3092 => x"87",
          3093 => x"54",
          3094 => x"bc",
          3095 => x"3f",
          3096 => x"33",
          3097 => x"2e",
          3098 => x"87",
          3099 => x"87",
          3100 => x"54",
          3101 => x"d8",
          3102 => x"3f",
          3103 => x"33",
          3104 => x"2e",
          3105 => x"87",
          3106 => x"87",
          3107 => x"54",
          3108 => x"f4",
          3109 => x"3f",
          3110 => x"33",
          3111 => x"2e",
          3112 => x"87",
          3113 => x"87",
          3114 => x"54",
          3115 => x"90",
          3116 => x"3f",
          3117 => x"33",
          3118 => x"2e",
          3119 => x"87",
          3120 => x"87",
          3121 => x"54",
          3122 => x"ac",
          3123 => x"3f",
          3124 => x"33",
          3125 => x"2e",
          3126 => x"88",
          3127 => x"81",
          3128 => x"8e",
          3129 => x"88",
          3130 => x"73",
          3131 => x"38",
          3132 => x"33",
          3133 => x"e8",
          3134 => x"3f",
          3135 => x"33",
          3136 => x"2e",
          3137 => x"88",
          3138 => x"81",
          3139 => x"8d",
          3140 => x"88",
          3141 => x"73",
          3142 => x"38",
          3143 => x"51",
          3144 => x"82",
          3145 => x"54",
          3146 => x"88",
          3147 => x"bc",
          3148 => x"3f",
          3149 => x"33",
          3150 => x"2e",
          3151 => x"f4",
          3152 => x"c3",
          3153 => x"a5",
          3154 => x"80",
          3155 => x"81",
          3156 => x"87",
          3157 => x"88",
          3158 => x"73",
          3159 => x"38",
          3160 => x"51",
          3161 => x"81",
          3162 => x"87",
          3163 => x"88",
          3164 => x"81",
          3165 => x"8c",
          3166 => x"88",
          3167 => x"81",
          3168 => x"8c",
          3169 => x"88",
          3170 => x"81",
          3171 => x"8c",
          3172 => x"f5",
          3173 => x"ef",
          3174 => x"8c",
          3175 => x"f5",
          3176 => x"c7",
          3177 => x"90",
          3178 => x"84",
          3179 => x"51",
          3180 => x"82",
          3181 => x"bd",
          3182 => x"76",
          3183 => x"54",
          3184 => x"08",
          3185 => x"a0",
          3186 => x"3f",
          3187 => x"33",
          3188 => x"2e",
          3189 => x"88",
          3190 => x"bd",
          3191 => x"75",
          3192 => x"3f",
          3193 => x"08",
          3194 => x"29",
          3195 => x"54",
          3196 => x"dc",
          3197 => x"f6",
          3198 => x"ef",
          3199 => x"9e",
          3200 => x"80",
          3201 => x"82",
          3202 => x"56",
          3203 => x"52",
          3204 => x"c7",
          3205 => x"dc",
          3206 => x"c0",
          3207 => x"31",
          3208 => x"8c",
          3209 => x"81",
          3210 => x"8b",
          3211 => x"85",
          3212 => x"d3",
          3213 => x"0d",
          3214 => x"0d",
          3215 => x"33",
          3216 => x"71",
          3217 => x"38",
          3218 => x"0b",
          3219 => x"d0",
          3220 => x"08",
          3221 => x"a4",
          3222 => x"81",
          3223 => x"97",
          3224 => x"b4",
          3225 => x"81",
          3226 => x"8b",
          3227 => x"c0",
          3228 => x"81",
          3229 => x"85",
          3230 => x"3d",
          3231 => x"88",
          3232 => x"80",
          3233 => x"96",
          3234 => x"82",
          3235 => x"87",
          3236 => x"0c",
          3237 => x"0d",
          3238 => x"08",
          3239 => x"a4",
          3240 => x"8c",
          3241 => x"8c",
          3242 => x"11",
          3243 => x"53",
          3244 => x"f8",
          3245 => x"70",
          3246 => x"0c",
          3247 => x"82",
          3248 => x"84",
          3249 => x"f9",
          3250 => x"7b",
          3251 => x"a0",
          3252 => x"08",
          3253 => x"90",
          3254 => x"58",
          3255 => x"53",
          3256 => x"ba",
          3257 => x"88",
          3258 => x"51",
          3259 => x"76",
          3260 => x"12",
          3261 => x"0c",
          3262 => x"0c",
          3263 => x"0c",
          3264 => x"0c",
          3265 => x"0c",
          3266 => x"0c",
          3267 => x"0c",
          3268 => x"0c",
          3269 => x"0c",
          3270 => x"0c",
          3271 => x"73",
          3272 => x"16",
          3273 => x"15",
          3274 => x"8c",
          3275 => x"3d",
          3276 => x"3d",
          3277 => x"11",
          3278 => x"08",
          3279 => x"71",
          3280 => x"09",
          3281 => x"38",
          3282 => x"70",
          3283 => x"70",
          3284 => x"81",
          3285 => x"84",
          3286 => x"84",
          3287 => x"88",
          3288 => x"8c",
          3289 => x"53",
          3290 => x"73",
          3291 => x"c4",
          3292 => x"0c",
          3293 => x"0b",
          3294 => x"72",
          3295 => x"0c",
          3296 => x"73",
          3297 => x"51",
          3298 => x"2e",
          3299 => x"b3",
          3300 => x"08",
          3301 => x"52",
          3302 => x"09",
          3303 => x"38",
          3304 => x"12",
          3305 => x"94",
          3306 => x"15",
          3307 => x"13",
          3308 => x"12",
          3309 => x"08",
          3310 => x"70",
          3311 => x"52",
          3312 => x"72",
          3313 => x"0c",
          3314 => x"04",
          3315 => x"79",
          3316 => x"76",
          3317 => x"b5",
          3318 => x"f0",
          3319 => x"c4",
          3320 => x"75",
          3321 => x"8f",
          3322 => x"08",
          3323 => x"c7",
          3324 => x"08",
          3325 => x"83",
          3326 => x"fc",
          3327 => x"70",
          3328 => x"91",
          3329 => x"dc",
          3330 => x"dc",
          3331 => x"82",
          3332 => x"07",
          3333 => x"8c",
          3334 => x"70",
          3335 => x"07",
          3336 => x"07",
          3337 => x"51",
          3338 => x"54",
          3339 => x"09",
          3340 => x"d9",
          3341 => x"76",
          3342 => x"80",
          3343 => x"0b",
          3344 => x"08",
          3345 => x"8c",
          3346 => x"05",
          3347 => x"c0",
          3348 => x"08",
          3349 => x"38",
          3350 => x"87",
          3351 => x"08",
          3352 => x"88",
          3353 => x"17",
          3354 => x"17",
          3355 => x"14",
          3356 => x"08",
          3357 => x"0c",
          3358 => x"fd",
          3359 => x"52",
          3360 => x"08",
          3361 => x"3f",
          3362 => x"08",
          3363 => x"8c",
          3364 => x"3d",
          3365 => x"3d",
          3366 => x"71",
          3367 => x"38",
          3368 => x"fd",
          3369 => x"3d",
          3370 => x"3d",
          3371 => x"05",
          3372 => x"8a",
          3373 => x"06",
          3374 => x"51",
          3375 => x"8c",
          3376 => x"71",
          3377 => x"38",
          3378 => x"82",
          3379 => x"81",
          3380 => x"f8",
          3381 => x"82",
          3382 => x"52",
          3383 => x"85",
          3384 => x"71",
          3385 => x"0d",
          3386 => x"0d",
          3387 => x"33",
          3388 => x"08",
          3389 => x"f0",
          3390 => x"ff",
          3391 => x"82",
          3392 => x"84",
          3393 => x"fd",
          3394 => x"54",
          3395 => x"81",
          3396 => x"53",
          3397 => x"8e",
          3398 => x"ff",
          3399 => x"14",
          3400 => x"3f",
          3401 => x"3d",
          3402 => x"3d",
          3403 => x"8c",
          3404 => x"82",
          3405 => x"56",
          3406 => x"70",
          3407 => x"53",
          3408 => x"2e",
          3409 => x"81",
          3410 => x"81",
          3411 => x"da",
          3412 => x"74",
          3413 => x"0c",
          3414 => x"04",
          3415 => x"66",
          3416 => x"78",
          3417 => x"5a",
          3418 => x"80",
          3419 => x"38",
          3420 => x"09",
          3421 => x"de",
          3422 => x"7a",
          3423 => x"5c",
          3424 => x"5b",
          3425 => x"09",
          3426 => x"38",
          3427 => x"39",
          3428 => x"09",
          3429 => x"38",
          3430 => x"70",
          3431 => x"33",
          3432 => x"2e",
          3433 => x"92",
          3434 => x"19",
          3435 => x"70",
          3436 => x"33",
          3437 => x"53",
          3438 => x"16",
          3439 => x"26",
          3440 => x"88",
          3441 => x"05",
          3442 => x"05",
          3443 => x"05",
          3444 => x"5b",
          3445 => x"80",
          3446 => x"30",
          3447 => x"80",
          3448 => x"cc",
          3449 => x"70",
          3450 => x"25",
          3451 => x"54",
          3452 => x"53",
          3453 => x"8c",
          3454 => x"07",
          3455 => x"05",
          3456 => x"5a",
          3457 => x"83",
          3458 => x"54",
          3459 => x"27",
          3460 => x"16",
          3461 => x"06",
          3462 => x"80",
          3463 => x"aa",
          3464 => x"cf",
          3465 => x"73",
          3466 => x"81",
          3467 => x"80",
          3468 => x"38",
          3469 => x"2e",
          3470 => x"81",
          3471 => x"80",
          3472 => x"8a",
          3473 => x"39",
          3474 => x"2e",
          3475 => x"73",
          3476 => x"8a",
          3477 => x"d3",
          3478 => x"80",
          3479 => x"80",
          3480 => x"ee",
          3481 => x"39",
          3482 => x"71",
          3483 => x"53",
          3484 => x"54",
          3485 => x"2e",
          3486 => x"15",
          3487 => x"33",
          3488 => x"72",
          3489 => x"81",
          3490 => x"39",
          3491 => x"56",
          3492 => x"27",
          3493 => x"51",
          3494 => x"75",
          3495 => x"72",
          3496 => x"38",
          3497 => x"df",
          3498 => x"16",
          3499 => x"7b",
          3500 => x"38",
          3501 => x"f2",
          3502 => x"77",
          3503 => x"12",
          3504 => x"53",
          3505 => x"5c",
          3506 => x"5c",
          3507 => x"5c",
          3508 => x"5c",
          3509 => x"51",
          3510 => x"fd",
          3511 => x"82",
          3512 => x"06",
          3513 => x"80",
          3514 => x"77",
          3515 => x"53",
          3516 => x"18",
          3517 => x"72",
          3518 => x"c4",
          3519 => x"70",
          3520 => x"25",
          3521 => x"55",
          3522 => x"8d",
          3523 => x"2e",
          3524 => x"30",
          3525 => x"5b",
          3526 => x"8f",
          3527 => x"7b",
          3528 => x"dc",
          3529 => x"8c",
          3530 => x"ff",
          3531 => x"75",
          3532 => x"a7",
          3533 => x"dc",
          3534 => x"74",
          3535 => x"a7",
          3536 => x"80",
          3537 => x"38",
          3538 => x"72",
          3539 => x"54",
          3540 => x"72",
          3541 => x"05",
          3542 => x"17",
          3543 => x"77",
          3544 => x"51",
          3545 => x"9f",
          3546 => x"72",
          3547 => x"79",
          3548 => x"81",
          3549 => x"72",
          3550 => x"38",
          3551 => x"05",
          3552 => x"ad",
          3553 => x"17",
          3554 => x"81",
          3555 => x"b0",
          3556 => x"38",
          3557 => x"81",
          3558 => x"06",
          3559 => x"9f",
          3560 => x"55",
          3561 => x"97",
          3562 => x"f9",
          3563 => x"81",
          3564 => x"8b",
          3565 => x"16",
          3566 => x"73",
          3567 => x"96",
          3568 => x"e0",
          3569 => x"17",
          3570 => x"33",
          3571 => x"f9",
          3572 => x"f2",
          3573 => x"16",
          3574 => x"7b",
          3575 => x"38",
          3576 => x"c6",
          3577 => x"96",
          3578 => x"fd",
          3579 => x"3d",
          3580 => x"05",
          3581 => x"52",
          3582 => x"e0",
          3583 => x"0d",
          3584 => x"0d",
          3585 => x"f8",
          3586 => x"88",
          3587 => x"51",
          3588 => x"82",
          3589 => x"53",
          3590 => x"80",
          3591 => x"f8",
          3592 => x"0d",
          3593 => x"0d",
          3594 => x"08",
          3595 => x"f0",
          3596 => x"88",
          3597 => x"52",
          3598 => x"3f",
          3599 => x"f0",
          3600 => x"0d",
          3601 => x"0d",
          3602 => x"8c",
          3603 => x"56",
          3604 => x"80",
          3605 => x"2e",
          3606 => x"82",
          3607 => x"52",
          3608 => x"8c",
          3609 => x"ff",
          3610 => x"80",
          3611 => x"38",
          3612 => x"b9",
          3613 => x"32",
          3614 => x"80",
          3615 => x"52",
          3616 => x"8b",
          3617 => x"2e",
          3618 => x"14",
          3619 => x"9f",
          3620 => x"38",
          3621 => x"73",
          3622 => x"38",
          3623 => x"72",
          3624 => x"14",
          3625 => x"f8",
          3626 => x"af",
          3627 => x"52",
          3628 => x"8a",
          3629 => x"3f",
          3630 => x"82",
          3631 => x"87",
          3632 => x"fe",
          3633 => x"8c",
          3634 => x"82",
          3635 => x"77",
          3636 => x"53",
          3637 => x"72",
          3638 => x"0c",
          3639 => x"04",
          3640 => x"7a",
          3641 => x"80",
          3642 => x"58",
          3643 => x"33",
          3644 => x"a0",
          3645 => x"06",
          3646 => x"13",
          3647 => x"39",
          3648 => x"09",
          3649 => x"38",
          3650 => x"11",
          3651 => x"08",
          3652 => x"54",
          3653 => x"2e",
          3654 => x"80",
          3655 => x"08",
          3656 => x"0c",
          3657 => x"33",
          3658 => x"80",
          3659 => x"38",
          3660 => x"80",
          3661 => x"38",
          3662 => x"57",
          3663 => x"0c",
          3664 => x"33",
          3665 => x"39",
          3666 => x"74",
          3667 => x"38",
          3668 => x"80",
          3669 => x"89",
          3670 => x"38",
          3671 => x"d0",
          3672 => x"55",
          3673 => x"80",
          3674 => x"39",
          3675 => x"d9",
          3676 => x"80",
          3677 => x"27",
          3678 => x"80",
          3679 => x"89",
          3680 => x"70",
          3681 => x"55",
          3682 => x"70",
          3683 => x"55",
          3684 => x"27",
          3685 => x"14",
          3686 => x"06",
          3687 => x"74",
          3688 => x"73",
          3689 => x"38",
          3690 => x"14",
          3691 => x"05",
          3692 => x"08",
          3693 => x"54",
          3694 => x"39",
          3695 => x"84",
          3696 => x"55",
          3697 => x"81",
          3698 => x"8c",
          3699 => x"3d",
          3700 => x"3d",
          3701 => x"5a",
          3702 => x"7a",
          3703 => x"08",
          3704 => x"53",
          3705 => x"09",
          3706 => x"38",
          3707 => x"0c",
          3708 => x"ad",
          3709 => x"06",
          3710 => x"76",
          3711 => x"0c",
          3712 => x"33",
          3713 => x"73",
          3714 => x"81",
          3715 => x"38",
          3716 => x"05",
          3717 => x"08",
          3718 => x"53",
          3719 => x"2e",
          3720 => x"57",
          3721 => x"2e",
          3722 => x"39",
          3723 => x"13",
          3724 => x"08",
          3725 => x"53",
          3726 => x"55",
          3727 => x"80",
          3728 => x"14",
          3729 => x"88",
          3730 => x"27",
          3731 => x"eb",
          3732 => x"53",
          3733 => x"89",
          3734 => x"38",
          3735 => x"55",
          3736 => x"8a",
          3737 => x"a0",
          3738 => x"c2",
          3739 => x"74",
          3740 => x"e0",
          3741 => x"ff",
          3742 => x"d0",
          3743 => x"ff",
          3744 => x"90",
          3745 => x"38",
          3746 => x"81",
          3747 => x"53",
          3748 => x"ca",
          3749 => x"27",
          3750 => x"77",
          3751 => x"08",
          3752 => x"0c",
          3753 => x"33",
          3754 => x"ff",
          3755 => x"80",
          3756 => x"74",
          3757 => x"79",
          3758 => x"74",
          3759 => x"0c",
          3760 => x"04",
          3761 => x"76",
          3762 => x"98",
          3763 => x"2b",
          3764 => x"72",
          3765 => x"82",
          3766 => x"51",
          3767 => x"80",
          3768 => x"dc",
          3769 => x"53",
          3770 => x"9c",
          3771 => x"d8",
          3772 => x"02",
          3773 => x"05",
          3774 => x"52",
          3775 => x"72",
          3776 => x"06",
          3777 => x"53",
          3778 => x"dc",
          3779 => x"0d",
          3780 => x"0d",
          3781 => x"05",
          3782 => x"71",
          3783 => x"53",
          3784 => x"9f",
          3785 => x"f3",
          3786 => x"51",
          3787 => x"88",
          3788 => x"3f",
          3789 => x"05",
          3790 => x"34",
          3791 => x"06",
          3792 => x"76",
          3793 => x"3f",
          3794 => x"86",
          3795 => x"f6",
          3796 => x"02",
          3797 => x"05",
          3798 => x"05",
          3799 => x"82",
          3800 => x"70",
          3801 => x"88",
          3802 => x"08",
          3803 => x"5a",
          3804 => x"80",
          3805 => x"74",
          3806 => x"3f",
          3807 => x"33",
          3808 => x"82",
          3809 => x"81",
          3810 => x"58",
          3811 => x"bc",
          3812 => x"dc",
          3813 => x"82",
          3814 => x"70",
          3815 => x"88",
          3816 => x"08",
          3817 => x"74",
          3818 => x"38",
          3819 => x"52",
          3820 => x"9f",
          3821 => x"a8",
          3822 => x"55",
          3823 => x"a8",
          3824 => x"ff",
          3825 => x"75",
          3826 => x"80",
          3827 => x"a8",
          3828 => x"2e",
          3829 => x"89",
          3830 => x"75",
          3831 => x"38",
          3832 => x"33",
          3833 => x"38",
          3834 => x"05",
          3835 => x"78",
          3836 => x"80",
          3837 => x"82",
          3838 => x"52",
          3839 => x"fd",
          3840 => x"89",
          3841 => x"80",
          3842 => x"8c",
          3843 => x"dc",
          3844 => x"57",
          3845 => x"89",
          3846 => x"80",
          3847 => x"82",
          3848 => x"80",
          3849 => x"89",
          3850 => x"80",
          3851 => x"3d",
          3852 => x"80",
          3853 => x"82",
          3854 => x"80",
          3855 => x"75",
          3856 => x"3f",
          3857 => x"08",
          3858 => x"82",
          3859 => x"25",
          3860 => x"8c",
          3861 => x"05",
          3862 => x"55",
          3863 => x"75",
          3864 => x"81",
          3865 => x"f0",
          3866 => x"ff",
          3867 => x"2e",
          3868 => x"ff",
          3869 => x"3d",
          3870 => x"3d",
          3871 => x"08",
          3872 => x"5a",
          3873 => x"58",
          3874 => x"82",
          3875 => x"51",
          3876 => x"3f",
          3877 => x"08",
          3878 => x"ff",
          3879 => x"a4",
          3880 => x"80",
          3881 => x"3d",
          3882 => x"80",
          3883 => x"82",
          3884 => x"80",
          3885 => x"75",
          3886 => x"3f",
          3887 => x"08",
          3888 => x"55",
          3889 => x"8c",
          3890 => x"8e",
          3891 => x"dc",
          3892 => x"70",
          3893 => x"80",
          3894 => x"09",
          3895 => x"72",
          3896 => x"51",
          3897 => x"77",
          3898 => x"73",
          3899 => x"82",
          3900 => x"8c",
          3901 => x"51",
          3902 => x"3f",
          3903 => x"08",
          3904 => x"38",
          3905 => x"51",
          3906 => x"78",
          3907 => x"81",
          3908 => x"75",
          3909 => x"d5",
          3910 => x"51",
          3911 => x"ab",
          3912 => x"82",
          3913 => x"74",
          3914 => x"77",
          3915 => x"0c",
          3916 => x"04",
          3917 => x"7c",
          3918 => x"71",
          3919 => x"59",
          3920 => x"a0",
          3921 => x"06",
          3922 => x"33",
          3923 => x"77",
          3924 => x"38",
          3925 => x"5b",
          3926 => x"56",
          3927 => x"a0",
          3928 => x"06",
          3929 => x"75",
          3930 => x"80",
          3931 => x"29",
          3932 => x"05",
          3933 => x"55",
          3934 => x"82",
          3935 => x"53",
          3936 => x"08",
          3937 => x"3f",
          3938 => x"08",
          3939 => x"84",
          3940 => x"74",
          3941 => x"38",
          3942 => x"88",
          3943 => x"fc",
          3944 => x"39",
          3945 => x"8c",
          3946 => x"53",
          3947 => x"f6",
          3948 => x"8c",
          3949 => x"2e",
          3950 => x"53",
          3951 => x"51",
          3952 => x"82",
          3953 => x"81",
          3954 => x"74",
          3955 => x"54",
          3956 => x"14",
          3957 => x"06",
          3958 => x"74",
          3959 => x"38",
          3960 => x"82",
          3961 => x"8c",
          3962 => x"d3",
          3963 => x"3d",
          3964 => x"05",
          3965 => x"33",
          3966 => x"0b",
          3967 => x"82",
          3968 => x"5b",
          3969 => x"08",
          3970 => x"82",
          3971 => x"54",
          3972 => x"38",
          3973 => x"b4",
          3974 => x"dc",
          3975 => x"a4",
          3976 => x"dc",
          3977 => x"80",
          3978 => x"53",
          3979 => x"08",
          3980 => x"dc",
          3981 => x"ed",
          3982 => x"dc",
          3983 => x"8b",
          3984 => x"a8",
          3985 => x"3f",
          3986 => x"82",
          3987 => x"53",
          3988 => x"90",
          3989 => x"54",
          3990 => x"3f",
          3991 => x"08",
          3992 => x"dc",
          3993 => x"09",
          3994 => x"c1",
          3995 => x"dc",
          3996 => x"fa",
          3997 => x"dc",
          3998 => x"0b",
          3999 => x"08",
          4000 => x"82",
          4001 => x"ff",
          4002 => x"55",
          4003 => x"34",
          4004 => x"81",
          4005 => x"75",
          4006 => x"3f",
          4007 => x"09",
          4008 => x"a7",
          4009 => x"81",
          4010 => x"a0",
          4011 => x"5d",
          4012 => x"82",
          4013 => x"98",
          4014 => x"2c",
          4015 => x"ff",
          4016 => x"78",
          4017 => x"82",
          4018 => x"70",
          4019 => x"98",
          4020 => x"fc",
          4021 => x"2b",
          4022 => x"71",
          4023 => x"70",
          4024 => x"f8",
          4025 => x"08",
          4026 => x"51",
          4027 => x"59",
          4028 => x"5d",
          4029 => x"73",
          4030 => x"e9",
          4031 => x"27",
          4032 => x"81",
          4033 => x"81",
          4034 => x"70",
          4035 => x"55",
          4036 => x"80",
          4037 => x"53",
          4038 => x"51",
          4039 => x"82",
          4040 => x"81",
          4041 => x"73",
          4042 => x"38",
          4043 => x"fc",
          4044 => x"b1",
          4045 => x"80",
          4046 => x"80",
          4047 => x"98",
          4048 => x"ff",
          4049 => x"55",
          4050 => x"97",
          4051 => x"74",
          4052 => x"f6",
          4053 => x"8c",
          4054 => x"ff",
          4055 => x"cc",
          4056 => x"80",
          4057 => x"2e",
          4058 => x"81",
          4059 => x"82",
          4060 => x"74",
          4061 => x"98",
          4062 => x"fc",
          4063 => x"2b",
          4064 => x"70",
          4065 => x"82",
          4066 => x"dc",
          4067 => x"51",
          4068 => x"58",
          4069 => x"77",
          4070 => x"06",
          4071 => x"81",
          4072 => x"08",
          4073 => x"0b",
          4074 => x"34",
          4075 => x"8c",
          4076 => x"39",
          4077 => x"80",
          4078 => x"8c",
          4079 => x"af",
          4080 => x"7d",
          4081 => x"73",
          4082 => x"e1",
          4083 => x"29",
          4084 => x"05",
          4085 => x"04",
          4086 => x"33",
          4087 => x"2e",
          4088 => x"82",
          4089 => x"55",
          4090 => x"ab",
          4091 => x"2b",
          4092 => x"51",
          4093 => x"24",
          4094 => x"1a",
          4095 => x"81",
          4096 => x"81",
          4097 => x"81",
          4098 => x"70",
          4099 => x"8d",
          4100 => x"51",
          4101 => x"82",
          4102 => x"81",
          4103 => x"74",
          4104 => x"34",
          4105 => x"ae",
          4106 => x"34",
          4107 => x"33",
          4108 => x"27",
          4109 => x"14",
          4110 => x"8d",
          4111 => x"8d",
          4112 => x"81",
          4113 => x"81",
          4114 => x"70",
          4115 => x"8d",
          4116 => x"51",
          4117 => x"77",
          4118 => x"74",
          4119 => x"52",
          4120 => x"3f",
          4121 => x"0a",
          4122 => x"0a",
          4123 => x"2c",
          4124 => x"33",
          4125 => x"73",
          4126 => x"38",
          4127 => x"33",
          4128 => x"70",
          4129 => x"8d",
          4130 => x"51",
          4131 => x"77",
          4132 => x"38",
          4133 => x"92",
          4134 => x"80",
          4135 => x"80",
          4136 => x"98",
          4137 => x"84",
          4138 => x"55",
          4139 => x"e4",
          4140 => x"39",
          4141 => x"33",
          4142 => x"06",
          4143 => x"80",
          4144 => x"38",
          4145 => x"33",
          4146 => x"73",
          4147 => x"34",
          4148 => x"73",
          4149 => x"34",
          4150 => x"ce",
          4151 => x"88",
          4152 => x"2b",
          4153 => x"82",
          4154 => x"57",
          4155 => x"74",
          4156 => x"38",
          4157 => x"81",
          4158 => x"34",
          4159 => x"e7",
          4160 => x"81",
          4161 => x"81",
          4162 => x"70",
          4163 => x"8d",
          4164 => x"51",
          4165 => x"24",
          4166 => x"51",
          4167 => x"82",
          4168 => x"70",
          4169 => x"98",
          4170 => x"84",
          4171 => x"56",
          4172 => x"24",
          4173 => x"88",
          4174 => x"3f",
          4175 => x"0a",
          4176 => x"0a",
          4177 => x"2c",
          4178 => x"33",
          4179 => x"75",
          4180 => x"38",
          4181 => x"82",
          4182 => x"7a",
          4183 => x"74",
          4184 => x"e6",
          4185 => x"8d",
          4186 => x"51",
          4187 => x"82",
          4188 => x"81",
          4189 => x"73",
          4190 => x"8d",
          4191 => x"73",
          4192 => x"c9",
          4193 => x"73",
          4194 => x"f3",
          4195 => x"bd",
          4196 => x"34",
          4197 => x"82",
          4198 => x"54",
          4199 => x"fa",
          4200 => x"51",
          4201 => x"82",
          4202 => x"ff",
          4203 => x"82",
          4204 => x"73",
          4205 => x"54",
          4206 => x"8d",
          4207 => x"8d",
          4208 => x"55",
          4209 => x"f9",
          4210 => x"14",
          4211 => x"8d",
          4212 => x"98",
          4213 => x"2c",
          4214 => x"06",
          4215 => x"74",
          4216 => x"38",
          4217 => x"81",
          4218 => x"34",
          4219 => x"e5",
          4220 => x"81",
          4221 => x"81",
          4222 => x"70",
          4223 => x"8d",
          4224 => x"51",
          4225 => x"24",
          4226 => x"51",
          4227 => x"82",
          4228 => x"70",
          4229 => x"98",
          4230 => x"84",
          4231 => x"56",
          4232 => x"24",
          4233 => x"88",
          4234 => x"3f",
          4235 => x"0a",
          4236 => x"0a",
          4237 => x"2c",
          4238 => x"33",
          4239 => x"75",
          4240 => x"38",
          4241 => x"82",
          4242 => x"70",
          4243 => x"82",
          4244 => x"59",
          4245 => x"77",
          4246 => x"38",
          4247 => x"73",
          4248 => x"34",
          4249 => x"33",
          4250 => x"be",
          4251 => x"88",
          4252 => x"ff",
          4253 => x"84",
          4254 => x"54",
          4255 => x"dc",
          4256 => x"39",
          4257 => x"82",
          4258 => x"55",
          4259 => x"a4",
          4260 => x"cb",
          4261 => x"8c",
          4262 => x"8d",
          4263 => x"8c",
          4264 => x"ff",
          4265 => x"53",
          4266 => x"51",
          4267 => x"93",
          4268 => x"39",
          4269 => x"82",
          4270 => x"fc",
          4271 => x"54",
          4272 => x"a5",
          4273 => x"cb",
          4274 => x"8c",
          4275 => x"8d",
          4276 => x"8c",
          4277 => x"ff",
          4278 => x"53",
          4279 => x"51",
          4280 => x"ff",
          4281 => x"de",
          4282 => x"55",
          4283 => x"f7",
          4284 => x"51",
          4285 => x"80",
          4286 => x"93",
          4287 => x"06",
          4288 => x"88",
          4289 => x"74",
          4290 => x"38",
          4291 => x"de",
          4292 => x"39",
          4293 => x"82",
          4294 => x"84",
          4295 => x"54",
          4296 => x"a9",
          4297 => x"ca",
          4298 => x"8c",
          4299 => x"8d",
          4300 => x"8c",
          4301 => x"ff",
          4302 => x"53",
          4303 => x"51",
          4304 => x"81",
          4305 => x"81",
          4306 => x"a8",
          4307 => x"55",
          4308 => x"f6",
          4309 => x"51",
          4310 => x"82",
          4311 => x"82",
          4312 => x"82",
          4313 => x"81",
          4314 => x"05",
          4315 => x"79",
          4316 => x"3f",
          4317 => x"53",
          4318 => x"33",
          4319 => x"ef",
          4320 => x"a9",
          4321 => x"88",
          4322 => x"ff",
          4323 => x"84",
          4324 => x"54",
          4325 => x"f6",
          4326 => x"14",
          4327 => x"8d",
          4328 => x"1a",
          4329 => x"54",
          4330 => x"f6",
          4331 => x"8d",
          4332 => x"73",
          4333 => x"f5",
          4334 => x"e1",
          4335 => x"8d",
          4336 => x"05",
          4337 => x"8d",
          4338 => x"e1",
          4339 => x"82",
          4340 => x"80",
          4341 => x"84",
          4342 => x"8c",
          4343 => x"3d",
          4344 => x"3d",
          4345 => x"05",
          4346 => x"52",
          4347 => x"87",
          4348 => x"c4",
          4349 => x"71",
          4350 => x"0c",
          4351 => x"04",
          4352 => x"02",
          4353 => x"02",
          4354 => x"05",
          4355 => x"83",
          4356 => x"26",
          4357 => x"72",
          4358 => x"c0",
          4359 => x"53",
          4360 => x"74",
          4361 => x"38",
          4362 => x"73",
          4363 => x"c0",
          4364 => x"51",
          4365 => x"85",
          4366 => x"98",
          4367 => x"52",
          4368 => x"82",
          4369 => x"70",
          4370 => x"38",
          4371 => x"8c",
          4372 => x"ec",
          4373 => x"fc",
          4374 => x"52",
          4375 => x"87",
          4376 => x"08",
          4377 => x"2e",
          4378 => x"82",
          4379 => x"34",
          4380 => x"13",
          4381 => x"82",
          4382 => x"86",
          4383 => x"f3",
          4384 => x"62",
          4385 => x"05",
          4386 => x"57",
          4387 => x"83",
          4388 => x"fe",
          4389 => x"8c",
          4390 => x"06",
          4391 => x"71",
          4392 => x"71",
          4393 => x"2b",
          4394 => x"80",
          4395 => x"92",
          4396 => x"c0",
          4397 => x"41",
          4398 => x"5a",
          4399 => x"87",
          4400 => x"0c",
          4401 => x"84",
          4402 => x"08",
          4403 => x"70",
          4404 => x"53",
          4405 => x"2e",
          4406 => x"08",
          4407 => x"70",
          4408 => x"34",
          4409 => x"80",
          4410 => x"53",
          4411 => x"2e",
          4412 => x"53",
          4413 => x"26",
          4414 => x"80",
          4415 => x"87",
          4416 => x"08",
          4417 => x"38",
          4418 => x"8c",
          4419 => x"80",
          4420 => x"78",
          4421 => x"99",
          4422 => x"0c",
          4423 => x"8c",
          4424 => x"08",
          4425 => x"51",
          4426 => x"38",
          4427 => x"8d",
          4428 => x"17",
          4429 => x"81",
          4430 => x"53",
          4431 => x"2e",
          4432 => x"fc",
          4433 => x"52",
          4434 => x"7d",
          4435 => x"ed",
          4436 => x"80",
          4437 => x"71",
          4438 => x"38",
          4439 => x"53",
          4440 => x"dc",
          4441 => x"0d",
          4442 => x"0d",
          4443 => x"02",
          4444 => x"05",
          4445 => x"58",
          4446 => x"80",
          4447 => x"fc",
          4448 => x"8c",
          4449 => x"06",
          4450 => x"71",
          4451 => x"81",
          4452 => x"38",
          4453 => x"2b",
          4454 => x"80",
          4455 => x"92",
          4456 => x"c0",
          4457 => x"40",
          4458 => x"5a",
          4459 => x"c0",
          4460 => x"76",
          4461 => x"76",
          4462 => x"75",
          4463 => x"2a",
          4464 => x"51",
          4465 => x"80",
          4466 => x"7a",
          4467 => x"5c",
          4468 => x"81",
          4469 => x"81",
          4470 => x"06",
          4471 => x"80",
          4472 => x"87",
          4473 => x"08",
          4474 => x"38",
          4475 => x"8c",
          4476 => x"80",
          4477 => x"77",
          4478 => x"99",
          4479 => x"0c",
          4480 => x"8c",
          4481 => x"08",
          4482 => x"51",
          4483 => x"38",
          4484 => x"8d",
          4485 => x"70",
          4486 => x"84",
          4487 => x"5b",
          4488 => x"2e",
          4489 => x"fc",
          4490 => x"52",
          4491 => x"7d",
          4492 => x"f8",
          4493 => x"80",
          4494 => x"71",
          4495 => x"38",
          4496 => x"53",
          4497 => x"dc",
          4498 => x"0d",
          4499 => x"0d",
          4500 => x"05",
          4501 => x"02",
          4502 => x"05",
          4503 => x"54",
          4504 => x"fe",
          4505 => x"dc",
          4506 => x"53",
          4507 => x"80",
          4508 => x"0b",
          4509 => x"8c",
          4510 => x"71",
          4511 => x"dc",
          4512 => x"24",
          4513 => x"84",
          4514 => x"92",
          4515 => x"54",
          4516 => x"8d",
          4517 => x"39",
          4518 => x"80",
          4519 => x"cb",
          4520 => x"70",
          4521 => x"81",
          4522 => x"52",
          4523 => x"8a",
          4524 => x"98",
          4525 => x"71",
          4526 => x"c0",
          4527 => x"52",
          4528 => x"81",
          4529 => x"c0",
          4530 => x"53",
          4531 => x"82",
          4532 => x"71",
          4533 => x"39",
          4534 => x"39",
          4535 => x"77",
          4536 => x"81",
          4537 => x"72",
          4538 => x"84",
          4539 => x"73",
          4540 => x"0c",
          4541 => x"04",
          4542 => x"74",
          4543 => x"71",
          4544 => x"2b",
          4545 => x"dc",
          4546 => x"84",
          4547 => x"fd",
          4548 => x"83",
          4549 => x"12",
          4550 => x"2b",
          4551 => x"07",
          4552 => x"70",
          4553 => x"2b",
          4554 => x"07",
          4555 => x"0c",
          4556 => x"56",
          4557 => x"3d",
          4558 => x"3d",
          4559 => x"84",
          4560 => x"22",
          4561 => x"72",
          4562 => x"54",
          4563 => x"2a",
          4564 => x"34",
          4565 => x"04",
          4566 => x"73",
          4567 => x"70",
          4568 => x"05",
          4569 => x"88",
          4570 => x"72",
          4571 => x"54",
          4572 => x"2a",
          4573 => x"70",
          4574 => x"34",
          4575 => x"51",
          4576 => x"83",
          4577 => x"fe",
          4578 => x"75",
          4579 => x"51",
          4580 => x"92",
          4581 => x"81",
          4582 => x"73",
          4583 => x"55",
          4584 => x"51",
          4585 => x"3d",
          4586 => x"3d",
          4587 => x"76",
          4588 => x"72",
          4589 => x"05",
          4590 => x"11",
          4591 => x"38",
          4592 => x"04",
          4593 => x"78",
          4594 => x"56",
          4595 => x"81",
          4596 => x"74",
          4597 => x"56",
          4598 => x"31",
          4599 => x"52",
          4600 => x"80",
          4601 => x"71",
          4602 => x"38",
          4603 => x"dc",
          4604 => x"0d",
          4605 => x"0d",
          4606 => x"51",
          4607 => x"73",
          4608 => x"81",
          4609 => x"33",
          4610 => x"38",
          4611 => x"8c",
          4612 => x"3d",
          4613 => x"0b",
          4614 => x"0c",
          4615 => x"82",
          4616 => x"04",
          4617 => x"7b",
          4618 => x"83",
          4619 => x"5a",
          4620 => x"80",
          4621 => x"54",
          4622 => x"53",
          4623 => x"53",
          4624 => x"52",
          4625 => x"3f",
          4626 => x"08",
          4627 => x"81",
          4628 => x"82",
          4629 => x"83",
          4630 => x"16",
          4631 => x"18",
          4632 => x"18",
          4633 => x"58",
          4634 => x"9f",
          4635 => x"33",
          4636 => x"2e",
          4637 => x"93",
          4638 => x"76",
          4639 => x"52",
          4640 => x"51",
          4641 => x"83",
          4642 => x"79",
          4643 => x"0c",
          4644 => x"04",
          4645 => x"78",
          4646 => x"80",
          4647 => x"17",
          4648 => x"38",
          4649 => x"fc",
          4650 => x"dc",
          4651 => x"8c",
          4652 => x"38",
          4653 => x"53",
          4654 => x"81",
          4655 => x"f7",
          4656 => x"8c",
          4657 => x"2e",
          4658 => x"55",
          4659 => x"b0",
          4660 => x"82",
          4661 => x"88",
          4662 => x"f8",
          4663 => x"70",
          4664 => x"c0",
          4665 => x"dc",
          4666 => x"8c",
          4667 => x"91",
          4668 => x"55",
          4669 => x"09",
          4670 => x"f0",
          4671 => x"33",
          4672 => x"2e",
          4673 => x"80",
          4674 => x"80",
          4675 => x"dc",
          4676 => x"17",
          4677 => x"fd",
          4678 => x"d4",
          4679 => x"b2",
          4680 => x"96",
          4681 => x"85",
          4682 => x"75",
          4683 => x"3f",
          4684 => x"e4",
          4685 => x"98",
          4686 => x"9c",
          4687 => x"08",
          4688 => x"17",
          4689 => x"3f",
          4690 => x"52",
          4691 => x"51",
          4692 => x"a0",
          4693 => x"05",
          4694 => x"0c",
          4695 => x"75",
          4696 => x"33",
          4697 => x"3f",
          4698 => x"34",
          4699 => x"52",
          4700 => x"51",
          4701 => x"82",
          4702 => x"80",
          4703 => x"81",
          4704 => x"8c",
          4705 => x"3d",
          4706 => x"3d",
          4707 => x"1a",
          4708 => x"fe",
          4709 => x"54",
          4710 => x"73",
          4711 => x"8a",
          4712 => x"71",
          4713 => x"08",
          4714 => x"75",
          4715 => x"0c",
          4716 => x"04",
          4717 => x"7a",
          4718 => x"56",
          4719 => x"77",
          4720 => x"38",
          4721 => x"08",
          4722 => x"38",
          4723 => x"54",
          4724 => x"2e",
          4725 => x"72",
          4726 => x"38",
          4727 => x"8d",
          4728 => x"39",
          4729 => x"81",
          4730 => x"b6",
          4731 => x"2a",
          4732 => x"2a",
          4733 => x"05",
          4734 => x"55",
          4735 => x"82",
          4736 => x"81",
          4737 => x"83",
          4738 => x"b4",
          4739 => x"17",
          4740 => x"a4",
          4741 => x"55",
          4742 => x"57",
          4743 => x"3f",
          4744 => x"08",
          4745 => x"74",
          4746 => x"14",
          4747 => x"70",
          4748 => x"07",
          4749 => x"71",
          4750 => x"52",
          4751 => x"72",
          4752 => x"75",
          4753 => x"58",
          4754 => x"76",
          4755 => x"15",
          4756 => x"73",
          4757 => x"3f",
          4758 => x"08",
          4759 => x"76",
          4760 => x"06",
          4761 => x"05",
          4762 => x"3f",
          4763 => x"08",
          4764 => x"06",
          4765 => x"76",
          4766 => x"15",
          4767 => x"73",
          4768 => x"3f",
          4769 => x"08",
          4770 => x"82",
          4771 => x"06",
          4772 => x"05",
          4773 => x"3f",
          4774 => x"08",
          4775 => x"58",
          4776 => x"58",
          4777 => x"dc",
          4778 => x"0d",
          4779 => x"0d",
          4780 => x"5a",
          4781 => x"59",
          4782 => x"82",
          4783 => x"98",
          4784 => x"82",
          4785 => x"33",
          4786 => x"2e",
          4787 => x"72",
          4788 => x"38",
          4789 => x"8d",
          4790 => x"39",
          4791 => x"81",
          4792 => x"f7",
          4793 => x"2a",
          4794 => x"2a",
          4795 => x"05",
          4796 => x"55",
          4797 => x"82",
          4798 => x"59",
          4799 => x"08",
          4800 => x"74",
          4801 => x"16",
          4802 => x"16",
          4803 => x"59",
          4804 => x"53",
          4805 => x"8f",
          4806 => x"2b",
          4807 => x"74",
          4808 => x"71",
          4809 => x"72",
          4810 => x"0b",
          4811 => x"74",
          4812 => x"17",
          4813 => x"75",
          4814 => x"3f",
          4815 => x"08",
          4816 => x"dc",
          4817 => x"38",
          4818 => x"06",
          4819 => x"78",
          4820 => x"54",
          4821 => x"77",
          4822 => x"33",
          4823 => x"71",
          4824 => x"51",
          4825 => x"34",
          4826 => x"76",
          4827 => x"17",
          4828 => x"75",
          4829 => x"3f",
          4830 => x"08",
          4831 => x"dc",
          4832 => x"38",
          4833 => x"ff",
          4834 => x"10",
          4835 => x"76",
          4836 => x"51",
          4837 => x"be",
          4838 => x"2a",
          4839 => x"05",
          4840 => x"f9",
          4841 => x"8c",
          4842 => x"82",
          4843 => x"ab",
          4844 => x"0a",
          4845 => x"2b",
          4846 => x"70",
          4847 => x"70",
          4848 => x"54",
          4849 => x"82",
          4850 => x"8f",
          4851 => x"07",
          4852 => x"f7",
          4853 => x"0b",
          4854 => x"78",
          4855 => x"0c",
          4856 => x"04",
          4857 => x"7a",
          4858 => x"08",
          4859 => x"59",
          4860 => x"a4",
          4861 => x"17",
          4862 => x"38",
          4863 => x"aa",
          4864 => x"73",
          4865 => x"fd",
          4866 => x"8c",
          4867 => x"82",
          4868 => x"80",
          4869 => x"39",
          4870 => x"eb",
          4871 => x"80",
          4872 => x"8c",
          4873 => x"80",
          4874 => x"52",
          4875 => x"84",
          4876 => x"dc",
          4877 => x"8c",
          4878 => x"2e",
          4879 => x"82",
          4880 => x"81",
          4881 => x"82",
          4882 => x"ff",
          4883 => x"80",
          4884 => x"75",
          4885 => x"3f",
          4886 => x"08",
          4887 => x"16",
          4888 => x"90",
          4889 => x"55",
          4890 => x"27",
          4891 => x"15",
          4892 => x"84",
          4893 => x"07",
          4894 => x"17",
          4895 => x"76",
          4896 => x"a6",
          4897 => x"73",
          4898 => x"0c",
          4899 => x"04",
          4900 => x"7c",
          4901 => x"59",
          4902 => x"95",
          4903 => x"08",
          4904 => x"2e",
          4905 => x"17",
          4906 => x"b2",
          4907 => x"ae",
          4908 => x"7a",
          4909 => x"3f",
          4910 => x"82",
          4911 => x"27",
          4912 => x"82",
          4913 => x"55",
          4914 => x"08",
          4915 => x"d2",
          4916 => x"08",
          4917 => x"08",
          4918 => x"38",
          4919 => x"17",
          4920 => x"54",
          4921 => x"82",
          4922 => x"7a",
          4923 => x"06",
          4924 => x"81",
          4925 => x"17",
          4926 => x"83",
          4927 => x"75",
          4928 => x"f9",
          4929 => x"59",
          4930 => x"08",
          4931 => x"81",
          4932 => x"82",
          4933 => x"59",
          4934 => x"08",
          4935 => x"70",
          4936 => x"25",
          4937 => x"82",
          4938 => x"54",
          4939 => x"55",
          4940 => x"38",
          4941 => x"08",
          4942 => x"38",
          4943 => x"54",
          4944 => x"90",
          4945 => x"18",
          4946 => x"38",
          4947 => x"39",
          4948 => x"38",
          4949 => x"16",
          4950 => x"08",
          4951 => x"38",
          4952 => x"78",
          4953 => x"38",
          4954 => x"51",
          4955 => x"82",
          4956 => x"80",
          4957 => x"80",
          4958 => x"dc",
          4959 => x"09",
          4960 => x"38",
          4961 => x"08",
          4962 => x"dc",
          4963 => x"30",
          4964 => x"80",
          4965 => x"07",
          4966 => x"55",
          4967 => x"38",
          4968 => x"09",
          4969 => x"ae",
          4970 => x"80",
          4971 => x"53",
          4972 => x"51",
          4973 => x"82",
          4974 => x"82",
          4975 => x"30",
          4976 => x"dc",
          4977 => x"25",
          4978 => x"79",
          4979 => x"38",
          4980 => x"8f",
          4981 => x"79",
          4982 => x"f9",
          4983 => x"8c",
          4984 => x"74",
          4985 => x"8c",
          4986 => x"17",
          4987 => x"90",
          4988 => x"54",
          4989 => x"86",
          4990 => x"90",
          4991 => x"17",
          4992 => x"54",
          4993 => x"34",
          4994 => x"56",
          4995 => x"90",
          4996 => x"80",
          4997 => x"82",
          4998 => x"55",
          4999 => x"56",
          5000 => x"82",
          5001 => x"8c",
          5002 => x"f8",
          5003 => x"70",
          5004 => x"f0",
          5005 => x"dc",
          5006 => x"56",
          5007 => x"08",
          5008 => x"7b",
          5009 => x"f6",
          5010 => x"8c",
          5011 => x"8c",
          5012 => x"17",
          5013 => x"80",
          5014 => x"b4",
          5015 => x"57",
          5016 => x"77",
          5017 => x"81",
          5018 => x"15",
          5019 => x"78",
          5020 => x"81",
          5021 => x"53",
          5022 => x"15",
          5023 => x"e9",
          5024 => x"dc",
          5025 => x"df",
          5026 => x"22",
          5027 => x"30",
          5028 => x"70",
          5029 => x"51",
          5030 => x"82",
          5031 => x"8a",
          5032 => x"f8",
          5033 => x"7c",
          5034 => x"56",
          5035 => x"80",
          5036 => x"f1",
          5037 => x"06",
          5038 => x"e9",
          5039 => x"18",
          5040 => x"08",
          5041 => x"38",
          5042 => x"82",
          5043 => x"38",
          5044 => x"54",
          5045 => x"74",
          5046 => x"82",
          5047 => x"22",
          5048 => x"79",
          5049 => x"38",
          5050 => x"98",
          5051 => x"cd",
          5052 => x"22",
          5053 => x"54",
          5054 => x"26",
          5055 => x"52",
          5056 => x"b0",
          5057 => x"dc",
          5058 => x"8c",
          5059 => x"2e",
          5060 => x"0b",
          5061 => x"08",
          5062 => x"98",
          5063 => x"8c",
          5064 => x"85",
          5065 => x"bd",
          5066 => x"31",
          5067 => x"73",
          5068 => x"f4",
          5069 => x"8c",
          5070 => x"18",
          5071 => x"18",
          5072 => x"08",
          5073 => x"72",
          5074 => x"38",
          5075 => x"58",
          5076 => x"89",
          5077 => x"18",
          5078 => x"ff",
          5079 => x"05",
          5080 => x"80",
          5081 => x"8c",
          5082 => x"3d",
          5083 => x"3d",
          5084 => x"08",
          5085 => x"a0",
          5086 => x"54",
          5087 => x"77",
          5088 => x"80",
          5089 => x"0c",
          5090 => x"53",
          5091 => x"80",
          5092 => x"38",
          5093 => x"06",
          5094 => x"b5",
          5095 => x"98",
          5096 => x"14",
          5097 => x"92",
          5098 => x"2a",
          5099 => x"56",
          5100 => x"26",
          5101 => x"80",
          5102 => x"16",
          5103 => x"77",
          5104 => x"53",
          5105 => x"38",
          5106 => x"51",
          5107 => x"82",
          5108 => x"53",
          5109 => x"0b",
          5110 => x"08",
          5111 => x"38",
          5112 => x"8c",
          5113 => x"2e",
          5114 => x"98",
          5115 => x"8c",
          5116 => x"80",
          5117 => x"8a",
          5118 => x"15",
          5119 => x"80",
          5120 => x"14",
          5121 => x"51",
          5122 => x"82",
          5123 => x"53",
          5124 => x"8c",
          5125 => x"2e",
          5126 => x"82",
          5127 => x"dc",
          5128 => x"ba",
          5129 => x"82",
          5130 => x"ff",
          5131 => x"82",
          5132 => x"52",
          5133 => x"f3",
          5134 => x"dc",
          5135 => x"72",
          5136 => x"72",
          5137 => x"f2",
          5138 => x"8c",
          5139 => x"15",
          5140 => x"15",
          5141 => x"b4",
          5142 => x"0c",
          5143 => x"82",
          5144 => x"8a",
          5145 => x"f7",
          5146 => x"7d",
          5147 => x"5b",
          5148 => x"76",
          5149 => x"3f",
          5150 => x"08",
          5151 => x"dc",
          5152 => x"38",
          5153 => x"08",
          5154 => x"08",
          5155 => x"f0",
          5156 => x"8c",
          5157 => x"82",
          5158 => x"80",
          5159 => x"8c",
          5160 => x"18",
          5161 => x"51",
          5162 => x"81",
          5163 => x"81",
          5164 => x"81",
          5165 => x"dc",
          5166 => x"83",
          5167 => x"77",
          5168 => x"72",
          5169 => x"38",
          5170 => x"75",
          5171 => x"81",
          5172 => x"a5",
          5173 => x"dc",
          5174 => x"52",
          5175 => x"8e",
          5176 => x"dc",
          5177 => x"8c",
          5178 => x"2e",
          5179 => x"73",
          5180 => x"81",
          5181 => x"87",
          5182 => x"8c",
          5183 => x"3d",
          5184 => x"3d",
          5185 => x"11",
          5186 => x"ec",
          5187 => x"dc",
          5188 => x"ff",
          5189 => x"33",
          5190 => x"71",
          5191 => x"81",
          5192 => x"94",
          5193 => x"d0",
          5194 => x"dc",
          5195 => x"73",
          5196 => x"82",
          5197 => x"85",
          5198 => x"fc",
          5199 => x"79",
          5200 => x"ff",
          5201 => x"12",
          5202 => x"eb",
          5203 => x"70",
          5204 => x"72",
          5205 => x"81",
          5206 => x"73",
          5207 => x"94",
          5208 => x"d6",
          5209 => x"0d",
          5210 => x"0d",
          5211 => x"55",
          5212 => x"5a",
          5213 => x"08",
          5214 => x"8a",
          5215 => x"08",
          5216 => x"ee",
          5217 => x"8c",
          5218 => x"82",
          5219 => x"80",
          5220 => x"15",
          5221 => x"55",
          5222 => x"38",
          5223 => x"e6",
          5224 => x"33",
          5225 => x"70",
          5226 => x"58",
          5227 => x"86",
          5228 => x"8c",
          5229 => x"73",
          5230 => x"83",
          5231 => x"73",
          5232 => x"38",
          5233 => x"06",
          5234 => x"80",
          5235 => x"75",
          5236 => x"38",
          5237 => x"08",
          5238 => x"54",
          5239 => x"2e",
          5240 => x"83",
          5241 => x"73",
          5242 => x"38",
          5243 => x"51",
          5244 => x"82",
          5245 => x"58",
          5246 => x"08",
          5247 => x"15",
          5248 => x"38",
          5249 => x"0b",
          5250 => x"77",
          5251 => x"0c",
          5252 => x"04",
          5253 => x"77",
          5254 => x"54",
          5255 => x"51",
          5256 => x"82",
          5257 => x"55",
          5258 => x"08",
          5259 => x"14",
          5260 => x"51",
          5261 => x"82",
          5262 => x"55",
          5263 => x"08",
          5264 => x"53",
          5265 => x"08",
          5266 => x"08",
          5267 => x"3f",
          5268 => x"14",
          5269 => x"08",
          5270 => x"3f",
          5271 => x"17",
          5272 => x"8c",
          5273 => x"3d",
          5274 => x"3d",
          5275 => x"08",
          5276 => x"54",
          5277 => x"53",
          5278 => x"82",
          5279 => x"8d",
          5280 => x"08",
          5281 => x"34",
          5282 => x"15",
          5283 => x"0d",
          5284 => x"0d",
          5285 => x"57",
          5286 => x"17",
          5287 => x"08",
          5288 => x"82",
          5289 => x"89",
          5290 => x"55",
          5291 => x"14",
          5292 => x"16",
          5293 => x"71",
          5294 => x"38",
          5295 => x"09",
          5296 => x"38",
          5297 => x"73",
          5298 => x"81",
          5299 => x"ae",
          5300 => x"05",
          5301 => x"15",
          5302 => x"70",
          5303 => x"34",
          5304 => x"8a",
          5305 => x"38",
          5306 => x"05",
          5307 => x"81",
          5308 => x"17",
          5309 => x"12",
          5310 => x"34",
          5311 => x"9c",
          5312 => x"e8",
          5313 => x"8c",
          5314 => x"0c",
          5315 => x"e7",
          5316 => x"8c",
          5317 => x"17",
          5318 => x"51",
          5319 => x"82",
          5320 => x"84",
          5321 => x"3d",
          5322 => x"3d",
          5323 => x"08",
          5324 => x"61",
          5325 => x"55",
          5326 => x"2e",
          5327 => x"55",
          5328 => x"2e",
          5329 => x"80",
          5330 => x"94",
          5331 => x"1c",
          5332 => x"81",
          5333 => x"61",
          5334 => x"56",
          5335 => x"2e",
          5336 => x"83",
          5337 => x"73",
          5338 => x"70",
          5339 => x"25",
          5340 => x"51",
          5341 => x"38",
          5342 => x"0c",
          5343 => x"51",
          5344 => x"26",
          5345 => x"80",
          5346 => x"34",
          5347 => x"51",
          5348 => x"82",
          5349 => x"55",
          5350 => x"91",
          5351 => x"1d",
          5352 => x"8b",
          5353 => x"79",
          5354 => x"3f",
          5355 => x"57",
          5356 => x"55",
          5357 => x"2e",
          5358 => x"80",
          5359 => x"18",
          5360 => x"1a",
          5361 => x"70",
          5362 => x"2a",
          5363 => x"07",
          5364 => x"5a",
          5365 => x"8c",
          5366 => x"54",
          5367 => x"81",
          5368 => x"39",
          5369 => x"70",
          5370 => x"2a",
          5371 => x"75",
          5372 => x"8c",
          5373 => x"2e",
          5374 => x"a0",
          5375 => x"38",
          5376 => x"0c",
          5377 => x"76",
          5378 => x"38",
          5379 => x"b8",
          5380 => x"70",
          5381 => x"5a",
          5382 => x"76",
          5383 => x"38",
          5384 => x"70",
          5385 => x"dc",
          5386 => x"72",
          5387 => x"80",
          5388 => x"51",
          5389 => x"73",
          5390 => x"38",
          5391 => x"18",
          5392 => x"1a",
          5393 => x"55",
          5394 => x"2e",
          5395 => x"83",
          5396 => x"73",
          5397 => x"70",
          5398 => x"25",
          5399 => x"51",
          5400 => x"38",
          5401 => x"75",
          5402 => x"81",
          5403 => x"81",
          5404 => x"27",
          5405 => x"73",
          5406 => x"38",
          5407 => x"70",
          5408 => x"32",
          5409 => x"80",
          5410 => x"2a",
          5411 => x"56",
          5412 => x"81",
          5413 => x"57",
          5414 => x"f5",
          5415 => x"2b",
          5416 => x"25",
          5417 => x"80",
          5418 => x"fa",
          5419 => x"57",
          5420 => x"e6",
          5421 => x"8c",
          5422 => x"2e",
          5423 => x"18",
          5424 => x"1a",
          5425 => x"56",
          5426 => x"3f",
          5427 => x"08",
          5428 => x"e8",
          5429 => x"54",
          5430 => x"80",
          5431 => x"17",
          5432 => x"34",
          5433 => x"11",
          5434 => x"74",
          5435 => x"75",
          5436 => x"8c",
          5437 => x"3f",
          5438 => x"08",
          5439 => x"9f",
          5440 => x"99",
          5441 => x"e0",
          5442 => x"ff",
          5443 => x"79",
          5444 => x"74",
          5445 => x"57",
          5446 => x"77",
          5447 => x"76",
          5448 => x"38",
          5449 => x"73",
          5450 => x"09",
          5451 => x"38",
          5452 => x"84",
          5453 => x"27",
          5454 => x"39",
          5455 => x"f2",
          5456 => x"80",
          5457 => x"54",
          5458 => x"34",
          5459 => x"58",
          5460 => x"f2",
          5461 => x"8c",
          5462 => x"82",
          5463 => x"80",
          5464 => x"1b",
          5465 => x"51",
          5466 => x"82",
          5467 => x"56",
          5468 => x"08",
          5469 => x"9c",
          5470 => x"33",
          5471 => x"80",
          5472 => x"38",
          5473 => x"bf",
          5474 => x"86",
          5475 => x"15",
          5476 => x"2a",
          5477 => x"51",
          5478 => x"92",
          5479 => x"79",
          5480 => x"e4",
          5481 => x"8c",
          5482 => x"2e",
          5483 => x"52",
          5484 => x"ba",
          5485 => x"39",
          5486 => x"33",
          5487 => x"80",
          5488 => x"74",
          5489 => x"81",
          5490 => x"38",
          5491 => x"70",
          5492 => x"82",
          5493 => x"54",
          5494 => x"96",
          5495 => x"06",
          5496 => x"2e",
          5497 => x"ff",
          5498 => x"1c",
          5499 => x"80",
          5500 => x"81",
          5501 => x"ba",
          5502 => x"b6",
          5503 => x"2a",
          5504 => x"51",
          5505 => x"38",
          5506 => x"70",
          5507 => x"81",
          5508 => x"55",
          5509 => x"e1",
          5510 => x"08",
          5511 => x"1d",
          5512 => x"7c",
          5513 => x"3f",
          5514 => x"08",
          5515 => x"fa",
          5516 => x"82",
          5517 => x"8f",
          5518 => x"f6",
          5519 => x"5b",
          5520 => x"70",
          5521 => x"59",
          5522 => x"73",
          5523 => x"c6",
          5524 => x"81",
          5525 => x"70",
          5526 => x"52",
          5527 => x"8d",
          5528 => x"38",
          5529 => x"09",
          5530 => x"a5",
          5531 => x"d0",
          5532 => x"ff",
          5533 => x"53",
          5534 => x"91",
          5535 => x"73",
          5536 => x"d0",
          5537 => x"71",
          5538 => x"f7",
          5539 => x"81",
          5540 => x"55",
          5541 => x"55",
          5542 => x"81",
          5543 => x"74",
          5544 => x"56",
          5545 => x"12",
          5546 => x"70",
          5547 => x"38",
          5548 => x"81",
          5549 => x"51",
          5550 => x"51",
          5551 => x"89",
          5552 => x"70",
          5553 => x"53",
          5554 => x"70",
          5555 => x"51",
          5556 => x"09",
          5557 => x"38",
          5558 => x"38",
          5559 => x"77",
          5560 => x"70",
          5561 => x"2a",
          5562 => x"07",
          5563 => x"51",
          5564 => x"8f",
          5565 => x"84",
          5566 => x"83",
          5567 => x"94",
          5568 => x"74",
          5569 => x"38",
          5570 => x"0c",
          5571 => x"86",
          5572 => x"a0",
          5573 => x"82",
          5574 => x"8c",
          5575 => x"fa",
          5576 => x"56",
          5577 => x"17",
          5578 => x"b0",
          5579 => x"52",
          5580 => x"e0",
          5581 => x"82",
          5582 => x"81",
          5583 => x"b2",
          5584 => x"b4",
          5585 => x"dc",
          5586 => x"ff",
          5587 => x"55",
          5588 => x"d5",
          5589 => x"06",
          5590 => x"80",
          5591 => x"33",
          5592 => x"81",
          5593 => x"81",
          5594 => x"81",
          5595 => x"eb",
          5596 => x"70",
          5597 => x"07",
          5598 => x"73",
          5599 => x"81",
          5600 => x"81",
          5601 => x"83",
          5602 => x"9c",
          5603 => x"16",
          5604 => x"3f",
          5605 => x"08",
          5606 => x"dc",
          5607 => x"9d",
          5608 => x"81",
          5609 => x"81",
          5610 => x"e0",
          5611 => x"8c",
          5612 => x"82",
          5613 => x"80",
          5614 => x"82",
          5615 => x"8c",
          5616 => x"3d",
          5617 => x"3d",
          5618 => x"84",
          5619 => x"05",
          5620 => x"80",
          5621 => x"51",
          5622 => x"82",
          5623 => x"58",
          5624 => x"0b",
          5625 => x"08",
          5626 => x"38",
          5627 => x"08",
          5628 => x"8d",
          5629 => x"08",
          5630 => x"56",
          5631 => x"86",
          5632 => x"75",
          5633 => x"fe",
          5634 => x"54",
          5635 => x"2e",
          5636 => x"14",
          5637 => x"ca",
          5638 => x"dc",
          5639 => x"06",
          5640 => x"54",
          5641 => x"38",
          5642 => x"86",
          5643 => x"82",
          5644 => x"06",
          5645 => x"56",
          5646 => x"38",
          5647 => x"80",
          5648 => x"81",
          5649 => x"52",
          5650 => x"51",
          5651 => x"82",
          5652 => x"81",
          5653 => x"81",
          5654 => x"83",
          5655 => x"87",
          5656 => x"2e",
          5657 => x"82",
          5658 => x"06",
          5659 => x"56",
          5660 => x"38",
          5661 => x"74",
          5662 => x"a3",
          5663 => x"dc",
          5664 => x"06",
          5665 => x"2e",
          5666 => x"80",
          5667 => x"3d",
          5668 => x"83",
          5669 => x"15",
          5670 => x"53",
          5671 => x"8d",
          5672 => x"15",
          5673 => x"3f",
          5674 => x"08",
          5675 => x"70",
          5676 => x"0c",
          5677 => x"16",
          5678 => x"80",
          5679 => x"80",
          5680 => x"54",
          5681 => x"84",
          5682 => x"5b",
          5683 => x"80",
          5684 => x"7a",
          5685 => x"fc",
          5686 => x"8c",
          5687 => x"ff",
          5688 => x"77",
          5689 => x"81",
          5690 => x"76",
          5691 => x"81",
          5692 => x"2e",
          5693 => x"8d",
          5694 => x"26",
          5695 => x"bf",
          5696 => x"f4",
          5697 => x"dc",
          5698 => x"ff",
          5699 => x"84",
          5700 => x"81",
          5701 => x"38",
          5702 => x"51",
          5703 => x"82",
          5704 => x"83",
          5705 => x"58",
          5706 => x"80",
          5707 => x"db",
          5708 => x"8c",
          5709 => x"77",
          5710 => x"80",
          5711 => x"82",
          5712 => x"c4",
          5713 => x"11",
          5714 => x"06",
          5715 => x"8d",
          5716 => x"26",
          5717 => x"74",
          5718 => x"78",
          5719 => x"c1",
          5720 => x"59",
          5721 => x"15",
          5722 => x"2e",
          5723 => x"13",
          5724 => x"72",
          5725 => x"38",
          5726 => x"eb",
          5727 => x"14",
          5728 => x"3f",
          5729 => x"08",
          5730 => x"dc",
          5731 => x"23",
          5732 => x"57",
          5733 => x"83",
          5734 => x"c7",
          5735 => x"d8",
          5736 => x"dc",
          5737 => x"ff",
          5738 => x"8d",
          5739 => x"14",
          5740 => x"3f",
          5741 => x"08",
          5742 => x"14",
          5743 => x"3f",
          5744 => x"08",
          5745 => x"06",
          5746 => x"72",
          5747 => x"97",
          5748 => x"22",
          5749 => x"84",
          5750 => x"5a",
          5751 => x"83",
          5752 => x"14",
          5753 => x"79",
          5754 => x"96",
          5755 => x"8c",
          5756 => x"82",
          5757 => x"80",
          5758 => x"38",
          5759 => x"08",
          5760 => x"ff",
          5761 => x"38",
          5762 => x"83",
          5763 => x"83",
          5764 => x"74",
          5765 => x"85",
          5766 => x"89",
          5767 => x"76",
          5768 => x"c3",
          5769 => x"70",
          5770 => x"7b",
          5771 => x"73",
          5772 => x"17",
          5773 => x"ac",
          5774 => x"55",
          5775 => x"09",
          5776 => x"38",
          5777 => x"51",
          5778 => x"82",
          5779 => x"83",
          5780 => x"53",
          5781 => x"82",
          5782 => x"82",
          5783 => x"e0",
          5784 => x"ab",
          5785 => x"dc",
          5786 => x"0c",
          5787 => x"53",
          5788 => x"56",
          5789 => x"81",
          5790 => x"13",
          5791 => x"74",
          5792 => x"82",
          5793 => x"74",
          5794 => x"81",
          5795 => x"06",
          5796 => x"83",
          5797 => x"2a",
          5798 => x"72",
          5799 => x"26",
          5800 => x"ff",
          5801 => x"0c",
          5802 => x"15",
          5803 => x"0b",
          5804 => x"76",
          5805 => x"81",
          5806 => x"38",
          5807 => x"51",
          5808 => x"82",
          5809 => x"83",
          5810 => x"53",
          5811 => x"09",
          5812 => x"f9",
          5813 => x"52",
          5814 => x"b8",
          5815 => x"dc",
          5816 => x"38",
          5817 => x"08",
          5818 => x"84",
          5819 => x"d8",
          5820 => x"8c",
          5821 => x"ff",
          5822 => x"72",
          5823 => x"2e",
          5824 => x"80",
          5825 => x"14",
          5826 => x"3f",
          5827 => x"08",
          5828 => x"a4",
          5829 => x"81",
          5830 => x"84",
          5831 => x"d7",
          5832 => x"8c",
          5833 => x"8a",
          5834 => x"2e",
          5835 => x"9d",
          5836 => x"14",
          5837 => x"3f",
          5838 => x"08",
          5839 => x"84",
          5840 => x"d7",
          5841 => x"8c",
          5842 => x"15",
          5843 => x"34",
          5844 => x"22",
          5845 => x"72",
          5846 => x"23",
          5847 => x"23",
          5848 => x"15",
          5849 => x"75",
          5850 => x"0c",
          5851 => x"04",
          5852 => x"77",
          5853 => x"73",
          5854 => x"38",
          5855 => x"72",
          5856 => x"38",
          5857 => x"71",
          5858 => x"38",
          5859 => x"84",
          5860 => x"52",
          5861 => x"09",
          5862 => x"38",
          5863 => x"51",
          5864 => x"82",
          5865 => x"81",
          5866 => x"88",
          5867 => x"08",
          5868 => x"39",
          5869 => x"73",
          5870 => x"74",
          5871 => x"0c",
          5872 => x"04",
          5873 => x"02",
          5874 => x"7a",
          5875 => x"fc",
          5876 => x"f4",
          5877 => x"54",
          5878 => x"8c",
          5879 => x"bc",
          5880 => x"dc",
          5881 => x"82",
          5882 => x"70",
          5883 => x"73",
          5884 => x"38",
          5885 => x"78",
          5886 => x"2e",
          5887 => x"74",
          5888 => x"0c",
          5889 => x"80",
          5890 => x"80",
          5891 => x"70",
          5892 => x"51",
          5893 => x"82",
          5894 => x"54",
          5895 => x"dc",
          5896 => x"0d",
          5897 => x"0d",
          5898 => x"05",
          5899 => x"33",
          5900 => x"54",
          5901 => x"84",
          5902 => x"bf",
          5903 => x"98",
          5904 => x"53",
          5905 => x"05",
          5906 => x"fa",
          5907 => x"dc",
          5908 => x"8c",
          5909 => x"a4",
          5910 => x"68",
          5911 => x"70",
          5912 => x"c6",
          5913 => x"dc",
          5914 => x"8c",
          5915 => x"38",
          5916 => x"05",
          5917 => x"2b",
          5918 => x"80",
          5919 => x"86",
          5920 => x"06",
          5921 => x"2e",
          5922 => x"74",
          5923 => x"38",
          5924 => x"09",
          5925 => x"38",
          5926 => x"f8",
          5927 => x"dc",
          5928 => x"39",
          5929 => x"33",
          5930 => x"73",
          5931 => x"77",
          5932 => x"81",
          5933 => x"73",
          5934 => x"38",
          5935 => x"bc",
          5936 => x"07",
          5937 => x"b4",
          5938 => x"2a",
          5939 => x"51",
          5940 => x"2e",
          5941 => x"62",
          5942 => x"e8",
          5943 => x"8c",
          5944 => x"82",
          5945 => x"52",
          5946 => x"51",
          5947 => x"62",
          5948 => x"8b",
          5949 => x"53",
          5950 => x"51",
          5951 => x"80",
          5952 => x"05",
          5953 => x"3f",
          5954 => x"0b",
          5955 => x"75",
          5956 => x"f1",
          5957 => x"11",
          5958 => x"80",
          5959 => x"97",
          5960 => x"51",
          5961 => x"82",
          5962 => x"55",
          5963 => x"08",
          5964 => x"b7",
          5965 => x"c4",
          5966 => x"05",
          5967 => x"2a",
          5968 => x"51",
          5969 => x"80",
          5970 => x"84",
          5971 => x"39",
          5972 => x"70",
          5973 => x"54",
          5974 => x"a9",
          5975 => x"06",
          5976 => x"2e",
          5977 => x"55",
          5978 => x"73",
          5979 => x"d6",
          5980 => x"8c",
          5981 => x"ff",
          5982 => x"0c",
          5983 => x"8c",
          5984 => x"f8",
          5985 => x"2a",
          5986 => x"51",
          5987 => x"2e",
          5988 => x"80",
          5989 => x"7a",
          5990 => x"a0",
          5991 => x"a4",
          5992 => x"53",
          5993 => x"e6",
          5994 => x"8c",
          5995 => x"8c",
          5996 => x"1b",
          5997 => x"05",
          5998 => x"d3",
          5999 => x"dc",
          6000 => x"dc",
          6001 => x"0c",
          6002 => x"56",
          6003 => x"84",
          6004 => x"90",
          6005 => x"0b",
          6006 => x"80",
          6007 => x"0c",
          6008 => x"1a",
          6009 => x"2a",
          6010 => x"51",
          6011 => x"2e",
          6012 => x"82",
          6013 => x"80",
          6014 => x"38",
          6015 => x"08",
          6016 => x"8a",
          6017 => x"89",
          6018 => x"59",
          6019 => x"76",
          6020 => x"d7",
          6021 => x"8c",
          6022 => x"82",
          6023 => x"81",
          6024 => x"82",
          6025 => x"dc",
          6026 => x"09",
          6027 => x"38",
          6028 => x"78",
          6029 => x"30",
          6030 => x"80",
          6031 => x"77",
          6032 => x"38",
          6033 => x"06",
          6034 => x"c3",
          6035 => x"1a",
          6036 => x"38",
          6037 => x"06",
          6038 => x"2e",
          6039 => x"52",
          6040 => x"a6",
          6041 => x"dc",
          6042 => x"82",
          6043 => x"75",
          6044 => x"8c",
          6045 => x"9c",
          6046 => x"39",
          6047 => x"74",
          6048 => x"8c",
          6049 => x"3d",
          6050 => x"3d",
          6051 => x"65",
          6052 => x"5d",
          6053 => x"0c",
          6054 => x"05",
          6055 => x"f9",
          6056 => x"8c",
          6057 => x"82",
          6058 => x"8a",
          6059 => x"33",
          6060 => x"2e",
          6061 => x"56",
          6062 => x"90",
          6063 => x"06",
          6064 => x"74",
          6065 => x"b6",
          6066 => x"82",
          6067 => x"34",
          6068 => x"aa",
          6069 => x"91",
          6070 => x"56",
          6071 => x"8c",
          6072 => x"1a",
          6073 => x"74",
          6074 => x"38",
          6075 => x"80",
          6076 => x"38",
          6077 => x"70",
          6078 => x"56",
          6079 => x"b2",
          6080 => x"11",
          6081 => x"77",
          6082 => x"5b",
          6083 => x"38",
          6084 => x"88",
          6085 => x"8f",
          6086 => x"08",
          6087 => x"d5",
          6088 => x"8c",
          6089 => x"81",
          6090 => x"9f",
          6091 => x"2e",
          6092 => x"74",
          6093 => x"98",
          6094 => x"7e",
          6095 => x"3f",
          6096 => x"08",
          6097 => x"83",
          6098 => x"dc",
          6099 => x"89",
          6100 => x"77",
          6101 => x"d6",
          6102 => x"7f",
          6103 => x"58",
          6104 => x"75",
          6105 => x"75",
          6106 => x"77",
          6107 => x"7c",
          6108 => x"33",
          6109 => x"3f",
          6110 => x"08",
          6111 => x"7e",
          6112 => x"56",
          6113 => x"2e",
          6114 => x"16",
          6115 => x"55",
          6116 => x"94",
          6117 => x"53",
          6118 => x"b0",
          6119 => x"31",
          6120 => x"05",
          6121 => x"3f",
          6122 => x"56",
          6123 => x"9c",
          6124 => x"19",
          6125 => x"06",
          6126 => x"31",
          6127 => x"76",
          6128 => x"7b",
          6129 => x"08",
          6130 => x"d1",
          6131 => x"8c",
          6132 => x"81",
          6133 => x"94",
          6134 => x"ff",
          6135 => x"05",
          6136 => x"cf",
          6137 => x"76",
          6138 => x"17",
          6139 => x"1e",
          6140 => x"18",
          6141 => x"5e",
          6142 => x"39",
          6143 => x"82",
          6144 => x"90",
          6145 => x"f2",
          6146 => x"63",
          6147 => x"40",
          6148 => x"7e",
          6149 => x"fc",
          6150 => x"51",
          6151 => x"82",
          6152 => x"55",
          6153 => x"08",
          6154 => x"18",
          6155 => x"80",
          6156 => x"74",
          6157 => x"39",
          6158 => x"70",
          6159 => x"81",
          6160 => x"56",
          6161 => x"80",
          6162 => x"38",
          6163 => x"0b",
          6164 => x"82",
          6165 => x"39",
          6166 => x"19",
          6167 => x"83",
          6168 => x"18",
          6169 => x"56",
          6170 => x"27",
          6171 => x"09",
          6172 => x"2e",
          6173 => x"94",
          6174 => x"83",
          6175 => x"56",
          6176 => x"38",
          6177 => x"22",
          6178 => x"89",
          6179 => x"55",
          6180 => x"75",
          6181 => x"18",
          6182 => x"9c",
          6183 => x"85",
          6184 => x"08",
          6185 => x"d7",
          6186 => x"8c",
          6187 => x"82",
          6188 => x"80",
          6189 => x"38",
          6190 => x"ff",
          6191 => x"ff",
          6192 => x"38",
          6193 => x"0c",
          6194 => x"85",
          6195 => x"19",
          6196 => x"b0",
          6197 => x"19",
          6198 => x"81",
          6199 => x"74",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"98",
          6203 => x"7e",
          6204 => x"3f",
          6205 => x"08",
          6206 => x"d2",
          6207 => x"dc",
          6208 => x"89",
          6209 => x"78",
          6210 => x"d5",
          6211 => x"7f",
          6212 => x"58",
          6213 => x"75",
          6214 => x"75",
          6215 => x"78",
          6216 => x"7c",
          6217 => x"33",
          6218 => x"3f",
          6219 => x"08",
          6220 => x"7e",
          6221 => x"78",
          6222 => x"74",
          6223 => x"38",
          6224 => x"b0",
          6225 => x"31",
          6226 => x"05",
          6227 => x"51",
          6228 => x"7e",
          6229 => x"83",
          6230 => x"89",
          6231 => x"db",
          6232 => x"08",
          6233 => x"26",
          6234 => x"51",
          6235 => x"82",
          6236 => x"fd",
          6237 => x"77",
          6238 => x"55",
          6239 => x"0c",
          6240 => x"83",
          6241 => x"80",
          6242 => x"55",
          6243 => x"83",
          6244 => x"9c",
          6245 => x"7e",
          6246 => x"3f",
          6247 => x"08",
          6248 => x"75",
          6249 => x"94",
          6250 => x"ff",
          6251 => x"05",
          6252 => x"3f",
          6253 => x"0b",
          6254 => x"7b",
          6255 => x"08",
          6256 => x"76",
          6257 => x"08",
          6258 => x"1c",
          6259 => x"08",
          6260 => x"5c",
          6261 => x"83",
          6262 => x"74",
          6263 => x"fd",
          6264 => x"18",
          6265 => x"07",
          6266 => x"19",
          6267 => x"75",
          6268 => x"0c",
          6269 => x"04",
          6270 => x"7a",
          6271 => x"05",
          6272 => x"56",
          6273 => x"82",
          6274 => x"57",
          6275 => x"08",
          6276 => x"90",
          6277 => x"86",
          6278 => x"06",
          6279 => x"73",
          6280 => x"e9",
          6281 => x"08",
          6282 => x"cc",
          6283 => x"8c",
          6284 => x"82",
          6285 => x"80",
          6286 => x"16",
          6287 => x"33",
          6288 => x"55",
          6289 => x"34",
          6290 => x"53",
          6291 => x"08",
          6292 => x"3f",
          6293 => x"52",
          6294 => x"c9",
          6295 => x"88",
          6296 => x"96",
          6297 => x"f0",
          6298 => x"92",
          6299 => x"ca",
          6300 => x"81",
          6301 => x"34",
          6302 => x"df",
          6303 => x"dc",
          6304 => x"33",
          6305 => x"55",
          6306 => x"17",
          6307 => x"8c",
          6308 => x"3d",
          6309 => x"3d",
          6310 => x"52",
          6311 => x"3f",
          6312 => x"08",
          6313 => x"dc",
          6314 => x"86",
          6315 => x"52",
          6316 => x"bc",
          6317 => x"dc",
          6318 => x"8c",
          6319 => x"38",
          6320 => x"08",
          6321 => x"82",
          6322 => x"86",
          6323 => x"ff",
          6324 => x"3d",
          6325 => x"3f",
          6326 => x"0b",
          6327 => x"08",
          6328 => x"82",
          6329 => x"82",
          6330 => x"80",
          6331 => x"8c",
          6332 => x"3d",
          6333 => x"3d",
          6334 => x"93",
          6335 => x"52",
          6336 => x"e9",
          6337 => x"8c",
          6338 => x"82",
          6339 => x"80",
          6340 => x"58",
          6341 => x"3d",
          6342 => x"e0",
          6343 => x"8c",
          6344 => x"82",
          6345 => x"bc",
          6346 => x"c7",
          6347 => x"98",
          6348 => x"73",
          6349 => x"38",
          6350 => x"12",
          6351 => x"39",
          6352 => x"33",
          6353 => x"70",
          6354 => x"55",
          6355 => x"2e",
          6356 => x"7f",
          6357 => x"54",
          6358 => x"82",
          6359 => x"94",
          6360 => x"39",
          6361 => x"08",
          6362 => x"81",
          6363 => x"85",
          6364 => x"8c",
          6365 => x"3d",
          6366 => x"3d",
          6367 => x"5b",
          6368 => x"34",
          6369 => x"3d",
          6370 => x"52",
          6371 => x"e8",
          6372 => x"8c",
          6373 => x"82",
          6374 => x"82",
          6375 => x"43",
          6376 => x"11",
          6377 => x"58",
          6378 => x"80",
          6379 => x"38",
          6380 => x"3d",
          6381 => x"d5",
          6382 => x"8c",
          6383 => x"82",
          6384 => x"82",
          6385 => x"52",
          6386 => x"c8",
          6387 => x"dc",
          6388 => x"8c",
          6389 => x"c1",
          6390 => x"7b",
          6391 => x"3f",
          6392 => x"08",
          6393 => x"74",
          6394 => x"3f",
          6395 => x"08",
          6396 => x"dc",
          6397 => x"38",
          6398 => x"51",
          6399 => x"82",
          6400 => x"57",
          6401 => x"08",
          6402 => x"52",
          6403 => x"f2",
          6404 => x"8c",
          6405 => x"a6",
          6406 => x"74",
          6407 => x"3f",
          6408 => x"08",
          6409 => x"dc",
          6410 => x"cc",
          6411 => x"2e",
          6412 => x"86",
          6413 => x"81",
          6414 => x"81",
          6415 => x"3d",
          6416 => x"52",
          6417 => x"c9",
          6418 => x"3d",
          6419 => x"11",
          6420 => x"5a",
          6421 => x"2e",
          6422 => x"b9",
          6423 => x"16",
          6424 => x"33",
          6425 => x"73",
          6426 => x"16",
          6427 => x"26",
          6428 => x"75",
          6429 => x"38",
          6430 => x"05",
          6431 => x"6f",
          6432 => x"ff",
          6433 => x"55",
          6434 => x"74",
          6435 => x"38",
          6436 => x"11",
          6437 => x"74",
          6438 => x"39",
          6439 => x"09",
          6440 => x"38",
          6441 => x"11",
          6442 => x"74",
          6443 => x"82",
          6444 => x"70",
          6445 => x"fa",
          6446 => x"08",
          6447 => x"5c",
          6448 => x"73",
          6449 => x"38",
          6450 => x"1a",
          6451 => x"55",
          6452 => x"38",
          6453 => x"73",
          6454 => x"38",
          6455 => x"76",
          6456 => x"74",
          6457 => x"33",
          6458 => x"05",
          6459 => x"15",
          6460 => x"ba",
          6461 => x"05",
          6462 => x"ff",
          6463 => x"06",
          6464 => x"57",
          6465 => x"18",
          6466 => x"54",
          6467 => x"70",
          6468 => x"34",
          6469 => x"ee",
          6470 => x"34",
          6471 => x"dc",
          6472 => x"0d",
          6473 => x"0d",
          6474 => x"3d",
          6475 => x"71",
          6476 => x"ec",
          6477 => x"8c",
          6478 => x"82",
          6479 => x"82",
          6480 => x"15",
          6481 => x"82",
          6482 => x"15",
          6483 => x"76",
          6484 => x"90",
          6485 => x"81",
          6486 => x"06",
          6487 => x"72",
          6488 => x"56",
          6489 => x"54",
          6490 => x"17",
          6491 => x"78",
          6492 => x"38",
          6493 => x"22",
          6494 => x"59",
          6495 => x"78",
          6496 => x"76",
          6497 => x"51",
          6498 => x"3f",
          6499 => x"08",
          6500 => x"54",
          6501 => x"53",
          6502 => x"3f",
          6503 => x"08",
          6504 => x"38",
          6505 => x"75",
          6506 => x"18",
          6507 => x"31",
          6508 => x"57",
          6509 => x"b1",
          6510 => x"08",
          6511 => x"38",
          6512 => x"51",
          6513 => x"82",
          6514 => x"54",
          6515 => x"08",
          6516 => x"9a",
          6517 => x"dc",
          6518 => x"81",
          6519 => x"8c",
          6520 => x"16",
          6521 => x"16",
          6522 => x"2e",
          6523 => x"76",
          6524 => x"dc",
          6525 => x"31",
          6526 => x"18",
          6527 => x"90",
          6528 => x"81",
          6529 => x"06",
          6530 => x"56",
          6531 => x"9a",
          6532 => x"74",
          6533 => x"3f",
          6534 => x"08",
          6535 => x"dc",
          6536 => x"82",
          6537 => x"56",
          6538 => x"52",
          6539 => x"84",
          6540 => x"dc",
          6541 => x"ff",
          6542 => x"81",
          6543 => x"38",
          6544 => x"98",
          6545 => x"a6",
          6546 => x"16",
          6547 => x"39",
          6548 => x"16",
          6549 => x"75",
          6550 => x"53",
          6551 => x"aa",
          6552 => x"79",
          6553 => x"3f",
          6554 => x"08",
          6555 => x"0b",
          6556 => x"82",
          6557 => x"39",
          6558 => x"16",
          6559 => x"bb",
          6560 => x"2a",
          6561 => x"08",
          6562 => x"15",
          6563 => x"15",
          6564 => x"90",
          6565 => x"16",
          6566 => x"33",
          6567 => x"53",
          6568 => x"34",
          6569 => x"06",
          6570 => x"2e",
          6571 => x"9c",
          6572 => x"85",
          6573 => x"16",
          6574 => x"72",
          6575 => x"0c",
          6576 => x"04",
          6577 => x"79",
          6578 => x"75",
          6579 => x"8a",
          6580 => x"89",
          6581 => x"52",
          6582 => x"05",
          6583 => x"3f",
          6584 => x"08",
          6585 => x"dc",
          6586 => x"38",
          6587 => x"7a",
          6588 => x"d8",
          6589 => x"8c",
          6590 => x"82",
          6591 => x"80",
          6592 => x"16",
          6593 => x"2b",
          6594 => x"74",
          6595 => x"86",
          6596 => x"84",
          6597 => x"06",
          6598 => x"73",
          6599 => x"38",
          6600 => x"52",
          6601 => x"da",
          6602 => x"dc",
          6603 => x"0c",
          6604 => x"14",
          6605 => x"23",
          6606 => x"51",
          6607 => x"82",
          6608 => x"55",
          6609 => x"09",
          6610 => x"38",
          6611 => x"39",
          6612 => x"84",
          6613 => x"0c",
          6614 => x"82",
          6615 => x"89",
          6616 => x"fc",
          6617 => x"87",
          6618 => x"53",
          6619 => x"e7",
          6620 => x"8c",
          6621 => x"38",
          6622 => x"08",
          6623 => x"3d",
          6624 => x"3d",
          6625 => x"89",
          6626 => x"54",
          6627 => x"54",
          6628 => x"82",
          6629 => x"53",
          6630 => x"08",
          6631 => x"74",
          6632 => x"8c",
          6633 => x"73",
          6634 => x"3f",
          6635 => x"08",
          6636 => x"39",
          6637 => x"08",
          6638 => x"d3",
          6639 => x"8c",
          6640 => x"82",
          6641 => x"84",
          6642 => x"06",
          6643 => x"53",
          6644 => x"8c",
          6645 => x"38",
          6646 => x"51",
          6647 => x"72",
          6648 => x"cf",
          6649 => x"8c",
          6650 => x"32",
          6651 => x"72",
          6652 => x"70",
          6653 => x"08",
          6654 => x"54",
          6655 => x"8c",
          6656 => x"3d",
          6657 => x"3d",
          6658 => x"80",
          6659 => x"70",
          6660 => x"52",
          6661 => x"3f",
          6662 => x"08",
          6663 => x"dc",
          6664 => x"64",
          6665 => x"d6",
          6666 => x"8c",
          6667 => x"82",
          6668 => x"a0",
          6669 => x"cb",
          6670 => x"98",
          6671 => x"73",
          6672 => x"38",
          6673 => x"39",
          6674 => x"88",
          6675 => x"75",
          6676 => x"3f",
          6677 => x"dc",
          6678 => x"0d",
          6679 => x"0d",
          6680 => x"5c",
          6681 => x"3d",
          6682 => x"93",
          6683 => x"d6",
          6684 => x"dc",
          6685 => x"8c",
          6686 => x"80",
          6687 => x"0c",
          6688 => x"11",
          6689 => x"90",
          6690 => x"56",
          6691 => x"74",
          6692 => x"75",
          6693 => x"e4",
          6694 => x"81",
          6695 => x"5b",
          6696 => x"82",
          6697 => x"75",
          6698 => x"73",
          6699 => x"81",
          6700 => x"82",
          6701 => x"76",
          6702 => x"f0",
          6703 => x"f4",
          6704 => x"dc",
          6705 => x"d1",
          6706 => x"dc",
          6707 => x"ce",
          6708 => x"dc",
          6709 => x"82",
          6710 => x"07",
          6711 => x"05",
          6712 => x"53",
          6713 => x"98",
          6714 => x"26",
          6715 => x"f9",
          6716 => x"08",
          6717 => x"08",
          6718 => x"98",
          6719 => x"81",
          6720 => x"58",
          6721 => x"3f",
          6722 => x"08",
          6723 => x"dc",
          6724 => x"38",
          6725 => x"77",
          6726 => x"5d",
          6727 => x"74",
          6728 => x"81",
          6729 => x"b4",
          6730 => x"bb",
          6731 => x"8c",
          6732 => x"ff",
          6733 => x"30",
          6734 => x"1b",
          6735 => x"5b",
          6736 => x"39",
          6737 => x"ff",
          6738 => x"82",
          6739 => x"f0",
          6740 => x"30",
          6741 => x"1b",
          6742 => x"5b",
          6743 => x"83",
          6744 => x"58",
          6745 => x"92",
          6746 => x"0c",
          6747 => x"12",
          6748 => x"33",
          6749 => x"54",
          6750 => x"34",
          6751 => x"dc",
          6752 => x"0d",
          6753 => x"0d",
          6754 => x"fc",
          6755 => x"52",
          6756 => x"3f",
          6757 => x"08",
          6758 => x"dc",
          6759 => x"38",
          6760 => x"56",
          6761 => x"38",
          6762 => x"70",
          6763 => x"81",
          6764 => x"55",
          6765 => x"80",
          6766 => x"38",
          6767 => x"54",
          6768 => x"08",
          6769 => x"38",
          6770 => x"82",
          6771 => x"53",
          6772 => x"52",
          6773 => x"8c",
          6774 => x"dc",
          6775 => x"19",
          6776 => x"c9",
          6777 => x"08",
          6778 => x"ff",
          6779 => x"82",
          6780 => x"ff",
          6781 => x"06",
          6782 => x"56",
          6783 => x"08",
          6784 => x"81",
          6785 => x"82",
          6786 => x"75",
          6787 => x"54",
          6788 => x"08",
          6789 => x"27",
          6790 => x"17",
          6791 => x"8c",
          6792 => x"76",
          6793 => x"3f",
          6794 => x"08",
          6795 => x"08",
          6796 => x"90",
          6797 => x"c0",
          6798 => x"90",
          6799 => x"80",
          6800 => x"75",
          6801 => x"75",
          6802 => x"8c",
          6803 => x"3d",
          6804 => x"3d",
          6805 => x"a0",
          6806 => x"05",
          6807 => x"51",
          6808 => x"82",
          6809 => x"55",
          6810 => x"08",
          6811 => x"78",
          6812 => x"08",
          6813 => x"70",
          6814 => x"ae",
          6815 => x"dc",
          6816 => x"8c",
          6817 => x"db",
          6818 => x"fb",
          6819 => x"85",
          6820 => x"06",
          6821 => x"86",
          6822 => x"c7",
          6823 => x"2b",
          6824 => x"24",
          6825 => x"02",
          6826 => x"33",
          6827 => x"58",
          6828 => x"76",
          6829 => x"6b",
          6830 => x"cc",
          6831 => x"8c",
          6832 => x"84",
          6833 => x"06",
          6834 => x"73",
          6835 => x"d4",
          6836 => x"82",
          6837 => x"94",
          6838 => x"81",
          6839 => x"5a",
          6840 => x"08",
          6841 => x"8a",
          6842 => x"54",
          6843 => x"82",
          6844 => x"55",
          6845 => x"08",
          6846 => x"82",
          6847 => x"52",
          6848 => x"e5",
          6849 => x"dc",
          6850 => x"8c",
          6851 => x"38",
          6852 => x"cf",
          6853 => x"dc",
          6854 => x"88",
          6855 => x"dc",
          6856 => x"38",
          6857 => x"c2",
          6858 => x"dc",
          6859 => x"dc",
          6860 => x"82",
          6861 => x"07",
          6862 => x"55",
          6863 => x"2e",
          6864 => x"80",
          6865 => x"80",
          6866 => x"77",
          6867 => x"3f",
          6868 => x"08",
          6869 => x"38",
          6870 => x"ba",
          6871 => x"8c",
          6872 => x"74",
          6873 => x"0c",
          6874 => x"04",
          6875 => x"82",
          6876 => x"c0",
          6877 => x"3d",
          6878 => x"3f",
          6879 => x"08",
          6880 => x"dc",
          6881 => x"38",
          6882 => x"52",
          6883 => x"52",
          6884 => x"3f",
          6885 => x"08",
          6886 => x"dc",
          6887 => x"88",
          6888 => x"39",
          6889 => x"08",
          6890 => x"81",
          6891 => x"38",
          6892 => x"05",
          6893 => x"2a",
          6894 => x"55",
          6895 => x"81",
          6896 => x"5a",
          6897 => x"3d",
          6898 => x"c1",
          6899 => x"8c",
          6900 => x"55",
          6901 => x"dc",
          6902 => x"87",
          6903 => x"dc",
          6904 => x"09",
          6905 => x"38",
          6906 => x"8c",
          6907 => x"2e",
          6908 => x"86",
          6909 => x"81",
          6910 => x"81",
          6911 => x"8c",
          6912 => x"78",
          6913 => x"3f",
          6914 => x"08",
          6915 => x"dc",
          6916 => x"38",
          6917 => x"52",
          6918 => x"ff",
          6919 => x"78",
          6920 => x"b4",
          6921 => x"54",
          6922 => x"15",
          6923 => x"b2",
          6924 => x"ca",
          6925 => x"b6",
          6926 => x"53",
          6927 => x"53",
          6928 => x"3f",
          6929 => x"b4",
          6930 => x"d4",
          6931 => x"b6",
          6932 => x"54",
          6933 => x"d5",
          6934 => x"53",
          6935 => x"11",
          6936 => x"d7",
          6937 => x"81",
          6938 => x"34",
          6939 => x"a4",
          6940 => x"dc",
          6941 => x"8c",
          6942 => x"38",
          6943 => x"0a",
          6944 => x"05",
          6945 => x"d0",
          6946 => x"64",
          6947 => x"c9",
          6948 => x"54",
          6949 => x"15",
          6950 => x"81",
          6951 => x"34",
          6952 => x"b8",
          6953 => x"8c",
          6954 => x"8b",
          6955 => x"75",
          6956 => x"ff",
          6957 => x"73",
          6958 => x"0c",
          6959 => x"04",
          6960 => x"a9",
          6961 => x"51",
          6962 => x"82",
          6963 => x"ff",
          6964 => x"a9",
          6965 => x"ee",
          6966 => x"dc",
          6967 => x"8c",
          6968 => x"d3",
          6969 => x"a9",
          6970 => x"9d",
          6971 => x"58",
          6972 => x"82",
          6973 => x"55",
          6974 => x"08",
          6975 => x"02",
          6976 => x"33",
          6977 => x"54",
          6978 => x"82",
          6979 => x"53",
          6980 => x"52",
          6981 => x"88",
          6982 => x"b4",
          6983 => x"53",
          6984 => x"3d",
          6985 => x"ff",
          6986 => x"aa",
          6987 => x"73",
          6988 => x"3f",
          6989 => x"08",
          6990 => x"dc",
          6991 => x"63",
          6992 => x"81",
          6993 => x"65",
          6994 => x"2e",
          6995 => x"55",
          6996 => x"82",
          6997 => x"84",
          6998 => x"06",
          6999 => x"73",
          7000 => x"3f",
          7001 => x"08",
          7002 => x"dc",
          7003 => x"38",
          7004 => x"53",
          7005 => x"95",
          7006 => x"16",
          7007 => x"87",
          7008 => x"05",
          7009 => x"34",
          7010 => x"70",
          7011 => x"81",
          7012 => x"55",
          7013 => x"74",
          7014 => x"73",
          7015 => x"78",
          7016 => x"83",
          7017 => x"16",
          7018 => x"2a",
          7019 => x"51",
          7020 => x"80",
          7021 => x"38",
          7022 => x"80",
          7023 => x"52",
          7024 => x"be",
          7025 => x"dc",
          7026 => x"51",
          7027 => x"3f",
          7028 => x"8c",
          7029 => x"2e",
          7030 => x"82",
          7031 => x"52",
          7032 => x"b5",
          7033 => x"8c",
          7034 => x"80",
          7035 => x"58",
          7036 => x"dc",
          7037 => x"38",
          7038 => x"54",
          7039 => x"09",
          7040 => x"38",
          7041 => x"52",
          7042 => x"af",
          7043 => x"81",
          7044 => x"34",
          7045 => x"8c",
          7046 => x"38",
          7047 => x"ca",
          7048 => x"dc",
          7049 => x"8c",
          7050 => x"38",
          7051 => x"b5",
          7052 => x"8c",
          7053 => x"74",
          7054 => x"0c",
          7055 => x"04",
          7056 => x"02",
          7057 => x"33",
          7058 => x"80",
          7059 => x"57",
          7060 => x"95",
          7061 => x"52",
          7062 => x"d2",
          7063 => x"8c",
          7064 => x"82",
          7065 => x"80",
          7066 => x"5a",
          7067 => x"3d",
          7068 => x"c9",
          7069 => x"8c",
          7070 => x"82",
          7071 => x"b8",
          7072 => x"cf",
          7073 => x"a0",
          7074 => x"55",
          7075 => x"75",
          7076 => x"71",
          7077 => x"33",
          7078 => x"74",
          7079 => x"57",
          7080 => x"8b",
          7081 => x"54",
          7082 => x"15",
          7083 => x"ff",
          7084 => x"82",
          7085 => x"55",
          7086 => x"dc",
          7087 => x"0d",
          7088 => x"0d",
          7089 => x"53",
          7090 => x"05",
          7091 => x"51",
          7092 => x"82",
          7093 => x"55",
          7094 => x"08",
          7095 => x"76",
          7096 => x"93",
          7097 => x"51",
          7098 => x"82",
          7099 => x"55",
          7100 => x"08",
          7101 => x"80",
          7102 => x"81",
          7103 => x"86",
          7104 => x"38",
          7105 => x"86",
          7106 => x"90",
          7107 => x"54",
          7108 => x"ff",
          7109 => x"76",
          7110 => x"83",
          7111 => x"51",
          7112 => x"3f",
          7113 => x"08",
          7114 => x"8c",
          7115 => x"3d",
          7116 => x"3d",
          7117 => x"5c",
          7118 => x"98",
          7119 => x"52",
          7120 => x"d1",
          7121 => x"8c",
          7122 => x"8c",
          7123 => x"70",
          7124 => x"08",
          7125 => x"51",
          7126 => x"80",
          7127 => x"38",
          7128 => x"06",
          7129 => x"80",
          7130 => x"38",
          7131 => x"5f",
          7132 => x"3d",
          7133 => x"ff",
          7134 => x"82",
          7135 => x"57",
          7136 => x"08",
          7137 => x"74",
          7138 => x"c3",
          7139 => x"8c",
          7140 => x"82",
          7141 => x"bf",
          7142 => x"dc",
          7143 => x"dc",
          7144 => x"59",
          7145 => x"81",
          7146 => x"56",
          7147 => x"33",
          7148 => x"16",
          7149 => x"27",
          7150 => x"56",
          7151 => x"80",
          7152 => x"80",
          7153 => x"ff",
          7154 => x"70",
          7155 => x"56",
          7156 => x"e8",
          7157 => x"76",
          7158 => x"81",
          7159 => x"80",
          7160 => x"57",
          7161 => x"78",
          7162 => x"51",
          7163 => x"2e",
          7164 => x"73",
          7165 => x"38",
          7166 => x"08",
          7167 => x"b1",
          7168 => x"8c",
          7169 => x"82",
          7170 => x"a7",
          7171 => x"33",
          7172 => x"c3",
          7173 => x"2e",
          7174 => x"e4",
          7175 => x"2e",
          7176 => x"56",
          7177 => x"05",
          7178 => x"e3",
          7179 => x"dc",
          7180 => x"76",
          7181 => x"0c",
          7182 => x"04",
          7183 => x"82",
          7184 => x"ff",
          7185 => x"9d",
          7186 => x"fa",
          7187 => x"dc",
          7188 => x"dc",
          7189 => x"82",
          7190 => x"83",
          7191 => x"53",
          7192 => x"3d",
          7193 => x"ff",
          7194 => x"73",
          7195 => x"70",
          7196 => x"52",
          7197 => x"9f",
          7198 => x"bc",
          7199 => x"74",
          7200 => x"6d",
          7201 => x"70",
          7202 => x"af",
          7203 => x"8c",
          7204 => x"2e",
          7205 => x"70",
          7206 => x"57",
          7207 => x"fd",
          7208 => x"dc",
          7209 => x"8d",
          7210 => x"2b",
          7211 => x"81",
          7212 => x"86",
          7213 => x"dc",
          7214 => x"9f",
          7215 => x"ff",
          7216 => x"54",
          7217 => x"8a",
          7218 => x"70",
          7219 => x"06",
          7220 => x"ff",
          7221 => x"38",
          7222 => x"15",
          7223 => x"80",
          7224 => x"74",
          7225 => x"ec",
          7226 => x"89",
          7227 => x"dc",
          7228 => x"81",
          7229 => x"88",
          7230 => x"26",
          7231 => x"39",
          7232 => x"86",
          7233 => x"81",
          7234 => x"ff",
          7235 => x"38",
          7236 => x"54",
          7237 => x"81",
          7238 => x"81",
          7239 => x"78",
          7240 => x"5a",
          7241 => x"6d",
          7242 => x"81",
          7243 => x"57",
          7244 => x"9f",
          7245 => x"38",
          7246 => x"54",
          7247 => x"81",
          7248 => x"b1",
          7249 => x"2e",
          7250 => x"a7",
          7251 => x"15",
          7252 => x"54",
          7253 => x"09",
          7254 => x"38",
          7255 => x"76",
          7256 => x"41",
          7257 => x"52",
          7258 => x"52",
          7259 => x"b3",
          7260 => x"dc",
          7261 => x"8c",
          7262 => x"f7",
          7263 => x"74",
          7264 => x"e5",
          7265 => x"dc",
          7266 => x"8c",
          7267 => x"38",
          7268 => x"38",
          7269 => x"74",
          7270 => x"39",
          7271 => x"08",
          7272 => x"81",
          7273 => x"38",
          7274 => x"74",
          7275 => x"38",
          7276 => x"51",
          7277 => x"3f",
          7278 => x"08",
          7279 => x"dc",
          7280 => x"a0",
          7281 => x"dc",
          7282 => x"51",
          7283 => x"3f",
          7284 => x"0b",
          7285 => x"8b",
          7286 => x"67",
          7287 => x"a7",
          7288 => x"81",
          7289 => x"34",
          7290 => x"ad",
          7291 => x"8c",
          7292 => x"73",
          7293 => x"8c",
          7294 => x"3d",
          7295 => x"3d",
          7296 => x"02",
          7297 => x"cb",
          7298 => x"3d",
          7299 => x"72",
          7300 => x"5a",
          7301 => x"82",
          7302 => x"58",
          7303 => x"08",
          7304 => x"91",
          7305 => x"77",
          7306 => x"7c",
          7307 => x"38",
          7308 => x"59",
          7309 => x"90",
          7310 => x"81",
          7311 => x"06",
          7312 => x"73",
          7313 => x"54",
          7314 => x"82",
          7315 => x"39",
          7316 => x"8b",
          7317 => x"11",
          7318 => x"2b",
          7319 => x"54",
          7320 => x"fe",
          7321 => x"ff",
          7322 => x"70",
          7323 => x"07",
          7324 => x"8c",
          7325 => x"8c",
          7326 => x"40",
          7327 => x"55",
          7328 => x"88",
          7329 => x"08",
          7330 => x"38",
          7331 => x"77",
          7332 => x"56",
          7333 => x"51",
          7334 => x"3f",
          7335 => x"55",
          7336 => x"08",
          7337 => x"38",
          7338 => x"8c",
          7339 => x"2e",
          7340 => x"82",
          7341 => x"ff",
          7342 => x"38",
          7343 => x"08",
          7344 => x"16",
          7345 => x"2e",
          7346 => x"87",
          7347 => x"74",
          7348 => x"74",
          7349 => x"81",
          7350 => x"38",
          7351 => x"ff",
          7352 => x"2e",
          7353 => x"7b",
          7354 => x"80",
          7355 => x"81",
          7356 => x"81",
          7357 => x"06",
          7358 => x"56",
          7359 => x"52",
          7360 => x"af",
          7361 => x"8c",
          7362 => x"82",
          7363 => x"80",
          7364 => x"81",
          7365 => x"56",
          7366 => x"d3",
          7367 => x"ff",
          7368 => x"7c",
          7369 => x"55",
          7370 => x"b3",
          7371 => x"1b",
          7372 => x"1b",
          7373 => x"33",
          7374 => x"54",
          7375 => x"34",
          7376 => x"fe",
          7377 => x"08",
          7378 => x"74",
          7379 => x"75",
          7380 => x"16",
          7381 => x"33",
          7382 => x"73",
          7383 => x"77",
          7384 => x"8c",
          7385 => x"3d",
          7386 => x"3d",
          7387 => x"02",
          7388 => x"eb",
          7389 => x"3d",
          7390 => x"59",
          7391 => x"8b",
          7392 => x"82",
          7393 => x"24",
          7394 => x"82",
          7395 => x"84",
          7396 => x"8c",
          7397 => x"51",
          7398 => x"2e",
          7399 => x"75",
          7400 => x"dc",
          7401 => x"06",
          7402 => x"7e",
          7403 => x"d0",
          7404 => x"dc",
          7405 => x"06",
          7406 => x"56",
          7407 => x"74",
          7408 => x"76",
          7409 => x"81",
          7410 => x"8a",
          7411 => x"b2",
          7412 => x"fc",
          7413 => x"52",
          7414 => x"a4",
          7415 => x"8c",
          7416 => x"38",
          7417 => x"80",
          7418 => x"74",
          7419 => x"26",
          7420 => x"15",
          7421 => x"74",
          7422 => x"38",
          7423 => x"80",
          7424 => x"84",
          7425 => x"92",
          7426 => x"80",
          7427 => x"38",
          7428 => x"06",
          7429 => x"2e",
          7430 => x"56",
          7431 => x"78",
          7432 => x"89",
          7433 => x"2b",
          7434 => x"43",
          7435 => x"38",
          7436 => x"30",
          7437 => x"77",
          7438 => x"91",
          7439 => x"c2",
          7440 => x"f8",
          7441 => x"52",
          7442 => x"a4",
          7443 => x"56",
          7444 => x"08",
          7445 => x"77",
          7446 => x"77",
          7447 => x"dc",
          7448 => x"45",
          7449 => x"bf",
          7450 => x"8e",
          7451 => x"26",
          7452 => x"74",
          7453 => x"48",
          7454 => x"75",
          7455 => x"38",
          7456 => x"81",
          7457 => x"fa",
          7458 => x"2a",
          7459 => x"56",
          7460 => x"2e",
          7461 => x"87",
          7462 => x"82",
          7463 => x"38",
          7464 => x"55",
          7465 => x"83",
          7466 => x"81",
          7467 => x"56",
          7468 => x"80",
          7469 => x"38",
          7470 => x"83",
          7471 => x"06",
          7472 => x"78",
          7473 => x"91",
          7474 => x"0b",
          7475 => x"22",
          7476 => x"80",
          7477 => x"74",
          7478 => x"38",
          7479 => x"56",
          7480 => x"17",
          7481 => x"57",
          7482 => x"2e",
          7483 => x"75",
          7484 => x"79",
          7485 => x"fe",
          7486 => x"82",
          7487 => x"84",
          7488 => x"05",
          7489 => x"5e",
          7490 => x"80",
          7491 => x"dc",
          7492 => x"8a",
          7493 => x"fd",
          7494 => x"75",
          7495 => x"38",
          7496 => x"78",
          7497 => x"8c",
          7498 => x"0b",
          7499 => x"22",
          7500 => x"80",
          7501 => x"74",
          7502 => x"38",
          7503 => x"56",
          7504 => x"17",
          7505 => x"57",
          7506 => x"2e",
          7507 => x"75",
          7508 => x"79",
          7509 => x"fe",
          7510 => x"82",
          7511 => x"10",
          7512 => x"82",
          7513 => x"9f",
          7514 => x"38",
          7515 => x"8c",
          7516 => x"82",
          7517 => x"05",
          7518 => x"2a",
          7519 => x"56",
          7520 => x"17",
          7521 => x"81",
          7522 => x"60",
          7523 => x"65",
          7524 => x"12",
          7525 => x"30",
          7526 => x"74",
          7527 => x"59",
          7528 => x"7d",
          7529 => x"81",
          7530 => x"76",
          7531 => x"41",
          7532 => x"76",
          7533 => x"90",
          7534 => x"62",
          7535 => x"51",
          7536 => x"26",
          7537 => x"75",
          7538 => x"31",
          7539 => x"65",
          7540 => x"fe",
          7541 => x"82",
          7542 => x"58",
          7543 => x"09",
          7544 => x"38",
          7545 => x"08",
          7546 => x"26",
          7547 => x"78",
          7548 => x"79",
          7549 => x"78",
          7550 => x"86",
          7551 => x"82",
          7552 => x"06",
          7553 => x"83",
          7554 => x"82",
          7555 => x"27",
          7556 => x"8f",
          7557 => x"55",
          7558 => x"26",
          7559 => x"59",
          7560 => x"62",
          7561 => x"74",
          7562 => x"38",
          7563 => x"88",
          7564 => x"dc",
          7565 => x"26",
          7566 => x"86",
          7567 => x"1a",
          7568 => x"79",
          7569 => x"38",
          7570 => x"80",
          7571 => x"2e",
          7572 => x"83",
          7573 => x"9f",
          7574 => x"8b",
          7575 => x"06",
          7576 => x"74",
          7577 => x"84",
          7578 => x"52",
          7579 => x"a2",
          7580 => x"53",
          7581 => x"52",
          7582 => x"a2",
          7583 => x"80",
          7584 => x"51",
          7585 => x"3f",
          7586 => x"34",
          7587 => x"ff",
          7588 => x"1b",
          7589 => x"a2",
          7590 => x"90",
          7591 => x"83",
          7592 => x"70",
          7593 => x"80",
          7594 => x"55",
          7595 => x"ff",
          7596 => x"66",
          7597 => x"ff",
          7598 => x"38",
          7599 => x"ff",
          7600 => x"1b",
          7601 => x"f2",
          7602 => x"74",
          7603 => x"51",
          7604 => x"3f",
          7605 => x"1c",
          7606 => x"98",
          7607 => x"a0",
          7608 => x"ff",
          7609 => x"51",
          7610 => x"3f",
          7611 => x"1b",
          7612 => x"e4",
          7613 => x"2e",
          7614 => x"80",
          7615 => x"88",
          7616 => x"80",
          7617 => x"ff",
          7618 => x"7c",
          7619 => x"51",
          7620 => x"3f",
          7621 => x"1b",
          7622 => x"bc",
          7623 => x"b0",
          7624 => x"a0",
          7625 => x"52",
          7626 => x"ff",
          7627 => x"ff",
          7628 => x"c0",
          7629 => x"0b",
          7630 => x"34",
          7631 => x"fa",
          7632 => x"c7",
          7633 => x"39",
          7634 => x"0a",
          7635 => x"51",
          7636 => x"3f",
          7637 => x"ff",
          7638 => x"1b",
          7639 => x"da",
          7640 => x"0b",
          7641 => x"a9",
          7642 => x"34",
          7643 => x"fa",
          7644 => x"1b",
          7645 => x"8f",
          7646 => x"d5",
          7647 => x"1b",
          7648 => x"ff",
          7649 => x"81",
          7650 => x"7a",
          7651 => x"ff",
          7652 => x"81",
          7653 => x"dc",
          7654 => x"38",
          7655 => x"09",
          7656 => x"ee",
          7657 => x"60",
          7658 => x"7a",
          7659 => x"ff",
          7660 => x"84",
          7661 => x"52",
          7662 => x"9f",
          7663 => x"8b",
          7664 => x"52",
          7665 => x"9f",
          7666 => x"8a",
          7667 => x"52",
          7668 => x"51",
          7669 => x"3f",
          7670 => x"83",
          7671 => x"ff",
          7672 => x"82",
          7673 => x"1b",
          7674 => x"ec",
          7675 => x"d5",
          7676 => x"ff",
          7677 => x"75",
          7678 => x"05",
          7679 => x"7e",
          7680 => x"e5",
          7681 => x"60",
          7682 => x"52",
          7683 => x"9a",
          7684 => x"53",
          7685 => x"51",
          7686 => x"3f",
          7687 => x"58",
          7688 => x"09",
          7689 => x"38",
          7690 => x"51",
          7691 => x"3f",
          7692 => x"1b",
          7693 => x"a0",
          7694 => x"52",
          7695 => x"91",
          7696 => x"ff",
          7697 => x"81",
          7698 => x"f8",
          7699 => x"7a",
          7700 => x"84",
          7701 => x"61",
          7702 => x"26",
          7703 => x"57",
          7704 => x"53",
          7705 => x"51",
          7706 => x"3f",
          7707 => x"08",
          7708 => x"84",
          7709 => x"8c",
          7710 => x"7a",
          7711 => x"aa",
          7712 => x"75",
          7713 => x"56",
          7714 => x"81",
          7715 => x"80",
          7716 => x"38",
          7717 => x"83",
          7718 => x"63",
          7719 => x"74",
          7720 => x"38",
          7721 => x"54",
          7722 => x"52",
          7723 => x"99",
          7724 => x"8c",
          7725 => x"c1",
          7726 => x"75",
          7727 => x"56",
          7728 => x"8c",
          7729 => x"2e",
          7730 => x"56",
          7731 => x"ff",
          7732 => x"84",
          7733 => x"2e",
          7734 => x"56",
          7735 => x"58",
          7736 => x"38",
          7737 => x"77",
          7738 => x"ff",
          7739 => x"82",
          7740 => x"78",
          7741 => x"c2",
          7742 => x"1b",
          7743 => x"34",
          7744 => x"16",
          7745 => x"82",
          7746 => x"83",
          7747 => x"84",
          7748 => x"67",
          7749 => x"fd",
          7750 => x"51",
          7751 => x"3f",
          7752 => x"16",
          7753 => x"dc",
          7754 => x"bf",
          7755 => x"86",
          7756 => x"8c",
          7757 => x"16",
          7758 => x"83",
          7759 => x"ff",
          7760 => x"66",
          7761 => x"1b",
          7762 => x"8c",
          7763 => x"77",
          7764 => x"7e",
          7765 => x"91",
          7766 => x"82",
          7767 => x"a2",
          7768 => x"80",
          7769 => x"ff",
          7770 => x"81",
          7771 => x"dc",
          7772 => x"89",
          7773 => x"8a",
          7774 => x"86",
          7775 => x"dc",
          7776 => x"82",
          7777 => x"99",
          7778 => x"f5",
          7779 => x"60",
          7780 => x"79",
          7781 => x"5a",
          7782 => x"78",
          7783 => x"8d",
          7784 => x"55",
          7785 => x"fc",
          7786 => x"51",
          7787 => x"7a",
          7788 => x"81",
          7789 => x"8c",
          7790 => x"74",
          7791 => x"38",
          7792 => x"81",
          7793 => x"81",
          7794 => x"8a",
          7795 => x"06",
          7796 => x"76",
          7797 => x"76",
          7798 => x"55",
          7799 => x"dc",
          7800 => x"0d",
          7801 => x"0d",
          7802 => x"05",
          7803 => x"59",
          7804 => x"2e",
          7805 => x"87",
          7806 => x"76",
          7807 => x"84",
          7808 => x"80",
          7809 => x"38",
          7810 => x"77",
          7811 => x"56",
          7812 => x"34",
          7813 => x"bb",
          7814 => x"38",
          7815 => x"05",
          7816 => x"8c",
          7817 => x"08",
          7818 => x"3f",
          7819 => x"70",
          7820 => x"07",
          7821 => x"30",
          7822 => x"56",
          7823 => x"0c",
          7824 => x"18",
          7825 => x"0d",
          7826 => x"0d",
          7827 => x"08",
          7828 => x"75",
          7829 => x"89",
          7830 => x"54",
          7831 => x"16",
          7832 => x"51",
          7833 => x"82",
          7834 => x"91",
          7835 => x"08",
          7836 => x"81",
          7837 => x"88",
          7838 => x"83",
          7839 => x"74",
          7840 => x"0c",
          7841 => x"04",
          7842 => x"75",
          7843 => x"53",
          7844 => x"51",
          7845 => x"3f",
          7846 => x"85",
          7847 => x"ea",
          7848 => x"80",
          7849 => x"6a",
          7850 => x"70",
          7851 => x"d8",
          7852 => x"72",
          7853 => x"3f",
          7854 => x"8d",
          7855 => x"0d",
          7856 => x"0d",
          7857 => x"70",
          7858 => x"74",
          7859 => x"e1",
          7860 => x"77",
          7861 => x"85",
          7862 => x"80",
          7863 => x"33",
          7864 => x"2e",
          7865 => x"86",
          7866 => x"55",
          7867 => x"57",
          7868 => x"82",
          7869 => x"70",
          7870 => x"fe",
          7871 => x"82",
          7872 => x"82",
          7873 => x"54",
          7874 => x"08",
          7875 => x"db",
          7876 => x"8c",
          7877 => x"38",
          7878 => x"54",
          7879 => x"ff",
          7880 => x"17",
          7881 => x"06",
          7882 => x"77",
          7883 => x"ff",
          7884 => x"8c",
          7885 => x"3d",
          7886 => x"3d",
          7887 => x"71",
          7888 => x"8e",
          7889 => x"29",
          7890 => x"05",
          7891 => x"04",
          7892 => x"51",
          7893 => x"81",
          7894 => x"80",
          7895 => x"fd",
          7896 => x"f2",
          7897 => x"fc",
          7898 => x"39",
          7899 => x"51",
          7900 => x"81",
          7901 => x"80",
          7902 => x"fe",
          7903 => x"d6",
          7904 => x"c0",
          7905 => x"39",
          7906 => x"51",
          7907 => x"81",
          7908 => x"80",
          7909 => x"ff",
          7910 => x"39",
          7911 => x"51",
          7912 => x"ff",
          7913 => x"39",
          7914 => x"51",
          7915 => x"ff",
          7916 => x"39",
          7917 => x"51",
          7918 => x"80",
          7919 => x"39",
          7920 => x"51",
          7921 => x"80",
          7922 => x"39",
          7923 => x"51",
          7924 => x"81",
          7925 => x"f2",
          7926 => x"3d",
          7927 => x"3d",
          7928 => x"56",
          7929 => x"e7",
          7930 => x"74",
          7931 => x"e8",
          7932 => x"39",
          7933 => x"74",
          7934 => x"df",
          7935 => x"dc",
          7936 => x"51",
          7937 => x"3f",
          7938 => x"08",
          7939 => x"75",
          7940 => x"90",
          7941 => x"d3",
          7942 => x"0d",
          7943 => x"0d",
          7944 => x"05",
          7945 => x"33",
          7946 => x"68",
          7947 => x"7a",
          7948 => x"51",
          7949 => x"78",
          7950 => x"ff",
          7951 => x"81",
          7952 => x"07",
          7953 => x"06",
          7954 => x"56",
          7955 => x"38",
          7956 => x"52",
          7957 => x"52",
          7958 => x"c9",
          7959 => x"dc",
          7960 => x"8c",
          7961 => x"38",
          7962 => x"08",
          7963 => x"88",
          7964 => x"dc",
          7965 => x"3d",
          7966 => x"84",
          7967 => x"52",
          7968 => x"86",
          7969 => x"dc",
          7970 => x"8c",
          7971 => x"38",
          7972 => x"80",
          7973 => x"74",
          7974 => x"59",
          7975 => x"96",
          7976 => x"51",
          7977 => x"76",
          7978 => x"07",
          7979 => x"30",
          7980 => x"72",
          7981 => x"51",
          7982 => x"2e",
          7983 => x"81",
          7984 => x"c0",
          7985 => x"52",
          7986 => x"92",
          7987 => x"75",
          7988 => x"0c",
          7989 => x"04",
          7990 => x"7b",
          7991 => x"b3",
          7992 => x"58",
          7993 => x"53",
          7994 => x"51",
          7995 => x"82",
          7996 => x"a4",
          7997 => x"2e",
          7998 => x"81",
          7999 => x"98",
          8000 => x"7f",
          8001 => x"dc",
          8002 => x"7d",
          8003 => x"82",
          8004 => x"57",
          8005 => x"04",
          8006 => x"dc",
          8007 => x"0d",
          8008 => x"0d",
          8009 => x"02",
          8010 => x"cf",
          8011 => x"73",
          8012 => x"5f",
          8013 => x"5e",
          8014 => x"82",
          8015 => x"fe",
          8016 => x"82",
          8017 => x"fe",
          8018 => x"80",
          8019 => x"27",
          8020 => x"7b",
          8021 => x"38",
          8022 => x"a7",
          8023 => x"39",
          8024 => x"72",
          8025 => x"38",
          8026 => x"82",
          8027 => x"fe",
          8028 => x"89",
          8029 => x"d4",
          8030 => x"8b",
          8031 => x"55",
          8032 => x"74",
          8033 => x"7a",
          8034 => x"72",
          8035 => x"81",
          8036 => x"f4",
          8037 => x"39",
          8038 => x"51",
          8039 => x"3f",
          8040 => x"a1",
          8041 => x"53",
          8042 => x"8e",
          8043 => x"52",
          8044 => x"51",
          8045 => x"3f",
          8046 => x"81",
          8047 => x"ee",
          8048 => x"15",
          8049 => x"fe",
          8050 => x"ff",
          8051 => x"81",
          8052 => x"ee",
          8053 => x"55",
          8054 => x"bc",
          8055 => x"70",
          8056 => x"80",
          8057 => x"27",
          8058 => x"56",
          8059 => x"74",
          8060 => x"81",
          8061 => x"06",
          8062 => x"06",
          8063 => x"80",
          8064 => x"73",
          8065 => x"85",
          8066 => x"83",
          8067 => x"fe",
          8068 => x"81",
          8069 => x"39",
          8070 => x"51",
          8071 => x"3f",
          8072 => x"1c",
          8073 => x"de",
          8074 => x"8c",
          8075 => x"2b",
          8076 => x"51",
          8077 => x"2e",
          8078 => x"ab",
          8079 => x"be",
          8080 => x"dc",
          8081 => x"70",
          8082 => x"a0",
          8083 => x"72",
          8084 => x"30",
          8085 => x"73",
          8086 => x"51",
          8087 => x"57",
          8088 => x"73",
          8089 => x"76",
          8090 => x"81",
          8091 => x"80",
          8092 => x"7c",
          8093 => x"78",
          8094 => x"38",
          8095 => x"82",
          8096 => x"8f",
          8097 => x"fc",
          8098 => x"9b",
          8099 => x"81",
          8100 => x"81",
          8101 => x"fe",
          8102 => x"82",
          8103 => x"51",
          8104 => x"3f",
          8105 => x"54",
          8106 => x"53",
          8107 => x"33",
          8108 => x"94",
          8109 => x"b3",
          8110 => x"2e",
          8111 => x"e2",
          8112 => x"3d",
          8113 => x"3d",
          8114 => x"96",
          8115 => x"fe",
          8116 => x"81",
          8117 => x"ba",
          8118 => x"b0",
          8119 => x"b2",
          8120 => x"fe",
          8121 => x"72",
          8122 => x"81",
          8123 => x"71",
          8124 => x"38",
          8125 => x"d9",
          8126 => x"82",
          8127 => x"db",
          8128 => x"51",
          8129 => x"3f",
          8130 => x"70",
          8131 => x"52",
          8132 => x"95",
          8133 => x"fe",
          8134 => x"82",
          8135 => x"fe",
          8136 => x"80",
          8137 => x"ea",
          8138 => x"2a",
          8139 => x"51",
          8140 => x"2e",
          8141 => x"51",
          8142 => x"3f",
          8143 => x"51",
          8144 => x"3f",
          8145 => x"d8",
          8146 => x"84",
          8147 => x"06",
          8148 => x"80",
          8149 => x"81",
          8150 => x"b6",
          8151 => x"80",
          8152 => x"ae",
          8153 => x"fe",
          8154 => x"72",
          8155 => x"81",
          8156 => x"71",
          8157 => x"38",
          8158 => x"d8",
          8159 => x"83",
          8160 => x"da",
          8161 => x"51",
          8162 => x"3f",
          8163 => x"70",
          8164 => x"52",
          8165 => x"95",
          8166 => x"fe",
          8167 => x"82",
          8168 => x"fe",
          8169 => x"80",
          8170 => x"e6",
          8171 => x"2a",
          8172 => x"51",
          8173 => x"2e",
          8174 => x"51",
          8175 => x"3f",
          8176 => x"51",
          8177 => x"3f",
          8178 => x"d7",
          8179 => x"88",
          8180 => x"06",
          8181 => x"80",
          8182 => x"81",
          8183 => x"b2",
          8184 => x"d0",
          8185 => x"aa",
          8186 => x"fe",
          8187 => x"fe",
          8188 => x"84",
          8189 => x"fb",
          8190 => x"02",
          8191 => x"05",
          8192 => x"56",
          8193 => x"75",
          8194 => x"e2",
          8195 => x"c8",
          8196 => x"a7",
          8197 => x"82",
          8198 => x"82",
          8199 => x"ff",
          8200 => x"82",
          8201 => x"30",
          8202 => x"dc",
          8203 => x"25",
          8204 => x"51",
          8205 => x"82",
          8206 => x"82",
          8207 => x"54",
          8208 => x"09",
          8209 => x"38",
          8210 => x"53",
          8211 => x"51",
          8212 => x"82",
          8213 => x"80",
          8214 => x"82",
          8215 => x"51",
          8216 => x"3f",
          8217 => x"a3",
          8218 => x"aa",
          8219 => x"82",
          8220 => x"82",
          8221 => x"54",
          8222 => x"09",
          8223 => x"38",
          8224 => x"51",
          8225 => x"3f",
          8226 => x"8c",
          8227 => x"3d",
          8228 => x"3d",
          8229 => x"71",
          8230 => x"0c",
          8231 => x"52",
          8232 => x"86",
          8233 => x"8c",
          8234 => x"ff",
          8235 => x"7d",
          8236 => x"06",
          8237 => x"84",
          8238 => x"3d",
          8239 => x"fe",
          8240 => x"7c",
          8241 => x"82",
          8242 => x"ff",
          8243 => x"82",
          8244 => x"7d",
          8245 => x"82",
          8246 => x"8d",
          8247 => x"70",
          8248 => x"84",
          8249 => x"e8",
          8250 => x"3d",
          8251 => x"80",
          8252 => x"51",
          8253 => x"b4",
          8254 => x"05",
          8255 => x"3f",
          8256 => x"08",
          8257 => x"90",
          8258 => x"78",
          8259 => x"87",
          8260 => x"80",
          8261 => x"38",
          8262 => x"81",
          8263 => x"bd",
          8264 => x"78",
          8265 => x"ba",
          8266 => x"2e",
          8267 => x"8a",
          8268 => x"80",
          8269 => x"a1",
          8270 => x"c0",
          8271 => x"38",
          8272 => x"82",
          8273 => x"d2",
          8274 => x"f9",
          8275 => x"38",
          8276 => x"24",
          8277 => x"80",
          8278 => x"98",
          8279 => x"f8",
          8280 => x"38",
          8281 => x"78",
          8282 => x"8a",
          8283 => x"81",
          8284 => x"38",
          8285 => x"2e",
          8286 => x"8a",
          8287 => x"81",
          8288 => x"8f",
          8289 => x"39",
          8290 => x"80",
          8291 => x"84",
          8292 => x"ee",
          8293 => x"8c",
          8294 => x"2e",
          8295 => x"b4",
          8296 => x"11",
          8297 => x"05",
          8298 => x"b4",
          8299 => x"dc",
          8300 => x"fe",
          8301 => x"3d",
          8302 => x"53",
          8303 => x"51",
          8304 => x"3f",
          8305 => x"08",
          8306 => x"8c",
          8307 => x"82",
          8308 => x"fe",
          8309 => x"63",
          8310 => x"79",
          8311 => x"f2",
          8312 => x"78",
          8313 => x"05",
          8314 => x"7a",
          8315 => x"81",
          8316 => x"3d",
          8317 => x"53",
          8318 => x"51",
          8319 => x"3f",
          8320 => x"08",
          8321 => x"da",
          8322 => x"fe",
          8323 => x"ff",
          8324 => x"fe",
          8325 => x"82",
          8326 => x"80",
          8327 => x"38",
          8328 => x"f8",
          8329 => x"84",
          8330 => x"ed",
          8331 => x"8c",
          8332 => x"2e",
          8333 => x"82",
          8334 => x"fe",
          8335 => x"63",
          8336 => x"27",
          8337 => x"61",
          8338 => x"81",
          8339 => x"79",
          8340 => x"05",
          8341 => x"b4",
          8342 => x"11",
          8343 => x"05",
          8344 => x"fc",
          8345 => x"dc",
          8346 => x"fc",
          8347 => x"3d",
          8348 => x"53",
          8349 => x"51",
          8350 => x"3f",
          8351 => x"08",
          8352 => x"de",
          8353 => x"fe",
          8354 => x"ff",
          8355 => x"fe",
          8356 => x"82",
          8357 => x"80",
          8358 => x"38",
          8359 => x"51",
          8360 => x"3f",
          8361 => x"63",
          8362 => x"61",
          8363 => x"33",
          8364 => x"78",
          8365 => x"38",
          8366 => x"54",
          8367 => x"79",
          8368 => x"8c",
          8369 => x"a3",
          8370 => x"62",
          8371 => x"5a",
          8372 => x"85",
          8373 => x"bd",
          8374 => x"ff",
          8375 => x"ff",
          8376 => x"fe",
          8377 => x"82",
          8378 => x"80",
          8379 => x"88",
          8380 => x"78",
          8381 => x"38",
          8382 => x"08",
          8383 => x"39",
          8384 => x"33",
          8385 => x"2e",
          8386 => x"87",
          8387 => x"bc",
          8388 => x"a2",
          8389 => x"80",
          8390 => x"82",
          8391 => x"44",
          8392 => x"88",
          8393 => x"78",
          8394 => x"38",
          8395 => x"08",
          8396 => x"82",
          8397 => x"59",
          8398 => x"88",
          8399 => x"f8",
          8400 => x"39",
          8401 => x"08",
          8402 => x"44",
          8403 => x"fc",
          8404 => x"84",
          8405 => x"eb",
          8406 => x"8c",
          8407 => x"de",
          8408 => x"a0",
          8409 => x"80",
          8410 => x"82",
          8411 => x"43",
          8412 => x"82",
          8413 => x"59",
          8414 => x"88",
          8415 => x"e4",
          8416 => x"39",
          8417 => x"33",
          8418 => x"2e",
          8419 => x"87",
          8420 => x"aa",
          8421 => x"a3",
          8422 => x"80",
          8423 => x"82",
          8424 => x"43",
          8425 => x"88",
          8426 => x"78",
          8427 => x"38",
          8428 => x"08",
          8429 => x"82",
          8430 => x"88",
          8431 => x"3d",
          8432 => x"53",
          8433 => x"51",
          8434 => x"3f",
          8435 => x"08",
          8436 => x"38",
          8437 => x"5c",
          8438 => x"83",
          8439 => x"7a",
          8440 => x"30",
          8441 => x"9f",
          8442 => x"06",
          8443 => x"5a",
          8444 => x"88",
          8445 => x"2e",
          8446 => x"42",
          8447 => x"51",
          8448 => x"3f",
          8449 => x"54",
          8450 => x"52",
          8451 => x"91",
          8452 => x"b8",
          8453 => x"ef",
          8454 => x"39",
          8455 => x"80",
          8456 => x"84",
          8457 => x"e9",
          8458 => x"8c",
          8459 => x"2e",
          8460 => x"b4",
          8461 => x"11",
          8462 => x"05",
          8463 => x"a0",
          8464 => x"dc",
          8465 => x"a5",
          8466 => x"02",
          8467 => x"33",
          8468 => x"81",
          8469 => x"3d",
          8470 => x"53",
          8471 => x"51",
          8472 => x"3f",
          8473 => x"08",
          8474 => x"f6",
          8475 => x"33",
          8476 => x"85",
          8477 => x"e6",
          8478 => x"f8",
          8479 => x"fe",
          8480 => x"79",
          8481 => x"59",
          8482 => x"f8",
          8483 => x"79",
          8484 => x"b4",
          8485 => x"11",
          8486 => x"05",
          8487 => x"c0",
          8488 => x"dc",
          8489 => x"91",
          8490 => x"02",
          8491 => x"33",
          8492 => x"81",
          8493 => x"b5",
          8494 => x"d0",
          8495 => x"c7",
          8496 => x"39",
          8497 => x"f4",
          8498 => x"84",
          8499 => x"ea",
          8500 => x"8c",
          8501 => x"2e",
          8502 => x"b4",
          8503 => x"11",
          8504 => x"05",
          8505 => x"ea",
          8506 => x"dc",
          8507 => x"a6",
          8508 => x"02",
          8509 => x"79",
          8510 => x"5b",
          8511 => x"b4",
          8512 => x"11",
          8513 => x"05",
          8514 => x"c6",
          8515 => x"dc",
          8516 => x"f7",
          8517 => x"70",
          8518 => x"82",
          8519 => x"fe",
          8520 => x"80",
          8521 => x"51",
          8522 => x"3f",
          8523 => x"33",
          8524 => x"2e",
          8525 => x"78",
          8526 => x"38",
          8527 => x"41",
          8528 => x"3d",
          8529 => x"53",
          8530 => x"51",
          8531 => x"3f",
          8532 => x"08",
          8533 => x"38",
          8534 => x"be",
          8535 => x"70",
          8536 => x"23",
          8537 => x"ae",
          8538 => x"d0",
          8539 => x"97",
          8540 => x"39",
          8541 => x"f4",
          8542 => x"84",
          8543 => x"e8",
          8544 => x"8c",
          8545 => x"2e",
          8546 => x"b4",
          8547 => x"11",
          8548 => x"05",
          8549 => x"ba",
          8550 => x"dc",
          8551 => x"a1",
          8552 => x"71",
          8553 => x"84",
          8554 => x"3d",
          8555 => x"53",
          8556 => x"51",
          8557 => x"3f",
          8558 => x"08",
          8559 => x"a2",
          8560 => x"08",
          8561 => x"85",
          8562 => x"e4",
          8563 => x"f8",
          8564 => x"fe",
          8565 => x"79",
          8566 => x"59",
          8567 => x"f6",
          8568 => x"79",
          8569 => x"b4",
          8570 => x"11",
          8571 => x"05",
          8572 => x"de",
          8573 => x"dc",
          8574 => x"8d",
          8575 => x"71",
          8576 => x"84",
          8577 => x"b9",
          8578 => x"d0",
          8579 => x"f7",
          8580 => x"39",
          8581 => x"80",
          8582 => x"84",
          8583 => x"e5",
          8584 => x"8c",
          8585 => x"2e",
          8586 => x"63",
          8587 => x"f0",
          8588 => x"b7",
          8589 => x"78",
          8590 => x"ff",
          8591 => x"ff",
          8592 => x"fe",
          8593 => x"82",
          8594 => x"80",
          8595 => x"38",
          8596 => x"86",
          8597 => x"e3",
          8598 => x"59",
          8599 => x"8c",
          8600 => x"2e",
          8601 => x"82",
          8602 => x"52",
          8603 => x"51",
          8604 => x"3f",
          8605 => x"82",
          8606 => x"fe",
          8607 => x"fe",
          8608 => x"f4",
          8609 => x"86",
          8610 => x"dc",
          8611 => x"59",
          8612 => x"fe",
          8613 => x"f4",
          8614 => x"45",
          8615 => x"78",
          8616 => x"be",
          8617 => x"06",
          8618 => x"2e",
          8619 => x"b4",
          8620 => x"05",
          8621 => x"8b",
          8622 => x"dc",
          8623 => x"5b",
          8624 => x"b2",
          8625 => x"24",
          8626 => x"81",
          8627 => x"80",
          8628 => x"83",
          8629 => x"80",
          8630 => x"86",
          8631 => x"55",
          8632 => x"54",
          8633 => x"86",
          8634 => x"3d",
          8635 => x"51",
          8636 => x"3f",
          8637 => x"87",
          8638 => x"3d",
          8639 => x"51",
          8640 => x"3f",
          8641 => x"55",
          8642 => x"54",
          8643 => x"87",
          8644 => x"3d",
          8645 => x"51",
          8646 => x"3f",
          8647 => x"54",
          8648 => x"87",
          8649 => x"3d",
          8650 => x"51",
          8651 => x"3f",
          8652 => x"58",
          8653 => x"57",
          8654 => x"55",
          8655 => x"80",
          8656 => x"80",
          8657 => x"3d",
          8658 => x"51",
          8659 => x"82",
          8660 => x"82",
          8661 => x"09",
          8662 => x"72",
          8663 => x"51",
          8664 => x"80",
          8665 => x"26",
          8666 => x"5a",
          8667 => x"59",
          8668 => x"8d",
          8669 => x"70",
          8670 => x"5c",
          8671 => x"c0",
          8672 => x"32",
          8673 => x"07",
          8674 => x"38",
          8675 => x"09",
          8676 => x"ce",
          8677 => x"a0",
          8678 => x"cf",
          8679 => x"39",
          8680 => x"80",
          8681 => x"a4",
          8682 => x"94",
          8683 => x"54",
          8684 => x"80",
          8685 => x"fe",
          8686 => x"82",
          8687 => x"90",
          8688 => x"55",
          8689 => x"80",
          8690 => x"fe",
          8691 => x"72",
          8692 => x"08",
          8693 => x"87",
          8694 => x"70",
          8695 => x"87",
          8696 => x"72",
          8697 => x"f3",
          8698 => x"dc",
          8699 => x"75",
          8700 => x"87",
          8701 => x"73",
          8702 => x"df",
          8703 => x"8c",
          8704 => x"75",
          8705 => x"83",
          8706 => x"94",
          8707 => x"80",
          8708 => x"c0",
          8709 => x"b7",
          8710 => x"8c",
          8711 => x"ad",
          8712 => x"f4",
          8713 => x"ae",
          8714 => x"d7",
          8715 => x"b0",
          8716 => x"d3",
          8717 => x"bc",
          8718 => x"cb",
          8719 => x"c6",
          8720 => x"ba",
          8721 => x"ec",
          8722 => x"c6",
          8723 => x"00",
          8724 => x"55",
          8725 => x"5b",
          8726 => x"61",
          8727 => x"67",
          8728 => x"6d",
          8729 => x"d8",
          8730 => x"b4",
          8731 => x"57",
          8732 => x"97",
          8733 => x"ba",
          8734 => x"47",
          8735 => x"ad",
          8736 => x"ad",
          8737 => x"84",
          8738 => x"fa",
          8739 => x"85",
          8740 => x"ae",
          8741 => x"cc",
          8742 => x"50",
          8743 => x"57",
          8744 => x"5e",
          8745 => x"65",
          8746 => x"6c",
          8747 => x"73",
          8748 => x"7a",
          8749 => x"81",
          8750 => x"88",
          8751 => x"8f",
          8752 => x"96",
          8753 => x"9c",
          8754 => x"a2",
          8755 => x"a8",
          8756 => x"ae",
          8757 => x"b4",
          8758 => x"ba",
          8759 => x"c0",
          8760 => x"c6",
          8761 => x"25",
          8762 => x"64",
          8763 => x"3a",
          8764 => x"25",
          8765 => x"64",
          8766 => x"00",
          8767 => x"20",
          8768 => x"66",
          8769 => x"72",
          8770 => x"6f",
          8771 => x"00",
          8772 => x"72",
          8773 => x"53",
          8774 => x"63",
          8775 => x"69",
          8776 => x"00",
          8777 => x"65",
          8778 => x"65",
          8779 => x"6d",
          8780 => x"6d",
          8781 => x"65",
          8782 => x"00",
          8783 => x"20",
          8784 => x"53",
          8785 => x"4d",
          8786 => x"25",
          8787 => x"3a",
          8788 => x"58",
          8789 => x"00",
          8790 => x"20",
          8791 => x"41",
          8792 => x"20",
          8793 => x"25",
          8794 => x"3a",
          8795 => x"58",
          8796 => x"00",
          8797 => x"20",
          8798 => x"4e",
          8799 => x"41",
          8800 => x"25",
          8801 => x"3a",
          8802 => x"58",
          8803 => x"00",
          8804 => x"20",
          8805 => x"4d",
          8806 => x"20",
          8807 => x"25",
          8808 => x"3a",
          8809 => x"58",
          8810 => x"00",
          8811 => x"20",
          8812 => x"20",
          8813 => x"20",
          8814 => x"25",
          8815 => x"3a",
          8816 => x"58",
          8817 => x"00",
          8818 => x"20",
          8819 => x"43",
          8820 => x"20",
          8821 => x"44",
          8822 => x"63",
          8823 => x"3d",
          8824 => x"64",
          8825 => x"00",
          8826 => x"20",
          8827 => x"45",
          8828 => x"20",
          8829 => x"54",
          8830 => x"72",
          8831 => x"3d",
          8832 => x"64",
          8833 => x"00",
          8834 => x"20",
          8835 => x"52",
          8836 => x"52",
          8837 => x"43",
          8838 => x"6e",
          8839 => x"3d",
          8840 => x"64",
          8841 => x"00",
          8842 => x"20",
          8843 => x"48",
          8844 => x"45",
          8845 => x"53",
          8846 => x"00",
          8847 => x"20",
          8848 => x"49",
          8849 => x"00",
          8850 => x"20",
          8851 => x"54",
          8852 => x"00",
          8853 => x"20",
          8854 => x"0a",
          8855 => x"00",
          8856 => x"20",
          8857 => x"0a",
          8858 => x"00",
          8859 => x"72",
          8860 => x"65",
          8861 => x"00",
          8862 => x"20",
          8863 => x"20",
          8864 => x"65",
          8865 => x"65",
          8866 => x"72",
          8867 => x"64",
          8868 => x"73",
          8869 => x"25",
          8870 => x"0a",
          8871 => x"00",
          8872 => x"20",
          8873 => x"20",
          8874 => x"6f",
          8875 => x"53",
          8876 => x"74",
          8877 => x"64",
          8878 => x"73",
          8879 => x"25",
          8880 => x"0a",
          8881 => x"00",
          8882 => x"20",
          8883 => x"63",
          8884 => x"74",
          8885 => x"20",
          8886 => x"72",
          8887 => x"20",
          8888 => x"20",
          8889 => x"25",
          8890 => x"0a",
          8891 => x"00",
          8892 => x"63",
          8893 => x"00",
          8894 => x"20",
          8895 => x"20",
          8896 => x"20",
          8897 => x"20",
          8898 => x"20",
          8899 => x"20",
          8900 => x"20",
          8901 => x"25",
          8902 => x"0a",
          8903 => x"00",
          8904 => x"20",
          8905 => x"74",
          8906 => x"43",
          8907 => x"6b",
          8908 => x"65",
          8909 => x"20",
          8910 => x"20",
          8911 => x"25",
          8912 => x"30",
          8913 => x"48",
          8914 => x"00",
          8915 => x"20",
          8916 => x"41",
          8917 => x"6c",
          8918 => x"20",
          8919 => x"71",
          8920 => x"20",
          8921 => x"20",
          8922 => x"25",
          8923 => x"30",
          8924 => x"48",
          8925 => x"00",
          8926 => x"20",
          8927 => x"68",
          8928 => x"65",
          8929 => x"52",
          8930 => x"43",
          8931 => x"6b",
          8932 => x"65",
          8933 => x"25",
          8934 => x"30",
          8935 => x"48",
          8936 => x"00",
          8937 => x"6c",
          8938 => x"00",
          8939 => x"69",
          8940 => x"00",
          8941 => x"78",
          8942 => x"00",
          8943 => x"00",
          8944 => x"6d",
          8945 => x"00",
          8946 => x"6e",
          8947 => x"00",
          8948 => x"74",
          8949 => x"2e",
          8950 => x"00",
          8951 => x"74",
          8952 => x"00",
          8953 => x"74",
          8954 => x"00",
          8955 => x"00",
          8956 => x"64",
          8957 => x"73",
          8958 => x"00",
          8959 => x"6c",
          8960 => x"74",
          8961 => x"65",
          8962 => x"20",
          8963 => x"20",
          8964 => x"74",
          8965 => x"20",
          8966 => x"65",
          8967 => x"20",
          8968 => x"2e",
          8969 => x"00",
          8970 => x"6e",
          8971 => x"6f",
          8972 => x"2f",
          8973 => x"61",
          8974 => x"68",
          8975 => x"6f",
          8976 => x"66",
          8977 => x"2c",
          8978 => x"73",
          8979 => x"69",
          8980 => x"0a",
          8981 => x"00",
          8982 => x"04",
          8983 => x"00",
          8984 => x"01",
          8985 => x"00",
          8986 => x"00",
          8987 => x"02",
          8988 => x"fc",
          8989 => x"00",
          8990 => x"03",
          8991 => x"f8",
          8992 => x"00",
          8993 => x"04",
          8994 => x"f4",
          8995 => x"00",
          8996 => x"05",
          8997 => x"f0",
          8998 => x"00",
          8999 => x"06",
          9000 => x"ec",
          9001 => x"00",
          9002 => x"07",
          9003 => x"e8",
          9004 => x"00",
          9005 => x"08",
          9006 => x"e4",
          9007 => x"00",
          9008 => x"09",
          9009 => x"e0",
          9010 => x"00",
          9011 => x"0a",
          9012 => x"dc",
          9013 => x"00",
          9014 => x"0b",
          9015 => x"00",
          9016 => x"00",
          9017 => x"00",
          9018 => x"00",
          9019 => x"7e",
          9020 => x"7e",
          9021 => x"7e",
          9022 => x"7e",
          9023 => x"7e",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"2c",
          9028 => x"3d",
          9029 => x"5d",
          9030 => x"00",
          9031 => x"00",
          9032 => x"33",
          9033 => x"00",
          9034 => x"4d",
          9035 => x"53",
          9036 => x"00",
          9037 => x"4e",
          9038 => x"20",
          9039 => x"46",
          9040 => x"32",
          9041 => x"00",
          9042 => x"4e",
          9043 => x"20",
          9044 => x"46",
          9045 => x"20",
          9046 => x"00",
          9047 => x"08",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"41",
          9052 => x"80",
          9053 => x"49",
          9054 => x"8f",
          9055 => x"4f",
          9056 => x"55",
          9057 => x"9b",
          9058 => x"9f",
          9059 => x"55",
          9060 => x"a7",
          9061 => x"ab",
          9062 => x"af",
          9063 => x"b3",
          9064 => x"b7",
          9065 => x"bb",
          9066 => x"bf",
          9067 => x"c3",
          9068 => x"c7",
          9069 => x"cb",
          9070 => x"cf",
          9071 => x"d3",
          9072 => x"d7",
          9073 => x"db",
          9074 => x"df",
          9075 => x"e3",
          9076 => x"e7",
          9077 => x"eb",
          9078 => x"ef",
          9079 => x"f3",
          9080 => x"f7",
          9081 => x"fb",
          9082 => x"ff",
          9083 => x"3b",
          9084 => x"2f",
          9085 => x"3a",
          9086 => x"7c",
          9087 => x"00",
          9088 => x"04",
          9089 => x"40",
          9090 => x"00",
          9091 => x"00",
          9092 => x"02",
          9093 => x"08",
          9094 => x"20",
          9095 => x"00",
          9096 => x"69",
          9097 => x"00",
          9098 => x"63",
          9099 => x"00",
          9100 => x"69",
          9101 => x"00",
          9102 => x"61",
          9103 => x"00",
          9104 => x"65",
          9105 => x"00",
          9106 => x"65",
          9107 => x"00",
          9108 => x"70",
          9109 => x"00",
          9110 => x"66",
          9111 => x"00",
          9112 => x"6d",
          9113 => x"00",
          9114 => x"00",
          9115 => x"00",
          9116 => x"00",
          9117 => x"00",
          9118 => x"00",
          9119 => x"00",
          9120 => x"00",
          9121 => x"6c",
          9122 => x"00",
          9123 => x"00",
          9124 => x"74",
          9125 => x"00",
          9126 => x"65",
          9127 => x"00",
          9128 => x"6f",
          9129 => x"00",
          9130 => x"74",
          9131 => x"00",
          9132 => x"73",
          9133 => x"00",
          9134 => x"73",
          9135 => x"00",
          9136 => x"6f",
          9137 => x"00",
          9138 => x"6b",
          9139 => x"72",
          9140 => x"00",
          9141 => x"65",
          9142 => x"6c",
          9143 => x"72",
          9144 => x"0a",
          9145 => x"00",
          9146 => x"6b",
          9147 => x"74",
          9148 => x"61",
          9149 => x"0a",
          9150 => x"00",
          9151 => x"66",
          9152 => x"20",
          9153 => x"6e",
          9154 => x"00",
          9155 => x"70",
          9156 => x"20",
          9157 => x"6e",
          9158 => x"00",
          9159 => x"61",
          9160 => x"20",
          9161 => x"65",
          9162 => x"65",
          9163 => x"00",
          9164 => x"65",
          9165 => x"64",
          9166 => x"65",
          9167 => x"00",
          9168 => x"65",
          9169 => x"72",
          9170 => x"79",
          9171 => x"69",
          9172 => x"2e",
          9173 => x"00",
          9174 => x"65",
          9175 => x"6e",
          9176 => x"20",
          9177 => x"61",
          9178 => x"2e",
          9179 => x"00",
          9180 => x"69",
          9181 => x"72",
          9182 => x"20",
          9183 => x"74",
          9184 => x"65",
          9185 => x"00",
          9186 => x"76",
          9187 => x"75",
          9188 => x"72",
          9189 => x"20",
          9190 => x"61",
          9191 => x"2e",
          9192 => x"00",
          9193 => x"6b",
          9194 => x"74",
          9195 => x"61",
          9196 => x"64",
          9197 => x"00",
          9198 => x"63",
          9199 => x"61",
          9200 => x"6c",
          9201 => x"69",
          9202 => x"79",
          9203 => x"6d",
          9204 => x"75",
          9205 => x"6f",
          9206 => x"69",
          9207 => x"0a",
          9208 => x"00",
          9209 => x"6d",
          9210 => x"61",
          9211 => x"74",
          9212 => x"0a",
          9213 => x"00",
          9214 => x"65",
          9215 => x"2c",
          9216 => x"65",
          9217 => x"69",
          9218 => x"63",
          9219 => x"65",
          9220 => x"64",
          9221 => x"00",
          9222 => x"65",
          9223 => x"20",
          9224 => x"6b",
          9225 => x"0a",
          9226 => x"00",
          9227 => x"75",
          9228 => x"63",
          9229 => x"74",
          9230 => x"6d",
          9231 => x"2e",
          9232 => x"00",
          9233 => x"20",
          9234 => x"79",
          9235 => x"65",
          9236 => x"69",
          9237 => x"2e",
          9238 => x"00",
          9239 => x"61",
          9240 => x"65",
          9241 => x"69",
          9242 => x"72",
          9243 => x"74",
          9244 => x"00",
          9245 => x"63",
          9246 => x"2e",
          9247 => x"00",
          9248 => x"6e",
          9249 => x"20",
          9250 => x"6f",
          9251 => x"00",
          9252 => x"75",
          9253 => x"74",
          9254 => x"25",
          9255 => x"74",
          9256 => x"75",
          9257 => x"74",
          9258 => x"73",
          9259 => x"0a",
          9260 => x"00",
          9261 => x"64",
          9262 => x"00",
          9263 => x"58",
          9264 => x"00",
          9265 => x"00",
          9266 => x"58",
          9267 => x"00",
          9268 => x"20",
          9269 => x"20",
          9270 => x"00",
          9271 => x"58",
          9272 => x"00",
          9273 => x"00",
          9274 => x"00",
          9275 => x"00",
          9276 => x"00",
          9277 => x"20",
          9278 => x"28",
          9279 => x"00",
          9280 => x"30",
          9281 => x"30",
          9282 => x"00",
          9283 => x"30",
          9284 => x"00",
          9285 => x"55",
          9286 => x"65",
          9287 => x"30",
          9288 => x"20",
          9289 => x"25",
          9290 => x"2a",
          9291 => x"00",
          9292 => x"20",
          9293 => x"65",
          9294 => x"70",
          9295 => x"61",
          9296 => x"65",
          9297 => x"00",
          9298 => x"65",
          9299 => x"6e",
          9300 => x"72",
          9301 => x"0a",
          9302 => x"00",
          9303 => x"20",
          9304 => x"65",
          9305 => x"70",
          9306 => x"00",
          9307 => x"54",
          9308 => x"44",
          9309 => x"74",
          9310 => x"75",
          9311 => x"00",
          9312 => x"54",
          9313 => x"52",
          9314 => x"74",
          9315 => x"75",
          9316 => x"00",
          9317 => x"54",
          9318 => x"58",
          9319 => x"74",
          9320 => x"75",
          9321 => x"00",
          9322 => x"54",
          9323 => x"58",
          9324 => x"74",
          9325 => x"75",
          9326 => x"00",
          9327 => x"54",
          9328 => x"58",
          9329 => x"74",
          9330 => x"75",
          9331 => x"00",
          9332 => x"54",
          9333 => x"58",
          9334 => x"74",
          9335 => x"75",
          9336 => x"00",
          9337 => x"74",
          9338 => x"20",
          9339 => x"74",
          9340 => x"72",
          9341 => x"0a",
          9342 => x"00",
          9343 => x"62",
          9344 => x"67",
          9345 => x"6d",
          9346 => x"2e",
          9347 => x"00",
          9348 => x"6f",
          9349 => x"63",
          9350 => x"74",
          9351 => x"00",
          9352 => x"00",
          9353 => x"6c",
          9354 => x"74",
          9355 => x"6e",
          9356 => x"61",
          9357 => x"65",
          9358 => x"20",
          9359 => x"64",
          9360 => x"20",
          9361 => x"61",
          9362 => x"69",
          9363 => x"20",
          9364 => x"75",
          9365 => x"79",
          9366 => x"00",
          9367 => x"00",
          9368 => x"61",
          9369 => x"67",
          9370 => x"2e",
          9371 => x"00",
          9372 => x"79",
          9373 => x"2e",
          9374 => x"00",
          9375 => x"70",
          9376 => x"6e",
          9377 => x"2e",
          9378 => x"00",
          9379 => x"6c",
          9380 => x"30",
          9381 => x"2d",
          9382 => x"38",
          9383 => x"25",
          9384 => x"29",
          9385 => x"00",
          9386 => x"70",
          9387 => x"6d",
          9388 => x"0a",
          9389 => x"00",
          9390 => x"6d",
          9391 => x"74",
          9392 => x"00",
          9393 => x"58",
          9394 => x"32",
          9395 => x"00",
          9396 => x"0a",
          9397 => x"00",
          9398 => x"58",
          9399 => x"34",
          9400 => x"00",
          9401 => x"58",
          9402 => x"38",
          9403 => x"00",
          9404 => x"63",
          9405 => x"6e",
          9406 => x"6f",
          9407 => x"40",
          9408 => x"38",
          9409 => x"2e",
          9410 => x"00",
          9411 => x"6c",
          9412 => x"20",
          9413 => x"65",
          9414 => x"25",
          9415 => x"20",
          9416 => x"0a",
          9417 => x"00",
          9418 => x"6c",
          9419 => x"74",
          9420 => x"65",
          9421 => x"6f",
          9422 => x"28",
          9423 => x"2e",
          9424 => x"00",
          9425 => x"74",
          9426 => x"69",
          9427 => x"61",
          9428 => x"69",
          9429 => x"69",
          9430 => x"2e",
          9431 => x"00",
          9432 => x"64",
          9433 => x"62",
          9434 => x"69",
          9435 => x"2e",
          9436 => x"00",
          9437 => x"00",
          9438 => x"00",
          9439 => x"5c",
          9440 => x"25",
          9441 => x"73",
          9442 => x"00",
          9443 => x"5c",
          9444 => x"25",
          9445 => x"00",
          9446 => x"5c",
          9447 => x"00",
          9448 => x"20",
          9449 => x"6d",
          9450 => x"2e",
          9451 => x"00",
          9452 => x"6e",
          9453 => x"2e",
          9454 => x"00",
          9455 => x"62",
          9456 => x"67",
          9457 => x"74",
          9458 => x"75",
          9459 => x"2e",
          9460 => x"00",
          9461 => x"00",
          9462 => x"00",
          9463 => x"ff",
          9464 => x"00",
          9465 => x"ff",
          9466 => x"00",
          9467 => x"ff",
          9468 => x"00",
          9469 => x"00",
          9470 => x"00",
          9471 => x"ff",
          9472 => x"00",
          9473 => x"00",
          9474 => x"00",
          9475 => x"00",
          9476 => x"00",
          9477 => x"00",
          9478 => x"00",
          9479 => x"00",
          9480 => x"01",
          9481 => x"01",
          9482 => x"01",
          9483 => x"00",
          9484 => x"00",
          9485 => x"02",
          9486 => x"00",
          9487 => x"34",
          9488 => x"34",
          9489 => x"34",
          9490 => x"34",
          9491 => x"d0",
          9492 => x"00",
          9493 => x"00",
          9494 => x"00",
          9495 => x"00",
          9496 => x"00",
          9497 => x"00",
          9498 => x"00",
          9499 => x"00",
          9500 => x"00",
          9501 => x"00",
          9502 => x"00",
          9503 => x"00",
          9504 => x"00",
          9505 => x"00",
          9506 => x"00",
          9507 => x"00",
          9508 => x"00",
          9509 => x"00",
          9510 => x"00",
          9511 => x"00",
          9512 => x"00",
          9513 => x"00",
          9514 => x"00",
          9515 => x"dc",
          9516 => x"00",
          9517 => x"e4",
          9518 => x"00",
          9519 => x"ec",
          9520 => x"00",
          9521 => x"00",
          9522 => x"00",
          9523 => x"20",
          9524 => x"00",
          9525 => x"00",
          9526 => x"00",
          9527 => x"28",
          9528 => x"00",
          9529 => x"00",
          9530 => x"00",
          9531 => x"30",
          9532 => x"00",
          9533 => x"00",
          9534 => x"00",
          9535 => x"38",
          9536 => x"00",
          9537 => x"00",
          9538 => x"00",
          9539 => x"40",
          9540 => x"00",
          9541 => x"00",
          9542 => x"00",
          9543 => x"48",
          9544 => x"00",
          9545 => x"00",
          9546 => x"00",
          9547 => x"50",
          9548 => x"00",
          9549 => x"00",
          9550 => x"00",
          9551 => x"58",
          9552 => x"00",
          9553 => x"00",
          9554 => x"00",
          9555 => x"60",
          9556 => x"00",
          9557 => x"00",
          9558 => x"00",
          9559 => x"68",
          9560 => x"00",
          9561 => x"00",
          9562 => x"00",
          9563 => x"6c",
          9564 => x"00",
          9565 => x"00",
          9566 => x"00",
          9567 => x"70",
          9568 => x"00",
          9569 => x"00",
          9570 => x"00",
          9571 => x"74",
          9572 => x"00",
          9573 => x"00",
          9574 => x"00",
          9575 => x"78",
          9576 => x"00",
          9577 => x"00",
          9578 => x"00",
          9579 => x"7c",
          9580 => x"00",
          9581 => x"00",
          9582 => x"00",
          9583 => x"80",
          9584 => x"00",
          9585 => x"00",
          9586 => x"00",
          9587 => x"84",
          9588 => x"00",
          9589 => x"00",
          9590 => x"00",
          9591 => x"8c",
          9592 => x"00",
          9593 => x"00",
          9594 => x"00",
          9595 => x"90",
          9596 => x"00",
          9597 => x"00",
          9598 => x"00",
          9599 => x"98",
          9600 => x"00",
          9601 => x"00",
          9602 => x"00",
          9603 => x"a0",
          9604 => x"00",
          9605 => x"00",
          9606 => x"00",
          9607 => x"a8",
          9608 => x"00",
          9609 => x"00",
          9610 => x"00",
          9611 => x"b0",
          9612 => x"00",
          9613 => x"00",
          9614 => x"00",
          9615 => x"b8",
          9616 => x"00",
          9617 => x"00",
          9618 => x"00",
          9619 => x"c0",
          9620 => x"00",
          9621 => x"00",
          9622 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"70",
           281 => x"8e",
           282 => x"70",
           283 => x"0c",
           284 => x"88",
           285 => x"fe",
           286 => x"04",
           287 => x"00",
           288 => x"00",
           289 => x"08",
           290 => x"fd",
           291 => x"53",
           292 => x"05",
           293 => x"08",
           294 => x"51",
           295 => x"88",
           296 => x"0c",
           297 => x"0d",
           298 => x"94",
           299 => x"0c",
           300 => x"81",
           301 => x"8c",
           302 => x"94",
           303 => x"08",
           304 => x"3f",
           305 => x"88",
           306 => x"3d",
           307 => x"04",
           308 => x"94",
           309 => x"0d",
           310 => x"08",
           311 => x"94",
           312 => x"08",
           313 => x"38",
           314 => x"05",
           315 => x"08",
           316 => x"80",
           317 => x"f4",
           318 => x"08",
           319 => x"88",
           320 => x"94",
           321 => x"0c",
           322 => x"05",
           323 => x"fc",
           324 => x"08",
           325 => x"80",
           326 => x"94",
           327 => x"08",
           328 => x"8c",
           329 => x"0b",
           330 => x"05",
           331 => x"fc",
           332 => x"38",
           333 => x"08",
           334 => x"94",
           335 => x"08",
           336 => x"05",
           337 => x"94",
           338 => x"08",
           339 => x"88",
           340 => x"81",
           341 => x"08",
           342 => x"f8",
           343 => x"94",
           344 => x"08",
           345 => x"38",
           346 => x"05",
           347 => x"08",
           348 => x"94",
           349 => x"08",
           350 => x"54",
           351 => x"94",
           352 => x"08",
           353 => x"fb",
           354 => x"0b",
           355 => x"05",
           356 => x"88",
           357 => x"25",
           358 => x"08",
           359 => x"30",
           360 => x"05",
           361 => x"94",
           362 => x"0c",
           363 => x"05",
           364 => x"8c",
           365 => x"8c",
           366 => x"94",
           367 => x"0c",
           368 => x"08",
           369 => x"52",
           370 => x"05",
           371 => x"3f",
           372 => x"94",
           373 => x"0c",
           374 => x"fc",
           375 => x"2e",
           376 => x"08",
           377 => x"30",
           378 => x"05",
           379 => x"f8",
           380 => x"88",
           381 => x"3d",
           382 => x"04",
           383 => x"94",
           384 => x"0d",
           385 => x"08",
           386 => x"80",
           387 => x"f8",
           388 => x"08",
           389 => x"94",
           390 => x"08",
           391 => x"94",
           392 => x"08",
           393 => x"38",
           394 => x"08",
           395 => x"24",
           396 => x"08",
           397 => x"10",
           398 => x"05",
           399 => x"fc",
           400 => x"94",
           401 => x"0c",
           402 => x"08",
           403 => x"80",
           404 => x"38",
           405 => x"05",
           406 => x"88",
           407 => x"a1",
           408 => x"88",
           409 => x"08",
           410 => x"31",
           411 => x"05",
           412 => x"f8",
           413 => x"08",
           414 => x"07",
           415 => x"05",
           416 => x"fc",
           417 => x"2a",
           418 => x"05",
           419 => x"8c",
           420 => x"2a",
           421 => x"05",
           422 => x"39",
           423 => x"05",
           424 => x"8f",
           425 => x"88",
           426 => x"94",
           427 => x"0c",
           428 => x"94",
           429 => x"08",
           430 => x"f4",
           431 => x"94",
           432 => x"08",
           433 => x"3d",
           434 => x"04",
           435 => x"81",
           436 => x"c0",
           437 => x"81",
           438 => x"92",
           439 => x"0b",
           440 => x"8c",
           441 => x"92",
           442 => x"82",
           443 => x"70",
           444 => x"38",
           445 => x"8c",
           446 => x"e9",
           447 => x"92",
           448 => x"80",
           449 => x"71",
           450 => x"c0",
           451 => x"51",
           452 => x"88",
           453 => x"0b",
           454 => x"34",
           455 => x"9f",
           456 => x"0c",
           457 => x"04",
           458 => x"78",
           459 => x"58",
           460 => x"0b",
           461 => x"f0",
           462 => x"52",
           463 => x"70",
           464 => x"81",
           465 => x"38",
           466 => x"c0",
           467 => x"79",
           468 => x"80",
           469 => x"87",
           470 => x"0c",
           471 => x"8c",
           472 => x"2a",
           473 => x"51",
           474 => x"80",
           475 => x"87",
           476 => x"08",
           477 => x"06",
           478 => x"52",
           479 => x"80",
           480 => x"70",
           481 => x"38",
           482 => x"81",
           483 => x"ff",
           484 => x"15",
           485 => x"06",
           486 => x"2e",
           487 => x"c0",
           488 => x"51",
           489 => x"38",
           490 => x"8c",
           491 => x"95",
           492 => x"87",
           493 => x"0c",
           494 => x"8c",
           495 => x"06",
           496 => x"f4",
           497 => x"fc",
           498 => x"52",
           499 => x"2e",
           500 => x"8f",
           501 => x"98",
           502 => x"70",
           503 => x"81",
           504 => x"81",
           505 => x"0c",
           506 => x"04",
           507 => x"74",
           508 => x"71",
           509 => x"2b",
           510 => x"53",
           511 => x"0d",
           512 => x"0d",
           513 => x"33",
           514 => x"71",
           515 => x"88",
           516 => x"14",
           517 => x"07",
           518 => x"33",
           519 => x"0c",
           520 => x"56",
           521 => x"3d",
           522 => x"3d",
           523 => x"0b",
           524 => x"08",
           525 => x"77",
           526 => x"38",
           527 => x"08",
           528 => x"38",
           529 => x"74",
           530 => x"38",
           531 => x"ae",
           532 => x"39",
           533 => x"10",
           534 => x"53",
           535 => x"8c",
           536 => x"52",
           537 => x"52",
           538 => x"3f",
           539 => x"38",
           540 => x"f8",
           541 => x"83",
           542 => x"55",
           543 => x"54",
           544 => x"83",
           545 => x"76",
           546 => x"17",
           547 => x"88",
           548 => x"55",
           549 => x"88",
           550 => x"74",
           551 => x"3f",
           552 => x"0a",
           553 => x"39",
           554 => x"88",
           555 => x"0d",
           556 => x"0d",
           557 => x"9f",
           558 => x"19",
           559 => x"fe",
           560 => x"54",
           561 => x"73",
           562 => x"82",
           563 => x"71",
           564 => x"08",
           565 => x"75",
           566 => x"3d",
           567 => x"3d",
           568 => x"80",
           569 => x"0b",
           570 => x"70",
           571 => x"53",
           572 => x"09",
           573 => x"38",
           574 => x"fd",
           575 => x"08",
           576 => x"9a",
           577 => x"e4",
           578 => x"83",
           579 => x"73",
           580 => x"85",
           581 => x"fc",
           582 => x"0b",
           583 => x"f4",
           584 => x"80",
           585 => x"15",
           586 => x"81",
           587 => x"88",
           588 => x"26",
           589 => x"52",
           590 => x"90",
           591 => x"52",
           592 => x"09",
           593 => x"38",
           594 => x"53",
           595 => x"0c",
           596 => x"8b",
           597 => x"fe",
           598 => x"08",
           599 => x"90",
           600 => x"71",
           601 => x"80",
           602 => x"0c",
           603 => x"04",
           604 => x"78",
           605 => x"9f",
           606 => x"22",
           607 => x"83",
           608 => x"57",
           609 => x"73",
           610 => x"38",
           611 => x"53",
           612 => x"83",
           613 => x"39",
           614 => x"52",
           615 => x"38",
           616 => x"16",
           617 => x"08",
           618 => x"38",
           619 => x"17",
           620 => x"73",
           621 => x"38",
           622 => x"16",
           623 => x"74",
           624 => x"52",
           625 => x"72",
           626 => x"3f",
           627 => x"88",
           628 => x"38",
           629 => x"08",
           630 => x"27",
           631 => x"08",
           632 => x"88",
           633 => x"c9",
           634 => x"90",
           635 => x"75",
           636 => x"71",
           637 => x"3d",
           638 => x"3d",
           639 => x"64",
           640 => x"75",
           641 => x"a0",
           642 => x"06",
           643 => x"16",
           644 => x"ef",
           645 => x"33",
           646 => x"af",
           647 => x"06",
           648 => x"16",
           649 => x"88",
           650 => x"70",
           651 => x"74",
           652 => x"38",
           653 => x"df",
           654 => x"56",
           655 => x"82",
           656 => x"3d",
           657 => x"70",
           658 => x"8a",
           659 => x"70",
           660 => x"34",
           661 => x"74",
           662 => x"81",
           663 => x"80",
           664 => x"88",
           665 => x"5a",
           666 => x"70",
           667 => x"60",
           668 => x"70",
           669 => x"30",
           670 => x"71",
           671 => x"51",
           672 => x"53",
           673 => x"74",
           674 => x"76",
           675 => x"81",
           676 => x"81",
           677 => x"27",
           678 => x"74",
           679 => x"38",
           680 => x"70",
           681 => x"32",
           682 => x"73",
           683 => x"53",
           684 => x"56",
           685 => x"88",
           686 => x"ff",
           687 => x"81",
           688 => x"ff",
           689 => x"53",
           690 => x"76",
           691 => x"98",
           692 => x"7f",
           693 => x"76",
           694 => x"38",
           695 => x"8b",
           696 => x"51",
           697 => x"88",
           698 => x"38",
           699 => x"22",
           700 => x"83",
           701 => x"55",
           702 => x"52",
           703 => x"a8",
           704 => x"57",
           705 => x"fb",
           706 => x"55",
           707 => x"80",
           708 => x"1d",
           709 => x"2a",
           710 => x"51",
           711 => x"b2",
           712 => x"84",
           713 => x"08",
           714 => x"58",
           715 => x"77",
           716 => x"38",
           717 => x"05",
           718 => x"70",
           719 => x"33",
           720 => x"52",
           721 => x"80",
           722 => x"86",
           723 => x"2e",
           724 => x"51",
           725 => x"ff",
           726 => x"08",
           727 => x"b4",
           728 => x"76",
           729 => x"08",
           730 => x"51",
           731 => x"38",
           732 => x"70",
           733 => x"81",
           734 => x"56",
           735 => x"83",
           736 => x"81",
           737 => x"7c",
           738 => x"3f",
           739 => x"1d",
           740 => x"39",
           741 => x"90",
           742 => x"f9",
           743 => x"7b",
           744 => x"54",
           745 => x"77",
           746 => x"f6",
           747 => x"56",
           748 => x"e7",
           749 => x"f8",
           750 => x"08",
           751 => x"06",
           752 => x"74",
           753 => x"2e",
           754 => x"80",
           755 => x"54",
           756 => x"52",
           757 => x"d0",
           758 => x"56",
           759 => x"38",
           760 => x"88",
           761 => x"83",
           762 => x"55",
           763 => x"c6",
           764 => x"82",
           765 => x"53",
           766 => x"51",
           767 => x"88",
           768 => x"08",
           769 => x"51",
           770 => x"88",
           771 => x"ff",
           772 => x"81",
           773 => x"83",
           774 => x"75",
           775 => x"3d",
           776 => x"3d",
           777 => x"80",
           778 => x"0b",
           779 => x"f5",
           780 => x"08",
           781 => x"82",
           782 => x"f2",
           783 => x"53",
           784 => x"53",
           785 => x"d3",
           786 => x"81",
           787 => x"76",
           788 => x"81",
           789 => x"90",
           790 => x"53",
           791 => x"51",
           792 => x"88",
           793 => x"8d",
           794 => x"74",
           795 => x"38",
           796 => x"05",
           797 => x"3f",
           798 => x"08",
           799 => x"5a",
           800 => x"88",
           801 => x"06",
           802 => x"2e",
           803 => x"86",
           804 => x"82",
           805 => x"80",
           806 => x"86",
           807 => x"39",
           808 => x"53",
           809 => x"51",
           810 => x"81",
           811 => x"81",
           812 => x"3d",
           813 => x"f6",
           814 => x"08",
           815 => x"06",
           816 => x"38",
           817 => x"05",
           818 => x"3f",
           819 => x"02",
           820 => x"78",
           821 => x"88",
           822 => x"70",
           823 => x"5b",
           824 => x"88",
           825 => x"ff",
           826 => x"8c",
           827 => x"3d",
           828 => x"34",
           829 => x"05",
           830 => x"3f",
           831 => x"1a",
           832 => x"e2",
           833 => x"e4",
           834 => x"83",
           835 => x"56",
           836 => x"95",
           837 => x"51",
           838 => x"88",
           839 => x"51",
           840 => x"88",
           841 => x"ff",
           842 => x"31",
           843 => x"1b",
           844 => x"2a",
           845 => x"56",
           846 => x"55",
           847 => x"55",
           848 => x"88",
           849 => x"70",
           850 => x"88",
           851 => x"05",
           852 => x"83",
           853 => x"83",
           854 => x"83",
           855 => x"27",
           856 => x"57",
           857 => x"56",
           858 => x"80",
           859 => x"79",
           860 => x"2e",
           861 => x"90",
           862 => x"fb",
           863 => x"81",
           864 => x"90",
           865 => x"39",
           866 => x"18",
           867 => x"79",
           868 => x"06",
           869 => x"19",
           870 => x"05",
           871 => x"55",
           872 => x"1a",
           873 => x"0b",
           874 => x"0c",
           875 => x"88",
           876 => x"0d",
           877 => x"0d",
           878 => x"9f",
           879 => x"85",
           880 => x"2e",
           881 => x"80",
           882 => x"34",
           883 => x"11",
           884 => x"89",
           885 => x"57",
           886 => x"f8",
           887 => x"08",
           888 => x"80",
           889 => x"3d",
           890 => x"80",
           891 => x"02",
           892 => x"70",
           893 => x"81",
           894 => x"57",
           895 => x"85",
           896 => x"a1",
           897 => x"f5",
           898 => x"08",
           899 => x"98",
           900 => x"51",
           901 => x"88",
           902 => x"0c",
           903 => x"0c",
           904 => x"16",
           905 => x"0c",
           906 => x"04",
           907 => x"7d",
           908 => x"0b",
           909 => x"08",
           910 => x"58",
           911 => x"85",
           912 => x"2e",
           913 => x"81",
           914 => x"06",
           915 => x"74",
           916 => x"c3",
           917 => x"74",
           918 => x"86",
           919 => x"81",
           920 => x"57",
           921 => x"9c",
           922 => x"17",
           923 => x"74",
           924 => x"38",
           925 => x"80",
           926 => x"38",
           927 => x"70",
           928 => x"56",
           929 => x"c7",
           930 => x"33",
           931 => x"89",
           932 => x"81",
           933 => x"55",
           934 => x"76",
           935 => x"16",
           936 => x"39",
           937 => x"51",
           938 => x"88",
           939 => x"75",
           940 => x"38",
           941 => x"0c",
           942 => x"51",
           943 => x"88",
           944 => x"08",
           945 => x"8f",
           946 => x"1a",
           947 => x"98",
           948 => x"ff",
           949 => x"71",
           950 => x"77",
           951 => x"38",
           952 => x"54",
           953 => x"83",
           954 => x"a8",
           955 => x"78",
           956 => x"3f",
           957 => x"e5",
           958 => x"08",
           959 => x"0c",
           960 => x"7b",
           961 => x"0c",
           962 => x"2e",
           963 => x"74",
           964 => x"e2",
           965 => x"76",
           966 => x"3d",
           967 => x"3d",
           968 => x"94",
           969 => x"87",
           970 => x"73",
           971 => x"3f",
           972 => x"2b",
           973 => x"8c",
           974 => x"87",
           975 => x"74",
           976 => x"3f",
           977 => x"07",
           978 => x"8c",
           979 => x"94",
           980 => x"87",
           981 => x"73",
           982 => x"3f",
           983 => x"2b",
           984 => x"9c",
           985 => x"87",
           986 => x"74",
           987 => x"3f",
           988 => x"07",
           989 => x"9c",
           990 => x"83",
           991 => x"94",
           992 => x"80",
           993 => x"c0",
           994 => x"9f",
           995 => x"92",
           996 => x"b8",
           997 => x"51",
           998 => x"88",
           999 => x"a0",
          1000 => x"08",
          1001 => x"88",
          1002 => x"3d",
          1003 => x"84",
          1004 => x"51",
          1005 => x"88",
          1006 => x"75",
          1007 => x"2e",
          1008 => x"15",
          1009 => x"a0",
          1010 => x"04",
          1011 => x"39",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"00",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"4e",
          1018 => x"4f",
          1019 => x"00",
          1020 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"bb",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"0b",
          2058 => x"84",
          2059 => x"0b",
          2060 => x"0b",
          2061 => x"a3",
          2062 => x"0b",
          2063 => x"0b",
          2064 => x"c3",
          2065 => x"0b",
          2066 => x"0b",
          2067 => x"e3",
          2068 => x"0b",
          2069 => x"0b",
          2070 => x"83",
          2071 => x"0b",
          2072 => x"0b",
          2073 => x"a3",
          2074 => x"0b",
          2075 => x"0b",
          2076 => x"c3",
          2077 => x"0b",
          2078 => x"0b",
          2079 => x"e2",
          2080 => x"0b",
          2081 => x"0b",
          2082 => x"80",
          2083 => x"0b",
          2084 => x"0b",
          2085 => x"9e",
          2086 => x"0b",
          2087 => x"0b",
          2088 => x"be",
          2089 => x"0b",
          2090 => x"0b",
          2091 => x"de",
          2092 => x"0b",
          2093 => x"0b",
          2094 => x"fe",
          2095 => x"0b",
          2096 => x"0b",
          2097 => x"9e",
          2098 => x"0b",
          2099 => x"0b",
          2100 => x"be",
          2101 => x"0b",
          2102 => x"0b",
          2103 => x"de",
          2104 => x"0b",
          2105 => x"0b",
          2106 => x"fe",
          2107 => x"0b",
          2108 => x"0b",
          2109 => x"9e",
          2110 => x"0b",
          2111 => x"0b",
          2112 => x"be",
          2113 => x"0b",
          2114 => x"0b",
          2115 => x"de",
          2116 => x"0b",
          2117 => x"0b",
          2118 => x"fe",
          2119 => x"0b",
          2120 => x"0b",
          2121 => x"9e",
          2122 => x"0b",
          2123 => x"0b",
          2124 => x"be",
          2125 => x"0b",
          2126 => x"0b",
          2127 => x"de",
          2128 => x"0b",
          2129 => x"0b",
          2130 => x"fe",
          2131 => x"0b",
          2132 => x"0b",
          2133 => x"9c",
          2134 => x"0b",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"e8",
          2178 => x"2d",
          2179 => x"08",
          2180 => x"04",
          2181 => x"0c",
          2182 => x"2d",
          2183 => x"08",
          2184 => x"04",
          2185 => x"0c",
          2186 => x"2d",
          2187 => x"08",
          2188 => x"04",
          2189 => x"0c",
          2190 => x"2d",
          2191 => x"08",
          2192 => x"04",
          2193 => x"0c",
          2194 => x"2d",
          2195 => x"08",
          2196 => x"04",
          2197 => x"0c",
          2198 => x"2d",
          2199 => x"08",
          2200 => x"04",
          2201 => x"0c",
          2202 => x"2d",
          2203 => x"08",
          2204 => x"04",
          2205 => x"0c",
          2206 => x"2d",
          2207 => x"08",
          2208 => x"04",
          2209 => x"0c",
          2210 => x"2d",
          2211 => x"08",
          2212 => x"04",
          2213 => x"0c",
          2214 => x"2d",
          2215 => x"08",
          2216 => x"04",
          2217 => x"0c",
          2218 => x"2d",
          2219 => x"08",
          2220 => x"04",
          2221 => x"0c",
          2222 => x"2d",
          2223 => x"08",
          2224 => x"04",
          2225 => x"0c",
          2226 => x"2d",
          2227 => x"08",
          2228 => x"04",
          2229 => x"0c",
          2230 => x"82",
          2231 => x"83",
          2232 => x"82",
          2233 => x"ba",
          2234 => x"8c",
          2235 => x"80",
          2236 => x"8c",
          2237 => x"9a",
          2238 => x"e8",
          2239 => x"90",
          2240 => x"e8",
          2241 => x"2d",
          2242 => x"08",
          2243 => x"04",
          2244 => x"0c",
          2245 => x"82",
          2246 => x"83",
          2247 => x"82",
          2248 => x"81",
          2249 => x"82",
          2250 => x"83",
          2251 => x"82",
          2252 => x"81",
          2253 => x"82",
          2254 => x"83",
          2255 => x"82",
          2256 => x"81",
          2257 => x"82",
          2258 => x"83",
          2259 => x"82",
          2260 => x"81",
          2261 => x"82",
          2262 => x"83",
          2263 => x"82",
          2264 => x"81",
          2265 => x"82",
          2266 => x"83",
          2267 => x"82",
          2268 => x"81",
          2269 => x"82",
          2270 => x"83",
          2271 => x"82",
          2272 => x"81",
          2273 => x"82",
          2274 => x"83",
          2275 => x"82",
          2276 => x"81",
          2277 => x"82",
          2278 => x"83",
          2279 => x"82",
          2280 => x"81",
          2281 => x"82",
          2282 => x"83",
          2283 => x"82",
          2284 => x"81",
          2285 => x"82",
          2286 => x"83",
          2287 => x"82",
          2288 => x"81",
          2289 => x"82",
          2290 => x"83",
          2291 => x"82",
          2292 => x"81",
          2293 => x"82",
          2294 => x"83",
          2295 => x"82",
          2296 => x"81",
          2297 => x"82",
          2298 => x"83",
          2299 => x"82",
          2300 => x"81",
          2301 => x"82",
          2302 => x"83",
          2303 => x"82",
          2304 => x"81",
          2305 => x"82",
          2306 => x"83",
          2307 => x"82",
          2308 => x"81",
          2309 => x"82",
          2310 => x"83",
          2311 => x"82",
          2312 => x"81",
          2313 => x"82",
          2314 => x"83",
          2315 => x"82",
          2316 => x"81",
          2317 => x"82",
          2318 => x"83",
          2319 => x"82",
          2320 => x"81",
          2321 => x"82",
          2322 => x"83",
          2323 => x"82",
          2324 => x"81",
          2325 => x"82",
          2326 => x"83",
          2327 => x"82",
          2328 => x"81",
          2329 => x"82",
          2330 => x"83",
          2331 => x"82",
          2332 => x"81",
          2333 => x"82",
          2334 => x"83",
          2335 => x"82",
          2336 => x"81",
          2337 => x"82",
          2338 => x"83",
          2339 => x"82",
          2340 => x"81",
          2341 => x"82",
          2342 => x"83",
          2343 => x"82",
          2344 => x"81",
          2345 => x"82",
          2346 => x"83",
          2347 => x"82",
          2348 => x"81",
          2349 => x"82",
          2350 => x"83",
          2351 => x"82",
          2352 => x"81",
          2353 => x"82",
          2354 => x"83",
          2355 => x"82",
          2356 => x"80",
          2357 => x"82",
          2358 => x"83",
          2359 => x"82",
          2360 => x"80",
          2361 => x"82",
          2362 => x"83",
          2363 => x"82",
          2364 => x"80",
          2365 => x"82",
          2366 => x"83",
          2367 => x"82",
          2368 => x"b3",
          2369 => x"8c",
          2370 => x"80",
          2371 => x"8c",
          2372 => x"a5",
          2373 => x"e8",
          2374 => x"90",
          2375 => x"e8",
          2376 => x"2d",
          2377 => x"08",
          2378 => x"04",
          2379 => x"0c",
          2380 => x"2d",
          2381 => x"08",
          2382 => x"04",
          2383 => x"70",
          2384 => x"27",
          2385 => x"71",
          2386 => x"53",
          2387 => x"0b",
          2388 => x"a4",
          2389 => x"ef",
          2390 => x"04",
          2391 => x"08",
          2392 => x"e8",
          2393 => x"0d",
          2394 => x"8c",
          2395 => x"05",
          2396 => x"8c",
          2397 => x"05",
          2398 => x"c5",
          2399 => x"dc",
          2400 => x"8c",
          2401 => x"85",
          2402 => x"8c",
          2403 => x"82",
          2404 => x"02",
          2405 => x"0c",
          2406 => x"81",
          2407 => x"e8",
          2408 => x"08",
          2409 => x"e8",
          2410 => x"08",
          2411 => x"82",
          2412 => x"70",
          2413 => x"0c",
          2414 => x"0d",
          2415 => x"0c",
          2416 => x"e8",
          2417 => x"8c",
          2418 => x"3d",
          2419 => x"82",
          2420 => x"fc",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"8c",
          2425 => x"8c",
          2426 => x"05",
          2427 => x"38",
          2428 => x"08",
          2429 => x"80",
          2430 => x"80",
          2431 => x"e8",
          2432 => x"08",
          2433 => x"82",
          2434 => x"8c",
          2435 => x"82",
          2436 => x"8c",
          2437 => x"8c",
          2438 => x"05",
          2439 => x"8c",
          2440 => x"05",
          2441 => x"39",
          2442 => x"08",
          2443 => x"80",
          2444 => x"38",
          2445 => x"08",
          2446 => x"82",
          2447 => x"88",
          2448 => x"ad",
          2449 => x"e8",
          2450 => x"08",
          2451 => x"08",
          2452 => x"31",
          2453 => x"08",
          2454 => x"82",
          2455 => x"f8",
          2456 => x"8c",
          2457 => x"05",
          2458 => x"8c",
          2459 => x"05",
          2460 => x"e8",
          2461 => x"08",
          2462 => x"8c",
          2463 => x"05",
          2464 => x"e8",
          2465 => x"08",
          2466 => x"8c",
          2467 => x"05",
          2468 => x"39",
          2469 => x"08",
          2470 => x"80",
          2471 => x"82",
          2472 => x"88",
          2473 => x"82",
          2474 => x"f4",
          2475 => x"91",
          2476 => x"e8",
          2477 => x"08",
          2478 => x"e8",
          2479 => x"0c",
          2480 => x"e8",
          2481 => x"08",
          2482 => x"0c",
          2483 => x"82",
          2484 => x"04",
          2485 => x"76",
          2486 => x"55",
          2487 => x"8f",
          2488 => x"38",
          2489 => x"83",
          2490 => x"80",
          2491 => x"ff",
          2492 => x"ff",
          2493 => x"72",
          2494 => x"54",
          2495 => x"81",
          2496 => x"ff",
          2497 => x"ff",
          2498 => x"06",
          2499 => x"82",
          2500 => x"86",
          2501 => x"74",
          2502 => x"84",
          2503 => x"71",
          2504 => x"53",
          2505 => x"84",
          2506 => x"71",
          2507 => x"53",
          2508 => x"84",
          2509 => x"71",
          2510 => x"53",
          2511 => x"84",
          2512 => x"71",
          2513 => x"53",
          2514 => x"52",
          2515 => x"c9",
          2516 => x"27",
          2517 => x"70",
          2518 => x"08",
          2519 => x"05",
          2520 => x"12",
          2521 => x"26",
          2522 => x"54",
          2523 => x"fc",
          2524 => x"79",
          2525 => x"05",
          2526 => x"57",
          2527 => x"83",
          2528 => x"38",
          2529 => x"51",
          2530 => x"a4",
          2531 => x"52",
          2532 => x"93",
          2533 => x"70",
          2534 => x"34",
          2535 => x"71",
          2536 => x"81",
          2537 => x"74",
          2538 => x"0c",
          2539 => x"04",
          2540 => x"2b",
          2541 => x"71",
          2542 => x"51",
          2543 => x"72",
          2544 => x"72",
          2545 => x"05",
          2546 => x"71",
          2547 => x"53",
          2548 => x"70",
          2549 => x"0c",
          2550 => x"84",
          2551 => x"f0",
          2552 => x"8f",
          2553 => x"83",
          2554 => x"38",
          2555 => x"84",
          2556 => x"fc",
          2557 => x"83",
          2558 => x"70",
          2559 => x"39",
          2560 => x"76",
          2561 => x"73",
          2562 => x"54",
          2563 => x"70",
          2564 => x"71",
          2565 => x"09",
          2566 => x"fd",
          2567 => x"70",
          2568 => x"81",
          2569 => x"51",
          2570 => x"70",
          2571 => x"14",
          2572 => x"84",
          2573 => x"70",
          2574 => x"70",
          2575 => x"ff",
          2576 => x"f8",
          2577 => x"80",
          2578 => x"53",
          2579 => x"80",
          2580 => x"73",
          2581 => x"81",
          2582 => x"51",
          2583 => x"81",
          2584 => x"70",
          2585 => x"82",
          2586 => x"86",
          2587 => x"fd",
          2588 => x"70",
          2589 => x"53",
          2590 => x"b8",
          2591 => x"08",
          2592 => x"fb",
          2593 => x"06",
          2594 => x"82",
          2595 => x"51",
          2596 => x"70",
          2597 => x"13",
          2598 => x"09",
          2599 => x"ff",
          2600 => x"f8",
          2601 => x"80",
          2602 => x"52",
          2603 => x"2e",
          2604 => x"52",
          2605 => x"70",
          2606 => x"38",
          2607 => x"33",
          2608 => x"f8",
          2609 => x"31",
          2610 => x"0c",
          2611 => x"04",
          2612 => x"78",
          2613 => x"54",
          2614 => x"72",
          2615 => x"d9",
          2616 => x"07",
          2617 => x"70",
          2618 => x"d6",
          2619 => x"53",
          2620 => x"b1",
          2621 => x"74",
          2622 => x"74",
          2623 => x"81",
          2624 => x"72",
          2625 => x"89",
          2626 => x"ff",
          2627 => x"80",
          2628 => x"38",
          2629 => x"15",
          2630 => x"55",
          2631 => x"2e",
          2632 => x"d1",
          2633 => x"74",
          2634 => x"70",
          2635 => x"75",
          2636 => x"71",
          2637 => x"52",
          2638 => x"8c",
          2639 => x"3d",
          2640 => x"74",
          2641 => x"73",
          2642 => x"71",
          2643 => x"2e",
          2644 => x"76",
          2645 => x"95",
          2646 => x"53",
          2647 => x"b1",
          2648 => x"70",
          2649 => x"fd",
          2650 => x"70",
          2651 => x"81",
          2652 => x"51",
          2653 => x"38",
          2654 => x"17",
          2655 => x"73",
          2656 => x"74",
          2657 => x"2e",
          2658 => x"76",
          2659 => x"dd",
          2660 => x"82",
          2661 => x"88",
          2662 => x"fe",
          2663 => x"52",
          2664 => x"88",
          2665 => x"86",
          2666 => x"dc",
          2667 => x"06",
          2668 => x"14",
          2669 => x"80",
          2670 => x"71",
          2671 => x"0c",
          2672 => x"04",
          2673 => x"77",
          2674 => x"53",
          2675 => x"80",
          2676 => x"38",
          2677 => x"70",
          2678 => x"81",
          2679 => x"81",
          2680 => x"39",
          2681 => x"39",
          2682 => x"80",
          2683 => x"81",
          2684 => x"55",
          2685 => x"2e",
          2686 => x"55",
          2687 => x"84",
          2688 => x"38",
          2689 => x"06",
          2690 => x"2e",
          2691 => x"88",
          2692 => x"70",
          2693 => x"34",
          2694 => x"71",
          2695 => x"8c",
          2696 => x"3d",
          2697 => x"3d",
          2698 => x"72",
          2699 => x"91",
          2700 => x"fc",
          2701 => x"51",
          2702 => x"82",
          2703 => x"85",
          2704 => x"83",
          2705 => x"72",
          2706 => x"0c",
          2707 => x"04",
          2708 => x"76",
          2709 => x"ff",
          2710 => x"81",
          2711 => x"26",
          2712 => x"83",
          2713 => x"05",
          2714 => x"70",
          2715 => x"8a",
          2716 => x"33",
          2717 => x"70",
          2718 => x"fe",
          2719 => x"33",
          2720 => x"70",
          2721 => x"f2",
          2722 => x"33",
          2723 => x"70",
          2724 => x"e6",
          2725 => x"22",
          2726 => x"74",
          2727 => x"80",
          2728 => x"13",
          2729 => x"52",
          2730 => x"26",
          2731 => x"81",
          2732 => x"98",
          2733 => x"22",
          2734 => x"bc",
          2735 => x"33",
          2736 => x"b8",
          2737 => x"33",
          2738 => x"b4",
          2739 => x"33",
          2740 => x"b0",
          2741 => x"33",
          2742 => x"ac",
          2743 => x"33",
          2744 => x"a8",
          2745 => x"c0",
          2746 => x"73",
          2747 => x"a0",
          2748 => x"87",
          2749 => x"0c",
          2750 => x"82",
          2751 => x"86",
          2752 => x"f3",
          2753 => x"5b",
          2754 => x"9c",
          2755 => x"0c",
          2756 => x"bc",
          2757 => x"7b",
          2758 => x"98",
          2759 => x"79",
          2760 => x"87",
          2761 => x"08",
          2762 => x"1c",
          2763 => x"98",
          2764 => x"79",
          2765 => x"87",
          2766 => x"08",
          2767 => x"1c",
          2768 => x"98",
          2769 => x"79",
          2770 => x"87",
          2771 => x"08",
          2772 => x"1c",
          2773 => x"98",
          2774 => x"79",
          2775 => x"80",
          2776 => x"83",
          2777 => x"59",
          2778 => x"ff",
          2779 => x"1b",
          2780 => x"1b",
          2781 => x"1b",
          2782 => x"1b",
          2783 => x"1b",
          2784 => x"83",
          2785 => x"52",
          2786 => x"51",
          2787 => x"8f",
          2788 => x"ff",
          2789 => x"8f",
          2790 => x"30",
          2791 => x"51",
          2792 => x"0b",
          2793 => x"d4",
          2794 => x"0d",
          2795 => x"0d",
          2796 => x"82",
          2797 => x"70",
          2798 => x"57",
          2799 => x"c0",
          2800 => x"74",
          2801 => x"38",
          2802 => x"94",
          2803 => x"70",
          2804 => x"81",
          2805 => x"52",
          2806 => x"8c",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"38",
          2810 => x"70",
          2811 => x"51",
          2812 => x"8d",
          2813 => x"2a",
          2814 => x"51",
          2815 => x"be",
          2816 => x"ff",
          2817 => x"c0",
          2818 => x"70",
          2819 => x"38",
          2820 => x"90",
          2821 => x"0c",
          2822 => x"dc",
          2823 => x"0d",
          2824 => x"0d",
          2825 => x"33",
          2826 => x"87",
          2827 => x"81",
          2828 => x"55",
          2829 => x"94",
          2830 => x"80",
          2831 => x"87",
          2832 => x"51",
          2833 => x"96",
          2834 => x"06",
          2835 => x"70",
          2836 => x"38",
          2837 => x"70",
          2838 => x"51",
          2839 => x"72",
          2840 => x"81",
          2841 => x"70",
          2842 => x"38",
          2843 => x"70",
          2844 => x"51",
          2845 => x"38",
          2846 => x"06",
          2847 => x"94",
          2848 => x"80",
          2849 => x"87",
          2850 => x"52",
          2851 => x"87",
          2852 => x"f9",
          2853 => x"54",
          2854 => x"70",
          2855 => x"53",
          2856 => x"77",
          2857 => x"38",
          2858 => x"06",
          2859 => x"0b",
          2860 => x"33",
          2861 => x"06",
          2862 => x"58",
          2863 => x"84",
          2864 => x"2e",
          2865 => x"c0",
          2866 => x"70",
          2867 => x"2a",
          2868 => x"53",
          2869 => x"80",
          2870 => x"71",
          2871 => x"81",
          2872 => x"70",
          2873 => x"81",
          2874 => x"06",
          2875 => x"80",
          2876 => x"71",
          2877 => x"81",
          2878 => x"70",
          2879 => x"74",
          2880 => x"51",
          2881 => x"80",
          2882 => x"2e",
          2883 => x"c0",
          2884 => x"77",
          2885 => x"17",
          2886 => x"81",
          2887 => x"53",
          2888 => x"84",
          2889 => x"8c",
          2890 => x"3d",
          2891 => x"3d",
          2892 => x"82",
          2893 => x"70",
          2894 => x"54",
          2895 => x"94",
          2896 => x"80",
          2897 => x"87",
          2898 => x"51",
          2899 => x"82",
          2900 => x"06",
          2901 => x"70",
          2902 => x"38",
          2903 => x"06",
          2904 => x"94",
          2905 => x"80",
          2906 => x"87",
          2907 => x"52",
          2908 => x"81",
          2909 => x"8c",
          2910 => x"84",
          2911 => x"fe",
          2912 => x"0b",
          2913 => x"33",
          2914 => x"06",
          2915 => x"c0",
          2916 => x"70",
          2917 => x"38",
          2918 => x"94",
          2919 => x"70",
          2920 => x"81",
          2921 => x"51",
          2922 => x"80",
          2923 => x"72",
          2924 => x"51",
          2925 => x"80",
          2926 => x"2e",
          2927 => x"c0",
          2928 => x"71",
          2929 => x"2b",
          2930 => x"51",
          2931 => x"82",
          2932 => x"84",
          2933 => x"ff",
          2934 => x"c0",
          2935 => x"70",
          2936 => x"06",
          2937 => x"80",
          2938 => x"38",
          2939 => x"a4",
          2940 => x"d8",
          2941 => x"9e",
          2942 => x"87",
          2943 => x"c0",
          2944 => x"82",
          2945 => x"87",
          2946 => x"08",
          2947 => x"0c",
          2948 => x"9c",
          2949 => x"e8",
          2950 => x"9e",
          2951 => x"87",
          2952 => x"c0",
          2953 => x"82",
          2954 => x"87",
          2955 => x"08",
          2956 => x"0c",
          2957 => x"b4",
          2958 => x"f8",
          2959 => x"9e",
          2960 => x"87",
          2961 => x"c0",
          2962 => x"82",
          2963 => x"87",
          2964 => x"08",
          2965 => x"0c",
          2966 => x"c4",
          2967 => x"88",
          2968 => x"9e",
          2969 => x"70",
          2970 => x"23",
          2971 => x"84",
          2972 => x"90",
          2973 => x"9e",
          2974 => x"88",
          2975 => x"c0",
          2976 => x"82",
          2977 => x"81",
          2978 => x"9c",
          2979 => x"87",
          2980 => x"08",
          2981 => x"0a",
          2982 => x"52",
          2983 => x"83",
          2984 => x"71",
          2985 => x"34",
          2986 => x"c0",
          2987 => x"70",
          2988 => x"06",
          2989 => x"70",
          2990 => x"38",
          2991 => x"82",
          2992 => x"80",
          2993 => x"9e",
          2994 => x"90",
          2995 => x"51",
          2996 => x"80",
          2997 => x"81",
          2998 => x"88",
          2999 => x"0b",
          3000 => x"90",
          3001 => x"80",
          3002 => x"52",
          3003 => x"2e",
          3004 => x"52",
          3005 => x"a0",
          3006 => x"87",
          3007 => x"08",
          3008 => x"80",
          3009 => x"52",
          3010 => x"83",
          3011 => x"71",
          3012 => x"34",
          3013 => x"c0",
          3014 => x"70",
          3015 => x"06",
          3016 => x"70",
          3017 => x"38",
          3018 => x"82",
          3019 => x"80",
          3020 => x"9e",
          3021 => x"84",
          3022 => x"51",
          3023 => x"80",
          3024 => x"81",
          3025 => x"88",
          3026 => x"0b",
          3027 => x"90",
          3028 => x"80",
          3029 => x"52",
          3030 => x"2e",
          3031 => x"52",
          3032 => x"a4",
          3033 => x"87",
          3034 => x"08",
          3035 => x"80",
          3036 => x"52",
          3037 => x"83",
          3038 => x"71",
          3039 => x"34",
          3040 => x"c0",
          3041 => x"70",
          3042 => x"06",
          3043 => x"70",
          3044 => x"38",
          3045 => x"82",
          3046 => x"80",
          3047 => x"9e",
          3048 => x"a0",
          3049 => x"52",
          3050 => x"2e",
          3051 => x"52",
          3052 => x"a7",
          3053 => x"9e",
          3054 => x"98",
          3055 => x"8a",
          3056 => x"51",
          3057 => x"a8",
          3058 => x"87",
          3059 => x"08",
          3060 => x"06",
          3061 => x"70",
          3062 => x"38",
          3063 => x"82",
          3064 => x"87",
          3065 => x"08",
          3066 => x"06",
          3067 => x"51",
          3068 => x"82",
          3069 => x"80",
          3070 => x"9e",
          3071 => x"88",
          3072 => x"52",
          3073 => x"83",
          3074 => x"71",
          3075 => x"34",
          3076 => x"90",
          3077 => x"06",
          3078 => x"82",
          3079 => x"83",
          3080 => x"fb",
          3081 => x"f1",
          3082 => x"dc",
          3083 => x"9c",
          3084 => x"80",
          3085 => x"81",
          3086 => x"89",
          3087 => x"f2",
          3088 => x"c4",
          3089 => x"9e",
          3090 => x"80",
          3091 => x"82",
          3092 => x"82",
          3093 => x"11",
          3094 => x"f2",
          3095 => x"8c",
          3096 => x"a3",
          3097 => x"80",
          3098 => x"82",
          3099 => x"82",
          3100 => x"11",
          3101 => x"f2",
          3102 => x"f0",
          3103 => x"a0",
          3104 => x"80",
          3105 => x"82",
          3106 => x"82",
          3107 => x"11",
          3108 => x"f2",
          3109 => x"d4",
          3110 => x"a1",
          3111 => x"80",
          3112 => x"82",
          3113 => x"82",
          3114 => x"11",
          3115 => x"f3",
          3116 => x"b8",
          3117 => x"a2",
          3118 => x"80",
          3119 => x"82",
          3120 => x"82",
          3121 => x"11",
          3122 => x"f3",
          3123 => x"9c",
          3124 => x"a7",
          3125 => x"80",
          3126 => x"82",
          3127 => x"52",
          3128 => x"51",
          3129 => x"82",
          3130 => x"54",
          3131 => x"8d",
          3132 => x"ac",
          3133 => x"f3",
          3134 => x"f0",
          3135 => x"a9",
          3136 => x"80",
          3137 => x"82",
          3138 => x"52",
          3139 => x"51",
          3140 => x"82",
          3141 => x"54",
          3142 => x"88",
          3143 => x"a8",
          3144 => x"3f",
          3145 => x"33",
          3146 => x"2e",
          3147 => x"f4",
          3148 => x"d4",
          3149 => x"a4",
          3150 => x"80",
          3151 => x"81",
          3152 => x"87",
          3153 => x"88",
          3154 => x"73",
          3155 => x"38",
          3156 => x"51",
          3157 => x"82",
          3158 => x"54",
          3159 => x"88",
          3160 => x"e0",
          3161 => x"3f",
          3162 => x"51",
          3163 => x"82",
          3164 => x"52",
          3165 => x"51",
          3166 => x"82",
          3167 => x"52",
          3168 => x"51",
          3169 => x"82",
          3170 => x"52",
          3171 => x"51",
          3172 => x"81",
          3173 => x"86",
          3174 => x"88",
          3175 => x"81",
          3176 => x"8c",
          3177 => x"88",
          3178 => x"bd",
          3179 => x"75",
          3180 => x"3f",
          3181 => x"08",
          3182 => x"29",
          3183 => x"54",
          3184 => x"dc",
          3185 => x"f6",
          3186 => x"a0",
          3187 => x"a3",
          3188 => x"80",
          3189 => x"82",
          3190 => x"56",
          3191 => x"52",
          3192 => x"f8",
          3193 => x"dc",
          3194 => x"c0",
          3195 => x"31",
          3196 => x"8c",
          3197 => x"81",
          3198 => x"8b",
          3199 => x"88",
          3200 => x"73",
          3201 => x"38",
          3202 => x"08",
          3203 => x"c0",
          3204 => x"e6",
          3205 => x"8c",
          3206 => x"84",
          3207 => x"71",
          3208 => x"82",
          3209 => x"52",
          3210 => x"51",
          3211 => x"82",
          3212 => x"85",
          3213 => x"3d",
          3214 => x"3d",
          3215 => x"05",
          3216 => x"52",
          3217 => x"ac",
          3218 => x"29",
          3219 => x"f0",
          3220 => x"71",
          3221 => x"f7",
          3222 => x"39",
          3223 => x"51",
          3224 => x"f7",
          3225 => x"39",
          3226 => x"51",
          3227 => x"f7",
          3228 => x"39",
          3229 => x"51",
          3230 => x"84",
          3231 => x"71",
          3232 => x"04",
          3233 => x"c0",
          3234 => x"04",
          3235 => x"08",
          3236 => x"84",
          3237 => x"3d",
          3238 => x"ec",
          3239 => x"82",
          3240 => x"82",
          3241 => x"82",
          3242 => x"75",
          3243 => x"ff",
          3244 => x"b7",
          3245 => x"38",
          3246 => x"ec",
          3247 => x"72",
          3248 => x"0c",
          3249 => x"04",
          3250 => x"79",
          3251 => x"08",
          3252 => x"14",
          3253 => x"08",
          3254 => x"5a",
          3255 => x"57",
          3256 => x"26",
          3257 => x"13",
          3258 => x"53",
          3259 => x"0c",
          3260 => x"84",
          3261 => x"73",
          3262 => x"14",
          3263 => x"12",
          3264 => x"12",
          3265 => x"13",
          3266 => x"14",
          3267 => x"12",
          3268 => x"12",
          3269 => x"15",
          3270 => x"16",
          3271 => x"80",
          3272 => x"90",
          3273 => x"94",
          3274 => x"82",
          3275 => x"89",
          3276 => x"fc",
          3277 => x"8c",
          3278 => x"12",
          3279 => x"53",
          3280 => x"2e",
          3281 => x"a3",
          3282 => x"08",
          3283 => x"55",
          3284 => x"09",
          3285 => x"38",
          3286 => x"15",
          3287 => x"73",
          3288 => x"71",
          3289 => x"71",
          3290 => x"81",
          3291 => x"88",
          3292 => x"14",
          3293 => x"b4",
          3294 => x"0c",
          3295 => x"c4",
          3296 => x"08",
          3297 => x"0c",
          3298 => x"81",
          3299 => x"06",
          3300 => x"13",
          3301 => x"52",
          3302 => x"2e",
          3303 => x"a4",
          3304 => x"08",
          3305 => x"0c",
          3306 => x"90",
          3307 => x"90",
          3308 => x"94",
          3309 => x"14",
          3310 => x"08",
          3311 => x"0c",
          3312 => x"0c",
          3313 => x"dc",
          3314 => x"0d",
          3315 => x"0d",
          3316 => x"57",
          3317 => x"81",
          3318 => x"17",
          3319 => x"88",
          3320 => x"57",
          3321 => x"2e",
          3322 => x"16",
          3323 => x"80",
          3324 => x"16",
          3325 => x"39",
          3326 => x"17",
          3327 => x"06",
          3328 => x"fd",
          3329 => x"8c",
          3330 => x"8c",
          3331 => x"70",
          3332 => x"08",
          3333 => x"82",
          3334 => x"09",
          3335 => x"72",
          3336 => x"73",
          3337 => x"58",
          3338 => x"80",
          3339 => x"2e",
          3340 => x"80",
          3341 => x"39",
          3342 => x"51",
          3343 => x"81",
          3344 => x"dc",
          3345 => x"82",
          3346 => x"84",
          3347 => x"88",
          3348 => x"72",
          3349 => x"8c",
          3350 => x"26",
          3351 => x"13",
          3352 => x"39",
          3353 => x"88",
          3354 => x"8c",
          3355 => x"88",
          3356 => x"16",
          3357 => x"12",
          3358 => x"51",
          3359 => x"76",
          3360 => x"dc",
          3361 => x"c0",
          3362 => x"dc",
          3363 => x"82",
          3364 => x"89",
          3365 => x"ff",
          3366 => x"52",
          3367 => x"87",
          3368 => x"51",
          3369 => x"83",
          3370 => x"fe",
          3371 => x"93",
          3372 => x"72",
          3373 => x"81",
          3374 => x"8d",
          3375 => x"82",
          3376 => x"52",
          3377 => x"90",
          3378 => x"34",
          3379 => x"08",
          3380 => x"8c",
          3381 => x"39",
          3382 => x"08",
          3383 => x"2e",
          3384 => x"51",
          3385 => x"3d",
          3386 => x"3d",
          3387 => x"05",
          3388 => x"f0",
          3389 => x"8c",
          3390 => x"51",
          3391 => x"72",
          3392 => x"0c",
          3393 => x"04",
          3394 => x"75",
          3395 => x"70",
          3396 => x"53",
          3397 => x"2e",
          3398 => x"81",
          3399 => x"81",
          3400 => x"87",
          3401 => x"85",
          3402 => x"fc",
          3403 => x"82",
          3404 => x"78",
          3405 => x"0c",
          3406 => x"33",
          3407 => x"06",
          3408 => x"80",
          3409 => x"72",
          3410 => x"51",
          3411 => x"fe",
          3412 => x"39",
          3413 => x"f0",
          3414 => x"0d",
          3415 => x"0d",
          3416 => x"59",
          3417 => x"05",
          3418 => x"75",
          3419 => x"f8",
          3420 => x"2e",
          3421 => x"82",
          3422 => x"70",
          3423 => x"05",
          3424 => x"5b",
          3425 => x"2e",
          3426 => x"85",
          3427 => x"8b",
          3428 => x"2e",
          3429 => x"8a",
          3430 => x"78",
          3431 => x"5a",
          3432 => x"aa",
          3433 => x"06",
          3434 => x"84",
          3435 => x"7b",
          3436 => x"5d",
          3437 => x"59",
          3438 => x"d0",
          3439 => x"89",
          3440 => x"7a",
          3441 => x"10",
          3442 => x"d0",
          3443 => x"81",
          3444 => x"57",
          3445 => x"75",
          3446 => x"70",
          3447 => x"07",
          3448 => x"80",
          3449 => x"30",
          3450 => x"80",
          3451 => x"53",
          3452 => x"55",
          3453 => x"2e",
          3454 => x"84",
          3455 => x"81",
          3456 => x"57",
          3457 => x"2e",
          3458 => x"75",
          3459 => x"76",
          3460 => x"e0",
          3461 => x"ff",
          3462 => x"73",
          3463 => x"81",
          3464 => x"80",
          3465 => x"38",
          3466 => x"2e",
          3467 => x"73",
          3468 => x"8b",
          3469 => x"c2",
          3470 => x"38",
          3471 => x"73",
          3472 => x"81",
          3473 => x"8f",
          3474 => x"d5",
          3475 => x"38",
          3476 => x"24",
          3477 => x"80",
          3478 => x"38",
          3479 => x"73",
          3480 => x"80",
          3481 => x"ef",
          3482 => x"19",
          3483 => x"59",
          3484 => x"33",
          3485 => x"75",
          3486 => x"81",
          3487 => x"70",
          3488 => x"55",
          3489 => x"79",
          3490 => x"90",
          3491 => x"16",
          3492 => x"7b",
          3493 => x"a0",
          3494 => x"3f",
          3495 => x"53",
          3496 => x"e9",
          3497 => x"fc",
          3498 => x"81",
          3499 => x"72",
          3500 => x"b0",
          3501 => x"fb",
          3502 => x"39",
          3503 => x"83",
          3504 => x"59",
          3505 => x"82",
          3506 => x"88",
          3507 => x"8a",
          3508 => x"90",
          3509 => x"75",
          3510 => x"3f",
          3511 => x"79",
          3512 => x"81",
          3513 => x"72",
          3514 => x"38",
          3515 => x"59",
          3516 => x"84",
          3517 => x"58",
          3518 => x"80",
          3519 => x"30",
          3520 => x"80",
          3521 => x"55",
          3522 => x"25",
          3523 => x"80",
          3524 => x"74",
          3525 => x"07",
          3526 => x"0b",
          3527 => x"57",
          3528 => x"51",
          3529 => x"82",
          3530 => x"81",
          3531 => x"53",
          3532 => x"dc",
          3533 => x"8c",
          3534 => x"89",
          3535 => x"38",
          3536 => x"75",
          3537 => x"84",
          3538 => x"53",
          3539 => x"06",
          3540 => x"53",
          3541 => x"81",
          3542 => x"81",
          3543 => x"70",
          3544 => x"2a",
          3545 => x"76",
          3546 => x"38",
          3547 => x"38",
          3548 => x"70",
          3549 => x"53",
          3550 => x"8e",
          3551 => x"77",
          3552 => x"53",
          3553 => x"81",
          3554 => x"7a",
          3555 => x"55",
          3556 => x"83",
          3557 => x"79",
          3558 => x"81",
          3559 => x"72",
          3560 => x"17",
          3561 => x"27",
          3562 => x"51",
          3563 => x"75",
          3564 => x"72",
          3565 => x"81",
          3566 => x"7a",
          3567 => x"38",
          3568 => x"05",
          3569 => x"ff",
          3570 => x"70",
          3571 => x"57",
          3572 => x"76",
          3573 => x"81",
          3574 => x"72",
          3575 => x"84",
          3576 => x"f9",
          3577 => x"39",
          3578 => x"04",
          3579 => x"86",
          3580 => x"84",
          3581 => x"55",
          3582 => x"fa",
          3583 => x"3d",
          3584 => x"3d",
          3585 => x"8c",
          3586 => x"3d",
          3587 => x"75",
          3588 => x"3f",
          3589 => x"08",
          3590 => x"34",
          3591 => x"8c",
          3592 => x"3d",
          3593 => x"3d",
          3594 => x"f0",
          3595 => x"8c",
          3596 => x"3d",
          3597 => x"77",
          3598 => x"a1",
          3599 => x"8c",
          3600 => x"3d",
          3601 => x"3d",
          3602 => x"82",
          3603 => x"70",
          3604 => x"55",
          3605 => x"80",
          3606 => x"38",
          3607 => x"08",
          3608 => x"82",
          3609 => x"81",
          3610 => x"72",
          3611 => x"cb",
          3612 => x"2e",
          3613 => x"88",
          3614 => x"70",
          3615 => x"51",
          3616 => x"2e",
          3617 => x"80",
          3618 => x"ff",
          3619 => x"39",
          3620 => x"c8",
          3621 => x"52",
          3622 => x"c0",
          3623 => x"52",
          3624 => x"81",
          3625 => x"51",
          3626 => x"ff",
          3627 => x"15",
          3628 => x"34",
          3629 => x"f3",
          3630 => x"72",
          3631 => x"0c",
          3632 => x"04",
          3633 => x"82",
          3634 => x"75",
          3635 => x"0c",
          3636 => x"52",
          3637 => x"3f",
          3638 => x"f4",
          3639 => x"0d",
          3640 => x"0d",
          3641 => x"56",
          3642 => x"0c",
          3643 => x"70",
          3644 => x"73",
          3645 => x"81",
          3646 => x"81",
          3647 => x"ed",
          3648 => x"2e",
          3649 => x"8e",
          3650 => x"08",
          3651 => x"76",
          3652 => x"56",
          3653 => x"b0",
          3654 => x"06",
          3655 => x"75",
          3656 => x"76",
          3657 => x"70",
          3658 => x"73",
          3659 => x"8b",
          3660 => x"73",
          3661 => x"85",
          3662 => x"82",
          3663 => x"76",
          3664 => x"70",
          3665 => x"ac",
          3666 => x"a0",
          3667 => x"fa",
          3668 => x"53",
          3669 => x"57",
          3670 => x"98",
          3671 => x"39",
          3672 => x"80",
          3673 => x"26",
          3674 => x"86",
          3675 => x"80",
          3676 => x"57",
          3677 => x"74",
          3678 => x"38",
          3679 => x"27",
          3680 => x"14",
          3681 => x"06",
          3682 => x"14",
          3683 => x"06",
          3684 => x"74",
          3685 => x"f9",
          3686 => x"ff",
          3687 => x"89",
          3688 => x"38",
          3689 => x"c5",
          3690 => x"29",
          3691 => x"81",
          3692 => x"76",
          3693 => x"56",
          3694 => x"ba",
          3695 => x"2e",
          3696 => x"30",
          3697 => x"0c",
          3698 => x"82",
          3699 => x"8a",
          3700 => x"f8",
          3701 => x"7c",
          3702 => x"70",
          3703 => x"75",
          3704 => x"55",
          3705 => x"2e",
          3706 => x"87",
          3707 => x"76",
          3708 => x"73",
          3709 => x"81",
          3710 => x"81",
          3711 => x"77",
          3712 => x"70",
          3713 => x"58",
          3714 => x"09",
          3715 => x"c2",
          3716 => x"81",
          3717 => x"75",
          3718 => x"55",
          3719 => x"e2",
          3720 => x"90",
          3721 => x"f8",
          3722 => x"8f",
          3723 => x"81",
          3724 => x"75",
          3725 => x"55",
          3726 => x"81",
          3727 => x"27",
          3728 => x"d0",
          3729 => x"55",
          3730 => x"73",
          3731 => x"80",
          3732 => x"14",
          3733 => x"72",
          3734 => x"e0",
          3735 => x"80",
          3736 => x"39",
          3737 => x"55",
          3738 => x"80",
          3739 => x"e0",
          3740 => x"38",
          3741 => x"81",
          3742 => x"53",
          3743 => x"81",
          3744 => x"53",
          3745 => x"8e",
          3746 => x"70",
          3747 => x"55",
          3748 => x"27",
          3749 => x"77",
          3750 => x"74",
          3751 => x"76",
          3752 => x"77",
          3753 => x"70",
          3754 => x"55",
          3755 => x"77",
          3756 => x"38",
          3757 => x"74",
          3758 => x"55",
          3759 => x"dc",
          3760 => x"0d",
          3761 => x"0d",
          3762 => x"70",
          3763 => x"98",
          3764 => x"2c",
          3765 => x"70",
          3766 => x"53",
          3767 => x"51",
          3768 => x"f8",
          3769 => x"55",
          3770 => x"25",
          3771 => x"f8",
          3772 => x"12",
          3773 => x"97",
          3774 => x"33",
          3775 => x"70",
          3776 => x"81",
          3777 => x"81",
          3778 => x"8c",
          3779 => x"3d",
          3780 => x"3d",
          3781 => x"84",
          3782 => x"33",
          3783 => x"55",
          3784 => x"2e",
          3785 => x"51",
          3786 => x"a0",
          3787 => x"3f",
          3788 => x"f7",
          3789 => x"ff",
          3790 => x"73",
          3791 => x"ff",
          3792 => x"39",
          3793 => x"c0",
          3794 => x"34",
          3795 => x"04",
          3796 => x"7c",
          3797 => x"b7",
          3798 => x"88",
          3799 => x"33",
          3800 => x"33",
          3801 => x"82",
          3802 => x"70",
          3803 => x"59",
          3804 => x"74",
          3805 => x"38",
          3806 => x"9b",
          3807 => x"a8",
          3808 => x"29",
          3809 => x"05",
          3810 => x"54",
          3811 => x"f0",
          3812 => x"8c",
          3813 => x"0c",
          3814 => x"33",
          3815 => x"82",
          3816 => x"70",
          3817 => x"5a",
          3818 => x"a6",
          3819 => x"78",
          3820 => x"d6",
          3821 => x"89",
          3822 => x"05",
          3823 => x"89",
          3824 => x"81",
          3825 => x"93",
          3826 => x"38",
          3827 => x"89",
          3828 => x"80",
          3829 => x"82",
          3830 => x"56",
          3831 => x"ac",
          3832 => x"a0",
          3833 => x"a4",
          3834 => x"fc",
          3835 => x"53",
          3836 => x"51",
          3837 => x"3f",
          3838 => x"08",
          3839 => x"80",
          3840 => x"82",
          3841 => x"51",
          3842 => x"3f",
          3843 => x"04",
          3844 => x"81",
          3845 => x"82",
          3846 => x"51",
          3847 => x"3f",
          3848 => x"08",
          3849 => x"82",
          3850 => x"53",
          3851 => x"88",
          3852 => x"56",
          3853 => x"3f",
          3854 => x"08",
          3855 => x"38",
          3856 => x"ab",
          3857 => x"dc",
          3858 => x"0b",
          3859 => x"08",
          3860 => x"82",
          3861 => x"ff",
          3862 => x"55",
          3863 => x"34",
          3864 => x"52",
          3865 => x"f7",
          3866 => x"f6",
          3867 => x"ff",
          3868 => x"06",
          3869 => x"a6",
          3870 => x"d9",
          3871 => x"3d",
          3872 => x"08",
          3873 => x"70",
          3874 => x"52",
          3875 => x"08",
          3876 => x"92",
          3877 => x"dc",
          3878 => x"38",
          3879 => x"89",
          3880 => x"55",
          3881 => x"8b",
          3882 => x"56",
          3883 => x"3f",
          3884 => x"08",
          3885 => x"38",
          3886 => x"b3",
          3887 => x"dc",
          3888 => x"58",
          3889 => x"82",
          3890 => x"25",
          3891 => x"8c",
          3892 => x"05",
          3893 => x"55",
          3894 => x"74",
          3895 => x"70",
          3896 => x"2a",
          3897 => x"78",
          3898 => x"38",
          3899 => x"38",
          3900 => x"08",
          3901 => x"53",
          3902 => x"aa",
          3903 => x"dc",
          3904 => x"88",
          3905 => x"fc",
          3906 => x"3f",
          3907 => x"09",
          3908 => x"38",
          3909 => x"51",
          3910 => x"79",
          3911 => x"3f",
          3912 => x"54",
          3913 => x"08",
          3914 => x"58",
          3915 => x"dc",
          3916 => x"0d",
          3917 => x"0d",
          3918 => x"5c",
          3919 => x"57",
          3920 => x"73",
          3921 => x"81",
          3922 => x"78",
          3923 => x"56",
          3924 => x"98",
          3925 => x"70",
          3926 => x"33",
          3927 => x"73",
          3928 => x"81",
          3929 => x"75",
          3930 => x"38",
          3931 => x"88",
          3932 => x"ac",
          3933 => x"52",
          3934 => x"3f",
          3935 => x"08",
          3936 => x"74",
          3937 => x"c8",
          3938 => x"dc",
          3939 => x"38",
          3940 => x"55",
          3941 => x"88",
          3942 => x"2e",
          3943 => x"39",
          3944 => x"ab",
          3945 => x"5a",
          3946 => x"11",
          3947 => x"51",
          3948 => x"82",
          3949 => x"80",
          3950 => x"7a",
          3951 => x"77",
          3952 => x"3f",
          3953 => x"08",
          3954 => x"55",
          3955 => x"74",
          3956 => x"81",
          3957 => x"ff",
          3958 => x"82",
          3959 => x"8e",
          3960 => x"73",
          3961 => x"0c",
          3962 => x"04",
          3963 => x"b0",
          3964 => x"84",
          3965 => x"05",
          3966 => x"80",
          3967 => x"34",
          3968 => x"33",
          3969 => x"a4",
          3970 => x"38",
          3971 => x"33",
          3972 => x"9a",
          3973 => x"eb",
          3974 => x"8c",
          3975 => x"89",
          3976 => x"8c",
          3977 => x"2e",
          3978 => x"93",
          3979 => x"cc",
          3980 => x"8c",
          3981 => x"bb",
          3982 => x"8c",
          3983 => x"2e",
          3984 => x"f8",
          3985 => x"a4",
          3986 => x"39",
          3987 => x"08",
          3988 => x"52",
          3989 => x"52",
          3990 => x"b0",
          3991 => x"dc",
          3992 => x"8c",
          3993 => x"2e",
          3994 => x"80",
          3995 => x"8c",
          3996 => x"d3",
          3997 => x"8c",
          3998 => x"80",
          3999 => x"dc",
          4000 => x"38",
          4001 => x"08",
          4002 => x"17",
          4003 => x"74",
          4004 => x"74",
          4005 => x"52",
          4006 => x"b4",
          4007 => x"2e",
          4008 => x"ff",
          4009 => x"39",
          4010 => x"89",
          4011 => x"3d",
          4012 => x"3f",
          4013 => x"08",
          4014 => x"98",
          4015 => x"78",
          4016 => x"38",
          4017 => x"06",
          4018 => x"33",
          4019 => x"70",
          4020 => x"8c",
          4021 => x"98",
          4022 => x"2c",
          4023 => x"05",
          4024 => x"81",
          4025 => x"70",
          4026 => x"33",
          4027 => x"51",
          4028 => x"59",
          4029 => x"56",
          4030 => x"80",
          4031 => x"74",
          4032 => x"74",
          4033 => x"29",
          4034 => x"05",
          4035 => x"51",
          4036 => x"24",
          4037 => x"76",
          4038 => x"77",
          4039 => x"3f",
          4040 => x"08",
          4041 => x"54",
          4042 => x"d7",
          4043 => x"8c",
          4044 => x"56",
          4045 => x"81",
          4046 => x"81",
          4047 => x"70",
          4048 => x"81",
          4049 => x"51",
          4050 => x"26",
          4051 => x"53",
          4052 => x"51",
          4053 => x"82",
          4054 => x"81",
          4055 => x"73",
          4056 => x"39",
          4057 => x"80",
          4058 => x"38",
          4059 => x"74",
          4060 => x"34",
          4061 => x"70",
          4062 => x"8c",
          4063 => x"98",
          4064 => x"2c",
          4065 => x"70",
          4066 => x"f8",
          4067 => x"5e",
          4068 => x"57",
          4069 => x"74",
          4070 => x"81",
          4071 => x"38",
          4072 => x"14",
          4073 => x"80",
          4074 => x"80",
          4075 => x"82",
          4076 => x"92",
          4077 => x"8d",
          4078 => x"82",
          4079 => x"78",
          4080 => x"75",
          4081 => x"54",
          4082 => x"fd",
          4083 => x"84",
          4084 => x"e4",
          4085 => x"08",
          4086 => x"88",
          4087 => x"7e",
          4088 => x"38",
          4089 => x"33",
          4090 => x"27",
          4091 => x"98",
          4092 => x"2c",
          4093 => x"75",
          4094 => x"74",
          4095 => x"33",
          4096 => x"74",
          4097 => x"29",
          4098 => x"05",
          4099 => x"82",
          4100 => x"56",
          4101 => x"39",
          4102 => x"33",
          4103 => x"54",
          4104 => x"88",
          4105 => x"54",
          4106 => x"74",
          4107 => x"84",
          4108 => x"7e",
          4109 => x"81",
          4110 => x"82",
          4111 => x"82",
          4112 => x"70",
          4113 => x"29",
          4114 => x"05",
          4115 => x"82",
          4116 => x"5a",
          4117 => x"74",
          4118 => x"38",
          4119 => x"33",
          4120 => x"c7",
          4121 => x"80",
          4122 => x"80",
          4123 => x"98",
          4124 => x"84",
          4125 => x"55",
          4126 => x"e0",
          4127 => x"88",
          4128 => x"2b",
          4129 => x"82",
          4130 => x"5a",
          4131 => x"74",
          4132 => x"9a",
          4133 => x"e8",
          4134 => x"81",
          4135 => x"81",
          4136 => x"70",
          4137 => x"8d",
          4138 => x"51",
          4139 => x"24",
          4140 => x"fa",
          4141 => x"88",
          4142 => x"ff",
          4143 => x"73",
          4144 => x"ea",
          4145 => x"84",
          4146 => x"54",
          4147 => x"84",
          4148 => x"54",
          4149 => x"88",
          4150 => x"e7",
          4151 => x"8d",
          4152 => x"98",
          4153 => x"2c",
          4154 => x"33",
          4155 => x"57",
          4156 => x"a7",
          4157 => x"54",
          4158 => x"74",
          4159 => x"51",
          4160 => x"74",
          4161 => x"29",
          4162 => x"05",
          4163 => x"82",
          4164 => x"58",
          4165 => x"75",
          4166 => x"a0",
          4167 => x"3f",
          4168 => x"33",
          4169 => x"70",
          4170 => x"8d",
          4171 => x"51",
          4172 => x"74",
          4173 => x"38",
          4174 => x"ef",
          4175 => x"80",
          4176 => x"80",
          4177 => x"98",
          4178 => x"84",
          4179 => x"55",
          4180 => x"e4",
          4181 => x"39",
          4182 => x"33",
          4183 => x"80",
          4184 => x"51",
          4185 => x"82",
          4186 => x"79",
          4187 => x"3f",
          4188 => x"08",
          4189 => x"54",
          4190 => x"82",
          4191 => x"54",
          4192 => x"84",
          4193 => x"53",
          4194 => x"51",
          4195 => x"84",
          4196 => x"7a",
          4197 => x"39",
          4198 => x"33",
          4199 => x"2e",
          4200 => x"88",
          4201 => x"3f",
          4202 => x"33",
          4203 => x"73",
          4204 => x"34",
          4205 => x"06",
          4206 => x"82",
          4207 => x"82",
          4208 => x"55",
          4209 => x"2e",
          4210 => x"ff",
          4211 => x"82",
          4212 => x"74",
          4213 => x"98",
          4214 => x"ff",
          4215 => x"55",
          4216 => x"a7",
          4217 => x"54",
          4218 => x"74",
          4219 => x"51",
          4220 => x"74",
          4221 => x"29",
          4222 => x"05",
          4223 => x"82",
          4224 => x"58",
          4225 => x"75",
          4226 => x"a0",
          4227 => x"3f",
          4228 => x"33",
          4229 => x"70",
          4230 => x"8d",
          4231 => x"51",
          4232 => x"74",
          4233 => x"38",
          4234 => x"ff",
          4235 => x"80",
          4236 => x"80",
          4237 => x"98",
          4238 => x"84",
          4239 => x"55",
          4240 => x"e4",
          4241 => x"39",
          4242 => x"33",
          4243 => x"06",
          4244 => x"33",
          4245 => x"74",
          4246 => x"d2",
          4247 => x"54",
          4248 => x"88",
          4249 => x"70",
          4250 => x"e4",
          4251 => x"8d",
          4252 => x"81",
          4253 => x"8d",
          4254 => x"56",
          4255 => x"26",
          4256 => x"aa",
          4257 => x"38",
          4258 => x"08",
          4259 => x"2e",
          4260 => x"51",
          4261 => x"82",
          4262 => x"82",
          4263 => x"82",
          4264 => x"81",
          4265 => x"05",
          4266 => x"79",
          4267 => x"3f",
          4268 => x"c1",
          4269 => x"29",
          4270 => x"05",
          4271 => x"56",
          4272 => x"2e",
          4273 => x"51",
          4274 => x"82",
          4275 => x"82",
          4276 => x"82",
          4277 => x"81",
          4278 => x"05",
          4279 => x"79",
          4280 => x"3f",
          4281 => x"80",
          4282 => x"08",
          4283 => x"2e",
          4284 => x"74",
          4285 => x"3f",
          4286 => x"7a",
          4287 => x"81",
          4288 => x"82",
          4289 => x"55",
          4290 => x"89",
          4291 => x"ca",
          4292 => x"c8",
          4293 => x"29",
          4294 => x"05",
          4295 => x"56",
          4296 => x"2e",
          4297 => x"51",
          4298 => x"82",
          4299 => x"82",
          4300 => x"82",
          4301 => x"81",
          4302 => x"05",
          4303 => x"79",
          4304 => x"3f",
          4305 => x"73",
          4306 => x"5b",
          4307 => x"08",
          4308 => x"2e",
          4309 => x"74",
          4310 => x"3f",
          4311 => x"08",
          4312 => x"34",
          4313 => x"08",
          4314 => x"81",
          4315 => x"52",
          4316 => x"e0",
          4317 => x"88",
          4318 => x"84",
          4319 => x"51",
          4320 => x"f6",
          4321 => x"8d",
          4322 => x"81",
          4323 => x"8d",
          4324 => x"56",
          4325 => x"27",
          4326 => x"81",
          4327 => x"82",
          4328 => x"74",
          4329 => x"52",
          4330 => x"3f",
          4331 => x"82",
          4332 => x"54",
          4333 => x"f5",
          4334 => x"51",
          4335 => x"82",
          4336 => x"ff",
          4337 => x"82",
          4338 => x"f5",
          4339 => x"0b",
          4340 => x"34",
          4341 => x"8d",
          4342 => x"82",
          4343 => x"af",
          4344 => x"ff",
          4345 => x"8f",
          4346 => x"81",
          4347 => x"26",
          4348 => x"89",
          4349 => x"52",
          4350 => x"dc",
          4351 => x"0d",
          4352 => x"0d",
          4353 => x"33",
          4354 => x"9f",
          4355 => x"53",
          4356 => x"81",
          4357 => x"38",
          4358 => x"87",
          4359 => x"11",
          4360 => x"54",
          4361 => x"84",
          4362 => x"54",
          4363 => x"87",
          4364 => x"11",
          4365 => x"0c",
          4366 => x"c0",
          4367 => x"70",
          4368 => x"70",
          4369 => x"51",
          4370 => x"8a",
          4371 => x"98",
          4372 => x"70",
          4373 => x"08",
          4374 => x"06",
          4375 => x"38",
          4376 => x"8c",
          4377 => x"80",
          4378 => x"71",
          4379 => x"14",
          4380 => x"c4",
          4381 => x"70",
          4382 => x"0c",
          4383 => x"04",
          4384 => x"60",
          4385 => x"8c",
          4386 => x"33",
          4387 => x"5b",
          4388 => x"5a",
          4389 => x"82",
          4390 => x"81",
          4391 => x"52",
          4392 => x"38",
          4393 => x"84",
          4394 => x"92",
          4395 => x"c0",
          4396 => x"87",
          4397 => x"13",
          4398 => x"57",
          4399 => x"0b",
          4400 => x"8c",
          4401 => x"0c",
          4402 => x"75",
          4403 => x"2a",
          4404 => x"51",
          4405 => x"80",
          4406 => x"7b",
          4407 => x"7b",
          4408 => x"5d",
          4409 => x"59",
          4410 => x"06",
          4411 => x"73",
          4412 => x"81",
          4413 => x"ff",
          4414 => x"72",
          4415 => x"38",
          4416 => x"8c",
          4417 => x"c3",
          4418 => x"98",
          4419 => x"71",
          4420 => x"38",
          4421 => x"2e",
          4422 => x"76",
          4423 => x"92",
          4424 => x"72",
          4425 => x"06",
          4426 => x"f7",
          4427 => x"5a",
          4428 => x"80",
          4429 => x"70",
          4430 => x"5a",
          4431 => x"80",
          4432 => x"73",
          4433 => x"06",
          4434 => x"38",
          4435 => x"fe",
          4436 => x"fc",
          4437 => x"52",
          4438 => x"83",
          4439 => x"71",
          4440 => x"8c",
          4441 => x"3d",
          4442 => x"3d",
          4443 => x"64",
          4444 => x"bf",
          4445 => x"40",
          4446 => x"59",
          4447 => x"58",
          4448 => x"82",
          4449 => x"81",
          4450 => x"52",
          4451 => x"09",
          4452 => x"b1",
          4453 => x"84",
          4454 => x"92",
          4455 => x"c0",
          4456 => x"87",
          4457 => x"13",
          4458 => x"56",
          4459 => x"87",
          4460 => x"0c",
          4461 => x"82",
          4462 => x"58",
          4463 => x"84",
          4464 => x"06",
          4465 => x"71",
          4466 => x"38",
          4467 => x"05",
          4468 => x"0c",
          4469 => x"73",
          4470 => x"81",
          4471 => x"71",
          4472 => x"38",
          4473 => x"8c",
          4474 => x"d0",
          4475 => x"98",
          4476 => x"71",
          4477 => x"38",
          4478 => x"2e",
          4479 => x"76",
          4480 => x"92",
          4481 => x"72",
          4482 => x"06",
          4483 => x"f7",
          4484 => x"59",
          4485 => x"1a",
          4486 => x"06",
          4487 => x"59",
          4488 => x"80",
          4489 => x"73",
          4490 => x"06",
          4491 => x"38",
          4492 => x"fe",
          4493 => x"fc",
          4494 => x"52",
          4495 => x"83",
          4496 => x"71",
          4497 => x"8c",
          4498 => x"3d",
          4499 => x"3d",
          4500 => x"84",
          4501 => x"33",
          4502 => x"a7",
          4503 => x"54",
          4504 => x"fa",
          4505 => x"8c",
          4506 => x"06",
          4507 => x"72",
          4508 => x"85",
          4509 => x"98",
          4510 => x"56",
          4511 => x"80",
          4512 => x"76",
          4513 => x"74",
          4514 => x"c0",
          4515 => x"54",
          4516 => x"2e",
          4517 => x"d4",
          4518 => x"2e",
          4519 => x"80",
          4520 => x"08",
          4521 => x"70",
          4522 => x"51",
          4523 => x"2e",
          4524 => x"c0",
          4525 => x"52",
          4526 => x"87",
          4527 => x"08",
          4528 => x"38",
          4529 => x"87",
          4530 => x"14",
          4531 => x"70",
          4532 => x"52",
          4533 => x"96",
          4534 => x"92",
          4535 => x"0a",
          4536 => x"39",
          4537 => x"0c",
          4538 => x"39",
          4539 => x"54",
          4540 => x"dc",
          4541 => x"0d",
          4542 => x"0d",
          4543 => x"33",
          4544 => x"88",
          4545 => x"8c",
          4546 => x"51",
          4547 => x"04",
          4548 => x"75",
          4549 => x"82",
          4550 => x"90",
          4551 => x"2b",
          4552 => x"33",
          4553 => x"88",
          4554 => x"71",
          4555 => x"dc",
          4556 => x"54",
          4557 => x"85",
          4558 => x"ff",
          4559 => x"02",
          4560 => x"05",
          4561 => x"70",
          4562 => x"05",
          4563 => x"88",
          4564 => x"72",
          4565 => x"0d",
          4566 => x"0d",
          4567 => x"52",
          4568 => x"81",
          4569 => x"70",
          4570 => x"70",
          4571 => x"05",
          4572 => x"88",
          4573 => x"72",
          4574 => x"54",
          4575 => x"2a",
          4576 => x"34",
          4577 => x"04",
          4578 => x"76",
          4579 => x"54",
          4580 => x"2e",
          4581 => x"70",
          4582 => x"33",
          4583 => x"05",
          4584 => x"11",
          4585 => x"84",
          4586 => x"fe",
          4587 => x"77",
          4588 => x"53",
          4589 => x"81",
          4590 => x"ff",
          4591 => x"f4",
          4592 => x"0d",
          4593 => x"0d",
          4594 => x"56",
          4595 => x"70",
          4596 => x"33",
          4597 => x"05",
          4598 => x"71",
          4599 => x"56",
          4600 => x"72",
          4601 => x"38",
          4602 => x"e2",
          4603 => x"8c",
          4604 => x"3d",
          4605 => x"3d",
          4606 => x"54",
          4607 => x"71",
          4608 => x"38",
          4609 => x"70",
          4610 => x"f3",
          4611 => x"82",
          4612 => x"84",
          4613 => x"80",
          4614 => x"dc",
          4615 => x"0b",
          4616 => x"0c",
          4617 => x"0d",
          4618 => x"0b",
          4619 => x"56",
          4620 => x"2e",
          4621 => x"81",
          4622 => x"08",
          4623 => x"70",
          4624 => x"33",
          4625 => x"a2",
          4626 => x"dc",
          4627 => x"09",
          4628 => x"38",
          4629 => x"08",
          4630 => x"b0",
          4631 => x"a4",
          4632 => x"9c",
          4633 => x"56",
          4634 => x"27",
          4635 => x"16",
          4636 => x"82",
          4637 => x"06",
          4638 => x"54",
          4639 => x"78",
          4640 => x"33",
          4641 => x"3f",
          4642 => x"5a",
          4643 => x"dc",
          4644 => x"0d",
          4645 => x"0d",
          4646 => x"56",
          4647 => x"b0",
          4648 => x"af",
          4649 => x"fe",
          4650 => x"8c",
          4651 => x"82",
          4652 => x"9f",
          4653 => x"74",
          4654 => x"52",
          4655 => x"51",
          4656 => x"82",
          4657 => x"80",
          4658 => x"ff",
          4659 => x"74",
          4660 => x"76",
          4661 => x"0c",
          4662 => x"04",
          4663 => x"7a",
          4664 => x"fe",
          4665 => x"8c",
          4666 => x"82",
          4667 => x"81",
          4668 => x"33",
          4669 => x"2e",
          4670 => x"80",
          4671 => x"17",
          4672 => x"81",
          4673 => x"06",
          4674 => x"84",
          4675 => x"8c",
          4676 => x"b4",
          4677 => x"56",
          4678 => x"82",
          4679 => x"84",
          4680 => x"fc",
          4681 => x"8b",
          4682 => x"52",
          4683 => x"a9",
          4684 => x"85",
          4685 => x"84",
          4686 => x"fc",
          4687 => x"17",
          4688 => x"9c",
          4689 => x"91",
          4690 => x"08",
          4691 => x"17",
          4692 => x"3f",
          4693 => x"81",
          4694 => x"19",
          4695 => x"53",
          4696 => x"17",
          4697 => x"82",
          4698 => x"18",
          4699 => x"80",
          4700 => x"33",
          4701 => x"3f",
          4702 => x"08",
          4703 => x"38",
          4704 => x"82",
          4705 => x"8a",
          4706 => x"fb",
          4707 => x"fe",
          4708 => x"08",
          4709 => x"56",
          4710 => x"74",
          4711 => x"38",
          4712 => x"75",
          4713 => x"16",
          4714 => x"53",
          4715 => x"dc",
          4716 => x"0d",
          4717 => x"0d",
          4718 => x"08",
          4719 => x"81",
          4720 => x"df",
          4721 => x"15",
          4722 => x"d7",
          4723 => x"33",
          4724 => x"82",
          4725 => x"38",
          4726 => x"89",
          4727 => x"2e",
          4728 => x"bf",
          4729 => x"2e",
          4730 => x"81",
          4731 => x"81",
          4732 => x"89",
          4733 => x"08",
          4734 => x"52",
          4735 => x"3f",
          4736 => x"08",
          4737 => x"74",
          4738 => x"14",
          4739 => x"81",
          4740 => x"2a",
          4741 => x"05",
          4742 => x"57",
          4743 => x"f5",
          4744 => x"dc",
          4745 => x"38",
          4746 => x"06",
          4747 => x"33",
          4748 => x"78",
          4749 => x"06",
          4750 => x"5c",
          4751 => x"53",
          4752 => x"38",
          4753 => x"06",
          4754 => x"39",
          4755 => x"a4",
          4756 => x"52",
          4757 => x"bd",
          4758 => x"dc",
          4759 => x"38",
          4760 => x"fe",
          4761 => x"b4",
          4762 => x"8d",
          4763 => x"dc",
          4764 => x"ff",
          4765 => x"39",
          4766 => x"a4",
          4767 => x"52",
          4768 => x"91",
          4769 => x"dc",
          4770 => x"76",
          4771 => x"fc",
          4772 => x"b4",
          4773 => x"f8",
          4774 => x"dc",
          4775 => x"06",
          4776 => x"81",
          4777 => x"8c",
          4778 => x"3d",
          4779 => x"3d",
          4780 => x"7e",
          4781 => x"82",
          4782 => x"27",
          4783 => x"76",
          4784 => x"27",
          4785 => x"75",
          4786 => x"79",
          4787 => x"38",
          4788 => x"89",
          4789 => x"2e",
          4790 => x"80",
          4791 => x"2e",
          4792 => x"81",
          4793 => x"81",
          4794 => x"89",
          4795 => x"08",
          4796 => x"52",
          4797 => x"3f",
          4798 => x"08",
          4799 => x"dc",
          4800 => x"38",
          4801 => x"06",
          4802 => x"81",
          4803 => x"06",
          4804 => x"77",
          4805 => x"2e",
          4806 => x"84",
          4807 => x"06",
          4808 => x"06",
          4809 => x"53",
          4810 => x"81",
          4811 => x"34",
          4812 => x"a4",
          4813 => x"52",
          4814 => x"d9",
          4815 => x"dc",
          4816 => x"8c",
          4817 => x"94",
          4818 => x"ff",
          4819 => x"05",
          4820 => x"54",
          4821 => x"38",
          4822 => x"74",
          4823 => x"06",
          4824 => x"07",
          4825 => x"74",
          4826 => x"39",
          4827 => x"a4",
          4828 => x"52",
          4829 => x"9d",
          4830 => x"dc",
          4831 => x"8c",
          4832 => x"d8",
          4833 => x"ff",
          4834 => x"76",
          4835 => x"06",
          4836 => x"05",
          4837 => x"3f",
          4838 => x"87",
          4839 => x"08",
          4840 => x"51",
          4841 => x"82",
          4842 => x"59",
          4843 => x"08",
          4844 => x"f0",
          4845 => x"82",
          4846 => x"06",
          4847 => x"05",
          4848 => x"54",
          4849 => x"3f",
          4850 => x"08",
          4851 => x"74",
          4852 => x"51",
          4853 => x"81",
          4854 => x"34",
          4855 => x"dc",
          4856 => x"0d",
          4857 => x"0d",
          4858 => x"72",
          4859 => x"56",
          4860 => x"27",
          4861 => x"98",
          4862 => x"9d",
          4863 => x"2e",
          4864 => x"53",
          4865 => x"51",
          4866 => x"82",
          4867 => x"54",
          4868 => x"08",
          4869 => x"93",
          4870 => x"80",
          4871 => x"54",
          4872 => x"82",
          4873 => x"54",
          4874 => x"74",
          4875 => x"fb",
          4876 => x"8c",
          4877 => x"82",
          4878 => x"80",
          4879 => x"38",
          4880 => x"08",
          4881 => x"38",
          4882 => x"08",
          4883 => x"38",
          4884 => x"52",
          4885 => x"d6",
          4886 => x"dc",
          4887 => x"98",
          4888 => x"11",
          4889 => x"57",
          4890 => x"74",
          4891 => x"81",
          4892 => x"0c",
          4893 => x"81",
          4894 => x"84",
          4895 => x"55",
          4896 => x"ff",
          4897 => x"54",
          4898 => x"dc",
          4899 => x"0d",
          4900 => x"0d",
          4901 => x"08",
          4902 => x"79",
          4903 => x"17",
          4904 => x"80",
          4905 => x"98",
          4906 => x"26",
          4907 => x"58",
          4908 => x"52",
          4909 => x"fd",
          4910 => x"74",
          4911 => x"08",
          4912 => x"38",
          4913 => x"08",
          4914 => x"dc",
          4915 => x"82",
          4916 => x"17",
          4917 => x"dc",
          4918 => x"c7",
          4919 => x"90",
          4920 => x"56",
          4921 => x"2e",
          4922 => x"77",
          4923 => x"81",
          4924 => x"38",
          4925 => x"98",
          4926 => x"26",
          4927 => x"56",
          4928 => x"51",
          4929 => x"80",
          4930 => x"dc",
          4931 => x"09",
          4932 => x"38",
          4933 => x"08",
          4934 => x"dc",
          4935 => x"30",
          4936 => x"80",
          4937 => x"07",
          4938 => x"08",
          4939 => x"55",
          4940 => x"ef",
          4941 => x"dc",
          4942 => x"95",
          4943 => x"08",
          4944 => x"27",
          4945 => x"98",
          4946 => x"89",
          4947 => x"85",
          4948 => x"db",
          4949 => x"81",
          4950 => x"17",
          4951 => x"89",
          4952 => x"75",
          4953 => x"ac",
          4954 => x"7a",
          4955 => x"3f",
          4956 => x"08",
          4957 => x"38",
          4958 => x"8c",
          4959 => x"2e",
          4960 => x"86",
          4961 => x"dc",
          4962 => x"8c",
          4963 => x"70",
          4964 => x"07",
          4965 => x"7c",
          4966 => x"55",
          4967 => x"f8",
          4968 => x"2e",
          4969 => x"ff",
          4970 => x"55",
          4971 => x"ff",
          4972 => x"76",
          4973 => x"3f",
          4974 => x"08",
          4975 => x"08",
          4976 => x"8c",
          4977 => x"80",
          4978 => x"55",
          4979 => x"94",
          4980 => x"2e",
          4981 => x"53",
          4982 => x"51",
          4983 => x"82",
          4984 => x"55",
          4985 => x"75",
          4986 => x"98",
          4987 => x"05",
          4988 => x"56",
          4989 => x"26",
          4990 => x"15",
          4991 => x"84",
          4992 => x"07",
          4993 => x"18",
          4994 => x"ff",
          4995 => x"2e",
          4996 => x"39",
          4997 => x"39",
          4998 => x"08",
          4999 => x"81",
          5000 => x"74",
          5001 => x"0c",
          5002 => x"04",
          5003 => x"7a",
          5004 => x"f3",
          5005 => x"8c",
          5006 => x"81",
          5007 => x"dc",
          5008 => x"38",
          5009 => x"51",
          5010 => x"82",
          5011 => x"82",
          5012 => x"b0",
          5013 => x"84",
          5014 => x"52",
          5015 => x"52",
          5016 => x"3f",
          5017 => x"39",
          5018 => x"8a",
          5019 => x"75",
          5020 => x"38",
          5021 => x"19",
          5022 => x"81",
          5023 => x"ed",
          5024 => x"8c",
          5025 => x"2e",
          5026 => x"15",
          5027 => x"70",
          5028 => x"07",
          5029 => x"53",
          5030 => x"75",
          5031 => x"0c",
          5032 => x"04",
          5033 => x"7a",
          5034 => x"58",
          5035 => x"f0",
          5036 => x"80",
          5037 => x"9f",
          5038 => x"80",
          5039 => x"90",
          5040 => x"17",
          5041 => x"aa",
          5042 => x"53",
          5043 => x"88",
          5044 => x"08",
          5045 => x"38",
          5046 => x"53",
          5047 => x"17",
          5048 => x"72",
          5049 => x"fe",
          5050 => x"08",
          5051 => x"80",
          5052 => x"16",
          5053 => x"2b",
          5054 => x"75",
          5055 => x"73",
          5056 => x"f5",
          5057 => x"8c",
          5058 => x"82",
          5059 => x"ff",
          5060 => x"81",
          5061 => x"dc",
          5062 => x"38",
          5063 => x"82",
          5064 => x"26",
          5065 => x"58",
          5066 => x"73",
          5067 => x"39",
          5068 => x"51",
          5069 => x"82",
          5070 => x"98",
          5071 => x"94",
          5072 => x"17",
          5073 => x"58",
          5074 => x"9a",
          5075 => x"81",
          5076 => x"74",
          5077 => x"98",
          5078 => x"83",
          5079 => x"b4",
          5080 => x"0c",
          5081 => x"82",
          5082 => x"8a",
          5083 => x"f8",
          5084 => x"70",
          5085 => x"08",
          5086 => x"57",
          5087 => x"0a",
          5088 => x"38",
          5089 => x"15",
          5090 => x"08",
          5091 => x"72",
          5092 => x"cb",
          5093 => x"ff",
          5094 => x"81",
          5095 => x"13",
          5096 => x"94",
          5097 => x"74",
          5098 => x"85",
          5099 => x"22",
          5100 => x"73",
          5101 => x"38",
          5102 => x"8a",
          5103 => x"05",
          5104 => x"06",
          5105 => x"8a",
          5106 => x"73",
          5107 => x"3f",
          5108 => x"08",
          5109 => x"81",
          5110 => x"dc",
          5111 => x"ff",
          5112 => x"82",
          5113 => x"ff",
          5114 => x"38",
          5115 => x"82",
          5116 => x"26",
          5117 => x"7b",
          5118 => x"98",
          5119 => x"55",
          5120 => x"94",
          5121 => x"73",
          5122 => x"3f",
          5123 => x"08",
          5124 => x"82",
          5125 => x"80",
          5126 => x"38",
          5127 => x"8c",
          5128 => x"2e",
          5129 => x"55",
          5130 => x"08",
          5131 => x"38",
          5132 => x"08",
          5133 => x"fb",
          5134 => x"8c",
          5135 => x"38",
          5136 => x"0c",
          5137 => x"51",
          5138 => x"82",
          5139 => x"98",
          5140 => x"90",
          5141 => x"16",
          5142 => x"15",
          5143 => x"74",
          5144 => x"0c",
          5145 => x"04",
          5146 => x"7b",
          5147 => x"5b",
          5148 => x"52",
          5149 => x"ac",
          5150 => x"dc",
          5151 => x"8c",
          5152 => x"ec",
          5153 => x"dc",
          5154 => x"17",
          5155 => x"51",
          5156 => x"82",
          5157 => x"54",
          5158 => x"08",
          5159 => x"82",
          5160 => x"9c",
          5161 => x"33",
          5162 => x"72",
          5163 => x"09",
          5164 => x"38",
          5165 => x"8c",
          5166 => x"72",
          5167 => x"55",
          5168 => x"53",
          5169 => x"8e",
          5170 => x"56",
          5171 => x"09",
          5172 => x"38",
          5173 => x"8c",
          5174 => x"81",
          5175 => x"fd",
          5176 => x"8c",
          5177 => x"82",
          5178 => x"80",
          5179 => x"38",
          5180 => x"09",
          5181 => x"38",
          5182 => x"82",
          5183 => x"8b",
          5184 => x"fd",
          5185 => x"9a",
          5186 => x"eb",
          5187 => x"8c",
          5188 => x"ff",
          5189 => x"70",
          5190 => x"53",
          5191 => x"09",
          5192 => x"38",
          5193 => x"eb",
          5194 => x"8c",
          5195 => x"2b",
          5196 => x"72",
          5197 => x"0c",
          5198 => x"04",
          5199 => x"77",
          5200 => x"ff",
          5201 => x"9a",
          5202 => x"55",
          5203 => x"76",
          5204 => x"53",
          5205 => x"09",
          5206 => x"38",
          5207 => x"52",
          5208 => x"eb",
          5209 => x"3d",
          5210 => x"3d",
          5211 => x"5b",
          5212 => x"08",
          5213 => x"15",
          5214 => x"81",
          5215 => x"15",
          5216 => x"51",
          5217 => x"82",
          5218 => x"58",
          5219 => x"08",
          5220 => x"9c",
          5221 => x"33",
          5222 => x"86",
          5223 => x"80",
          5224 => x"13",
          5225 => x"06",
          5226 => x"06",
          5227 => x"72",
          5228 => x"82",
          5229 => x"53",
          5230 => x"2e",
          5231 => x"53",
          5232 => x"a9",
          5233 => x"74",
          5234 => x"72",
          5235 => x"38",
          5236 => x"99",
          5237 => x"dc",
          5238 => x"06",
          5239 => x"88",
          5240 => x"06",
          5241 => x"54",
          5242 => x"a0",
          5243 => x"74",
          5244 => x"3f",
          5245 => x"08",
          5246 => x"dc",
          5247 => x"98",
          5248 => x"fa",
          5249 => x"80",
          5250 => x"0c",
          5251 => x"dc",
          5252 => x"0d",
          5253 => x"0d",
          5254 => x"57",
          5255 => x"73",
          5256 => x"3f",
          5257 => x"08",
          5258 => x"dc",
          5259 => x"98",
          5260 => x"75",
          5261 => x"3f",
          5262 => x"08",
          5263 => x"dc",
          5264 => x"a0",
          5265 => x"dc",
          5266 => x"14",
          5267 => x"db",
          5268 => x"a0",
          5269 => x"14",
          5270 => x"ac",
          5271 => x"83",
          5272 => x"82",
          5273 => x"87",
          5274 => x"fd",
          5275 => x"70",
          5276 => x"08",
          5277 => x"55",
          5278 => x"3f",
          5279 => x"08",
          5280 => x"13",
          5281 => x"73",
          5282 => x"83",
          5283 => x"3d",
          5284 => x"3d",
          5285 => x"57",
          5286 => x"89",
          5287 => x"17",
          5288 => x"81",
          5289 => x"70",
          5290 => x"55",
          5291 => x"08",
          5292 => x"81",
          5293 => x"52",
          5294 => x"a8",
          5295 => x"2e",
          5296 => x"84",
          5297 => x"52",
          5298 => x"09",
          5299 => x"38",
          5300 => x"81",
          5301 => x"81",
          5302 => x"73",
          5303 => x"55",
          5304 => x"55",
          5305 => x"c5",
          5306 => x"88",
          5307 => x"0b",
          5308 => x"9c",
          5309 => x"8b",
          5310 => x"17",
          5311 => x"08",
          5312 => x"52",
          5313 => x"82",
          5314 => x"76",
          5315 => x"51",
          5316 => x"82",
          5317 => x"86",
          5318 => x"12",
          5319 => x"3f",
          5320 => x"08",
          5321 => x"88",
          5322 => x"f3",
          5323 => x"70",
          5324 => x"80",
          5325 => x"51",
          5326 => x"af",
          5327 => x"81",
          5328 => x"dc",
          5329 => x"74",
          5330 => x"38",
          5331 => x"88",
          5332 => x"39",
          5333 => x"80",
          5334 => x"56",
          5335 => x"af",
          5336 => x"06",
          5337 => x"56",
          5338 => x"32",
          5339 => x"80",
          5340 => x"51",
          5341 => x"dc",
          5342 => x"1c",
          5343 => x"33",
          5344 => x"9f",
          5345 => x"ff",
          5346 => x"1c",
          5347 => x"7a",
          5348 => x"3f",
          5349 => x"08",
          5350 => x"39",
          5351 => x"a0",
          5352 => x"5e",
          5353 => x"52",
          5354 => x"ff",
          5355 => x"59",
          5356 => x"33",
          5357 => x"ae",
          5358 => x"06",
          5359 => x"78",
          5360 => x"81",
          5361 => x"32",
          5362 => x"9f",
          5363 => x"26",
          5364 => x"53",
          5365 => x"73",
          5366 => x"17",
          5367 => x"34",
          5368 => x"db",
          5369 => x"32",
          5370 => x"9f",
          5371 => x"54",
          5372 => x"2e",
          5373 => x"80",
          5374 => x"75",
          5375 => x"bd",
          5376 => x"7e",
          5377 => x"a0",
          5378 => x"bd",
          5379 => x"82",
          5380 => x"18",
          5381 => x"1a",
          5382 => x"a0",
          5383 => x"fc",
          5384 => x"32",
          5385 => x"80",
          5386 => x"30",
          5387 => x"71",
          5388 => x"51",
          5389 => x"55",
          5390 => x"ac",
          5391 => x"81",
          5392 => x"78",
          5393 => x"51",
          5394 => x"af",
          5395 => x"06",
          5396 => x"55",
          5397 => x"32",
          5398 => x"80",
          5399 => x"51",
          5400 => x"db",
          5401 => x"39",
          5402 => x"09",
          5403 => x"38",
          5404 => x"7c",
          5405 => x"54",
          5406 => x"a2",
          5407 => x"32",
          5408 => x"ae",
          5409 => x"72",
          5410 => x"9f",
          5411 => x"51",
          5412 => x"74",
          5413 => x"88",
          5414 => x"fe",
          5415 => x"98",
          5416 => x"80",
          5417 => x"75",
          5418 => x"81",
          5419 => x"33",
          5420 => x"51",
          5421 => x"82",
          5422 => x"80",
          5423 => x"78",
          5424 => x"81",
          5425 => x"5a",
          5426 => x"d2",
          5427 => x"dc",
          5428 => x"80",
          5429 => x"1c",
          5430 => x"27",
          5431 => x"79",
          5432 => x"74",
          5433 => x"7a",
          5434 => x"74",
          5435 => x"39",
          5436 => x"fa",
          5437 => x"fe",
          5438 => x"dc",
          5439 => x"ff",
          5440 => x"73",
          5441 => x"38",
          5442 => x"81",
          5443 => x"54",
          5444 => x"75",
          5445 => x"17",
          5446 => x"39",
          5447 => x"0c",
          5448 => x"99",
          5449 => x"54",
          5450 => x"2e",
          5451 => x"84",
          5452 => x"34",
          5453 => x"76",
          5454 => x"8b",
          5455 => x"81",
          5456 => x"56",
          5457 => x"80",
          5458 => x"1b",
          5459 => x"08",
          5460 => x"51",
          5461 => x"82",
          5462 => x"56",
          5463 => x"08",
          5464 => x"98",
          5465 => x"76",
          5466 => x"3f",
          5467 => x"08",
          5468 => x"dc",
          5469 => x"38",
          5470 => x"70",
          5471 => x"73",
          5472 => x"be",
          5473 => x"33",
          5474 => x"73",
          5475 => x"8b",
          5476 => x"83",
          5477 => x"06",
          5478 => x"73",
          5479 => x"53",
          5480 => x"51",
          5481 => x"82",
          5482 => x"80",
          5483 => x"75",
          5484 => x"f3",
          5485 => x"9f",
          5486 => x"1c",
          5487 => x"74",
          5488 => x"38",
          5489 => x"09",
          5490 => x"e7",
          5491 => x"2a",
          5492 => x"77",
          5493 => x"51",
          5494 => x"2e",
          5495 => x"81",
          5496 => x"80",
          5497 => x"38",
          5498 => x"ab",
          5499 => x"55",
          5500 => x"75",
          5501 => x"73",
          5502 => x"55",
          5503 => x"82",
          5504 => x"06",
          5505 => x"ab",
          5506 => x"33",
          5507 => x"70",
          5508 => x"55",
          5509 => x"2e",
          5510 => x"1b",
          5511 => x"06",
          5512 => x"52",
          5513 => x"db",
          5514 => x"dc",
          5515 => x"0c",
          5516 => x"74",
          5517 => x"0c",
          5518 => x"04",
          5519 => x"7c",
          5520 => x"08",
          5521 => x"55",
          5522 => x"59",
          5523 => x"81",
          5524 => x"70",
          5525 => x"33",
          5526 => x"52",
          5527 => x"2e",
          5528 => x"ee",
          5529 => x"2e",
          5530 => x"81",
          5531 => x"33",
          5532 => x"81",
          5533 => x"52",
          5534 => x"26",
          5535 => x"14",
          5536 => x"06",
          5537 => x"52",
          5538 => x"80",
          5539 => x"0b",
          5540 => x"59",
          5541 => x"7a",
          5542 => x"70",
          5543 => x"33",
          5544 => x"05",
          5545 => x"9f",
          5546 => x"53",
          5547 => x"89",
          5548 => x"70",
          5549 => x"54",
          5550 => x"12",
          5551 => x"26",
          5552 => x"12",
          5553 => x"06",
          5554 => x"30",
          5555 => x"51",
          5556 => x"2e",
          5557 => x"85",
          5558 => x"be",
          5559 => x"74",
          5560 => x"30",
          5561 => x"9f",
          5562 => x"2a",
          5563 => x"54",
          5564 => x"2e",
          5565 => x"15",
          5566 => x"55",
          5567 => x"ff",
          5568 => x"39",
          5569 => x"86",
          5570 => x"7c",
          5571 => x"51",
          5572 => x"8d",
          5573 => x"70",
          5574 => x"0c",
          5575 => x"04",
          5576 => x"78",
          5577 => x"83",
          5578 => x"0b",
          5579 => x"79",
          5580 => x"e2",
          5581 => x"55",
          5582 => x"08",
          5583 => x"84",
          5584 => x"df",
          5585 => x"8c",
          5586 => x"ff",
          5587 => x"83",
          5588 => x"d4",
          5589 => x"81",
          5590 => x"38",
          5591 => x"17",
          5592 => x"74",
          5593 => x"09",
          5594 => x"38",
          5595 => x"81",
          5596 => x"30",
          5597 => x"79",
          5598 => x"54",
          5599 => x"74",
          5600 => x"09",
          5601 => x"38",
          5602 => x"fa",
          5603 => x"ea",
          5604 => x"b1",
          5605 => x"dc",
          5606 => x"8c",
          5607 => x"2e",
          5608 => x"53",
          5609 => x"52",
          5610 => x"51",
          5611 => x"82",
          5612 => x"55",
          5613 => x"08",
          5614 => x"38",
          5615 => x"82",
          5616 => x"88",
          5617 => x"f2",
          5618 => x"02",
          5619 => x"cb",
          5620 => x"55",
          5621 => x"60",
          5622 => x"3f",
          5623 => x"08",
          5624 => x"80",
          5625 => x"dc",
          5626 => x"fc",
          5627 => x"dc",
          5628 => x"82",
          5629 => x"70",
          5630 => x"8c",
          5631 => x"2e",
          5632 => x"73",
          5633 => x"81",
          5634 => x"33",
          5635 => x"80",
          5636 => x"81",
          5637 => x"d7",
          5638 => x"8c",
          5639 => x"ff",
          5640 => x"06",
          5641 => x"98",
          5642 => x"2e",
          5643 => x"74",
          5644 => x"81",
          5645 => x"8a",
          5646 => x"ac",
          5647 => x"39",
          5648 => x"77",
          5649 => x"81",
          5650 => x"33",
          5651 => x"3f",
          5652 => x"08",
          5653 => x"70",
          5654 => x"55",
          5655 => x"86",
          5656 => x"80",
          5657 => x"74",
          5658 => x"81",
          5659 => x"8a",
          5660 => x"f4",
          5661 => x"53",
          5662 => x"fd",
          5663 => x"8c",
          5664 => x"ff",
          5665 => x"82",
          5666 => x"06",
          5667 => x"8c",
          5668 => x"58",
          5669 => x"f6",
          5670 => x"58",
          5671 => x"2e",
          5672 => x"fa",
          5673 => x"e8",
          5674 => x"dc",
          5675 => x"78",
          5676 => x"5a",
          5677 => x"90",
          5678 => x"75",
          5679 => x"38",
          5680 => x"3d",
          5681 => x"70",
          5682 => x"08",
          5683 => x"7a",
          5684 => x"38",
          5685 => x"51",
          5686 => x"82",
          5687 => x"81",
          5688 => x"81",
          5689 => x"38",
          5690 => x"83",
          5691 => x"38",
          5692 => x"84",
          5693 => x"38",
          5694 => x"81",
          5695 => x"38",
          5696 => x"db",
          5697 => x"8c",
          5698 => x"ff",
          5699 => x"72",
          5700 => x"09",
          5701 => x"d0",
          5702 => x"14",
          5703 => x"3f",
          5704 => x"08",
          5705 => x"06",
          5706 => x"38",
          5707 => x"51",
          5708 => x"82",
          5709 => x"58",
          5710 => x"0c",
          5711 => x"33",
          5712 => x"80",
          5713 => x"ff",
          5714 => x"ff",
          5715 => x"55",
          5716 => x"81",
          5717 => x"38",
          5718 => x"06",
          5719 => x"80",
          5720 => x"52",
          5721 => x"8a",
          5722 => x"80",
          5723 => x"ff",
          5724 => x"53",
          5725 => x"86",
          5726 => x"83",
          5727 => x"c5",
          5728 => x"f5",
          5729 => x"dc",
          5730 => x"8c",
          5731 => x"15",
          5732 => x"06",
          5733 => x"76",
          5734 => x"80",
          5735 => x"da",
          5736 => x"8c",
          5737 => x"ff",
          5738 => x"74",
          5739 => x"d4",
          5740 => x"dc",
          5741 => x"dc",
          5742 => x"c2",
          5743 => x"b9",
          5744 => x"dc",
          5745 => x"ff",
          5746 => x"56",
          5747 => x"83",
          5748 => x"14",
          5749 => x"71",
          5750 => x"5a",
          5751 => x"26",
          5752 => x"8a",
          5753 => x"74",
          5754 => x"ff",
          5755 => x"82",
          5756 => x"55",
          5757 => x"08",
          5758 => x"ec",
          5759 => x"dc",
          5760 => x"ff",
          5761 => x"83",
          5762 => x"74",
          5763 => x"26",
          5764 => x"57",
          5765 => x"26",
          5766 => x"57",
          5767 => x"56",
          5768 => x"82",
          5769 => x"15",
          5770 => x"0c",
          5771 => x"0c",
          5772 => x"a4",
          5773 => x"1d",
          5774 => x"54",
          5775 => x"2e",
          5776 => x"af",
          5777 => x"14",
          5778 => x"3f",
          5779 => x"08",
          5780 => x"06",
          5781 => x"72",
          5782 => x"79",
          5783 => x"80",
          5784 => x"d9",
          5785 => x"8c",
          5786 => x"15",
          5787 => x"2b",
          5788 => x"8d",
          5789 => x"2e",
          5790 => x"77",
          5791 => x"0c",
          5792 => x"76",
          5793 => x"38",
          5794 => x"70",
          5795 => x"81",
          5796 => x"53",
          5797 => x"89",
          5798 => x"56",
          5799 => x"08",
          5800 => x"38",
          5801 => x"15",
          5802 => x"8c",
          5803 => x"80",
          5804 => x"34",
          5805 => x"09",
          5806 => x"92",
          5807 => x"14",
          5808 => x"3f",
          5809 => x"08",
          5810 => x"06",
          5811 => x"2e",
          5812 => x"80",
          5813 => x"1b",
          5814 => x"db",
          5815 => x"8c",
          5816 => x"ea",
          5817 => x"dc",
          5818 => x"34",
          5819 => x"51",
          5820 => x"82",
          5821 => x"83",
          5822 => x"53",
          5823 => x"d5",
          5824 => x"06",
          5825 => x"b4",
          5826 => x"84",
          5827 => x"dc",
          5828 => x"85",
          5829 => x"09",
          5830 => x"38",
          5831 => x"51",
          5832 => x"82",
          5833 => x"86",
          5834 => x"f2",
          5835 => x"06",
          5836 => x"9c",
          5837 => x"d8",
          5838 => x"dc",
          5839 => x"0c",
          5840 => x"51",
          5841 => x"82",
          5842 => x"8c",
          5843 => x"74",
          5844 => x"9c",
          5845 => x"53",
          5846 => x"9c",
          5847 => x"15",
          5848 => x"94",
          5849 => x"56",
          5850 => x"dc",
          5851 => x"0d",
          5852 => x"0d",
          5853 => x"55",
          5854 => x"b9",
          5855 => x"53",
          5856 => x"b1",
          5857 => x"52",
          5858 => x"a9",
          5859 => x"22",
          5860 => x"57",
          5861 => x"2e",
          5862 => x"99",
          5863 => x"33",
          5864 => x"3f",
          5865 => x"08",
          5866 => x"71",
          5867 => x"74",
          5868 => x"83",
          5869 => x"78",
          5870 => x"52",
          5871 => x"dc",
          5872 => x"0d",
          5873 => x"0d",
          5874 => x"33",
          5875 => x"3d",
          5876 => x"56",
          5877 => x"8b",
          5878 => x"82",
          5879 => x"24",
          5880 => x"8c",
          5881 => x"29",
          5882 => x"05",
          5883 => x"55",
          5884 => x"84",
          5885 => x"34",
          5886 => x"80",
          5887 => x"80",
          5888 => x"75",
          5889 => x"75",
          5890 => x"38",
          5891 => x"3d",
          5892 => x"05",
          5893 => x"3f",
          5894 => x"08",
          5895 => x"8c",
          5896 => x"3d",
          5897 => x"3d",
          5898 => x"84",
          5899 => x"05",
          5900 => x"89",
          5901 => x"2e",
          5902 => x"77",
          5903 => x"54",
          5904 => x"05",
          5905 => x"84",
          5906 => x"f6",
          5907 => x"8c",
          5908 => x"82",
          5909 => x"84",
          5910 => x"5c",
          5911 => x"3d",
          5912 => x"ed",
          5913 => x"8c",
          5914 => x"82",
          5915 => x"92",
          5916 => x"d7",
          5917 => x"98",
          5918 => x"73",
          5919 => x"38",
          5920 => x"9c",
          5921 => x"80",
          5922 => x"38",
          5923 => x"95",
          5924 => x"2e",
          5925 => x"aa",
          5926 => x"ea",
          5927 => x"8c",
          5928 => x"9e",
          5929 => x"05",
          5930 => x"54",
          5931 => x"38",
          5932 => x"70",
          5933 => x"54",
          5934 => x"8e",
          5935 => x"83",
          5936 => x"88",
          5937 => x"83",
          5938 => x"83",
          5939 => x"06",
          5940 => x"80",
          5941 => x"38",
          5942 => x"51",
          5943 => x"82",
          5944 => x"56",
          5945 => x"0a",
          5946 => x"05",
          5947 => x"3f",
          5948 => x"0b",
          5949 => x"80",
          5950 => x"7a",
          5951 => x"3f",
          5952 => x"9c",
          5953 => x"d1",
          5954 => x"81",
          5955 => x"34",
          5956 => x"80",
          5957 => x"b0",
          5958 => x"54",
          5959 => x"52",
          5960 => x"05",
          5961 => x"3f",
          5962 => x"08",
          5963 => x"dc",
          5964 => x"38",
          5965 => x"82",
          5966 => x"b2",
          5967 => x"84",
          5968 => x"06",
          5969 => x"73",
          5970 => x"38",
          5971 => x"ad",
          5972 => x"2a",
          5973 => x"51",
          5974 => x"2e",
          5975 => x"81",
          5976 => x"80",
          5977 => x"87",
          5978 => x"39",
          5979 => x"51",
          5980 => x"82",
          5981 => x"7b",
          5982 => x"12",
          5983 => x"82",
          5984 => x"81",
          5985 => x"83",
          5986 => x"06",
          5987 => x"80",
          5988 => x"77",
          5989 => x"58",
          5990 => x"08",
          5991 => x"63",
          5992 => x"63",
          5993 => x"57",
          5994 => x"82",
          5995 => x"82",
          5996 => x"88",
          5997 => x"9c",
          5998 => x"d2",
          5999 => x"8c",
          6000 => x"8c",
          6001 => x"1b",
          6002 => x"0c",
          6003 => x"22",
          6004 => x"77",
          6005 => x"80",
          6006 => x"34",
          6007 => x"1a",
          6008 => x"94",
          6009 => x"85",
          6010 => x"06",
          6011 => x"80",
          6012 => x"38",
          6013 => x"08",
          6014 => x"84",
          6015 => x"dc",
          6016 => x"0c",
          6017 => x"70",
          6018 => x"52",
          6019 => x"39",
          6020 => x"51",
          6021 => x"82",
          6022 => x"57",
          6023 => x"08",
          6024 => x"38",
          6025 => x"8c",
          6026 => x"2e",
          6027 => x"83",
          6028 => x"75",
          6029 => x"74",
          6030 => x"07",
          6031 => x"54",
          6032 => x"8a",
          6033 => x"75",
          6034 => x"73",
          6035 => x"98",
          6036 => x"a9",
          6037 => x"ff",
          6038 => x"80",
          6039 => x"76",
          6040 => x"d6",
          6041 => x"8c",
          6042 => x"38",
          6043 => x"39",
          6044 => x"82",
          6045 => x"05",
          6046 => x"84",
          6047 => x"0c",
          6048 => x"82",
          6049 => x"97",
          6050 => x"f2",
          6051 => x"63",
          6052 => x"40",
          6053 => x"7e",
          6054 => x"fc",
          6055 => x"51",
          6056 => x"82",
          6057 => x"55",
          6058 => x"08",
          6059 => x"19",
          6060 => x"80",
          6061 => x"74",
          6062 => x"39",
          6063 => x"81",
          6064 => x"56",
          6065 => x"82",
          6066 => x"39",
          6067 => x"1a",
          6068 => x"82",
          6069 => x"0b",
          6070 => x"81",
          6071 => x"39",
          6072 => x"94",
          6073 => x"55",
          6074 => x"83",
          6075 => x"7b",
          6076 => x"89",
          6077 => x"08",
          6078 => x"06",
          6079 => x"81",
          6080 => x"8a",
          6081 => x"05",
          6082 => x"06",
          6083 => x"a8",
          6084 => x"38",
          6085 => x"55",
          6086 => x"19",
          6087 => x"51",
          6088 => x"82",
          6089 => x"55",
          6090 => x"ff",
          6091 => x"ff",
          6092 => x"38",
          6093 => x"0c",
          6094 => x"52",
          6095 => x"cb",
          6096 => x"dc",
          6097 => x"ff",
          6098 => x"8c",
          6099 => x"7c",
          6100 => x"57",
          6101 => x"80",
          6102 => x"1a",
          6103 => x"22",
          6104 => x"75",
          6105 => x"38",
          6106 => x"58",
          6107 => x"53",
          6108 => x"1b",
          6109 => x"88",
          6110 => x"dc",
          6111 => x"38",
          6112 => x"33",
          6113 => x"80",
          6114 => x"b0",
          6115 => x"31",
          6116 => x"27",
          6117 => x"80",
          6118 => x"52",
          6119 => x"77",
          6120 => x"7d",
          6121 => x"e0",
          6122 => x"2b",
          6123 => x"76",
          6124 => x"94",
          6125 => x"ff",
          6126 => x"71",
          6127 => x"7b",
          6128 => x"38",
          6129 => x"19",
          6130 => x"51",
          6131 => x"82",
          6132 => x"fe",
          6133 => x"53",
          6134 => x"83",
          6135 => x"b4",
          6136 => x"51",
          6137 => x"7b",
          6138 => x"08",
          6139 => x"76",
          6140 => x"08",
          6141 => x"0c",
          6142 => x"f3",
          6143 => x"75",
          6144 => x"0c",
          6145 => x"04",
          6146 => x"60",
          6147 => x"40",
          6148 => x"80",
          6149 => x"3d",
          6150 => x"77",
          6151 => x"3f",
          6152 => x"08",
          6153 => x"dc",
          6154 => x"91",
          6155 => x"74",
          6156 => x"38",
          6157 => x"b8",
          6158 => x"33",
          6159 => x"70",
          6160 => x"56",
          6161 => x"74",
          6162 => x"a4",
          6163 => x"82",
          6164 => x"34",
          6165 => x"98",
          6166 => x"91",
          6167 => x"56",
          6168 => x"94",
          6169 => x"11",
          6170 => x"76",
          6171 => x"75",
          6172 => x"80",
          6173 => x"38",
          6174 => x"70",
          6175 => x"56",
          6176 => x"fd",
          6177 => x"11",
          6178 => x"77",
          6179 => x"5c",
          6180 => x"38",
          6181 => x"88",
          6182 => x"74",
          6183 => x"52",
          6184 => x"18",
          6185 => x"51",
          6186 => x"82",
          6187 => x"55",
          6188 => x"08",
          6189 => x"ab",
          6190 => x"2e",
          6191 => x"74",
          6192 => x"95",
          6193 => x"19",
          6194 => x"08",
          6195 => x"88",
          6196 => x"55",
          6197 => x"9c",
          6198 => x"09",
          6199 => x"38",
          6200 => x"c1",
          6201 => x"dc",
          6202 => x"38",
          6203 => x"52",
          6204 => x"97",
          6205 => x"dc",
          6206 => x"fe",
          6207 => x"8c",
          6208 => x"7c",
          6209 => x"57",
          6210 => x"80",
          6211 => x"1b",
          6212 => x"22",
          6213 => x"75",
          6214 => x"38",
          6215 => x"59",
          6216 => x"53",
          6217 => x"1a",
          6218 => x"be",
          6219 => x"dc",
          6220 => x"38",
          6221 => x"08",
          6222 => x"56",
          6223 => x"9b",
          6224 => x"53",
          6225 => x"77",
          6226 => x"7d",
          6227 => x"16",
          6228 => x"3f",
          6229 => x"0b",
          6230 => x"78",
          6231 => x"80",
          6232 => x"18",
          6233 => x"08",
          6234 => x"7e",
          6235 => x"3f",
          6236 => x"08",
          6237 => x"7e",
          6238 => x"0c",
          6239 => x"19",
          6240 => x"08",
          6241 => x"84",
          6242 => x"57",
          6243 => x"27",
          6244 => x"56",
          6245 => x"52",
          6246 => x"f9",
          6247 => x"dc",
          6248 => x"38",
          6249 => x"52",
          6250 => x"83",
          6251 => x"b4",
          6252 => x"d4",
          6253 => x"81",
          6254 => x"34",
          6255 => x"7e",
          6256 => x"0c",
          6257 => x"1a",
          6258 => x"94",
          6259 => x"1b",
          6260 => x"5e",
          6261 => x"27",
          6262 => x"55",
          6263 => x"0c",
          6264 => x"90",
          6265 => x"c0",
          6266 => x"90",
          6267 => x"56",
          6268 => x"dc",
          6269 => x"0d",
          6270 => x"0d",
          6271 => x"fc",
          6272 => x"52",
          6273 => x"3f",
          6274 => x"08",
          6275 => x"dc",
          6276 => x"38",
          6277 => x"70",
          6278 => x"81",
          6279 => x"55",
          6280 => x"80",
          6281 => x"16",
          6282 => x"51",
          6283 => x"82",
          6284 => x"57",
          6285 => x"08",
          6286 => x"a4",
          6287 => x"11",
          6288 => x"55",
          6289 => x"16",
          6290 => x"08",
          6291 => x"75",
          6292 => x"e8",
          6293 => x"08",
          6294 => x"51",
          6295 => x"82",
          6296 => x"52",
          6297 => x"c9",
          6298 => x"52",
          6299 => x"c9",
          6300 => x"54",
          6301 => x"15",
          6302 => x"cc",
          6303 => x"8c",
          6304 => x"17",
          6305 => x"06",
          6306 => x"90",
          6307 => x"82",
          6308 => x"8a",
          6309 => x"fc",
          6310 => x"70",
          6311 => x"d9",
          6312 => x"dc",
          6313 => x"8c",
          6314 => x"38",
          6315 => x"05",
          6316 => x"f1",
          6317 => x"8c",
          6318 => x"82",
          6319 => x"87",
          6320 => x"dc",
          6321 => x"72",
          6322 => x"0c",
          6323 => x"04",
          6324 => x"84",
          6325 => x"e4",
          6326 => x"80",
          6327 => x"dc",
          6328 => x"38",
          6329 => x"08",
          6330 => x"34",
          6331 => x"82",
          6332 => x"83",
          6333 => x"ef",
          6334 => x"53",
          6335 => x"05",
          6336 => x"51",
          6337 => x"82",
          6338 => x"55",
          6339 => x"08",
          6340 => x"76",
          6341 => x"93",
          6342 => x"51",
          6343 => x"82",
          6344 => x"55",
          6345 => x"08",
          6346 => x"80",
          6347 => x"70",
          6348 => x"56",
          6349 => x"89",
          6350 => x"94",
          6351 => x"b2",
          6352 => x"05",
          6353 => x"2a",
          6354 => x"51",
          6355 => x"80",
          6356 => x"76",
          6357 => x"52",
          6358 => x"3f",
          6359 => x"08",
          6360 => x"8e",
          6361 => x"dc",
          6362 => x"09",
          6363 => x"38",
          6364 => x"82",
          6365 => x"93",
          6366 => x"e4",
          6367 => x"6f",
          6368 => x"7a",
          6369 => x"9e",
          6370 => x"05",
          6371 => x"51",
          6372 => x"82",
          6373 => x"57",
          6374 => x"08",
          6375 => x"7b",
          6376 => x"94",
          6377 => x"55",
          6378 => x"73",
          6379 => x"ed",
          6380 => x"93",
          6381 => x"55",
          6382 => x"82",
          6383 => x"57",
          6384 => x"08",
          6385 => x"68",
          6386 => x"c9",
          6387 => x"8c",
          6388 => x"82",
          6389 => x"82",
          6390 => x"52",
          6391 => x"a3",
          6392 => x"dc",
          6393 => x"52",
          6394 => x"b8",
          6395 => x"dc",
          6396 => x"8c",
          6397 => x"a2",
          6398 => x"74",
          6399 => x"3f",
          6400 => x"08",
          6401 => x"dc",
          6402 => x"69",
          6403 => x"d9",
          6404 => x"82",
          6405 => x"2e",
          6406 => x"52",
          6407 => x"cf",
          6408 => x"dc",
          6409 => x"8c",
          6410 => x"2e",
          6411 => x"84",
          6412 => x"06",
          6413 => x"57",
          6414 => x"76",
          6415 => x"9e",
          6416 => x"05",
          6417 => x"dc",
          6418 => x"90",
          6419 => x"81",
          6420 => x"56",
          6421 => x"80",
          6422 => x"02",
          6423 => x"81",
          6424 => x"70",
          6425 => x"56",
          6426 => x"81",
          6427 => x"78",
          6428 => x"38",
          6429 => x"99",
          6430 => x"81",
          6431 => x"18",
          6432 => x"18",
          6433 => x"58",
          6434 => x"33",
          6435 => x"ee",
          6436 => x"6f",
          6437 => x"af",
          6438 => x"8d",
          6439 => x"2e",
          6440 => x"8a",
          6441 => x"6f",
          6442 => x"af",
          6443 => x"0b",
          6444 => x"33",
          6445 => x"81",
          6446 => x"70",
          6447 => x"52",
          6448 => x"56",
          6449 => x"8d",
          6450 => x"70",
          6451 => x"51",
          6452 => x"f5",
          6453 => x"54",
          6454 => x"a7",
          6455 => x"74",
          6456 => x"38",
          6457 => x"73",
          6458 => x"81",
          6459 => x"81",
          6460 => x"39",
          6461 => x"81",
          6462 => x"74",
          6463 => x"81",
          6464 => x"91",
          6465 => x"6e",
          6466 => x"59",
          6467 => x"7a",
          6468 => x"5c",
          6469 => x"26",
          6470 => x"7a",
          6471 => x"8c",
          6472 => x"3d",
          6473 => x"3d",
          6474 => x"8d",
          6475 => x"54",
          6476 => x"55",
          6477 => x"82",
          6478 => x"53",
          6479 => x"08",
          6480 => x"91",
          6481 => x"72",
          6482 => x"8c",
          6483 => x"73",
          6484 => x"38",
          6485 => x"70",
          6486 => x"81",
          6487 => x"57",
          6488 => x"73",
          6489 => x"08",
          6490 => x"94",
          6491 => x"75",
          6492 => x"97",
          6493 => x"11",
          6494 => x"2b",
          6495 => x"73",
          6496 => x"38",
          6497 => x"16",
          6498 => x"d0",
          6499 => x"dc",
          6500 => x"78",
          6501 => x"55",
          6502 => x"c0",
          6503 => x"dc",
          6504 => x"96",
          6505 => x"70",
          6506 => x"94",
          6507 => x"71",
          6508 => x"08",
          6509 => x"53",
          6510 => x"15",
          6511 => x"a6",
          6512 => x"74",
          6513 => x"3f",
          6514 => x"08",
          6515 => x"dc",
          6516 => x"81",
          6517 => x"8c",
          6518 => x"2e",
          6519 => x"82",
          6520 => x"88",
          6521 => x"98",
          6522 => x"80",
          6523 => x"38",
          6524 => x"80",
          6525 => x"77",
          6526 => x"08",
          6527 => x"0c",
          6528 => x"70",
          6529 => x"81",
          6530 => x"5a",
          6531 => x"2e",
          6532 => x"52",
          6533 => x"f9",
          6534 => x"dc",
          6535 => x"8c",
          6536 => x"38",
          6537 => x"08",
          6538 => x"73",
          6539 => x"c7",
          6540 => x"8c",
          6541 => x"73",
          6542 => x"38",
          6543 => x"af",
          6544 => x"73",
          6545 => x"27",
          6546 => x"98",
          6547 => x"a0",
          6548 => x"08",
          6549 => x"0c",
          6550 => x"06",
          6551 => x"2e",
          6552 => x"52",
          6553 => x"a3",
          6554 => x"dc",
          6555 => x"82",
          6556 => x"34",
          6557 => x"c4",
          6558 => x"91",
          6559 => x"53",
          6560 => x"89",
          6561 => x"dc",
          6562 => x"94",
          6563 => x"8c",
          6564 => x"27",
          6565 => x"8c",
          6566 => x"15",
          6567 => x"07",
          6568 => x"16",
          6569 => x"ff",
          6570 => x"80",
          6571 => x"77",
          6572 => x"2e",
          6573 => x"9c",
          6574 => x"53",
          6575 => x"dc",
          6576 => x"0d",
          6577 => x"0d",
          6578 => x"54",
          6579 => x"81",
          6580 => x"53",
          6581 => x"05",
          6582 => x"84",
          6583 => x"e7",
          6584 => x"dc",
          6585 => x"8c",
          6586 => x"ea",
          6587 => x"0c",
          6588 => x"51",
          6589 => x"82",
          6590 => x"55",
          6591 => x"08",
          6592 => x"ab",
          6593 => x"98",
          6594 => x"80",
          6595 => x"38",
          6596 => x"70",
          6597 => x"81",
          6598 => x"57",
          6599 => x"ad",
          6600 => x"08",
          6601 => x"d3",
          6602 => x"8c",
          6603 => x"17",
          6604 => x"86",
          6605 => x"17",
          6606 => x"75",
          6607 => x"3f",
          6608 => x"08",
          6609 => x"2e",
          6610 => x"85",
          6611 => x"86",
          6612 => x"2e",
          6613 => x"76",
          6614 => x"73",
          6615 => x"0c",
          6616 => x"04",
          6617 => x"76",
          6618 => x"05",
          6619 => x"53",
          6620 => x"82",
          6621 => x"87",
          6622 => x"dc",
          6623 => x"86",
          6624 => x"fb",
          6625 => x"79",
          6626 => x"05",
          6627 => x"56",
          6628 => x"3f",
          6629 => x"08",
          6630 => x"dc",
          6631 => x"38",
          6632 => x"82",
          6633 => x"52",
          6634 => x"f8",
          6635 => x"dc",
          6636 => x"ca",
          6637 => x"dc",
          6638 => x"51",
          6639 => x"82",
          6640 => x"53",
          6641 => x"08",
          6642 => x"81",
          6643 => x"80",
          6644 => x"82",
          6645 => x"a6",
          6646 => x"73",
          6647 => x"3f",
          6648 => x"51",
          6649 => x"82",
          6650 => x"84",
          6651 => x"70",
          6652 => x"2c",
          6653 => x"dc",
          6654 => x"51",
          6655 => x"82",
          6656 => x"87",
          6657 => x"ee",
          6658 => x"57",
          6659 => x"3d",
          6660 => x"3d",
          6661 => x"af",
          6662 => x"dc",
          6663 => x"8c",
          6664 => x"38",
          6665 => x"51",
          6666 => x"82",
          6667 => x"55",
          6668 => x"08",
          6669 => x"80",
          6670 => x"70",
          6671 => x"58",
          6672 => x"85",
          6673 => x"8d",
          6674 => x"2e",
          6675 => x"52",
          6676 => x"be",
          6677 => x"8c",
          6678 => x"3d",
          6679 => x"3d",
          6680 => x"55",
          6681 => x"92",
          6682 => x"52",
          6683 => x"de",
          6684 => x"8c",
          6685 => x"82",
          6686 => x"82",
          6687 => x"74",
          6688 => x"98",
          6689 => x"11",
          6690 => x"59",
          6691 => x"75",
          6692 => x"38",
          6693 => x"81",
          6694 => x"5b",
          6695 => x"82",
          6696 => x"39",
          6697 => x"08",
          6698 => x"59",
          6699 => x"09",
          6700 => x"38",
          6701 => x"57",
          6702 => x"3d",
          6703 => x"c1",
          6704 => x"8c",
          6705 => x"2e",
          6706 => x"8c",
          6707 => x"2e",
          6708 => x"8c",
          6709 => x"70",
          6710 => x"08",
          6711 => x"7a",
          6712 => x"7f",
          6713 => x"54",
          6714 => x"77",
          6715 => x"80",
          6716 => x"15",
          6717 => x"dc",
          6718 => x"75",
          6719 => x"52",
          6720 => x"52",
          6721 => x"8d",
          6722 => x"dc",
          6723 => x"8c",
          6724 => x"d6",
          6725 => x"33",
          6726 => x"1a",
          6727 => x"54",
          6728 => x"09",
          6729 => x"38",
          6730 => x"ff",
          6731 => x"82",
          6732 => x"83",
          6733 => x"70",
          6734 => x"25",
          6735 => x"59",
          6736 => x"9b",
          6737 => x"51",
          6738 => x"3f",
          6739 => x"08",
          6740 => x"70",
          6741 => x"25",
          6742 => x"59",
          6743 => x"75",
          6744 => x"7a",
          6745 => x"ff",
          6746 => x"7c",
          6747 => x"90",
          6748 => x"11",
          6749 => x"56",
          6750 => x"15",
          6751 => x"8c",
          6752 => x"3d",
          6753 => x"3d",
          6754 => x"3d",
          6755 => x"70",
          6756 => x"dd",
          6757 => x"dc",
          6758 => x"8c",
          6759 => x"a8",
          6760 => x"33",
          6761 => x"a0",
          6762 => x"33",
          6763 => x"70",
          6764 => x"55",
          6765 => x"73",
          6766 => x"8e",
          6767 => x"08",
          6768 => x"18",
          6769 => x"80",
          6770 => x"38",
          6771 => x"08",
          6772 => x"08",
          6773 => x"c4",
          6774 => x"8c",
          6775 => x"88",
          6776 => x"80",
          6777 => x"17",
          6778 => x"51",
          6779 => x"3f",
          6780 => x"08",
          6781 => x"81",
          6782 => x"81",
          6783 => x"dc",
          6784 => x"09",
          6785 => x"38",
          6786 => x"39",
          6787 => x"77",
          6788 => x"dc",
          6789 => x"08",
          6790 => x"98",
          6791 => x"82",
          6792 => x"52",
          6793 => x"bd",
          6794 => x"dc",
          6795 => x"17",
          6796 => x"0c",
          6797 => x"80",
          6798 => x"73",
          6799 => x"75",
          6800 => x"38",
          6801 => x"34",
          6802 => x"82",
          6803 => x"89",
          6804 => x"e2",
          6805 => x"53",
          6806 => x"a4",
          6807 => x"3d",
          6808 => x"3f",
          6809 => x"08",
          6810 => x"dc",
          6811 => x"38",
          6812 => x"3d",
          6813 => x"3d",
          6814 => x"d1",
          6815 => x"8c",
          6816 => x"82",
          6817 => x"81",
          6818 => x"80",
          6819 => x"70",
          6820 => x"81",
          6821 => x"56",
          6822 => x"81",
          6823 => x"98",
          6824 => x"74",
          6825 => x"38",
          6826 => x"05",
          6827 => x"06",
          6828 => x"55",
          6829 => x"38",
          6830 => x"51",
          6831 => x"82",
          6832 => x"74",
          6833 => x"81",
          6834 => x"56",
          6835 => x"80",
          6836 => x"54",
          6837 => x"08",
          6838 => x"2e",
          6839 => x"73",
          6840 => x"dc",
          6841 => x"52",
          6842 => x"52",
          6843 => x"3f",
          6844 => x"08",
          6845 => x"dc",
          6846 => x"38",
          6847 => x"08",
          6848 => x"cc",
          6849 => x"8c",
          6850 => x"82",
          6851 => x"86",
          6852 => x"80",
          6853 => x"8c",
          6854 => x"2e",
          6855 => x"8c",
          6856 => x"c0",
          6857 => x"ce",
          6858 => x"8c",
          6859 => x"8c",
          6860 => x"70",
          6861 => x"08",
          6862 => x"51",
          6863 => x"80",
          6864 => x"73",
          6865 => x"38",
          6866 => x"52",
          6867 => x"95",
          6868 => x"dc",
          6869 => x"8c",
          6870 => x"ff",
          6871 => x"82",
          6872 => x"55",
          6873 => x"dc",
          6874 => x"0d",
          6875 => x"0d",
          6876 => x"3d",
          6877 => x"9a",
          6878 => x"cb",
          6879 => x"dc",
          6880 => x"8c",
          6881 => x"b0",
          6882 => x"69",
          6883 => x"70",
          6884 => x"97",
          6885 => x"dc",
          6886 => x"8c",
          6887 => x"38",
          6888 => x"94",
          6889 => x"dc",
          6890 => x"09",
          6891 => x"88",
          6892 => x"df",
          6893 => x"85",
          6894 => x"51",
          6895 => x"74",
          6896 => x"78",
          6897 => x"8a",
          6898 => x"57",
          6899 => x"82",
          6900 => x"75",
          6901 => x"8c",
          6902 => x"38",
          6903 => x"8c",
          6904 => x"2e",
          6905 => x"83",
          6906 => x"82",
          6907 => x"ff",
          6908 => x"06",
          6909 => x"54",
          6910 => x"73",
          6911 => x"82",
          6912 => x"52",
          6913 => x"a4",
          6914 => x"dc",
          6915 => x"8c",
          6916 => x"9a",
          6917 => x"a0",
          6918 => x"51",
          6919 => x"3f",
          6920 => x"0b",
          6921 => x"78",
          6922 => x"bf",
          6923 => x"88",
          6924 => x"80",
          6925 => x"ff",
          6926 => x"75",
          6927 => x"11",
          6928 => x"f8",
          6929 => x"78",
          6930 => x"80",
          6931 => x"ff",
          6932 => x"78",
          6933 => x"80",
          6934 => x"7f",
          6935 => x"d4",
          6936 => x"c9",
          6937 => x"54",
          6938 => x"15",
          6939 => x"cb",
          6940 => x"8c",
          6941 => x"82",
          6942 => x"b2",
          6943 => x"b2",
          6944 => x"96",
          6945 => x"b5",
          6946 => x"53",
          6947 => x"51",
          6948 => x"64",
          6949 => x"8b",
          6950 => x"54",
          6951 => x"15",
          6952 => x"ff",
          6953 => x"82",
          6954 => x"54",
          6955 => x"53",
          6956 => x"51",
          6957 => x"3f",
          6958 => x"dc",
          6959 => x"0d",
          6960 => x"0d",
          6961 => x"05",
          6962 => x"3f",
          6963 => x"3d",
          6964 => x"52",
          6965 => x"d5",
          6966 => x"8c",
          6967 => x"82",
          6968 => x"82",
          6969 => x"4d",
          6970 => x"52",
          6971 => x"52",
          6972 => x"3f",
          6973 => x"08",
          6974 => x"dc",
          6975 => x"38",
          6976 => x"05",
          6977 => x"06",
          6978 => x"73",
          6979 => x"a0",
          6980 => x"08",
          6981 => x"ff",
          6982 => x"ff",
          6983 => x"ac",
          6984 => x"92",
          6985 => x"54",
          6986 => x"3f",
          6987 => x"52",
          6988 => x"f7",
          6989 => x"dc",
          6990 => x"8c",
          6991 => x"38",
          6992 => x"09",
          6993 => x"38",
          6994 => x"08",
          6995 => x"88",
          6996 => x"39",
          6997 => x"08",
          6998 => x"81",
          6999 => x"38",
          7000 => x"b1",
          7001 => x"dc",
          7002 => x"8c",
          7003 => x"c8",
          7004 => x"93",
          7005 => x"ff",
          7006 => x"8d",
          7007 => x"b4",
          7008 => x"af",
          7009 => x"17",
          7010 => x"33",
          7011 => x"70",
          7012 => x"55",
          7013 => x"38",
          7014 => x"54",
          7015 => x"34",
          7016 => x"0b",
          7017 => x"8b",
          7018 => x"84",
          7019 => x"06",
          7020 => x"73",
          7021 => x"e5",
          7022 => x"2e",
          7023 => x"75",
          7024 => x"c6",
          7025 => x"8c",
          7026 => x"78",
          7027 => x"bb",
          7028 => x"82",
          7029 => x"80",
          7030 => x"38",
          7031 => x"08",
          7032 => x"ff",
          7033 => x"82",
          7034 => x"79",
          7035 => x"58",
          7036 => x"8c",
          7037 => x"c0",
          7038 => x"33",
          7039 => x"2e",
          7040 => x"99",
          7041 => x"75",
          7042 => x"c6",
          7043 => x"54",
          7044 => x"15",
          7045 => x"82",
          7046 => x"9c",
          7047 => x"c8",
          7048 => x"8c",
          7049 => x"82",
          7050 => x"8c",
          7051 => x"ff",
          7052 => x"82",
          7053 => x"55",
          7054 => x"dc",
          7055 => x"0d",
          7056 => x"0d",
          7057 => x"05",
          7058 => x"05",
          7059 => x"33",
          7060 => x"53",
          7061 => x"05",
          7062 => x"51",
          7063 => x"82",
          7064 => x"55",
          7065 => x"08",
          7066 => x"78",
          7067 => x"95",
          7068 => x"51",
          7069 => x"82",
          7070 => x"55",
          7071 => x"08",
          7072 => x"80",
          7073 => x"81",
          7074 => x"86",
          7075 => x"38",
          7076 => x"61",
          7077 => x"12",
          7078 => x"7a",
          7079 => x"51",
          7080 => x"74",
          7081 => x"78",
          7082 => x"83",
          7083 => x"51",
          7084 => x"3f",
          7085 => x"08",
          7086 => x"8c",
          7087 => x"3d",
          7088 => x"3d",
          7089 => x"82",
          7090 => x"d0",
          7091 => x"3d",
          7092 => x"3f",
          7093 => x"08",
          7094 => x"dc",
          7095 => x"38",
          7096 => x"52",
          7097 => x"05",
          7098 => x"3f",
          7099 => x"08",
          7100 => x"dc",
          7101 => x"02",
          7102 => x"33",
          7103 => x"54",
          7104 => x"a6",
          7105 => x"22",
          7106 => x"71",
          7107 => x"53",
          7108 => x"51",
          7109 => x"3f",
          7110 => x"0b",
          7111 => x"76",
          7112 => x"b8",
          7113 => x"dc",
          7114 => x"82",
          7115 => x"93",
          7116 => x"ea",
          7117 => x"6b",
          7118 => x"53",
          7119 => x"05",
          7120 => x"51",
          7121 => x"82",
          7122 => x"82",
          7123 => x"30",
          7124 => x"dc",
          7125 => x"25",
          7126 => x"79",
          7127 => x"85",
          7128 => x"75",
          7129 => x"73",
          7130 => x"f9",
          7131 => x"80",
          7132 => x"8d",
          7133 => x"54",
          7134 => x"3f",
          7135 => x"08",
          7136 => x"dc",
          7137 => x"38",
          7138 => x"51",
          7139 => x"82",
          7140 => x"57",
          7141 => x"08",
          7142 => x"8c",
          7143 => x"8c",
          7144 => x"5b",
          7145 => x"18",
          7146 => x"18",
          7147 => x"74",
          7148 => x"81",
          7149 => x"78",
          7150 => x"8b",
          7151 => x"54",
          7152 => x"75",
          7153 => x"38",
          7154 => x"1b",
          7155 => x"55",
          7156 => x"2e",
          7157 => x"39",
          7158 => x"09",
          7159 => x"38",
          7160 => x"80",
          7161 => x"70",
          7162 => x"25",
          7163 => x"80",
          7164 => x"38",
          7165 => x"bc",
          7166 => x"11",
          7167 => x"ff",
          7168 => x"82",
          7169 => x"57",
          7170 => x"08",
          7171 => x"70",
          7172 => x"80",
          7173 => x"83",
          7174 => x"80",
          7175 => x"84",
          7176 => x"a7",
          7177 => x"b4",
          7178 => x"ad",
          7179 => x"8c",
          7180 => x"0c",
          7181 => x"dc",
          7182 => x"0d",
          7183 => x"0d",
          7184 => x"3d",
          7185 => x"52",
          7186 => x"ce",
          7187 => x"8c",
          7188 => x"8c",
          7189 => x"54",
          7190 => x"08",
          7191 => x"8b",
          7192 => x"8b",
          7193 => x"59",
          7194 => x"3f",
          7195 => x"33",
          7196 => x"06",
          7197 => x"57",
          7198 => x"81",
          7199 => x"58",
          7200 => x"06",
          7201 => x"4e",
          7202 => x"ff",
          7203 => x"82",
          7204 => x"80",
          7205 => x"6c",
          7206 => x"53",
          7207 => x"ae",
          7208 => x"8c",
          7209 => x"2e",
          7210 => x"88",
          7211 => x"6d",
          7212 => x"55",
          7213 => x"8c",
          7214 => x"ff",
          7215 => x"83",
          7216 => x"51",
          7217 => x"26",
          7218 => x"15",
          7219 => x"ff",
          7220 => x"80",
          7221 => x"87",
          7222 => x"ec",
          7223 => x"74",
          7224 => x"38",
          7225 => x"fb",
          7226 => x"ae",
          7227 => x"8c",
          7228 => x"38",
          7229 => x"27",
          7230 => x"89",
          7231 => x"8b",
          7232 => x"27",
          7233 => x"55",
          7234 => x"81",
          7235 => x"8f",
          7236 => x"2a",
          7237 => x"70",
          7238 => x"34",
          7239 => x"74",
          7240 => x"05",
          7241 => x"17",
          7242 => x"70",
          7243 => x"52",
          7244 => x"73",
          7245 => x"c8",
          7246 => x"33",
          7247 => x"73",
          7248 => x"81",
          7249 => x"80",
          7250 => x"02",
          7251 => x"76",
          7252 => x"51",
          7253 => x"2e",
          7254 => x"87",
          7255 => x"57",
          7256 => x"79",
          7257 => x"80",
          7258 => x"70",
          7259 => x"ba",
          7260 => x"8c",
          7261 => x"82",
          7262 => x"80",
          7263 => x"52",
          7264 => x"bf",
          7265 => x"8c",
          7266 => x"82",
          7267 => x"8d",
          7268 => x"c4",
          7269 => x"e5",
          7270 => x"c6",
          7271 => x"dc",
          7272 => x"09",
          7273 => x"cc",
          7274 => x"76",
          7275 => x"c4",
          7276 => x"74",
          7277 => x"b0",
          7278 => x"dc",
          7279 => x"8c",
          7280 => x"38",
          7281 => x"8c",
          7282 => x"67",
          7283 => x"db",
          7284 => x"88",
          7285 => x"34",
          7286 => x"52",
          7287 => x"ab",
          7288 => x"54",
          7289 => x"15",
          7290 => x"ff",
          7291 => x"82",
          7292 => x"54",
          7293 => x"82",
          7294 => x"9c",
          7295 => x"f2",
          7296 => x"62",
          7297 => x"80",
          7298 => x"93",
          7299 => x"55",
          7300 => x"5e",
          7301 => x"3f",
          7302 => x"08",
          7303 => x"dc",
          7304 => x"38",
          7305 => x"58",
          7306 => x"38",
          7307 => x"97",
          7308 => x"08",
          7309 => x"38",
          7310 => x"70",
          7311 => x"81",
          7312 => x"55",
          7313 => x"87",
          7314 => x"39",
          7315 => x"90",
          7316 => x"82",
          7317 => x"8a",
          7318 => x"89",
          7319 => x"7f",
          7320 => x"56",
          7321 => x"3f",
          7322 => x"06",
          7323 => x"72",
          7324 => x"82",
          7325 => x"05",
          7326 => x"7c",
          7327 => x"55",
          7328 => x"27",
          7329 => x"16",
          7330 => x"83",
          7331 => x"76",
          7332 => x"80",
          7333 => x"79",
          7334 => x"99",
          7335 => x"7f",
          7336 => x"14",
          7337 => x"83",
          7338 => x"82",
          7339 => x"81",
          7340 => x"38",
          7341 => x"08",
          7342 => x"95",
          7343 => x"dc",
          7344 => x"81",
          7345 => x"7b",
          7346 => x"06",
          7347 => x"39",
          7348 => x"56",
          7349 => x"09",
          7350 => x"b9",
          7351 => x"80",
          7352 => x"80",
          7353 => x"78",
          7354 => x"7a",
          7355 => x"38",
          7356 => x"73",
          7357 => x"81",
          7358 => x"ff",
          7359 => x"74",
          7360 => x"ff",
          7361 => x"82",
          7362 => x"58",
          7363 => x"08",
          7364 => x"74",
          7365 => x"16",
          7366 => x"73",
          7367 => x"39",
          7368 => x"7e",
          7369 => x"0c",
          7370 => x"2e",
          7371 => x"88",
          7372 => x"8c",
          7373 => x"1a",
          7374 => x"07",
          7375 => x"1b",
          7376 => x"08",
          7377 => x"16",
          7378 => x"75",
          7379 => x"38",
          7380 => x"90",
          7381 => x"15",
          7382 => x"54",
          7383 => x"34",
          7384 => x"82",
          7385 => x"90",
          7386 => x"e9",
          7387 => x"6d",
          7388 => x"80",
          7389 => x"9d",
          7390 => x"5c",
          7391 => x"3f",
          7392 => x"0b",
          7393 => x"08",
          7394 => x"38",
          7395 => x"08",
          7396 => x"8d",
          7397 => x"08",
          7398 => x"80",
          7399 => x"80",
          7400 => x"8c",
          7401 => x"ff",
          7402 => x"52",
          7403 => x"a0",
          7404 => x"8c",
          7405 => x"ff",
          7406 => x"06",
          7407 => x"56",
          7408 => x"38",
          7409 => x"70",
          7410 => x"55",
          7411 => x"8b",
          7412 => x"3d",
          7413 => x"83",
          7414 => x"ff",
          7415 => x"82",
          7416 => x"99",
          7417 => x"74",
          7418 => x"38",
          7419 => x"80",
          7420 => x"ff",
          7421 => x"55",
          7422 => x"83",
          7423 => x"78",
          7424 => x"38",
          7425 => x"26",
          7426 => x"81",
          7427 => x"8b",
          7428 => x"79",
          7429 => x"80",
          7430 => x"93",
          7431 => x"39",
          7432 => x"6e",
          7433 => x"89",
          7434 => x"48",
          7435 => x"83",
          7436 => x"61",
          7437 => x"25",
          7438 => x"55",
          7439 => x"8a",
          7440 => x"3d",
          7441 => x"81",
          7442 => x"ff",
          7443 => x"81",
          7444 => x"dc",
          7445 => x"38",
          7446 => x"70",
          7447 => x"8c",
          7448 => x"56",
          7449 => x"38",
          7450 => x"55",
          7451 => x"75",
          7452 => x"38",
          7453 => x"70",
          7454 => x"ff",
          7455 => x"83",
          7456 => x"78",
          7457 => x"89",
          7458 => x"81",
          7459 => x"06",
          7460 => x"80",
          7461 => x"77",
          7462 => x"74",
          7463 => x"8d",
          7464 => x"06",
          7465 => x"2e",
          7466 => x"77",
          7467 => x"93",
          7468 => x"74",
          7469 => x"cb",
          7470 => x"7d",
          7471 => x"81",
          7472 => x"38",
          7473 => x"66",
          7474 => x"81",
          7475 => x"90",
          7476 => x"74",
          7477 => x"38",
          7478 => x"98",
          7479 => x"90",
          7480 => x"82",
          7481 => x"57",
          7482 => x"80",
          7483 => x"76",
          7484 => x"38",
          7485 => x"51",
          7486 => x"3f",
          7487 => x"08",
          7488 => x"87",
          7489 => x"2a",
          7490 => x"5c",
          7491 => x"8c",
          7492 => x"80",
          7493 => x"44",
          7494 => x"0a",
          7495 => x"ec",
          7496 => x"39",
          7497 => x"66",
          7498 => x"81",
          7499 => x"80",
          7500 => x"74",
          7501 => x"38",
          7502 => x"98",
          7503 => x"80",
          7504 => x"82",
          7505 => x"57",
          7506 => x"80",
          7507 => x"76",
          7508 => x"38",
          7509 => x"51",
          7510 => x"3f",
          7511 => x"08",
          7512 => x"57",
          7513 => x"08",
          7514 => x"96",
          7515 => x"82",
          7516 => x"10",
          7517 => x"08",
          7518 => x"72",
          7519 => x"59",
          7520 => x"ff",
          7521 => x"5d",
          7522 => x"44",
          7523 => x"11",
          7524 => x"70",
          7525 => x"71",
          7526 => x"06",
          7527 => x"52",
          7528 => x"40",
          7529 => x"09",
          7530 => x"38",
          7531 => x"18",
          7532 => x"39",
          7533 => x"79",
          7534 => x"70",
          7535 => x"58",
          7536 => x"76",
          7537 => x"38",
          7538 => x"7d",
          7539 => x"70",
          7540 => x"55",
          7541 => x"3f",
          7542 => x"08",
          7543 => x"2e",
          7544 => x"9b",
          7545 => x"dc",
          7546 => x"f5",
          7547 => x"38",
          7548 => x"38",
          7549 => x"59",
          7550 => x"38",
          7551 => x"7d",
          7552 => x"81",
          7553 => x"38",
          7554 => x"0b",
          7555 => x"08",
          7556 => x"78",
          7557 => x"1a",
          7558 => x"c0",
          7559 => x"74",
          7560 => x"39",
          7561 => x"55",
          7562 => x"8f",
          7563 => x"fd",
          7564 => x"8c",
          7565 => x"f5",
          7566 => x"78",
          7567 => x"79",
          7568 => x"80",
          7569 => x"f1",
          7570 => x"39",
          7571 => x"81",
          7572 => x"06",
          7573 => x"55",
          7574 => x"27",
          7575 => x"81",
          7576 => x"56",
          7577 => x"38",
          7578 => x"80",
          7579 => x"ff",
          7580 => x"8b",
          7581 => x"a8",
          7582 => x"ff",
          7583 => x"84",
          7584 => x"1b",
          7585 => x"b3",
          7586 => x"1c",
          7587 => x"ff",
          7588 => x"8e",
          7589 => x"a1",
          7590 => x"0b",
          7591 => x"7d",
          7592 => x"30",
          7593 => x"84",
          7594 => x"51",
          7595 => x"51",
          7596 => x"3f",
          7597 => x"83",
          7598 => x"90",
          7599 => x"ff",
          7600 => x"93",
          7601 => x"a0",
          7602 => x"39",
          7603 => x"1b",
          7604 => x"85",
          7605 => x"95",
          7606 => x"52",
          7607 => x"ff",
          7608 => x"81",
          7609 => x"1b",
          7610 => x"cf",
          7611 => x"9c",
          7612 => x"a0",
          7613 => x"83",
          7614 => x"06",
          7615 => x"82",
          7616 => x"52",
          7617 => x"51",
          7618 => x"3f",
          7619 => x"1b",
          7620 => x"c5",
          7621 => x"ac",
          7622 => x"a0",
          7623 => x"52",
          7624 => x"ff",
          7625 => x"86",
          7626 => x"51",
          7627 => x"3f",
          7628 => x"80",
          7629 => x"a9",
          7630 => x"1c",
          7631 => x"81",
          7632 => x"80",
          7633 => x"ae",
          7634 => x"b2",
          7635 => x"1b",
          7636 => x"85",
          7637 => x"ff",
          7638 => x"96",
          7639 => x"9f",
          7640 => x"80",
          7641 => x"34",
          7642 => x"1c",
          7643 => x"81",
          7644 => x"ab",
          7645 => x"a0",
          7646 => x"d4",
          7647 => x"fe",
          7648 => x"59",
          7649 => x"3f",
          7650 => x"53",
          7651 => x"51",
          7652 => x"3f",
          7653 => x"8c",
          7654 => x"e7",
          7655 => x"2e",
          7656 => x"80",
          7657 => x"54",
          7658 => x"53",
          7659 => x"51",
          7660 => x"3f",
          7661 => x"80",
          7662 => x"ff",
          7663 => x"84",
          7664 => x"d2",
          7665 => x"ff",
          7666 => x"86",
          7667 => x"f2",
          7668 => x"1b",
          7669 => x"81",
          7670 => x"52",
          7671 => x"51",
          7672 => x"3f",
          7673 => x"ec",
          7674 => x"9e",
          7675 => x"d4",
          7676 => x"51",
          7677 => x"3f",
          7678 => x"87",
          7679 => x"52",
          7680 => x"9a",
          7681 => x"54",
          7682 => x"7a",
          7683 => x"ff",
          7684 => x"65",
          7685 => x"7a",
          7686 => x"8f",
          7687 => x"80",
          7688 => x"2e",
          7689 => x"9a",
          7690 => x"7a",
          7691 => x"a9",
          7692 => x"84",
          7693 => x"9e",
          7694 => x"0a",
          7695 => x"51",
          7696 => x"ff",
          7697 => x"7d",
          7698 => x"38",
          7699 => x"52",
          7700 => x"9e",
          7701 => x"55",
          7702 => x"62",
          7703 => x"74",
          7704 => x"75",
          7705 => x"7e",
          7706 => x"fe",
          7707 => x"dc",
          7708 => x"38",
          7709 => x"82",
          7710 => x"52",
          7711 => x"9e",
          7712 => x"16",
          7713 => x"56",
          7714 => x"38",
          7715 => x"77",
          7716 => x"8d",
          7717 => x"7d",
          7718 => x"38",
          7719 => x"57",
          7720 => x"83",
          7721 => x"76",
          7722 => x"7a",
          7723 => x"ff",
          7724 => x"82",
          7725 => x"81",
          7726 => x"16",
          7727 => x"56",
          7728 => x"38",
          7729 => x"83",
          7730 => x"86",
          7731 => x"ff",
          7732 => x"38",
          7733 => x"82",
          7734 => x"81",
          7735 => x"06",
          7736 => x"fe",
          7737 => x"53",
          7738 => x"51",
          7739 => x"3f",
          7740 => x"52",
          7741 => x"9c",
          7742 => x"be",
          7743 => x"75",
          7744 => x"81",
          7745 => x"0b",
          7746 => x"77",
          7747 => x"75",
          7748 => x"60",
          7749 => x"80",
          7750 => x"75",
          7751 => x"bc",
          7752 => x"85",
          7753 => x"8c",
          7754 => x"2a",
          7755 => x"75",
          7756 => x"82",
          7757 => x"87",
          7758 => x"52",
          7759 => x"51",
          7760 => x"3f",
          7761 => x"ca",
          7762 => x"9c",
          7763 => x"54",
          7764 => x"52",
          7765 => x"98",
          7766 => x"56",
          7767 => x"08",
          7768 => x"53",
          7769 => x"51",
          7770 => x"3f",
          7771 => x"8c",
          7772 => x"38",
          7773 => x"56",
          7774 => x"56",
          7775 => x"8c",
          7776 => x"75",
          7777 => x"0c",
          7778 => x"04",
          7779 => x"7d",
          7780 => x"80",
          7781 => x"05",
          7782 => x"76",
          7783 => x"38",
          7784 => x"11",
          7785 => x"53",
          7786 => x"79",
          7787 => x"3f",
          7788 => x"09",
          7789 => x"38",
          7790 => x"55",
          7791 => x"db",
          7792 => x"70",
          7793 => x"34",
          7794 => x"74",
          7795 => x"81",
          7796 => x"80",
          7797 => x"55",
          7798 => x"76",
          7799 => x"8c",
          7800 => x"3d",
          7801 => x"3d",
          7802 => x"84",
          7803 => x"33",
          7804 => x"8a",
          7805 => x"06",
          7806 => x"52",
          7807 => x"3f",
          7808 => x"56",
          7809 => x"be",
          7810 => x"08",
          7811 => x"05",
          7812 => x"75",
          7813 => x"56",
          7814 => x"a1",
          7815 => x"fc",
          7816 => x"53",
          7817 => x"76",
          7818 => x"dc",
          7819 => x"32",
          7820 => x"72",
          7821 => x"70",
          7822 => x"56",
          7823 => x"18",
          7824 => x"88",
          7825 => x"3d",
          7826 => x"3d",
          7827 => x"11",
          7828 => x"80",
          7829 => x"38",
          7830 => x"05",
          7831 => x"8c",
          7832 => x"08",
          7833 => x"3f",
          7834 => x"08",
          7835 => x"16",
          7836 => x"09",
          7837 => x"38",
          7838 => x"55",
          7839 => x"55",
          7840 => x"dc",
          7841 => x"0d",
          7842 => x"0d",
          7843 => x"cc",
          7844 => x"73",
          7845 => x"93",
          7846 => x"0c",
          7847 => x"04",
          7848 => x"02",
          7849 => x"33",
          7850 => x"3d",
          7851 => x"54",
          7852 => x"52",
          7853 => x"ae",
          7854 => x"ff",
          7855 => x"3d",
          7856 => x"3d",
          7857 => x"08",
          7858 => x"59",
          7859 => x"80",
          7860 => x"39",
          7861 => x"0c",
          7862 => x"54",
          7863 => x"74",
          7864 => x"a0",
          7865 => x"06",
          7866 => x"15",
          7867 => x"80",
          7868 => x"29",
          7869 => x"05",
          7870 => x"56",
          7871 => x"3f",
          7872 => x"08",
          7873 => x"08",
          7874 => x"76",
          7875 => x"fe",
          7876 => x"82",
          7877 => x"8b",
          7878 => x"33",
          7879 => x"2e",
          7880 => x"81",
          7881 => x"ff",
          7882 => x"98",
          7883 => x"38",
          7884 => x"82",
          7885 => x"8a",
          7886 => x"ff",
          7887 => x"52",
          7888 => x"81",
          7889 => x"84",
          7890 => x"94",
          7891 => x"08",
          7892 => x"c8",
          7893 => x"39",
          7894 => x"51",
          7895 => x"81",
          7896 => x"80",
          7897 => x"fd",
          7898 => x"eb",
          7899 => x"8c",
          7900 => x"39",
          7901 => x"51",
          7902 => x"81",
          7903 => x"80",
          7904 => x"fe",
          7905 => x"cf",
          7906 => x"d8",
          7907 => x"39",
          7908 => x"51",
          7909 => x"81",
          7910 => x"bb",
          7911 => x"a4",
          7912 => x"81",
          7913 => x"af",
          7914 => x"e4",
          7915 => x"81",
          7916 => x"a3",
          7917 => x"98",
          7918 => x"82",
          7919 => x"97",
          7920 => x"c4",
          7921 => x"82",
          7922 => x"8b",
          7923 => x"f4",
          7924 => x"82",
          7925 => x"fe",
          7926 => x"83",
          7927 => x"fb",
          7928 => x"79",
          7929 => x"87",
          7930 => x"38",
          7931 => x"87",
          7932 => x"91",
          7933 => x"52",
          7934 => x"d2",
          7935 => x"8c",
          7936 => x"75",
          7937 => x"d4",
          7938 => x"dc",
          7939 => x"53",
          7940 => x"81",
          7941 => x"f7",
          7942 => x"3d",
          7943 => x"3d",
          7944 => x"84",
          7945 => x"05",
          7946 => x"80",
          7947 => x"70",
          7948 => x"25",
          7949 => x"59",
          7950 => x"87",
          7951 => x"38",
          7952 => x"76",
          7953 => x"ff",
          7954 => x"93",
          7955 => x"80",
          7956 => x"76",
          7957 => x"70",
          7958 => x"bf",
          7959 => x"8c",
          7960 => x"82",
          7961 => x"b8",
          7962 => x"dc",
          7963 => x"98",
          7964 => x"8c",
          7965 => x"96",
          7966 => x"54",
          7967 => x"77",
          7968 => x"c4",
          7969 => x"8c",
          7970 => x"82",
          7971 => x"90",
          7972 => x"74",
          7973 => x"38",
          7974 => x"19",
          7975 => x"39",
          7976 => x"05",
          7977 => x"3f",
          7978 => x"78",
          7979 => x"7b",
          7980 => x"2a",
          7981 => x"57",
          7982 => x"80",
          7983 => x"82",
          7984 => x"87",
          7985 => x"08",
          7986 => x"fe",
          7987 => x"56",
          7988 => x"dc",
          7989 => x"0d",
          7990 => x"0d",
          7991 => x"05",
          7992 => x"57",
          7993 => x"80",
          7994 => x"79",
          7995 => x"3f",
          7996 => x"08",
          7997 => x"80",
          7998 => x"75",
          7999 => x"38",
          8000 => x"55",
          8001 => x"8c",
          8002 => x"52",
          8003 => x"2d",
          8004 => x"08",
          8005 => x"77",
          8006 => x"8c",
          8007 => x"3d",
          8008 => x"3d",
          8009 => x"63",
          8010 => x"80",
          8011 => x"73",
          8012 => x"41",
          8013 => x"5e",
          8014 => x"52",
          8015 => x"51",
          8016 => x"3f",
          8017 => x"51",
          8018 => x"3f",
          8019 => x"79",
          8020 => x"38",
          8021 => x"89",
          8022 => x"2e",
          8023 => x"c6",
          8024 => x"53",
          8025 => x"8e",
          8026 => x"52",
          8027 => x"51",
          8028 => x"3f",
          8029 => x"81",
          8030 => x"ef",
          8031 => x"15",
          8032 => x"39",
          8033 => x"72",
          8034 => x"38",
          8035 => x"82",
          8036 => x"fe",
          8037 => x"89",
          8038 => x"d0",
          8039 => x"e8",
          8040 => x"55",
          8041 => x"18",
          8042 => x"27",
          8043 => x"33",
          8044 => x"dc",
          8045 => x"b4",
          8046 => x"82",
          8047 => x"fe",
          8048 => x"81",
          8049 => x"51",
          8050 => x"3f",
          8051 => x"82",
          8052 => x"fe",
          8053 => x"80",
          8054 => x"27",
          8055 => x"18",
          8056 => x"53",
          8057 => x"7a",
          8058 => x"81",
          8059 => x"9f",
          8060 => x"38",
          8061 => x"73",
          8062 => x"ff",
          8063 => x"72",
          8064 => x"38",
          8065 => x"26",
          8066 => x"51",
          8067 => x"51",
          8068 => x"3f",
          8069 => x"c1",
          8070 => x"ec",
          8071 => x"e8",
          8072 => x"79",
          8073 => x"fe",
          8074 => x"82",
          8075 => x"98",
          8076 => x"2c",
          8077 => x"a0",
          8078 => x"06",
          8079 => x"de",
          8080 => x"8c",
          8081 => x"2b",
          8082 => x"70",
          8083 => x"30",
          8084 => x"70",
          8085 => x"07",
          8086 => x"06",
          8087 => x"59",
          8088 => x"80",
          8089 => x"38",
          8090 => x"09",
          8091 => x"38",
          8092 => x"39",
          8093 => x"72",
          8094 => x"be",
          8095 => x"72",
          8096 => x"0c",
          8097 => x"04",
          8098 => x"02",
          8099 => x"82",
          8100 => x"82",
          8101 => x"55",
          8102 => x"3f",
          8103 => x"22",
          8104 => x"96",
          8105 => x"80",
          8106 => x"8c",
          8107 => x"8d",
          8108 => x"82",
          8109 => x"f2",
          8110 => x"80",
          8111 => x"fe",
          8112 => x"86",
          8113 => x"fe",
          8114 => x"c0",
          8115 => x"53",
          8116 => x"3f",
          8117 => x"d9",
          8118 => x"82",
          8119 => x"db",
          8120 => x"51",
          8121 => x"3f",
          8122 => x"70",
          8123 => x"52",
          8124 => x"95",
          8125 => x"fe",
          8126 => x"82",
          8127 => x"fe",
          8128 => x"80",
          8129 => x"8b",
          8130 => x"2a",
          8131 => x"51",
          8132 => x"2e",
          8133 => x"51",
          8134 => x"3f",
          8135 => x"51",
          8136 => x"3f",
          8137 => x"d8",
          8138 => x"83",
          8139 => x"06",
          8140 => x"80",
          8141 => x"81",
          8142 => x"d7",
          8143 => x"ec",
          8144 => x"cf",
          8145 => x"fe",
          8146 => x"72",
          8147 => x"81",
          8148 => x"71",
          8149 => x"38",
          8150 => x"d8",
          8151 => x"83",
          8152 => x"da",
          8153 => x"51",
          8154 => x"3f",
          8155 => x"70",
          8156 => x"52",
          8157 => x"95",
          8158 => x"fe",
          8159 => x"82",
          8160 => x"fe",
          8161 => x"80",
          8162 => x"87",
          8163 => x"2a",
          8164 => x"51",
          8165 => x"2e",
          8166 => x"51",
          8167 => x"3f",
          8168 => x"51",
          8169 => x"3f",
          8170 => x"d7",
          8171 => x"87",
          8172 => x"06",
          8173 => x"80",
          8174 => x"81",
          8175 => x"d3",
          8176 => x"bc",
          8177 => x"cb",
          8178 => x"fe",
          8179 => x"72",
          8180 => x"81",
          8181 => x"71",
          8182 => x"38",
          8183 => x"d7",
          8184 => x"83",
          8185 => x"d9",
          8186 => x"51",
          8187 => x"3f",
          8188 => x"3f",
          8189 => x"04",
          8190 => x"77",
          8191 => x"a3",
          8192 => x"55",
          8193 => x"52",
          8194 => x"ce",
          8195 => x"89",
          8196 => x"73",
          8197 => x"53",
          8198 => x"52",
          8199 => x"51",
          8200 => x"3f",
          8201 => x"08",
          8202 => x"8c",
          8203 => x"80",
          8204 => x"31",
          8205 => x"73",
          8206 => x"34",
          8207 => x"33",
          8208 => x"2e",
          8209 => x"ac",
          8210 => x"f4",
          8211 => x"75",
          8212 => x"3f",
          8213 => x"08",
          8214 => x"38",
          8215 => x"08",
          8216 => x"a4",
          8217 => x"82",
          8218 => x"c4",
          8219 => x"0b",
          8220 => x"34",
          8221 => x"33",
          8222 => x"2e",
          8223 => x"89",
          8224 => x"75",
          8225 => x"e4",
          8226 => x"82",
          8227 => x"87",
          8228 => x"ce",
          8229 => x"70",
          8230 => x"f0",
          8231 => x"81",
          8232 => x"ff",
          8233 => x"82",
          8234 => x"81",
          8235 => x"78",
          8236 => x"81",
          8237 => x"82",
          8238 => x"96",
          8239 => x"59",
          8240 => x"3f",
          8241 => x"52",
          8242 => x"51",
          8243 => x"3f",
          8244 => x"08",
          8245 => x"38",
          8246 => x"51",
          8247 => x"81",
          8248 => x"82",
          8249 => x"fe",
          8250 => x"96",
          8251 => x"5a",
          8252 => x"79",
          8253 => x"3f",
          8254 => x"84",
          8255 => x"c2",
          8256 => x"dc",
          8257 => x"70",
          8258 => x"59",
          8259 => x"2e",
          8260 => x"78",
          8261 => x"b2",
          8262 => x"2e",
          8263 => x"78",
          8264 => x"38",
          8265 => x"ff",
          8266 => x"bc",
          8267 => x"38",
          8268 => x"78",
          8269 => x"83",
          8270 => x"80",
          8271 => x"dd",
          8272 => x"2e",
          8273 => x"8a",
          8274 => x"80",
          8275 => x"ea",
          8276 => x"f9",
          8277 => x"78",
          8278 => x"88",
          8279 => x"80",
          8280 => x"b1",
          8281 => x"39",
          8282 => x"2e",
          8283 => x"78",
          8284 => x"8b",
          8285 => x"82",
          8286 => x"38",
          8287 => x"78",
          8288 => x"8a",
          8289 => x"93",
          8290 => x"ff",
          8291 => x"ff",
          8292 => x"fe",
          8293 => x"82",
          8294 => x"80",
          8295 => x"38",
          8296 => x"fc",
          8297 => x"84",
          8298 => x"ee",
          8299 => x"8c",
          8300 => x"2e",
          8301 => x"b4",
          8302 => x"11",
          8303 => x"05",
          8304 => x"9d",
          8305 => x"dc",
          8306 => x"82",
          8307 => x"42",
          8308 => x"51",
          8309 => x"3f",
          8310 => x"5a",
          8311 => x"81",
          8312 => x"59",
          8313 => x"84",
          8314 => x"7a",
          8315 => x"38",
          8316 => x"b4",
          8317 => x"11",
          8318 => x"05",
          8319 => x"e1",
          8320 => x"dc",
          8321 => x"fd",
          8322 => x"3d",
          8323 => x"53",
          8324 => x"51",
          8325 => x"3f",
          8326 => x"08",
          8327 => x"c3",
          8328 => x"fe",
          8329 => x"ff",
          8330 => x"fe",
          8331 => x"82",
          8332 => x"80",
          8333 => x"38",
          8334 => x"51",
          8335 => x"3f",
          8336 => x"63",
          8337 => x"38",
          8338 => x"70",
          8339 => x"33",
          8340 => x"81",
          8341 => x"39",
          8342 => x"80",
          8343 => x"84",
          8344 => x"ec",
          8345 => x"8c",
          8346 => x"2e",
          8347 => x"b4",
          8348 => x"11",
          8349 => x"05",
          8350 => x"e5",
          8351 => x"dc",
          8352 => x"fc",
          8353 => x"3d",
          8354 => x"53",
          8355 => x"51",
          8356 => x"3f",
          8357 => x"08",
          8358 => x"c7",
          8359 => x"fc",
          8360 => x"e4",
          8361 => x"79",
          8362 => x"38",
          8363 => x"7b",
          8364 => x"5b",
          8365 => x"92",
          8366 => x"7a",
          8367 => x"53",
          8368 => x"85",
          8369 => x"ea",
          8370 => x"1a",
          8371 => x"43",
          8372 => x"82",
          8373 => x"82",
          8374 => x"3d",
          8375 => x"53",
          8376 => x"51",
          8377 => x"3f",
          8378 => x"08",
          8379 => x"82",
          8380 => x"59",
          8381 => x"89",
          8382 => x"d8",
          8383 => x"cd",
          8384 => x"a1",
          8385 => x"80",
          8386 => x"82",
          8387 => x"44",
          8388 => x"88",
          8389 => x"78",
          8390 => x"38",
          8391 => x"08",
          8392 => x"82",
          8393 => x"59",
          8394 => x"88",
          8395 => x"f0",
          8396 => x"39",
          8397 => x"33",
          8398 => x"2e",
          8399 => x"87",
          8400 => x"89",
          8401 => x"88",
          8402 => x"05",
          8403 => x"fe",
          8404 => x"ff",
          8405 => x"fe",
          8406 => x"82",
          8407 => x"80",
          8408 => x"88",
          8409 => x"78",
          8410 => x"38",
          8411 => x"08",
          8412 => x"39",
          8413 => x"33",
          8414 => x"2e",
          8415 => x"87",
          8416 => x"bb",
          8417 => x"a2",
          8418 => x"80",
          8419 => x"82",
          8420 => x"43",
          8421 => x"88",
          8422 => x"78",
          8423 => x"38",
          8424 => x"08",
          8425 => x"82",
          8426 => x"59",
          8427 => x"88",
          8428 => x"fc",
          8429 => x"39",
          8430 => x"08",
          8431 => x"b4",
          8432 => x"11",
          8433 => x"05",
          8434 => x"95",
          8435 => x"dc",
          8436 => x"a7",
          8437 => x"5c",
          8438 => x"2e",
          8439 => x"5c",
          8440 => x"70",
          8441 => x"07",
          8442 => x"7f",
          8443 => x"5a",
          8444 => x"2e",
          8445 => x"a0",
          8446 => x"88",
          8447 => x"a8",
          8448 => x"84",
          8449 => x"63",
          8450 => x"62",
          8451 => x"f2",
          8452 => x"85",
          8453 => x"e1",
          8454 => x"c7",
          8455 => x"ff",
          8456 => x"ff",
          8457 => x"fe",
          8458 => x"82",
          8459 => x"80",
          8460 => x"38",
          8461 => x"fc",
          8462 => x"84",
          8463 => x"e9",
          8464 => x"8c",
          8465 => x"2e",
          8466 => x"59",
          8467 => x"05",
          8468 => x"63",
          8469 => x"b4",
          8470 => x"11",
          8471 => x"05",
          8472 => x"fd",
          8473 => x"dc",
          8474 => x"f8",
          8475 => x"70",
          8476 => x"82",
          8477 => x"fe",
          8478 => x"80",
          8479 => x"51",
          8480 => x"3f",
          8481 => x"33",
          8482 => x"2e",
          8483 => x"9f",
          8484 => x"38",
          8485 => x"fc",
          8486 => x"84",
          8487 => x"e8",
          8488 => x"8c",
          8489 => x"2e",
          8490 => x"59",
          8491 => x"05",
          8492 => x"63",
          8493 => x"ff",
          8494 => x"85",
          8495 => x"e0",
          8496 => x"aa",
          8497 => x"fe",
          8498 => x"ff",
          8499 => x"fe",
          8500 => x"82",
          8501 => x"80",
          8502 => x"38",
          8503 => x"f0",
          8504 => x"84",
          8505 => x"e9",
          8506 => x"8c",
          8507 => x"2e",
          8508 => x"59",
          8509 => x"22",
          8510 => x"05",
          8511 => x"41",
          8512 => x"f0",
          8513 => x"84",
          8514 => x"e9",
          8515 => x"8c",
          8516 => x"38",
          8517 => x"60",
          8518 => x"52",
          8519 => x"51",
          8520 => x"3f",
          8521 => x"79",
          8522 => x"9a",
          8523 => x"79",
          8524 => x"ae",
          8525 => x"38",
          8526 => x"87",
          8527 => x"05",
          8528 => x"b4",
          8529 => x"11",
          8530 => x"05",
          8531 => x"83",
          8532 => x"dc",
          8533 => x"92",
          8534 => x"02",
          8535 => x"79",
          8536 => x"5b",
          8537 => x"ff",
          8538 => x"85",
          8539 => x"df",
          8540 => x"a3",
          8541 => x"fe",
          8542 => x"ff",
          8543 => x"fe",
          8544 => x"82",
          8545 => x"80",
          8546 => x"38",
          8547 => x"f0",
          8548 => x"84",
          8549 => x"e8",
          8550 => x"8c",
          8551 => x"2e",
          8552 => x"60",
          8553 => x"60",
          8554 => x"b4",
          8555 => x"11",
          8556 => x"05",
          8557 => x"9b",
          8558 => x"dc",
          8559 => x"f6",
          8560 => x"70",
          8561 => x"82",
          8562 => x"fe",
          8563 => x"80",
          8564 => x"51",
          8565 => x"3f",
          8566 => x"33",
          8567 => x"2e",
          8568 => x"9f",
          8569 => x"38",
          8570 => x"f0",
          8571 => x"84",
          8572 => x"e7",
          8573 => x"8c",
          8574 => x"2e",
          8575 => x"60",
          8576 => x"60",
          8577 => x"ff",
          8578 => x"85",
          8579 => x"dd",
          8580 => x"ae",
          8581 => x"ff",
          8582 => x"ff",
          8583 => x"fe",
          8584 => x"82",
          8585 => x"80",
          8586 => x"38",
          8587 => x"85",
          8588 => x"e3",
          8589 => x"59",
          8590 => x"3d",
          8591 => x"53",
          8592 => x"51",
          8593 => x"3f",
          8594 => x"08",
          8595 => x"93",
          8596 => x"82",
          8597 => x"fe",
          8598 => x"63",
          8599 => x"82",
          8600 => x"80",
          8601 => x"38",
          8602 => x"08",
          8603 => x"a8",
          8604 => x"f8",
          8605 => x"39",
          8606 => x"51",
          8607 => x"3f",
          8608 => x"3f",
          8609 => x"82",
          8610 => x"fe",
          8611 => x"80",
          8612 => x"39",
          8613 => x"3f",
          8614 => x"79",
          8615 => x"59",
          8616 => x"f4",
          8617 => x"7d",
          8618 => x"80",
          8619 => x"38",
          8620 => x"84",
          8621 => x"c6",
          8622 => x"8c",
          8623 => x"81",
          8624 => x"2e",
          8625 => x"82",
          8626 => x"7a",
          8627 => x"38",
          8628 => x"7a",
          8629 => x"38",
          8630 => x"82",
          8631 => x"7b",
          8632 => x"f8",
          8633 => x"82",
          8634 => x"b4",
          8635 => x"05",
          8636 => x"8e",
          8637 => x"82",
          8638 => x"b4",
          8639 => x"05",
          8640 => x"fe",
          8641 => x"7b",
          8642 => x"f8",
          8643 => x"82",
          8644 => x"b4",
          8645 => x"05",
          8646 => x"e6",
          8647 => x"7b",
          8648 => x"82",
          8649 => x"b4",
          8650 => x"05",
          8651 => x"d2",
          8652 => x"d8",
          8653 => x"a4",
          8654 => x"64",
          8655 => x"83",
          8656 => x"83",
          8657 => x"b4",
          8658 => x"05",
          8659 => x"3f",
          8660 => x"08",
          8661 => x"08",
          8662 => x"70",
          8663 => x"25",
          8664 => x"5f",
          8665 => x"83",
          8666 => x"81",
          8667 => x"06",
          8668 => x"2e",
          8669 => x"1b",
          8670 => x"06",
          8671 => x"fe",
          8672 => x"81",
          8673 => x"32",
          8674 => x"8a",
          8675 => x"2e",
          8676 => x"f2",
          8677 => x"87",
          8678 => x"e0",
          8679 => x"c3",
          8680 => x"0d",
          8681 => x"8d",
          8682 => x"c0",
          8683 => x"08",
          8684 => x"84",
          8685 => x"51",
          8686 => x"3f",
          8687 => x"08",
          8688 => x"08",
          8689 => x"84",
          8690 => x"51",
          8691 => x"3f",
          8692 => x"dc",
          8693 => x"0c",
          8694 => x"9c",
          8695 => x"55",
          8696 => x"52",
          8697 => x"ba",
          8698 => x"8c",
          8699 => x"2b",
          8700 => x"53",
          8701 => x"52",
          8702 => x"ba",
          8703 => x"82",
          8704 => x"07",
          8705 => x"80",
          8706 => x"c0",
          8707 => x"8c",
          8708 => x"87",
          8709 => x"0c",
          8710 => x"82",
          8711 => x"ba",
          8712 => x"8c",
          8713 => x"cb",
          8714 => x"d4",
          8715 => x"87",
          8716 => x"d9",
          8717 => x"87",
          8718 => x"d9",
          8719 => x"dd",
          8720 => x"d4",
          8721 => x"51",
          8722 => x"f0",
          8723 => x"04",
          8724 => x"22",
          8725 => x"22",
          8726 => x"22",
          8727 => x"22",
          8728 => x"22",
          8729 => x"2f",
          8730 => x"30",
          8731 => x"31",
          8732 => x"31",
          8733 => x"31",
          8734 => x"32",
          8735 => x"2e",
          8736 => x"2e",
          8737 => x"32",
          8738 => x"32",
          8739 => x"33",
          8740 => x"33",
          8741 => x"6b",
          8742 => x"6b",
          8743 => x"6b",
          8744 => x"6b",
          8745 => x"6b",
          8746 => x"6b",
          8747 => x"6b",
          8748 => x"6b",
          8749 => x"6b",
          8750 => x"6b",
          8751 => x"6b",
          8752 => x"6b",
          8753 => x"6b",
          8754 => x"6b",
          8755 => x"6b",
          8756 => x"6b",
          8757 => x"6b",
          8758 => x"6b",
          8759 => x"6b",
          8760 => x"6b",
          8761 => x"2f",
          8762 => x"25",
          8763 => x"64",
          8764 => x"3a",
          8765 => x"25",
          8766 => x"0a",
          8767 => x"43",
          8768 => x"6e",
          8769 => x"75",
          8770 => x"69",
          8771 => x"00",
          8772 => x"66",
          8773 => x"20",
          8774 => x"20",
          8775 => x"66",
          8776 => x"00",
          8777 => x"44",
          8778 => x"63",
          8779 => x"69",
          8780 => x"65",
          8781 => x"74",
          8782 => x"0a",
          8783 => x"20",
          8784 => x"20",
          8785 => x"41",
          8786 => x"28",
          8787 => x"58",
          8788 => x"38",
          8789 => x"0a",
          8790 => x"20",
          8791 => x"52",
          8792 => x"20",
          8793 => x"28",
          8794 => x"58",
          8795 => x"38",
          8796 => x"0a",
          8797 => x"20",
          8798 => x"53",
          8799 => x"52",
          8800 => x"28",
          8801 => x"58",
          8802 => x"38",
          8803 => x"0a",
          8804 => x"20",
          8805 => x"41",
          8806 => x"20",
          8807 => x"28",
          8808 => x"58",
          8809 => x"38",
          8810 => x"0a",
          8811 => x"20",
          8812 => x"4d",
          8813 => x"20",
          8814 => x"28",
          8815 => x"58",
          8816 => x"38",
          8817 => x"0a",
          8818 => x"20",
          8819 => x"20",
          8820 => x"44",
          8821 => x"28",
          8822 => x"69",
          8823 => x"20",
          8824 => x"32",
          8825 => x"0a",
          8826 => x"20",
          8827 => x"4d",
          8828 => x"20",
          8829 => x"28",
          8830 => x"65",
          8831 => x"20",
          8832 => x"32",
          8833 => x"0a",
          8834 => x"20",
          8835 => x"54",
          8836 => x"54",
          8837 => x"28",
          8838 => x"6e",
          8839 => x"73",
          8840 => x"32",
          8841 => x"0a",
          8842 => x"20",
          8843 => x"53",
          8844 => x"4e",
          8845 => x"55",
          8846 => x"00",
          8847 => x"20",
          8848 => x"20",
          8849 => x"0a",
          8850 => x"20",
          8851 => x"43",
          8852 => x"00",
          8853 => x"20",
          8854 => x"32",
          8855 => x"00",
          8856 => x"20",
          8857 => x"49",
          8858 => x"00",
          8859 => x"64",
          8860 => x"73",
          8861 => x"0a",
          8862 => x"20",
          8863 => x"55",
          8864 => x"73",
          8865 => x"56",
          8866 => x"6f",
          8867 => x"64",
          8868 => x"73",
          8869 => x"20",
          8870 => x"58",
          8871 => x"00",
          8872 => x"20",
          8873 => x"55",
          8874 => x"6d",
          8875 => x"20",
          8876 => x"72",
          8877 => x"64",
          8878 => x"73",
          8879 => x"20",
          8880 => x"58",
          8881 => x"00",
          8882 => x"20",
          8883 => x"61",
          8884 => x"53",
          8885 => x"74",
          8886 => x"64",
          8887 => x"73",
          8888 => x"20",
          8889 => x"20",
          8890 => x"58",
          8891 => x"00",
          8892 => x"73",
          8893 => x"00",
          8894 => x"20",
          8895 => x"55",
          8896 => x"20",
          8897 => x"20",
          8898 => x"20",
          8899 => x"20",
          8900 => x"20",
          8901 => x"20",
          8902 => x"58",
          8903 => x"00",
          8904 => x"20",
          8905 => x"73",
          8906 => x"20",
          8907 => x"63",
          8908 => x"72",
          8909 => x"20",
          8910 => x"20",
          8911 => x"20",
          8912 => x"25",
          8913 => x"4d",
          8914 => x"00",
          8915 => x"20",
          8916 => x"52",
          8917 => x"43",
          8918 => x"6b",
          8919 => x"65",
          8920 => x"20",
          8921 => x"20",
          8922 => x"20",
          8923 => x"25",
          8924 => x"4d",
          8925 => x"00",
          8926 => x"20",
          8927 => x"73",
          8928 => x"6e",
          8929 => x"44",
          8930 => x"20",
          8931 => x"63",
          8932 => x"72",
          8933 => x"20",
          8934 => x"25",
          8935 => x"4d",
          8936 => x"00",
          8937 => x"61",
          8938 => x"00",
          8939 => x"64",
          8940 => x"00",
          8941 => x"65",
          8942 => x"00",
          8943 => x"4f",
          8944 => x"4f",
          8945 => x"00",
          8946 => x"6b",
          8947 => x"6e",
          8948 => x"73",
          8949 => x"79",
          8950 => x"74",
          8951 => x"73",
          8952 => x"79",
          8953 => x"73",
          8954 => x"00",
          8955 => x"00",
          8956 => x"34",
          8957 => x"25",
          8958 => x"00",
          8959 => x"69",
          8960 => x"20",
          8961 => x"72",
          8962 => x"74",
          8963 => x"65",
          8964 => x"73",
          8965 => x"79",
          8966 => x"6c",
          8967 => x"6f",
          8968 => x"46",
          8969 => x"00",
          8970 => x"6e",
          8971 => x"20",
          8972 => x"6e",
          8973 => x"65",
          8974 => x"20",
          8975 => x"74",
          8976 => x"20",
          8977 => x"65",
          8978 => x"69",
          8979 => x"6c",
          8980 => x"2e",
          8981 => x"00",
          8982 => x"7d",
          8983 => x"00",
          8984 => x"00",
          8985 => x"7d",
          8986 => x"00",
          8987 => x"00",
          8988 => x"7c",
          8989 => x"00",
          8990 => x"00",
          8991 => x"7c",
          8992 => x"00",
          8993 => x"00",
          8994 => x"7c",
          8995 => x"00",
          8996 => x"00",
          8997 => x"7c",
          8998 => x"00",
          8999 => x"00",
          9000 => x"7c",
          9001 => x"00",
          9002 => x"00",
          9003 => x"7c",
          9004 => x"00",
          9005 => x"00",
          9006 => x"7c",
          9007 => x"00",
          9008 => x"00",
          9009 => x"7c",
          9010 => x"00",
          9011 => x"00",
          9012 => x"7c",
          9013 => x"00",
          9014 => x"00",
          9015 => x"44",
          9016 => x"43",
          9017 => x"42",
          9018 => x"41",
          9019 => x"36",
          9020 => x"35",
          9021 => x"34",
          9022 => x"33",
          9023 => x"31",
          9024 => x"00",
          9025 => x"00",
          9026 => x"00",
          9027 => x"2b",
          9028 => x"3c",
          9029 => x"5b",
          9030 => x"00",
          9031 => x"54",
          9032 => x"54",
          9033 => x"00",
          9034 => x"90",
          9035 => x"4f",
          9036 => x"30",
          9037 => x"20",
          9038 => x"45",
          9039 => x"20",
          9040 => x"33",
          9041 => x"20",
          9042 => x"20",
          9043 => x"45",
          9044 => x"20",
          9045 => x"20",
          9046 => x"20",
          9047 => x"7d",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"45",
          9052 => x"8f",
          9053 => x"45",
          9054 => x"8e",
          9055 => x"92",
          9056 => x"55",
          9057 => x"9a",
          9058 => x"9e",
          9059 => x"4f",
          9060 => x"a6",
          9061 => x"aa",
          9062 => x"ae",
          9063 => x"b2",
          9064 => x"b6",
          9065 => x"ba",
          9066 => x"be",
          9067 => x"c2",
          9068 => x"c6",
          9069 => x"ca",
          9070 => x"ce",
          9071 => x"d2",
          9072 => x"d6",
          9073 => x"da",
          9074 => x"de",
          9075 => x"e2",
          9076 => x"e6",
          9077 => x"ea",
          9078 => x"ee",
          9079 => x"f2",
          9080 => x"f6",
          9081 => x"fa",
          9082 => x"fe",
          9083 => x"2c",
          9084 => x"5d",
          9085 => x"2a",
          9086 => x"3f",
          9087 => x"00",
          9088 => x"00",
          9089 => x"00",
          9090 => x"02",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"6e",
          9097 => x"00",
          9098 => x"6f",
          9099 => x"00",
          9100 => x"6e",
          9101 => x"00",
          9102 => x"6f",
          9103 => x"00",
          9104 => x"78",
          9105 => x"00",
          9106 => x"6c",
          9107 => x"00",
          9108 => x"6f",
          9109 => x"00",
          9110 => x"69",
          9111 => x"00",
          9112 => x"75",
          9113 => x"00",
          9114 => x"62",
          9115 => x"68",
          9116 => x"77",
          9117 => x"64",
          9118 => x"65",
          9119 => x"64",
          9120 => x"65",
          9121 => x"6c",
          9122 => x"00",
          9123 => x"70",
          9124 => x"73",
          9125 => x"74",
          9126 => x"73",
          9127 => x"00",
          9128 => x"66",
          9129 => x"00",
          9130 => x"73",
          9131 => x"00",
          9132 => x"61",
          9133 => x"00",
          9134 => x"61",
          9135 => x"00",
          9136 => x"6c",
          9137 => x"00",
          9138 => x"73",
          9139 => x"72",
          9140 => x"0a",
          9141 => x"74",
          9142 => x"61",
          9143 => x"72",
          9144 => x"2e",
          9145 => x"00",
          9146 => x"73",
          9147 => x"6f",
          9148 => x"65",
          9149 => x"2e",
          9150 => x"00",
          9151 => x"20",
          9152 => x"65",
          9153 => x"75",
          9154 => x"0a",
          9155 => x"20",
          9156 => x"68",
          9157 => x"75",
          9158 => x"0a",
          9159 => x"76",
          9160 => x"64",
          9161 => x"6c",
          9162 => x"6d",
          9163 => x"00",
          9164 => x"63",
          9165 => x"20",
          9166 => x"69",
          9167 => x"0a",
          9168 => x"6c",
          9169 => x"6c",
          9170 => x"64",
          9171 => x"78",
          9172 => x"73",
          9173 => x"00",
          9174 => x"6c",
          9175 => x"61",
          9176 => x"65",
          9177 => x"76",
          9178 => x"64",
          9179 => x"00",
          9180 => x"20",
          9181 => x"77",
          9182 => x"65",
          9183 => x"6f",
          9184 => x"74",
          9185 => x"0a",
          9186 => x"69",
          9187 => x"6e",
          9188 => x"65",
          9189 => x"73",
          9190 => x"76",
          9191 => x"64",
          9192 => x"00",
          9193 => x"73",
          9194 => x"6f",
          9195 => x"6e",
          9196 => x"65",
          9197 => x"00",
          9198 => x"20",
          9199 => x"70",
          9200 => x"62",
          9201 => x"66",
          9202 => x"73",
          9203 => x"65",
          9204 => x"6f",
          9205 => x"20",
          9206 => x"64",
          9207 => x"2e",
          9208 => x"00",
          9209 => x"72",
          9210 => x"20",
          9211 => x"72",
          9212 => x"2e",
          9213 => x"00",
          9214 => x"6d",
          9215 => x"74",
          9216 => x"70",
          9217 => x"74",
          9218 => x"20",
          9219 => x"63",
          9220 => x"65",
          9221 => x"00",
          9222 => x"6c",
          9223 => x"73",
          9224 => x"63",
          9225 => x"2e",
          9226 => x"00",
          9227 => x"73",
          9228 => x"69",
          9229 => x"6e",
          9230 => x"65",
          9231 => x"79",
          9232 => x"00",
          9233 => x"6f",
          9234 => x"6e",
          9235 => x"70",
          9236 => x"66",
          9237 => x"73",
          9238 => x"00",
          9239 => x"72",
          9240 => x"74",
          9241 => x"20",
          9242 => x"6f",
          9243 => x"63",
          9244 => x"00",
          9245 => x"63",
          9246 => x"73",
          9247 => x"00",
          9248 => x"6b",
          9249 => x"6e",
          9250 => x"72",
          9251 => x"0a",
          9252 => x"6c",
          9253 => x"79",
          9254 => x"20",
          9255 => x"61",
          9256 => x"6c",
          9257 => x"79",
          9258 => x"2f",
          9259 => x"2e",
          9260 => x"00",
          9261 => x"61",
          9262 => x"00",
          9263 => x"38",
          9264 => x"00",
          9265 => x"20",
          9266 => x"34",
          9267 => x"00",
          9268 => x"20",
          9269 => x"20",
          9270 => x"00",
          9271 => x"32",
          9272 => x"00",
          9273 => x"00",
          9274 => x"00",
          9275 => x"0a",
          9276 => x"53",
          9277 => x"2a",
          9278 => x"20",
          9279 => x"00",
          9280 => x"2f",
          9281 => x"32",
          9282 => x"00",
          9283 => x"2e",
          9284 => x"00",
          9285 => x"50",
          9286 => x"72",
          9287 => x"25",
          9288 => x"29",
          9289 => x"20",
          9290 => x"2a",
          9291 => x"00",
          9292 => x"55",
          9293 => x"74",
          9294 => x"75",
          9295 => x"48",
          9296 => x"6c",
          9297 => x"00",
          9298 => x"6d",
          9299 => x"69",
          9300 => x"72",
          9301 => x"74",
          9302 => x"00",
          9303 => x"32",
          9304 => x"74",
          9305 => x"75",
          9306 => x"00",
          9307 => x"43",
          9308 => x"52",
          9309 => x"6e",
          9310 => x"72",
          9311 => x"0a",
          9312 => x"43",
          9313 => x"57",
          9314 => x"6e",
          9315 => x"72",
          9316 => x"0a",
          9317 => x"52",
          9318 => x"52",
          9319 => x"6e",
          9320 => x"72",
          9321 => x"0a",
          9322 => x"52",
          9323 => x"54",
          9324 => x"6e",
          9325 => x"72",
          9326 => x"0a",
          9327 => x"52",
          9328 => x"52",
          9329 => x"6e",
          9330 => x"72",
          9331 => x"0a",
          9332 => x"52",
          9333 => x"54",
          9334 => x"6e",
          9335 => x"72",
          9336 => x"0a",
          9337 => x"74",
          9338 => x"67",
          9339 => x"20",
          9340 => x"65",
          9341 => x"2e",
          9342 => x"00",
          9343 => x"61",
          9344 => x"6e",
          9345 => x"69",
          9346 => x"2e",
          9347 => x"00",
          9348 => x"74",
          9349 => x"65",
          9350 => x"61",
          9351 => x"00",
          9352 => x"00",
          9353 => x"69",
          9354 => x"20",
          9355 => x"69",
          9356 => x"69",
          9357 => x"73",
          9358 => x"64",
          9359 => x"72",
          9360 => x"2c",
          9361 => x"65",
          9362 => x"20",
          9363 => x"74",
          9364 => x"6e",
          9365 => x"6c",
          9366 => x"00",
          9367 => x"00",
          9368 => x"65",
          9369 => x"6e",
          9370 => x"2e",
          9371 => x"00",
          9372 => x"70",
          9373 => x"67",
          9374 => x"00",
          9375 => x"6d",
          9376 => x"69",
          9377 => x"2e",
          9378 => x"00",
          9379 => x"38",
          9380 => x"25",
          9381 => x"29",
          9382 => x"30",
          9383 => x"28",
          9384 => x"78",
          9385 => x"00",
          9386 => x"6d",
          9387 => x"65",
          9388 => x"79",
          9389 => x"00",
          9390 => x"6f",
          9391 => x"65",
          9392 => x"0a",
          9393 => x"38",
          9394 => x"30",
          9395 => x"00",
          9396 => x"3f",
          9397 => x"00",
          9398 => x"38",
          9399 => x"30",
          9400 => x"00",
          9401 => x"38",
          9402 => x"30",
          9403 => x"00",
          9404 => x"65",
          9405 => x"69",
          9406 => x"63",
          9407 => x"20",
          9408 => x"30",
          9409 => x"2e",
          9410 => x"00",
          9411 => x"6c",
          9412 => x"67",
          9413 => x"64",
          9414 => x"20",
          9415 => x"78",
          9416 => x"2e",
          9417 => x"00",
          9418 => x"6c",
          9419 => x"65",
          9420 => x"6e",
          9421 => x"63",
          9422 => x"20",
          9423 => x"29",
          9424 => x"00",
          9425 => x"73",
          9426 => x"74",
          9427 => x"20",
          9428 => x"6c",
          9429 => x"74",
          9430 => x"2e",
          9431 => x"00",
          9432 => x"6c",
          9433 => x"65",
          9434 => x"74",
          9435 => x"2e",
          9436 => x"00",
          9437 => x"55",
          9438 => x"6e",
          9439 => x"3a",
          9440 => x"5c",
          9441 => x"25",
          9442 => x"00",
          9443 => x"3a",
          9444 => x"5c",
          9445 => x"00",
          9446 => x"3a",
          9447 => x"00",
          9448 => x"64",
          9449 => x"6d",
          9450 => x"64",
          9451 => x"00",
          9452 => x"6e",
          9453 => x"67",
          9454 => x"0a",
          9455 => x"61",
          9456 => x"6e",
          9457 => x"6e",
          9458 => x"72",
          9459 => x"73",
          9460 => x"0a",
          9461 => x"00",
          9462 => x"00",
          9463 => x"7f",
          9464 => x"00",
          9465 => x"7f",
          9466 => x"00",
          9467 => x"7f",
          9468 => x"00",
          9469 => x"00",
          9470 => x"00",
          9471 => x"ff",
          9472 => x"00",
          9473 => x"00",
          9474 => x"78",
          9475 => x"00",
          9476 => x"e1",
          9477 => x"e1",
          9478 => x"e1",
          9479 => x"00",
          9480 => x"01",
          9481 => x"01",
          9482 => x"10",
          9483 => x"00",
          9484 => x"00",
          9485 => x"00",
          9486 => x"00",
          9487 => x"84",
          9488 => x"84",
          9489 => x"84",
          9490 => x"84",
          9491 => x"7b",
          9492 => x"00",
          9493 => x"00",
          9494 => x"00",
          9495 => x"00",
          9496 => x"00",
          9497 => x"00",
          9498 => x"00",
          9499 => x"00",
          9500 => x"00",
          9501 => x"00",
          9502 => x"00",
          9503 => x"00",
          9504 => x"00",
          9505 => x"00",
          9506 => x"00",
          9507 => x"00",
          9508 => x"00",
          9509 => x"00",
          9510 => x"00",
          9511 => x"00",
          9512 => x"00",
          9513 => x"00",
          9514 => x"00",
          9515 => x"7b",
          9516 => x"00",
          9517 => x"7b",
          9518 => x"00",
          9519 => x"7b",
          9520 => x"00",
          9521 => x"00",
          9522 => x"00",
          9523 => x"7e",
          9524 => x"01",
          9525 => x"00",
          9526 => x"00",
          9527 => x"7e",
          9528 => x"01",
          9529 => x"00",
          9530 => x"00",
          9531 => x"7e",
          9532 => x"03",
          9533 => x"00",
          9534 => x"00",
          9535 => x"7e",
          9536 => x"03",
          9537 => x"00",
          9538 => x"00",
          9539 => x"7e",
          9540 => x"03",
          9541 => x"00",
          9542 => x"00",
          9543 => x"7e",
          9544 => x"04",
          9545 => x"00",
          9546 => x"00",
          9547 => x"7e",
          9548 => x"04",
          9549 => x"00",
          9550 => x"00",
          9551 => x"7e",
          9552 => x"04",
          9553 => x"00",
          9554 => x"00",
          9555 => x"7e",
          9556 => x"04",
          9557 => x"00",
          9558 => x"00",
          9559 => x"7e",
          9560 => x"04",
          9561 => x"00",
          9562 => x"00",
          9563 => x"7e",
          9564 => x"04",
          9565 => x"00",
          9566 => x"00",
          9567 => x"7e",
          9568 => x"04",
          9569 => x"00",
          9570 => x"00",
          9571 => x"7e",
          9572 => x"05",
          9573 => x"00",
          9574 => x"00",
          9575 => x"7e",
          9576 => x"05",
          9577 => x"00",
          9578 => x"00",
          9579 => x"7e",
          9580 => x"05",
          9581 => x"00",
          9582 => x"00",
          9583 => x"7e",
          9584 => x"05",
          9585 => x"00",
          9586 => x"00",
          9587 => x"7e",
          9588 => x"07",
          9589 => x"00",
          9590 => x"00",
          9591 => x"7e",
          9592 => x"07",
          9593 => x"00",
          9594 => x"00",
          9595 => x"7e",
          9596 => x"08",
          9597 => x"00",
          9598 => x"00",
          9599 => x"7e",
          9600 => x"08",
          9601 => x"00",
          9602 => x"00",
          9603 => x"7e",
          9604 => x"08",
          9605 => x"00",
          9606 => x"00",
          9607 => x"7e",
          9608 => x"08",
          9609 => x"00",
          9610 => x"00",
          9611 => x"7e",
          9612 => x"09",
          9613 => x"00",
          9614 => x"00",
          9615 => x"7e",
          9616 => x"09",
          9617 => x"00",
          9618 => x"00",
          9619 => x"7e",
          9620 => x"09",
          9621 => x"00",
          9622 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"f4",
           281 => x"27",
           282 => x"71",
           283 => x"53",
           284 => x"0b",
           285 => x"88",
           286 => x"9d",
           287 => x"04",
           288 => x"04",
           289 => x"94",
           290 => x"0c",
           291 => x"80",
           292 => x"8c",
           293 => x"94",
           294 => x"08",
           295 => x"3f",
           296 => x"88",
           297 => x"3d",
           298 => x"04",
           299 => x"94",
           300 => x"0d",
           301 => x"08",
           302 => x"52",
           303 => x"05",
           304 => x"b9",
           305 => x"70",
           306 => x"85",
           307 => x"0c",
           308 => x"02",
           309 => x"3d",
           310 => x"94",
           311 => x"0c",
           312 => x"05",
           313 => x"ab",
           314 => x"88",
           315 => x"94",
           316 => x"0c",
           317 => x"08",
           318 => x"94",
           319 => x"08",
           320 => x"0b",
           321 => x"05",
           322 => x"f4",
           323 => x"08",
           324 => x"94",
           325 => x"08",
           326 => x"38",
           327 => x"05",
           328 => x"08",
           329 => x"80",
           330 => x"f0",
           331 => x"08",
           332 => x"88",
           333 => x"94",
           334 => x"0c",
           335 => x"05",
           336 => x"fc",
           337 => x"53",
           338 => x"05",
           339 => x"08",
           340 => x"51",
           341 => x"88",
           342 => x"08",
           343 => x"54",
           344 => x"05",
           345 => x"8c",
           346 => x"f8",
           347 => x"94",
           348 => x"0c",
           349 => x"05",
           350 => x"0c",
           351 => x"0d",
           352 => x"94",
           353 => x"0c",
           354 => x"80",
           355 => x"fc",
           356 => x"08",
           357 => x"80",
           358 => x"94",
           359 => x"08",
           360 => x"88",
           361 => x"0b",
           362 => x"05",
           363 => x"8c",
           364 => x"25",
           365 => x"08",
           366 => x"30",
           367 => x"05",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"ad",
           372 => x"70",
           373 => x"05",
           374 => x"08",
           375 => x"80",
           376 => x"94",
           377 => x"08",
           378 => x"f8",
           379 => x"08",
           380 => x"70",
           381 => x"87",
           382 => x"0c",
           383 => x"02",
           384 => x"3d",
           385 => x"94",
           386 => x"0c",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"05",
           391 => x"38",
           392 => x"05",
           393 => x"a3",
           394 => x"94",
           395 => x"08",
           396 => x"94",
           397 => x"08",
           398 => x"8c",
           399 => x"08",
           400 => x"10",
           401 => x"05",
           402 => x"94",
           403 => x"08",
           404 => x"c9",
           405 => x"8c",
           406 => x"08",
           407 => x"26",
           408 => x"08",
           409 => x"94",
           410 => x"08",
           411 => x"88",
           412 => x"08",
           413 => x"94",
           414 => x"08",
           415 => x"f8",
           416 => x"08",
           417 => x"81",
           418 => x"fc",
           419 => x"08",
           420 => x"81",
           421 => x"8c",
           422 => x"af",
           423 => x"90",
           424 => x"2e",
           425 => x"08",
           426 => x"70",
           427 => x"05",
           428 => x"39",
           429 => x"05",
           430 => x"08",
           431 => x"51",
           432 => x"05",
           433 => x"85",
           434 => x"0c",
           435 => x"0d",
           436 => x"87",
           437 => x"0c",
           438 => x"c0",
           439 => x"85",
           440 => x"98",
           441 => x"c0",
           442 => x"70",
           443 => x"51",
           444 => x"8a",
           445 => x"98",
           446 => x"70",
           447 => x"c0",
           448 => x"fc",
           449 => x"52",
           450 => x"87",
           451 => x"08",
           452 => x"2e",
           453 => x"0b",
           454 => x"f0",
           455 => x"0b",
           456 => x"88",
           457 => x"0d",
           458 => x"0d",
           459 => x"56",
           460 => x"0b",
           461 => x"9f",
           462 => x"06",
           463 => x"52",
           464 => x"09",
           465 => x"9e",
           466 => x"87",
           467 => x"0c",
           468 => x"92",
           469 => x"0b",
           470 => x"8c",
           471 => x"92",
           472 => x"85",
           473 => x"06",
           474 => x"70",
           475 => x"38",
           476 => x"84",
           477 => x"ff",
           478 => x"27",
           479 => x"73",
           480 => x"38",
           481 => x"8b",
           482 => x"70",
           483 => x"34",
           484 => x"81",
           485 => x"a2",
           486 => x"80",
           487 => x"87",
           488 => x"08",
           489 => x"b5",
           490 => x"98",
           491 => x"70",
           492 => x"0b",
           493 => x"8c",
           494 => x"92",
           495 => x"82",
           496 => x"70",
           497 => x"73",
           498 => x"06",
           499 => x"72",
           500 => x"06",
           501 => x"c0",
           502 => x"51",
           503 => x"09",
           504 => x"38",
           505 => x"88",
           506 => x"0d",
           507 => x"0d",
           508 => x"33",
           509 => x"88",
           510 => x"0c",
           511 => x"3d",
           512 => x"3d",
           513 => x"11",
           514 => x"33",
           515 => x"71",
           516 => x"81",
           517 => x"72",
           518 => x"75",
           519 => x"88",
           520 => x"54",
           521 => x"85",
           522 => x"f9",
           523 => x"0b",
           524 => x"f4",
           525 => x"81",
           526 => x"ed",
           527 => x"17",
           528 => x"e5",
           529 => x"55",
           530 => x"89",
           531 => x"2e",
           532 => x"d5",
           533 => x"76",
           534 => x"06",
           535 => x"2a",
           536 => x"05",
           537 => x"70",
           538 => x"bd",
           539 => x"b9",
           540 => x"fe",
           541 => x"08",
           542 => x"06",
           543 => x"84",
           544 => x"2b",
           545 => x"53",
           546 => x"8c",
           547 => x"52",
           548 => x"52",
           549 => x"3f",
           550 => x"38",
           551 => x"e2",
           552 => x"f0",
           553 => x"83",
           554 => x"74",
           555 => x"3d",
           556 => x"3d",
           557 => x"0b",
           558 => x"fe",
           559 => x"08",
           560 => x"56",
           561 => x"74",
           562 => x"38",
           563 => x"75",
           564 => x"16",
           565 => x"53",
           566 => x"87",
           567 => x"fd",
           568 => x"54",
           569 => x"0b",
           570 => x"08",
           571 => x"53",
           572 => x"2e",
           573 => x"8c",
           574 => x"51",
           575 => x"88",
           576 => x"53",
           577 => x"fd",
           578 => x"08",
           579 => x"06",
           580 => x"0c",
           581 => x"04",
           582 => x"76",
           583 => x"9f",
           584 => x"55",
           585 => x"88",
           586 => x"72",
           587 => x"38",
           588 => x"73",
           589 => x"81",
           590 => x"72",
           591 => x"33",
           592 => x"2e",
           593 => x"85",
           594 => x"08",
           595 => x"16",
           596 => x"2e",
           597 => x"51",
           598 => x"88",
           599 => x"39",
           600 => x"52",
           601 => x"0c",
           602 => x"88",
           603 => x"0d",
           604 => x"0d",
           605 => x"0b",
           606 => x"71",
           607 => x"70",
           608 => x"06",
           609 => x"55",
           610 => x"88",
           611 => x"08",
           612 => x"38",
           613 => x"dc",
           614 => x"06",
           615 => x"cf",
           616 => x"90",
           617 => x"15",
           618 => x"8f",
           619 => x"84",
           620 => x"52",
           621 => x"bc",
           622 => x"82",
           623 => x"05",
           624 => x"06",
           625 => x"38",
           626 => x"df",
           627 => x"71",
           628 => x"a0",
           629 => x"88",
           630 => x"08",
           631 => x"88",
           632 => x"0c",
           633 => x"fd",
           634 => x"08",
           635 => x"73",
           636 => x"52",
           637 => x"88",
           638 => x"f2",
           639 => x"62",
           640 => x"5c",
           641 => x"74",
           642 => x"81",
           643 => x"81",
           644 => x"56",
           645 => x"70",
           646 => x"74",
           647 => x"81",
           648 => x"81",
           649 => x"0b",
           650 => x"62",
           651 => x"55",
           652 => x"8f",
           653 => x"fd",
           654 => x"08",
           655 => x"34",
           656 => x"93",
           657 => x"08",
           658 => x"5f",
           659 => x"76",
           660 => x"58",
           661 => x"55",
           662 => x"09",
           663 => x"38",
           664 => x"5b",
           665 => x"5f",
           666 => x"1c",
           667 => x"06",
           668 => x"33",
           669 => x"70",
           670 => x"27",
           671 => x"07",
           672 => x"5b",
           673 => x"55",
           674 => x"38",
           675 => x"09",
           676 => x"38",
           677 => x"7a",
           678 => x"55",
           679 => x"9f",
           680 => x"32",
           681 => x"ae",
           682 => x"70",
           683 => x"2a",
           684 => x"51",
           685 => x"38",
           686 => x"5a",
           687 => x"77",
           688 => x"81",
           689 => x"1c",
           690 => x"55",
           691 => x"ff",
           692 => x"1e",
           693 => x"55",
           694 => x"83",
           695 => x"74",
           696 => x"7b",
           697 => x"3f",
           698 => x"ef",
           699 => x"7b",
           700 => x"2b",
           701 => x"54",
           702 => x"08",
           703 => x"f8",
           704 => x"08",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"8b",
           709 => x"83",
           710 => x"06",
           711 => x"74",
           712 => x"7d",
           713 => x"88",
           714 => x"5b",
           715 => x"58",
           716 => x"9a",
           717 => x"81",
           718 => x"79",
           719 => x"5b",
           720 => x"31",
           721 => x"75",
           722 => x"38",
           723 => x"80",
           724 => x"7b",
           725 => x"3f",
           726 => x"88",
           727 => x"08",
           728 => x"39",
           729 => x"1c",
           730 => x"33",
           731 => x"a5",
           732 => x"33",
           733 => x"70",
           734 => x"56",
           735 => x"38",
           736 => x"39",
           737 => x"39",
           738 => x"d3",
           739 => x"88",
           740 => x"af",
           741 => x"0c",
           742 => x"04",
           743 => x"79",
           744 => x"82",
           745 => x"53",
           746 => x"51",
           747 => x"83",
           748 => x"80",
           749 => x"51",
           750 => x"88",
           751 => x"ff",
           752 => x"56",
           753 => x"d5",
           754 => x"06",
           755 => x"75",
           756 => x"77",
           757 => x"f6",
           758 => x"08",
           759 => x"94",
           760 => x"f8",
           761 => x"08",
           762 => x"06",
           763 => x"82",
           764 => x"38",
           765 => x"d2",
           766 => x"76",
           767 => x"3f",
           768 => x"88",
           769 => x"76",
           770 => x"3f",
           771 => x"ff",
           772 => x"74",
           773 => x"2e",
           774 => x"56",
           775 => x"89",
           776 => x"ed",
           777 => x"59",
           778 => x"0b",
           779 => x"0c",
           780 => x"88",
           781 => x"55",
           782 => x"82",
           783 => x"75",
           784 => x"70",
           785 => x"fe",
           786 => x"08",
           787 => x"57",
           788 => x"09",
           789 => x"38",
           790 => x"be",
           791 => x"75",
           792 => x"3f",
           793 => x"38",
           794 => x"55",
           795 => x"ac",
           796 => x"e4",
           797 => x"8a",
           798 => x"88",
           799 => x"52",
           800 => x"3f",
           801 => x"ff",
           802 => x"83",
           803 => x"06",
           804 => x"56",
           805 => x"76",
           806 => x"38",
           807 => x"8f",
           808 => x"8d",
           809 => x"75",
           810 => x"3f",
           811 => x"08",
           812 => x"95",
           813 => x"51",
           814 => x"88",
           815 => x"ff",
           816 => x"8c",
           817 => x"f3",
           818 => x"b6",
           819 => x"58",
           820 => x"33",
           821 => x"02",
           822 => x"05",
           823 => x"59",
           824 => x"3f",
           825 => x"ff",
           826 => x"05",
           827 => x"8c",
           828 => x"1a",
           829 => x"e0",
           830 => x"f1",
           831 => x"84",
           832 => x"3d",
           833 => x"f5",
           834 => x"08",
           835 => x"06",
           836 => x"38",
           837 => x"05",
           838 => x"3f",
           839 => x"7a",
           840 => x"3f",
           841 => x"ff",
           842 => x"71",
           843 => x"84",
           844 => x"84",
           845 => x"33",
           846 => x"31",
           847 => x"51",
           848 => x"3f",
           849 => x"05",
           850 => x"0c",
           851 => x"8a",
           852 => x"74",
           853 => x"26",
           854 => x"57",
           855 => x"76",
           856 => x"83",
           857 => x"86",
           858 => x"2e",
           859 => x"76",
           860 => x"83",
           861 => x"06",
           862 => x"3d",
           863 => x"f5",
           864 => x"08",
           865 => x"88",
           866 => x"08",
           867 => x"0c",
           868 => x"ff",
           869 => x"08",
           870 => x"2a",
           871 => x"0c",
           872 => x"81",
           873 => x"0b",
           874 => x"f4",
           875 => x"75",
           876 => x"3d",
           877 => x"3d",
           878 => x"0b",
           879 => x"55",
           880 => x"80",
           881 => x"38",
           882 => x"16",
           883 => x"e0",
           884 => x"54",
           885 => x"54",
           886 => x"51",
           887 => x"88",
           888 => x"08",
           889 => x"88",
           890 => x"73",
           891 => x"38",
           892 => x"33",
           893 => x"70",
           894 => x"55",
           895 => x"2e",
           896 => x"54",
           897 => x"51",
           898 => x"88",
           899 => x"0c",
           900 => x"05",
           901 => x"3f",
           902 => x"16",
           903 => x"16",
           904 => x"81",
           905 => x"88",
           906 => x"0d",
           907 => x"0d",
           908 => x"0b",
           909 => x"f4",
           910 => x"5c",
           911 => x"0c",
           912 => x"80",
           913 => x"38",
           914 => x"81",
           915 => x"57",
           916 => x"81",
           917 => x"39",
           918 => x"34",
           919 => x"0b",
           920 => x"81",
           921 => x"39",
           922 => x"98",
           923 => x"55",
           924 => x"83",
           925 => x"77",
           926 => x"9a",
           927 => x"08",
           928 => x"06",
           929 => x"80",
           930 => x"16",
           931 => x"77",
           932 => x"70",
           933 => x"5b",
           934 => x"38",
           935 => x"a0",
           936 => x"8b",
           937 => x"08",
           938 => x"3f",
           939 => x"81",
           940 => x"aa",
           941 => x"17",
           942 => x"08",
           943 => x"3f",
           944 => x"88",
           945 => x"ff",
           946 => x"08",
           947 => x"0c",
           948 => x"83",
           949 => x"80",
           950 => x"55",
           951 => x"83",
           952 => x"74",
           953 => x"08",
           954 => x"53",
           955 => x"52",
           956 => x"b5",
           957 => x"fe",
           958 => x"16",
           959 => x"17",
           960 => x"31",
           961 => x"7c",
           962 => x"80",
           963 => x"38",
           964 => x"fe",
           965 => x"57",
           966 => x"8c",
           967 => x"fb",
           968 => x"c0",
           969 => x"54",
           970 => x"52",
           971 => x"d7",
           972 => x"90",
           973 => x"94",
           974 => x"54",
           975 => x"52",
           976 => x"c3",
           977 => x"08",
           978 => x"94",
           979 => x"c0",
           980 => x"54",
           981 => x"52",
           982 => x"ab",
           983 => x"90",
           984 => x"94",
           985 => x"54",
           986 => x"52",
           987 => x"97",
           988 => x"08",
           989 => x"94",
           990 => x"80",
           991 => x"c0",
           992 => x"8c",
           993 => x"87",
           994 => x"0c",
           995 => x"f9",
           996 => x"08",
           997 => x"e0",
           998 => x"3f",
           999 => x"38",
          1000 => x"88",
          1001 => x"98",
          1002 => x"87",
          1003 => x"53",
          1004 => x"74",
          1005 => x"3f",
          1006 => x"38",
          1007 => x"80",
          1008 => x"73",
          1009 => x"39",
          1010 => x"73",
          1011 => x"fb",
          1012 => x"ff",
          1013 => x"00",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"49",
          1018 => x"52",
          1019 => x"00",
          1020 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"aa",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"04",
          2058 => x"a4",
          2059 => x"0b",
          2060 => x"04",
          2061 => x"a4",
          2062 => x"0b",
          2063 => x"04",
          2064 => x"a4",
          2065 => x"0b",
          2066 => x"04",
          2067 => x"a4",
          2068 => x"0b",
          2069 => x"04",
          2070 => x"a5",
          2071 => x"0b",
          2072 => x"04",
          2073 => x"a5",
          2074 => x"0b",
          2075 => x"04",
          2076 => x"a5",
          2077 => x"0b",
          2078 => x"04",
          2079 => x"a5",
          2080 => x"0b",
          2081 => x"04",
          2082 => x"a6",
          2083 => x"0b",
          2084 => x"04",
          2085 => x"a6",
          2086 => x"0b",
          2087 => x"04",
          2088 => x"a6",
          2089 => x"0b",
          2090 => x"04",
          2091 => x"a6",
          2092 => x"0b",
          2093 => x"04",
          2094 => x"a6",
          2095 => x"0b",
          2096 => x"04",
          2097 => x"a7",
          2098 => x"0b",
          2099 => x"04",
          2100 => x"a7",
          2101 => x"0b",
          2102 => x"04",
          2103 => x"a7",
          2104 => x"0b",
          2105 => x"04",
          2106 => x"a7",
          2107 => x"0b",
          2108 => x"04",
          2109 => x"a8",
          2110 => x"0b",
          2111 => x"04",
          2112 => x"a8",
          2113 => x"0b",
          2114 => x"04",
          2115 => x"a8",
          2116 => x"0b",
          2117 => x"04",
          2118 => x"a8",
          2119 => x"0b",
          2120 => x"04",
          2121 => x"a9",
          2122 => x"0b",
          2123 => x"04",
          2124 => x"a9",
          2125 => x"0b",
          2126 => x"04",
          2127 => x"a9",
          2128 => x"0b",
          2129 => x"04",
          2130 => x"a9",
          2131 => x"0b",
          2132 => x"04",
          2133 => x"aa",
          2134 => x"0b",
          2135 => x"04",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"a4",
          2177 => x"8c",
          2178 => x"a0",
          2179 => x"e8",
          2180 => x"90",
          2181 => x"e8",
          2182 => x"aa",
          2183 => x"e8",
          2184 => x"90",
          2185 => x"e8",
          2186 => x"e9",
          2187 => x"e8",
          2188 => x"90",
          2189 => x"e8",
          2190 => x"87",
          2191 => x"e8",
          2192 => x"90",
          2193 => x"e8",
          2194 => x"c5",
          2195 => x"e8",
          2196 => x"90",
          2197 => x"e8",
          2198 => x"c3",
          2199 => x"e8",
          2200 => x"90",
          2201 => x"e8",
          2202 => x"aa",
          2203 => x"e8",
          2204 => x"90",
          2205 => x"e8",
          2206 => x"e0",
          2207 => x"e8",
          2208 => x"90",
          2209 => x"e8",
          2210 => x"d2",
          2211 => x"e8",
          2212 => x"90",
          2213 => x"e8",
          2214 => x"eb",
          2215 => x"e8",
          2216 => x"90",
          2217 => x"e8",
          2218 => x"dc",
          2219 => x"e8",
          2220 => x"90",
          2221 => x"e8",
          2222 => x"81",
          2223 => x"e8",
          2224 => x"90",
          2225 => x"e8",
          2226 => x"a5",
          2227 => x"e8",
          2228 => x"90",
          2229 => x"e8",
          2230 => x"2d",
          2231 => x"08",
          2232 => x"04",
          2233 => x"0c",
          2234 => x"82",
          2235 => x"83",
          2236 => x"82",
          2237 => x"b3",
          2238 => x"8c",
          2239 => x"80",
          2240 => x"8c",
          2241 => x"cf",
          2242 => x"e8",
          2243 => x"90",
          2244 => x"e8",
          2245 => x"2d",
          2246 => x"08",
          2247 => x"04",
          2248 => x"0c",
          2249 => x"2d",
          2250 => x"08",
          2251 => x"04",
          2252 => x"0c",
          2253 => x"2d",
          2254 => x"08",
          2255 => x"04",
          2256 => x"0c",
          2257 => x"2d",
          2258 => x"08",
          2259 => x"04",
          2260 => x"0c",
          2261 => x"2d",
          2262 => x"08",
          2263 => x"04",
          2264 => x"0c",
          2265 => x"2d",
          2266 => x"08",
          2267 => x"04",
          2268 => x"0c",
          2269 => x"2d",
          2270 => x"08",
          2271 => x"04",
          2272 => x"0c",
          2273 => x"2d",
          2274 => x"08",
          2275 => x"04",
          2276 => x"0c",
          2277 => x"2d",
          2278 => x"08",
          2279 => x"04",
          2280 => x"0c",
          2281 => x"2d",
          2282 => x"08",
          2283 => x"04",
          2284 => x"0c",
          2285 => x"2d",
          2286 => x"08",
          2287 => x"04",
          2288 => x"0c",
          2289 => x"2d",
          2290 => x"08",
          2291 => x"04",
          2292 => x"0c",
          2293 => x"2d",
          2294 => x"08",
          2295 => x"04",
          2296 => x"0c",
          2297 => x"2d",
          2298 => x"08",
          2299 => x"04",
          2300 => x"0c",
          2301 => x"2d",
          2302 => x"08",
          2303 => x"04",
          2304 => x"0c",
          2305 => x"2d",
          2306 => x"08",
          2307 => x"04",
          2308 => x"0c",
          2309 => x"2d",
          2310 => x"08",
          2311 => x"04",
          2312 => x"0c",
          2313 => x"2d",
          2314 => x"08",
          2315 => x"04",
          2316 => x"0c",
          2317 => x"2d",
          2318 => x"08",
          2319 => x"04",
          2320 => x"0c",
          2321 => x"2d",
          2322 => x"08",
          2323 => x"04",
          2324 => x"0c",
          2325 => x"2d",
          2326 => x"08",
          2327 => x"04",
          2328 => x"0c",
          2329 => x"2d",
          2330 => x"08",
          2331 => x"04",
          2332 => x"0c",
          2333 => x"2d",
          2334 => x"08",
          2335 => x"04",
          2336 => x"0c",
          2337 => x"2d",
          2338 => x"08",
          2339 => x"04",
          2340 => x"0c",
          2341 => x"2d",
          2342 => x"08",
          2343 => x"04",
          2344 => x"0c",
          2345 => x"2d",
          2346 => x"08",
          2347 => x"04",
          2348 => x"0c",
          2349 => x"2d",
          2350 => x"08",
          2351 => x"04",
          2352 => x"0c",
          2353 => x"2d",
          2354 => x"08",
          2355 => x"04",
          2356 => x"0c",
          2357 => x"2d",
          2358 => x"08",
          2359 => x"04",
          2360 => x"0c",
          2361 => x"2d",
          2362 => x"08",
          2363 => x"04",
          2364 => x"0c",
          2365 => x"2d",
          2366 => x"08",
          2367 => x"04",
          2368 => x"0c",
          2369 => x"82",
          2370 => x"83",
          2371 => x"82",
          2372 => x"b4",
          2373 => x"8c",
          2374 => x"80",
          2375 => x"8c",
          2376 => x"92",
          2377 => x"e8",
          2378 => x"90",
          2379 => x"e8",
          2380 => x"ba",
          2381 => x"e8",
          2382 => x"90",
          2383 => x"dc",
          2384 => x"9c",
          2385 => x"80",
          2386 => x"05",
          2387 => x"0b",
          2388 => x"04",
          2389 => x"81",
          2390 => x"3c",
          2391 => x"e8",
          2392 => x"8c",
          2393 => x"3d",
          2394 => x"82",
          2395 => x"8c",
          2396 => x"82",
          2397 => x"88",
          2398 => x"80",
          2399 => x"8c",
          2400 => x"82",
          2401 => x"54",
          2402 => x"82",
          2403 => x"04",
          2404 => x"08",
          2405 => x"e8",
          2406 => x"0d",
          2407 => x"8c",
          2408 => x"05",
          2409 => x"8c",
          2410 => x"05",
          2411 => x"3f",
          2412 => x"08",
          2413 => x"dc",
          2414 => x"3d",
          2415 => x"e8",
          2416 => x"8c",
          2417 => x"82",
          2418 => x"fd",
          2419 => x"0b",
          2420 => x"08",
          2421 => x"80",
          2422 => x"e8",
          2423 => x"0c",
          2424 => x"08",
          2425 => x"82",
          2426 => x"88",
          2427 => x"b9",
          2428 => x"e8",
          2429 => x"08",
          2430 => x"38",
          2431 => x"8c",
          2432 => x"05",
          2433 => x"38",
          2434 => x"08",
          2435 => x"10",
          2436 => x"08",
          2437 => x"82",
          2438 => x"fc",
          2439 => x"82",
          2440 => x"fc",
          2441 => x"b8",
          2442 => x"e8",
          2443 => x"08",
          2444 => x"e1",
          2445 => x"e8",
          2446 => x"08",
          2447 => x"08",
          2448 => x"26",
          2449 => x"8c",
          2450 => x"05",
          2451 => x"e8",
          2452 => x"08",
          2453 => x"e8",
          2454 => x"0c",
          2455 => x"08",
          2456 => x"82",
          2457 => x"fc",
          2458 => x"82",
          2459 => x"f8",
          2460 => x"8c",
          2461 => x"05",
          2462 => x"82",
          2463 => x"fc",
          2464 => x"8c",
          2465 => x"05",
          2466 => x"82",
          2467 => x"8c",
          2468 => x"95",
          2469 => x"e8",
          2470 => x"08",
          2471 => x"38",
          2472 => x"08",
          2473 => x"70",
          2474 => x"08",
          2475 => x"51",
          2476 => x"8c",
          2477 => x"05",
          2478 => x"8c",
          2479 => x"05",
          2480 => x"8c",
          2481 => x"05",
          2482 => x"dc",
          2483 => x"0d",
          2484 => x"0c",
          2485 => x"0d",
          2486 => x"7b",
          2487 => x"55",
          2488 => x"8c",
          2489 => x"07",
          2490 => x"70",
          2491 => x"38",
          2492 => x"71",
          2493 => x"38",
          2494 => x"05",
          2495 => x"70",
          2496 => x"34",
          2497 => x"71",
          2498 => x"81",
          2499 => x"74",
          2500 => x"0c",
          2501 => x"04",
          2502 => x"70",
          2503 => x"08",
          2504 => x"05",
          2505 => x"70",
          2506 => x"08",
          2507 => x"05",
          2508 => x"70",
          2509 => x"08",
          2510 => x"05",
          2511 => x"70",
          2512 => x"08",
          2513 => x"05",
          2514 => x"12",
          2515 => x"26",
          2516 => x"72",
          2517 => x"72",
          2518 => x"54",
          2519 => x"84",
          2520 => x"fc",
          2521 => x"83",
          2522 => x"70",
          2523 => x"39",
          2524 => x"76",
          2525 => x"8c",
          2526 => x"33",
          2527 => x"55",
          2528 => x"8a",
          2529 => x"06",
          2530 => x"2e",
          2531 => x"12",
          2532 => x"2e",
          2533 => x"73",
          2534 => x"55",
          2535 => x"52",
          2536 => x"09",
          2537 => x"38",
          2538 => x"dc",
          2539 => x"0d",
          2540 => x"88",
          2541 => x"70",
          2542 => x"07",
          2543 => x"8f",
          2544 => x"38",
          2545 => x"84",
          2546 => x"72",
          2547 => x"05",
          2548 => x"71",
          2549 => x"53",
          2550 => x"70",
          2551 => x"0c",
          2552 => x"71",
          2553 => x"38",
          2554 => x"90",
          2555 => x"70",
          2556 => x"0c",
          2557 => x"71",
          2558 => x"38",
          2559 => x"8e",
          2560 => x"0d",
          2561 => x"70",
          2562 => x"06",
          2563 => x"55",
          2564 => x"38",
          2565 => x"70",
          2566 => x"fb",
          2567 => x"06",
          2568 => x"82",
          2569 => x"51",
          2570 => x"54",
          2571 => x"84",
          2572 => x"70",
          2573 => x"0c",
          2574 => x"09",
          2575 => x"fd",
          2576 => x"70",
          2577 => x"81",
          2578 => x"51",
          2579 => x"70",
          2580 => x"38",
          2581 => x"70",
          2582 => x"33",
          2583 => x"70",
          2584 => x"34",
          2585 => x"74",
          2586 => x"0c",
          2587 => x"04",
          2588 => x"75",
          2589 => x"06",
          2590 => x"70",
          2591 => x"70",
          2592 => x"f7",
          2593 => x"12",
          2594 => x"84",
          2595 => x"06",
          2596 => x"53",
          2597 => x"84",
          2598 => x"70",
          2599 => x"fd",
          2600 => x"70",
          2601 => x"81",
          2602 => x"51",
          2603 => x"80",
          2604 => x"72",
          2605 => x"51",
          2606 => x"8a",
          2607 => x"70",
          2608 => x"70",
          2609 => x"74",
          2610 => x"dc",
          2611 => x"0d",
          2612 => x"0d",
          2613 => x"70",
          2614 => x"52",
          2615 => x"80",
          2616 => x"74",
          2617 => x"51",
          2618 => x"80",
          2619 => x"13",
          2620 => x"2e",
          2621 => x"33",
          2622 => x"51",
          2623 => x"09",
          2624 => x"38",
          2625 => x"81",
          2626 => x"81",
          2627 => x"70",
          2628 => x"fe",
          2629 => x"81",
          2630 => x"55",
          2631 => x"ff",
          2632 => x"06",
          2633 => x"33",
          2634 => x"51",
          2635 => x"06",
          2636 => x"06",
          2637 => x"51",
          2638 => x"82",
          2639 => x"88",
          2640 => x"71",
          2641 => x"83",
          2642 => x"38",
          2643 => x"08",
          2644 => x"74",
          2645 => x"ff",
          2646 => x"13",
          2647 => x"2e",
          2648 => x"08",
          2649 => x"fb",
          2650 => x"06",
          2651 => x"82",
          2652 => x"51",
          2653 => x"9a",
          2654 => x"84",
          2655 => x"83",
          2656 => x"38",
          2657 => x"08",
          2658 => x"74",
          2659 => x"fe",
          2660 => x"0b",
          2661 => x"0c",
          2662 => x"04",
          2663 => x"80",
          2664 => x"71",
          2665 => x"87",
          2666 => x"8c",
          2667 => x"ff",
          2668 => x"ff",
          2669 => x"72",
          2670 => x"38",
          2671 => x"dc",
          2672 => x"0d",
          2673 => x"0d",
          2674 => x"70",
          2675 => x"71",
          2676 => x"ca",
          2677 => x"51",
          2678 => x"09",
          2679 => x"38",
          2680 => x"f1",
          2681 => x"84",
          2682 => x"53",
          2683 => x"70",
          2684 => x"53",
          2685 => x"a0",
          2686 => x"81",
          2687 => x"2e",
          2688 => x"e5",
          2689 => x"ff",
          2690 => x"a0",
          2691 => x"06",
          2692 => x"73",
          2693 => x"55",
          2694 => x"0c",
          2695 => x"82",
          2696 => x"87",
          2697 => x"fc",
          2698 => x"53",
          2699 => x"2e",
          2700 => x"3d",
          2701 => x"72",
          2702 => x"3f",
          2703 => x"08",
          2704 => x"53",
          2705 => x"53",
          2706 => x"dc",
          2707 => x"0d",
          2708 => x"0d",
          2709 => x"33",
          2710 => x"53",
          2711 => x"8b",
          2712 => x"38",
          2713 => x"ff",
          2714 => x"52",
          2715 => x"81",
          2716 => x"13",
          2717 => x"52",
          2718 => x"80",
          2719 => x"13",
          2720 => x"52",
          2721 => x"80",
          2722 => x"13",
          2723 => x"52",
          2724 => x"80",
          2725 => x"13",
          2726 => x"52",
          2727 => x"26",
          2728 => x"8a",
          2729 => x"87",
          2730 => x"e7",
          2731 => x"38",
          2732 => x"c0",
          2733 => x"72",
          2734 => x"98",
          2735 => x"13",
          2736 => x"98",
          2737 => x"13",
          2738 => x"98",
          2739 => x"13",
          2740 => x"98",
          2741 => x"13",
          2742 => x"98",
          2743 => x"13",
          2744 => x"98",
          2745 => x"87",
          2746 => x"0c",
          2747 => x"98",
          2748 => x"0b",
          2749 => x"9c",
          2750 => x"71",
          2751 => x"0c",
          2752 => x"04",
          2753 => x"7f",
          2754 => x"98",
          2755 => x"7d",
          2756 => x"98",
          2757 => x"7d",
          2758 => x"c0",
          2759 => x"5a",
          2760 => x"34",
          2761 => x"b4",
          2762 => x"83",
          2763 => x"c0",
          2764 => x"5a",
          2765 => x"34",
          2766 => x"ac",
          2767 => x"85",
          2768 => x"c0",
          2769 => x"5a",
          2770 => x"34",
          2771 => x"a4",
          2772 => x"88",
          2773 => x"c0",
          2774 => x"5a",
          2775 => x"23",
          2776 => x"79",
          2777 => x"06",
          2778 => x"ff",
          2779 => x"86",
          2780 => x"85",
          2781 => x"84",
          2782 => x"83",
          2783 => x"82",
          2784 => x"7d",
          2785 => x"06",
          2786 => x"e4",
          2787 => x"3f",
          2788 => x"04",
          2789 => x"02",
          2790 => x"70",
          2791 => x"2a",
          2792 => x"70",
          2793 => x"87",
          2794 => x"3d",
          2795 => x"3d",
          2796 => x"0b",
          2797 => x"33",
          2798 => x"06",
          2799 => x"87",
          2800 => x"51",
          2801 => x"86",
          2802 => x"94",
          2803 => x"08",
          2804 => x"70",
          2805 => x"54",
          2806 => x"2e",
          2807 => x"91",
          2808 => x"06",
          2809 => x"d7",
          2810 => x"32",
          2811 => x"51",
          2812 => x"2e",
          2813 => x"93",
          2814 => x"06",
          2815 => x"ff",
          2816 => x"81",
          2817 => x"87",
          2818 => x"52",
          2819 => x"86",
          2820 => x"94",
          2821 => x"72",
          2822 => x"8c",
          2823 => x"3d",
          2824 => x"3d",
          2825 => x"05",
          2826 => x"82",
          2827 => x"70",
          2828 => x"57",
          2829 => x"c0",
          2830 => x"74",
          2831 => x"38",
          2832 => x"94",
          2833 => x"70",
          2834 => x"81",
          2835 => x"52",
          2836 => x"8c",
          2837 => x"2a",
          2838 => x"51",
          2839 => x"38",
          2840 => x"70",
          2841 => x"51",
          2842 => x"8d",
          2843 => x"2a",
          2844 => x"51",
          2845 => x"be",
          2846 => x"ff",
          2847 => x"c0",
          2848 => x"70",
          2849 => x"38",
          2850 => x"90",
          2851 => x"0c",
          2852 => x"04",
          2853 => x"79",
          2854 => x"33",
          2855 => x"06",
          2856 => x"70",
          2857 => x"fe",
          2858 => x"ff",
          2859 => x"0b",
          2860 => x"d4",
          2861 => x"ff",
          2862 => x"55",
          2863 => x"94",
          2864 => x"80",
          2865 => x"87",
          2866 => x"51",
          2867 => x"96",
          2868 => x"06",
          2869 => x"70",
          2870 => x"38",
          2871 => x"70",
          2872 => x"51",
          2873 => x"72",
          2874 => x"81",
          2875 => x"70",
          2876 => x"38",
          2877 => x"70",
          2878 => x"51",
          2879 => x"38",
          2880 => x"06",
          2881 => x"94",
          2882 => x"80",
          2883 => x"87",
          2884 => x"52",
          2885 => x"81",
          2886 => x"70",
          2887 => x"53",
          2888 => x"ff",
          2889 => x"82",
          2890 => x"89",
          2891 => x"fe",
          2892 => x"0b",
          2893 => x"33",
          2894 => x"06",
          2895 => x"c0",
          2896 => x"72",
          2897 => x"38",
          2898 => x"94",
          2899 => x"70",
          2900 => x"81",
          2901 => x"51",
          2902 => x"e2",
          2903 => x"ff",
          2904 => x"c0",
          2905 => x"70",
          2906 => x"38",
          2907 => x"90",
          2908 => x"70",
          2909 => x"82",
          2910 => x"51",
          2911 => x"04",
          2912 => x"0b",
          2913 => x"d4",
          2914 => x"ff",
          2915 => x"87",
          2916 => x"52",
          2917 => x"86",
          2918 => x"94",
          2919 => x"08",
          2920 => x"70",
          2921 => x"51",
          2922 => x"70",
          2923 => x"38",
          2924 => x"06",
          2925 => x"94",
          2926 => x"80",
          2927 => x"87",
          2928 => x"52",
          2929 => x"98",
          2930 => x"2c",
          2931 => x"71",
          2932 => x"0c",
          2933 => x"04",
          2934 => x"87",
          2935 => x"08",
          2936 => x"8a",
          2937 => x"70",
          2938 => x"b4",
          2939 => x"9e",
          2940 => x"87",
          2941 => x"c0",
          2942 => x"82",
          2943 => x"87",
          2944 => x"08",
          2945 => x"0c",
          2946 => x"98",
          2947 => x"e4",
          2948 => x"9e",
          2949 => x"87",
          2950 => x"c0",
          2951 => x"82",
          2952 => x"87",
          2953 => x"08",
          2954 => x"0c",
          2955 => x"b0",
          2956 => x"f4",
          2957 => x"9e",
          2958 => x"87",
          2959 => x"c0",
          2960 => x"82",
          2961 => x"87",
          2962 => x"08",
          2963 => x"0c",
          2964 => x"c0",
          2965 => x"84",
          2966 => x"9e",
          2967 => x"88",
          2968 => x"c0",
          2969 => x"51",
          2970 => x"8c",
          2971 => x"9e",
          2972 => x"88",
          2973 => x"c0",
          2974 => x"82",
          2975 => x"87",
          2976 => x"08",
          2977 => x"0c",
          2978 => x"88",
          2979 => x"0b",
          2980 => x"90",
          2981 => x"80",
          2982 => x"52",
          2983 => x"2e",
          2984 => x"52",
          2985 => x"9d",
          2986 => x"87",
          2987 => x"08",
          2988 => x"0a",
          2989 => x"52",
          2990 => x"83",
          2991 => x"71",
          2992 => x"34",
          2993 => x"c0",
          2994 => x"70",
          2995 => x"06",
          2996 => x"70",
          2997 => x"38",
          2998 => x"82",
          2999 => x"80",
          3000 => x"9e",
          3001 => x"88",
          3002 => x"51",
          3003 => x"80",
          3004 => x"81",
          3005 => x"88",
          3006 => x"0b",
          3007 => x"90",
          3008 => x"80",
          3009 => x"52",
          3010 => x"2e",
          3011 => x"52",
          3012 => x"a1",
          3013 => x"87",
          3014 => x"08",
          3015 => x"80",
          3016 => x"52",
          3017 => x"83",
          3018 => x"71",
          3019 => x"34",
          3020 => x"c0",
          3021 => x"70",
          3022 => x"06",
          3023 => x"70",
          3024 => x"38",
          3025 => x"82",
          3026 => x"80",
          3027 => x"9e",
          3028 => x"82",
          3029 => x"51",
          3030 => x"80",
          3031 => x"81",
          3032 => x"88",
          3033 => x"0b",
          3034 => x"90",
          3035 => x"80",
          3036 => x"52",
          3037 => x"2e",
          3038 => x"52",
          3039 => x"a5",
          3040 => x"87",
          3041 => x"08",
          3042 => x"80",
          3043 => x"52",
          3044 => x"83",
          3045 => x"71",
          3046 => x"34",
          3047 => x"c0",
          3048 => x"70",
          3049 => x"51",
          3050 => x"80",
          3051 => x"81",
          3052 => x"88",
          3053 => x"c0",
          3054 => x"70",
          3055 => x"70",
          3056 => x"51",
          3057 => x"88",
          3058 => x"0b",
          3059 => x"90",
          3060 => x"80",
          3061 => x"52",
          3062 => x"83",
          3063 => x"71",
          3064 => x"34",
          3065 => x"90",
          3066 => x"f0",
          3067 => x"2a",
          3068 => x"70",
          3069 => x"34",
          3070 => x"c0",
          3071 => x"70",
          3072 => x"52",
          3073 => x"2e",
          3074 => x"52",
          3075 => x"ab",
          3076 => x"9e",
          3077 => x"87",
          3078 => x"70",
          3079 => x"34",
          3080 => x"04",
          3081 => x"81",
          3082 => x"89",
          3083 => x"88",
          3084 => x"73",
          3085 => x"38",
          3086 => x"51",
          3087 => x"81",
          3088 => x"89",
          3089 => x"88",
          3090 => x"73",
          3091 => x"38",
          3092 => x"08",
          3093 => x"08",
          3094 => x"81",
          3095 => x"8f",
          3096 => x"88",
          3097 => x"73",
          3098 => x"38",
          3099 => x"08",
          3100 => x"08",
          3101 => x"81",
          3102 => x"8e",
          3103 => x"88",
          3104 => x"73",
          3105 => x"38",
          3106 => x"08",
          3107 => x"08",
          3108 => x"81",
          3109 => x"8e",
          3110 => x"88",
          3111 => x"73",
          3112 => x"38",
          3113 => x"08",
          3114 => x"08",
          3115 => x"81",
          3116 => x"8e",
          3117 => x"88",
          3118 => x"73",
          3119 => x"38",
          3120 => x"08",
          3121 => x"08",
          3122 => x"81",
          3123 => x"8e",
          3124 => x"88",
          3125 => x"73",
          3126 => x"38",
          3127 => x"33",
          3128 => x"c8",
          3129 => x"3f",
          3130 => x"33",
          3131 => x"2e",
          3132 => x"88",
          3133 => x"81",
          3134 => x"8d",
          3135 => x"88",
          3136 => x"73",
          3137 => x"38",
          3138 => x"33",
          3139 => x"88",
          3140 => x"3f",
          3141 => x"33",
          3142 => x"2e",
          3143 => x"f4",
          3144 => x"e5",
          3145 => x"9f",
          3146 => x"80",
          3147 => x"81",
          3148 => x"87",
          3149 => x"88",
          3150 => x"73",
          3151 => x"38",
          3152 => x"51",
          3153 => x"82",
          3154 => x"54",
          3155 => x"88",
          3156 => x"d4",
          3157 => x"3f",
          3158 => x"33",
          3159 => x"2e",
          3160 => x"f4",
          3161 => x"a1",
          3162 => x"ec",
          3163 => x"3f",
          3164 => x"08",
          3165 => x"f8",
          3166 => x"3f",
          3167 => x"08",
          3168 => x"a0",
          3169 => x"3f",
          3170 => x"08",
          3171 => x"c8",
          3172 => x"3f",
          3173 => x"51",
          3174 => x"82",
          3175 => x"52",
          3176 => x"51",
          3177 => x"82",
          3178 => x"56",
          3179 => x"52",
          3180 => x"a9",
          3181 => x"dc",
          3182 => x"c0",
          3183 => x"31",
          3184 => x"8c",
          3185 => x"81",
          3186 => x"8c",
          3187 => x"88",
          3188 => x"73",
          3189 => x"38",
          3190 => x"08",
          3191 => x"c0",
          3192 => x"e6",
          3193 => x"8c",
          3194 => x"84",
          3195 => x"71",
          3196 => x"82",
          3197 => x"52",
          3198 => x"51",
          3199 => x"82",
          3200 => x"54",
          3201 => x"a8",
          3202 => x"98",
          3203 => x"84",
          3204 => x"51",
          3205 => x"82",
          3206 => x"bd",
          3207 => x"76",
          3208 => x"54",
          3209 => x"08",
          3210 => x"f8",
          3211 => x"3f",
          3212 => x"51",
          3213 => x"87",
          3214 => x"fe",
          3215 => x"92",
          3216 => x"05",
          3217 => x"26",
          3218 => x"84",
          3219 => x"81",
          3220 => x"52",
          3221 => x"81",
          3222 => x"9d",
          3223 => x"ac",
          3224 => x"81",
          3225 => x"91",
          3226 => x"bc",
          3227 => x"81",
          3228 => x"85",
          3229 => x"c8",
          3230 => x"3f",
          3231 => x"04",
          3232 => x"0c",
          3233 => x"87",
          3234 => x"0c",
          3235 => x"b0",
          3236 => x"96",
          3237 => x"fe",
          3238 => x"8c",
          3239 => x"38",
          3240 => x"0b",
          3241 => x"0c",
          3242 => x"08",
          3243 => x"52",
          3244 => x"83",
          3245 => x"88",
          3246 => x"8c",
          3247 => x"53",
          3248 => x"dc",
          3249 => x"0d",
          3250 => x"0d",
          3251 => x"12",
          3252 => x"90",
          3253 => x"15",
          3254 => x"5e",
          3255 => x"59",
          3256 => x"77",
          3257 => x"75",
          3258 => x"08",
          3259 => x"71",
          3260 => x"31",
          3261 => x"80",
          3262 => x"84",
          3263 => x"8c",
          3264 => x"88",
          3265 => x"8c",
          3266 => x"88",
          3267 => x"90",
          3268 => x"94",
          3269 => x"94",
          3270 => x"90",
          3271 => x"39",
          3272 => x"73",
          3273 => x"74",
          3274 => x"77",
          3275 => x"0c",
          3276 => x"04",
          3277 => x"76",
          3278 => x"88",
          3279 => x"53",
          3280 => x"81",
          3281 => x"06",
          3282 => x"12",
          3283 => x"52",
          3284 => x"2e",
          3285 => x"94",
          3286 => x"08",
          3287 => x"0c",
          3288 => x"0c",
          3289 => x"0c",
          3290 => x"39",
          3291 => x"82",
          3292 => x"90",
          3293 => x"88",
          3294 => x"14",
          3295 => x"88",
          3296 => x"13",
          3297 => x"12",
          3298 => x"08",
          3299 => x"81",
          3300 => x"84",
          3301 => x"14",
          3302 => x"74",
          3303 => x"06",
          3304 => x"14",
          3305 => x"14",
          3306 => x"08",
          3307 => x"70",
          3308 => x"52",
          3309 => x"8c",
          3310 => x"15",
          3311 => x"13",
          3312 => x"12",
          3313 => x"8c",
          3314 => x"3d",
          3315 => x"3d",
          3316 => x"55",
          3317 => x"2e",
          3318 => x"9f",
          3319 => x"82",
          3320 => x"57",
          3321 => x"82",
          3322 => x"84",
          3323 => x"27",
          3324 => x"90",
          3325 => x"ed",
          3326 => x"ff",
          3327 => x"80",
          3328 => x"58",
          3329 => x"82",
          3330 => x"82",
          3331 => x"30",
          3332 => x"dc",
          3333 => x"25",
          3334 => x"08",
          3335 => x"70",
          3336 => x"25",
          3337 => x"58",
          3338 => x"56",
          3339 => x"74",
          3340 => x"06",
          3341 => x"88",
          3342 => x"75",
          3343 => x"39",
          3344 => x"8c",
          3345 => x"77",
          3346 => x"08",
          3347 => x"82",
          3348 => x"53",
          3349 => x"2e",
          3350 => x"73",
          3351 => x"8c",
          3352 => x"f0",
          3353 => x"08",
          3354 => x"72",
          3355 => x"75",
          3356 => x"88",
          3357 => x"8c",
          3358 => x"75",
          3359 => x"3f",
          3360 => x"8c",
          3361 => x"fc",
          3362 => x"8c",
          3363 => x"73",
          3364 => x"0c",
          3365 => x"04",
          3366 => x"73",
          3367 => x"2e",
          3368 => x"12",
          3369 => x"3f",
          3370 => x"04",
          3371 => x"02",
          3372 => x"53",
          3373 => x"09",
          3374 => x"38",
          3375 => x"3f",
          3376 => x"08",
          3377 => x"2e",
          3378 => x"72",
          3379 => x"f8",
          3380 => x"82",
          3381 => x"8f",
          3382 => x"f0",
          3383 => x"80",
          3384 => x"72",
          3385 => x"84",
          3386 => x"fe",
          3387 => x"97",
          3388 => x"8c",
          3389 => x"82",
          3390 => x"54",
          3391 => x"3f",
          3392 => x"f0",
          3393 => x"0d",
          3394 => x"0d",
          3395 => x"33",
          3396 => x"06",
          3397 => x"80",
          3398 => x"72",
          3399 => x"51",
          3400 => x"ff",
          3401 => x"39",
          3402 => x"04",
          3403 => x"77",
          3404 => x"08",
          3405 => x"f0",
          3406 => x"73",
          3407 => x"ff",
          3408 => x"71",
          3409 => x"38",
          3410 => x"06",
          3411 => x"54",
          3412 => x"e7",
          3413 => x"8c",
          3414 => x"3d",
          3415 => x"3d",
          3416 => x"59",
          3417 => x"81",
          3418 => x"56",
          3419 => x"84",
          3420 => x"a5",
          3421 => x"06",
          3422 => x"80",
          3423 => x"81",
          3424 => x"58",
          3425 => x"b0",
          3426 => x"06",
          3427 => x"5a",
          3428 => x"ad",
          3429 => x"06",
          3430 => x"5a",
          3431 => x"05",
          3432 => x"75",
          3433 => x"81",
          3434 => x"77",
          3435 => x"08",
          3436 => x"05",
          3437 => x"5d",
          3438 => x"39",
          3439 => x"72",
          3440 => x"38",
          3441 => x"7b",
          3442 => x"05",
          3443 => x"70",
          3444 => x"33",
          3445 => x"39",
          3446 => x"32",
          3447 => x"72",
          3448 => x"78",
          3449 => x"70",
          3450 => x"07",
          3451 => x"07",
          3452 => x"51",
          3453 => x"80",
          3454 => x"79",
          3455 => x"70",
          3456 => x"33",
          3457 => x"80",
          3458 => x"38",
          3459 => x"e0",
          3460 => x"38",
          3461 => x"81",
          3462 => x"53",
          3463 => x"2e",
          3464 => x"73",
          3465 => x"a2",
          3466 => x"c3",
          3467 => x"38",
          3468 => x"24",
          3469 => x"80",
          3470 => x"8c",
          3471 => x"39",
          3472 => x"2e",
          3473 => x"81",
          3474 => x"80",
          3475 => x"80",
          3476 => x"d5",
          3477 => x"73",
          3478 => x"8e",
          3479 => x"39",
          3480 => x"2e",
          3481 => x"80",
          3482 => x"84",
          3483 => x"56",
          3484 => x"74",
          3485 => x"72",
          3486 => x"38",
          3487 => x"15",
          3488 => x"54",
          3489 => x"38",
          3490 => x"56",
          3491 => x"81",
          3492 => x"72",
          3493 => x"38",
          3494 => x"90",
          3495 => x"06",
          3496 => x"2e",
          3497 => x"51",
          3498 => x"74",
          3499 => x"53",
          3500 => x"fd",
          3501 => x"51",
          3502 => x"ef",
          3503 => x"19",
          3504 => x"53",
          3505 => x"39",
          3506 => x"39",
          3507 => x"39",
          3508 => x"39",
          3509 => x"39",
          3510 => x"d0",
          3511 => x"39",
          3512 => x"70",
          3513 => x"53",
          3514 => x"88",
          3515 => x"19",
          3516 => x"39",
          3517 => x"54",
          3518 => x"74",
          3519 => x"70",
          3520 => x"07",
          3521 => x"55",
          3522 => x"80",
          3523 => x"72",
          3524 => x"38",
          3525 => x"90",
          3526 => x"80",
          3527 => x"5e",
          3528 => x"74",
          3529 => x"3f",
          3530 => x"08",
          3531 => x"7c",
          3532 => x"54",
          3533 => x"82",
          3534 => x"55",
          3535 => x"92",
          3536 => x"53",
          3537 => x"2e",
          3538 => x"14",
          3539 => x"ff",
          3540 => x"14",
          3541 => x"70",
          3542 => x"34",
          3543 => x"30",
          3544 => x"9f",
          3545 => x"57",
          3546 => x"85",
          3547 => x"b1",
          3548 => x"2a",
          3549 => x"51",
          3550 => x"2e",
          3551 => x"3d",
          3552 => x"05",
          3553 => x"34",
          3554 => x"76",
          3555 => x"54",
          3556 => x"72",
          3557 => x"54",
          3558 => x"70",
          3559 => x"56",
          3560 => x"81",
          3561 => x"7b",
          3562 => x"73",
          3563 => x"3f",
          3564 => x"53",
          3565 => x"74",
          3566 => x"53",
          3567 => x"eb",
          3568 => x"77",
          3569 => x"53",
          3570 => x"14",
          3571 => x"54",
          3572 => x"3f",
          3573 => x"74",
          3574 => x"53",
          3575 => x"fb",
          3576 => x"51",
          3577 => x"ef",
          3578 => x"0d",
          3579 => x"0d",
          3580 => x"70",
          3581 => x"08",
          3582 => x"51",
          3583 => x"85",
          3584 => x"fe",
          3585 => x"82",
          3586 => x"85",
          3587 => x"52",
          3588 => x"ca",
          3589 => x"f8",
          3590 => x"73",
          3591 => x"82",
          3592 => x"84",
          3593 => x"fd",
          3594 => x"8c",
          3595 => x"82",
          3596 => x"87",
          3597 => x"53",
          3598 => x"fa",
          3599 => x"82",
          3600 => x"85",
          3601 => x"fb",
          3602 => x"79",
          3603 => x"08",
          3604 => x"57",
          3605 => x"71",
          3606 => x"e0",
          3607 => x"f4",
          3608 => x"2d",
          3609 => x"08",
          3610 => x"53",
          3611 => x"80",
          3612 => x"8d",
          3613 => x"72",
          3614 => x"30",
          3615 => x"51",
          3616 => x"80",
          3617 => x"71",
          3618 => x"38",
          3619 => x"97",
          3620 => x"25",
          3621 => x"16",
          3622 => x"25",
          3623 => x"14",
          3624 => x"34",
          3625 => x"72",
          3626 => x"3f",
          3627 => x"73",
          3628 => x"72",
          3629 => x"f7",
          3630 => x"53",
          3631 => x"dc",
          3632 => x"0d",
          3633 => x"0d",
          3634 => x"08",
          3635 => x"f4",
          3636 => x"76",
          3637 => x"ef",
          3638 => x"8c",
          3639 => x"3d",
          3640 => x"3d",
          3641 => x"5a",
          3642 => x"7a",
          3643 => x"08",
          3644 => x"53",
          3645 => x"09",
          3646 => x"38",
          3647 => x"0c",
          3648 => x"ad",
          3649 => x"06",
          3650 => x"76",
          3651 => x"0c",
          3652 => x"33",
          3653 => x"73",
          3654 => x"81",
          3655 => x"38",
          3656 => x"05",
          3657 => x"08",
          3658 => x"53",
          3659 => x"2e",
          3660 => x"57",
          3661 => x"2e",
          3662 => x"39",
          3663 => x"13",
          3664 => x"08",
          3665 => x"53",
          3666 => x"55",
          3667 => x"80",
          3668 => x"14",
          3669 => x"88",
          3670 => x"27",
          3671 => x"eb",
          3672 => x"53",
          3673 => x"89",
          3674 => x"38",
          3675 => x"55",
          3676 => x"8a",
          3677 => x"a0",
          3678 => x"c2",
          3679 => x"74",
          3680 => x"e0",
          3681 => x"ff",
          3682 => x"d0",
          3683 => x"ff",
          3684 => x"90",
          3685 => x"38",
          3686 => x"81",
          3687 => x"53",
          3688 => x"ca",
          3689 => x"27",
          3690 => x"77",
          3691 => x"08",
          3692 => x"0c",
          3693 => x"33",
          3694 => x"ff",
          3695 => x"80",
          3696 => x"74",
          3697 => x"79",
          3698 => x"74",
          3699 => x"0c",
          3700 => x"04",
          3701 => x"7a",
          3702 => x"80",
          3703 => x"58",
          3704 => x"33",
          3705 => x"a0",
          3706 => x"06",
          3707 => x"13",
          3708 => x"39",
          3709 => x"09",
          3710 => x"38",
          3711 => x"11",
          3712 => x"08",
          3713 => x"54",
          3714 => x"2e",
          3715 => x"80",
          3716 => x"08",
          3717 => x"0c",
          3718 => x"33",
          3719 => x"80",
          3720 => x"38",
          3721 => x"80",
          3722 => x"38",
          3723 => x"57",
          3724 => x"0c",
          3725 => x"33",
          3726 => x"39",
          3727 => x"74",
          3728 => x"38",
          3729 => x"80",
          3730 => x"89",
          3731 => x"38",
          3732 => x"d0",
          3733 => x"55",
          3734 => x"80",
          3735 => x"39",
          3736 => x"d9",
          3737 => x"80",
          3738 => x"27",
          3739 => x"80",
          3740 => x"89",
          3741 => x"70",
          3742 => x"55",
          3743 => x"70",
          3744 => x"55",
          3745 => x"27",
          3746 => x"14",
          3747 => x"06",
          3748 => x"74",
          3749 => x"73",
          3750 => x"38",
          3751 => x"14",
          3752 => x"05",
          3753 => x"08",
          3754 => x"54",
          3755 => x"39",
          3756 => x"84",
          3757 => x"55",
          3758 => x"81",
          3759 => x"8c",
          3760 => x"3d",
          3761 => x"3d",
          3762 => x"2b",
          3763 => x"79",
          3764 => x"98",
          3765 => x"13",
          3766 => x"51",
          3767 => x"51",
          3768 => x"81",
          3769 => x"33",
          3770 => x"74",
          3771 => x"81",
          3772 => x"08",
          3773 => x"05",
          3774 => x"71",
          3775 => x"52",
          3776 => x"09",
          3777 => x"38",
          3778 => x"82",
          3779 => x"85",
          3780 => x"fc",
          3781 => x"02",
          3782 => x"05",
          3783 => x"54",
          3784 => x"80",
          3785 => x"88",
          3786 => x"3f",
          3787 => x"fc",
          3788 => x"f2",
          3789 => x"33",
          3790 => x"71",
          3791 => x"81",
          3792 => x"de",
          3793 => x"f3",
          3794 => x"73",
          3795 => x"0d",
          3796 => x"0d",
          3797 => x"05",
          3798 => x"02",
          3799 => x"05",
          3800 => x"a8",
          3801 => x"29",
          3802 => x"05",
          3803 => x"59",
          3804 => x"59",
          3805 => x"86",
          3806 => x"f2",
          3807 => x"89",
          3808 => x"84",
          3809 => x"d0",
          3810 => x"70",
          3811 => x"5a",
          3812 => x"82",
          3813 => x"75",
          3814 => x"a8",
          3815 => x"29",
          3816 => x"05",
          3817 => x"56",
          3818 => x"2e",
          3819 => x"53",
          3820 => x"51",
          3821 => x"82",
          3822 => x"81",
          3823 => x"82",
          3824 => x"74",
          3825 => x"55",
          3826 => x"87",
          3827 => x"82",
          3828 => x"77",
          3829 => x"38",
          3830 => x"08",
          3831 => x"2e",
          3832 => x"89",
          3833 => x"74",
          3834 => x"3d",
          3835 => x"76",
          3836 => x"75",
          3837 => x"91",
          3838 => x"a4",
          3839 => x"51",
          3840 => x"3f",
          3841 => x"08",
          3842 => x"ee",
          3843 => x"0d",
          3844 => x"0d",
          3845 => x"52",
          3846 => x"08",
          3847 => x"87",
          3848 => x"dc",
          3849 => x"38",
          3850 => x"08",
          3851 => x"52",
          3852 => x"52",
          3853 => x"d5",
          3854 => x"dc",
          3855 => x"b8",
          3856 => x"d8",
          3857 => x"8c",
          3858 => x"80",
          3859 => x"dc",
          3860 => x"38",
          3861 => x"08",
          3862 => x"17",
          3863 => x"74",
          3864 => x"76",
          3865 => x"81",
          3866 => x"57",
          3867 => x"74",
          3868 => x"81",
          3869 => x"38",
          3870 => x"04",
          3871 => x"aa",
          3872 => x"3d",
          3873 => x"81",
          3874 => x"80",
          3875 => x"a4",
          3876 => x"d1",
          3877 => x"8c",
          3878 => x"91",
          3879 => x"82",
          3880 => x"54",
          3881 => x"52",
          3882 => x"52",
          3883 => x"dd",
          3884 => x"dc",
          3885 => x"a4",
          3886 => x"d7",
          3887 => x"8c",
          3888 => x"18",
          3889 => x"0b",
          3890 => x"08",
          3891 => x"82",
          3892 => x"ff",
          3893 => x"55",
          3894 => x"34",
          3895 => x"30",
          3896 => x"9f",
          3897 => x"55",
          3898 => x"85",
          3899 => x"ad",
          3900 => x"a4",
          3901 => x"08",
          3902 => x"d0",
          3903 => x"8c",
          3904 => x"2e",
          3905 => x"f7",
          3906 => x"fd",
          3907 => x"2e",
          3908 => x"99",
          3909 => x"79",
          3910 => x"3f",
          3911 => x"d0",
          3912 => x"08",
          3913 => x"dc",
          3914 => x"80",
          3915 => x"8c",
          3916 => x"3d",
          3917 => x"3d",
          3918 => x"71",
          3919 => x"33",
          3920 => x"58",
          3921 => x"09",
          3922 => x"38",
          3923 => x"05",
          3924 => x"27",
          3925 => x"17",
          3926 => x"71",
          3927 => x"55",
          3928 => x"09",
          3929 => x"38",
          3930 => x"ea",
          3931 => x"73",
          3932 => x"89",
          3933 => x"08",
          3934 => x"f4",
          3935 => x"dc",
          3936 => x"52",
          3937 => x"d6",
          3938 => x"8c",
          3939 => x"c4",
          3940 => x"33",
          3941 => x"2e",
          3942 => x"82",
          3943 => x"b4",
          3944 => x"3f",
          3945 => x"1a",
          3946 => x"fc",
          3947 => x"05",
          3948 => x"3f",
          3949 => x"08",
          3950 => x"38",
          3951 => x"52",
          3952 => x"b8",
          3953 => x"dc",
          3954 => x"06",
          3955 => x"38",
          3956 => x"39",
          3957 => x"81",
          3958 => x"54",
          3959 => x"ff",
          3960 => x"54",
          3961 => x"dc",
          3962 => x"0d",
          3963 => x"0d",
          3964 => x"02",
          3965 => x"c3",
          3966 => x"5a",
          3967 => x"3d",
          3968 => x"a8",
          3969 => x"89",
          3970 => x"a3",
          3971 => x"a0",
          3972 => x"81",
          3973 => x"51",
          3974 => x"82",
          3975 => x"82",
          3976 => x"82",
          3977 => x"80",
          3978 => x"38",
          3979 => x"88",
          3980 => x"82",
          3981 => x"51",
          3982 => x"82",
          3983 => x"80",
          3984 => x"81",
          3985 => x"f3",
          3986 => x"e3",
          3987 => x"a4",
          3988 => x"f8",
          3989 => x"70",
          3990 => x"f6",
          3991 => x"8c",
          3992 => x"82",
          3993 => x"74",
          3994 => x"06",
          3995 => x"82",
          3996 => x"51",
          3997 => x"82",
          3998 => x"55",
          3999 => x"8c",
          4000 => x"9a",
          4001 => x"dc",
          4002 => x"70",
          4003 => x"80",
          4004 => x"53",
          4005 => x"06",
          4006 => x"f9",
          4007 => x"ff",
          4008 => x"06",
          4009 => x"87",
          4010 => x"82",
          4011 => x"8f",
          4012 => x"cc",
          4013 => x"dc",
          4014 => x"70",
          4015 => x"59",
          4016 => x"ee",
          4017 => x"ff",
          4018 => x"80",
          4019 => x"2b",
          4020 => x"82",
          4021 => x"70",
          4022 => x"97",
          4023 => x"2c",
          4024 => x"29",
          4025 => x"05",
          4026 => x"70",
          4027 => x"51",
          4028 => x"51",
          4029 => x"81",
          4030 => x"2e",
          4031 => x"77",
          4032 => x"38",
          4033 => x"0a",
          4034 => x"0a",
          4035 => x"2c",
          4036 => x"75",
          4037 => x"38",
          4038 => x"52",
          4039 => x"a6",
          4040 => x"dc",
          4041 => x"06",
          4042 => x"2e",
          4043 => x"82",
          4044 => x"81",
          4045 => x"74",
          4046 => x"29",
          4047 => x"05",
          4048 => x"70",
          4049 => x"56",
          4050 => x"8a",
          4051 => x"76",
          4052 => x"77",
          4053 => x"3f",
          4054 => x"08",
          4055 => x"54",
          4056 => x"d3",
          4057 => x"75",
          4058 => x"ca",
          4059 => x"55",
          4060 => x"80",
          4061 => x"2b",
          4062 => x"82",
          4063 => x"70",
          4064 => x"98",
          4065 => x"11",
          4066 => x"81",
          4067 => x"33",
          4068 => x"51",
          4069 => x"55",
          4070 => x"09",
          4071 => x"92",
          4072 => x"e0",
          4073 => x"0c",
          4074 => x"8d",
          4075 => x"0b",
          4076 => x"34",
          4077 => x"82",
          4078 => x"75",
          4079 => x"34",
          4080 => x"34",
          4081 => x"7e",
          4082 => x"26",
          4083 => x"73",
          4084 => x"f0",
          4085 => x"73",
          4086 => x"8d",
          4087 => x"73",
          4088 => x"cb",
          4089 => x"84",
          4090 => x"75",
          4091 => x"74",
          4092 => x"98",
          4093 => x"73",
          4094 => x"38",
          4095 => x"73",
          4096 => x"34",
          4097 => x"0a",
          4098 => x"0a",
          4099 => x"2c",
          4100 => x"33",
          4101 => x"df",
          4102 => x"88",
          4103 => x"56",
          4104 => x"8d",
          4105 => x"1a",
          4106 => x"33",
          4107 => x"8d",
          4108 => x"73",
          4109 => x"38",
          4110 => x"73",
          4111 => x"34",
          4112 => x"33",
          4113 => x"0a",
          4114 => x"0a",
          4115 => x"2c",
          4116 => x"33",
          4117 => x"56",
          4118 => x"a2",
          4119 => x"70",
          4120 => x"e8",
          4121 => x"81",
          4122 => x"81",
          4123 => x"70",
          4124 => x"8d",
          4125 => x"51",
          4126 => x"24",
          4127 => x"8d",
          4128 => x"98",
          4129 => x"2c",
          4130 => x"33",
          4131 => x"56",
          4132 => x"fc",
          4133 => x"51",
          4134 => x"74",
          4135 => x"29",
          4136 => x"05",
          4137 => x"82",
          4138 => x"56",
          4139 => x"75",
          4140 => x"fb",
          4141 => x"8d",
          4142 => x"81",
          4143 => x"55",
          4144 => x"fb",
          4145 => x"8d",
          4146 => x"05",
          4147 => x"8d",
          4148 => x"15",
          4149 => x"8d",
          4150 => x"51",
          4151 => x"82",
          4152 => x"70",
          4153 => x"98",
          4154 => x"84",
          4155 => x"56",
          4156 => x"25",
          4157 => x"1a",
          4158 => x"33",
          4159 => x"33",
          4160 => x"3f",
          4161 => x"0a",
          4162 => x"0a",
          4163 => x"2c",
          4164 => x"33",
          4165 => x"75",
          4166 => x"38",
          4167 => x"8c",
          4168 => x"88",
          4169 => x"2b",
          4170 => x"82",
          4171 => x"57",
          4172 => x"74",
          4173 => x"f7",
          4174 => x"e6",
          4175 => x"81",
          4176 => x"81",
          4177 => x"70",
          4178 => x"8d",
          4179 => x"51",
          4180 => x"25",
          4181 => x"d7",
          4182 => x"84",
          4183 => x"54",
          4184 => x"8a",
          4185 => x"3f",
          4186 => x"52",
          4187 => x"c6",
          4188 => x"dc",
          4189 => x"06",
          4190 => x"38",
          4191 => x"33",
          4192 => x"2e",
          4193 => x"81",
          4194 => x"79",
          4195 => x"3f",
          4196 => x"80",
          4197 => x"b7",
          4198 => x"88",
          4199 => x"80",
          4200 => x"38",
          4201 => x"84",
          4202 => x"88",
          4203 => x"54",
          4204 => x"88",
          4205 => x"ff",
          4206 => x"39",
          4207 => x"33",
          4208 => x"33",
          4209 => x"75",
          4210 => x"38",
          4211 => x"73",
          4212 => x"34",
          4213 => x"70",
          4214 => x"81",
          4215 => x"51",
          4216 => x"25",
          4217 => x"1a",
          4218 => x"33",
          4219 => x"33",
          4220 => x"3f",
          4221 => x"0a",
          4222 => x"0a",
          4223 => x"2c",
          4224 => x"33",
          4225 => x"75",
          4226 => x"38",
          4227 => x"9c",
          4228 => x"88",
          4229 => x"2b",
          4230 => x"82",
          4231 => x"57",
          4232 => x"74",
          4233 => x"87",
          4234 => x"e4",
          4235 => x"81",
          4236 => x"81",
          4237 => x"70",
          4238 => x"8d",
          4239 => x"51",
          4240 => x"25",
          4241 => x"e7",
          4242 => x"88",
          4243 => x"ff",
          4244 => x"84",
          4245 => x"54",
          4246 => x"f8",
          4247 => x"14",
          4248 => x"8d",
          4249 => x"1a",
          4250 => x"54",
          4251 => x"82",
          4252 => x"70",
          4253 => x"82",
          4254 => x"58",
          4255 => x"75",
          4256 => x"f8",
          4257 => x"ae",
          4258 => x"9c",
          4259 => x"80",
          4260 => x"74",
          4261 => x"3f",
          4262 => x"08",
          4263 => x"34",
          4264 => x"08",
          4265 => x"81",
          4266 => x"52",
          4267 => x"a5",
          4268 => x"81",
          4269 => x"84",
          4270 => x"d0",
          4271 => x"08",
          4272 => x"80",
          4273 => x"74",
          4274 => x"3f",
          4275 => x"08",
          4276 => x"34",
          4277 => x"08",
          4278 => x"81",
          4279 => x"52",
          4280 => x"f1",
          4281 => x"54",
          4282 => x"73",
          4283 => x"80",
          4284 => x"38",
          4285 => x"f8",
          4286 => x"39",
          4287 => x"09",
          4288 => x"38",
          4289 => x"08",
          4290 => x"2e",
          4291 => x"51",
          4292 => x"80",
          4293 => x"84",
          4294 => x"d0",
          4295 => x"08",
          4296 => x"80",
          4297 => x"74",
          4298 => x"3f",
          4299 => x"08",
          4300 => x"34",
          4301 => x"08",
          4302 => x"81",
          4303 => x"52",
          4304 => x"91",
          4305 => x"54",
          4306 => x"06",
          4307 => x"73",
          4308 => x"80",
          4309 => x"38",
          4310 => x"94",
          4311 => x"dc",
          4312 => x"84",
          4313 => x"dc",
          4314 => x"06",
          4315 => x"74",
          4316 => x"c6",
          4317 => x"8d",
          4318 => x"8d",
          4319 => x"79",
          4320 => x"3f",
          4321 => x"82",
          4322 => x"70",
          4323 => x"82",
          4324 => x"59",
          4325 => x"77",
          4326 => x"38",
          4327 => x"73",
          4328 => x"34",
          4329 => x"33",
          4330 => x"80",
          4331 => x"39",
          4332 => x"33",
          4333 => x"2e",
          4334 => x"88",
          4335 => x"3f",
          4336 => x"33",
          4337 => x"73",
          4338 => x"34",
          4339 => x"80",
          4340 => x"88",
          4341 => x"82",
          4342 => x"79",
          4343 => x"0c",
          4344 => x"04",
          4345 => x"02",
          4346 => x"51",
          4347 => x"72",
          4348 => x"82",
          4349 => x"33",
          4350 => x"8c",
          4351 => x"3d",
          4352 => x"3d",
          4353 => x"05",
          4354 => x"05",
          4355 => x"56",
          4356 => x"72",
          4357 => x"e0",
          4358 => x"2b",
          4359 => x"8c",
          4360 => x"88",
          4361 => x"2e",
          4362 => x"88",
          4363 => x"0c",
          4364 => x"8c",
          4365 => x"71",
          4366 => x"87",
          4367 => x"0c",
          4368 => x"08",
          4369 => x"51",
          4370 => x"2e",
          4371 => x"c0",
          4372 => x"51",
          4373 => x"71",
          4374 => x"80",
          4375 => x"92",
          4376 => x"98",
          4377 => x"70",
          4378 => x"38",
          4379 => x"c4",
          4380 => x"89",
          4381 => x"51",
          4382 => x"dc",
          4383 => x"0d",
          4384 => x"0d",
          4385 => x"02",
          4386 => x"05",
          4387 => x"58",
          4388 => x"52",
          4389 => x"3f",
          4390 => x"08",
          4391 => x"54",
          4392 => x"be",
          4393 => x"75",
          4394 => x"c0",
          4395 => x"87",
          4396 => x"12",
          4397 => x"84",
          4398 => x"40",
          4399 => x"85",
          4400 => x"98",
          4401 => x"7d",
          4402 => x"0c",
          4403 => x"85",
          4404 => x"06",
          4405 => x"71",
          4406 => x"38",
          4407 => x"71",
          4408 => x"05",
          4409 => x"19",
          4410 => x"a2",
          4411 => x"71",
          4412 => x"38",
          4413 => x"83",
          4414 => x"38",
          4415 => x"8a",
          4416 => x"98",
          4417 => x"71",
          4418 => x"c0",
          4419 => x"52",
          4420 => x"87",
          4421 => x"80",
          4422 => x"81",
          4423 => x"c0",
          4424 => x"53",
          4425 => x"82",
          4426 => x"71",
          4427 => x"1a",
          4428 => x"84",
          4429 => x"19",
          4430 => x"06",
          4431 => x"79",
          4432 => x"38",
          4433 => x"80",
          4434 => x"87",
          4435 => x"26",
          4436 => x"73",
          4437 => x"06",
          4438 => x"2e",
          4439 => x"52",
          4440 => x"82",
          4441 => x"8f",
          4442 => x"f3",
          4443 => x"62",
          4444 => x"05",
          4445 => x"57",
          4446 => x"83",
          4447 => x"52",
          4448 => x"3f",
          4449 => x"08",
          4450 => x"54",
          4451 => x"2e",
          4452 => x"81",
          4453 => x"74",
          4454 => x"c0",
          4455 => x"87",
          4456 => x"12",
          4457 => x"84",
          4458 => x"5f",
          4459 => x"0b",
          4460 => x"8c",
          4461 => x"0c",
          4462 => x"80",
          4463 => x"70",
          4464 => x"81",
          4465 => x"54",
          4466 => x"8c",
          4467 => x"81",
          4468 => x"7c",
          4469 => x"58",
          4470 => x"70",
          4471 => x"52",
          4472 => x"8a",
          4473 => x"98",
          4474 => x"71",
          4475 => x"c0",
          4476 => x"52",
          4477 => x"87",
          4478 => x"80",
          4479 => x"81",
          4480 => x"c0",
          4481 => x"53",
          4482 => x"82",
          4483 => x"71",
          4484 => x"19",
          4485 => x"81",
          4486 => x"ff",
          4487 => x"19",
          4488 => x"78",
          4489 => x"38",
          4490 => x"80",
          4491 => x"87",
          4492 => x"26",
          4493 => x"73",
          4494 => x"06",
          4495 => x"2e",
          4496 => x"52",
          4497 => x"82",
          4498 => x"8f",
          4499 => x"fa",
          4500 => x"02",
          4501 => x"05",
          4502 => x"05",
          4503 => x"71",
          4504 => x"57",
          4505 => x"82",
          4506 => x"81",
          4507 => x"54",
          4508 => x"38",
          4509 => x"c0",
          4510 => x"81",
          4511 => x"2e",
          4512 => x"71",
          4513 => x"38",
          4514 => x"87",
          4515 => x"11",
          4516 => x"80",
          4517 => x"80",
          4518 => x"83",
          4519 => x"38",
          4520 => x"72",
          4521 => x"2a",
          4522 => x"51",
          4523 => x"80",
          4524 => x"87",
          4525 => x"08",
          4526 => x"38",
          4527 => x"8c",
          4528 => x"96",
          4529 => x"0c",
          4530 => x"8c",
          4531 => x"08",
          4532 => x"51",
          4533 => x"38",
          4534 => x"56",
          4535 => x"80",
          4536 => x"85",
          4537 => x"77",
          4538 => x"83",
          4539 => x"75",
          4540 => x"8c",
          4541 => x"3d",
          4542 => x"3d",
          4543 => x"11",
          4544 => x"71",
          4545 => x"82",
          4546 => x"53",
          4547 => x"0d",
          4548 => x"0d",
          4549 => x"33",
          4550 => x"71",
          4551 => x"88",
          4552 => x"14",
          4553 => x"07",
          4554 => x"33",
          4555 => x"8c",
          4556 => x"53",
          4557 => x"52",
          4558 => x"04",
          4559 => x"73",
          4560 => x"92",
          4561 => x"52",
          4562 => x"81",
          4563 => x"70",
          4564 => x"70",
          4565 => x"3d",
          4566 => x"3d",
          4567 => x"52",
          4568 => x"70",
          4569 => x"34",
          4570 => x"51",
          4571 => x"81",
          4572 => x"70",
          4573 => x"70",
          4574 => x"05",
          4575 => x"88",
          4576 => x"72",
          4577 => x"0d",
          4578 => x"0d",
          4579 => x"54",
          4580 => x"80",
          4581 => x"71",
          4582 => x"53",
          4583 => x"81",
          4584 => x"ff",
          4585 => x"39",
          4586 => x"04",
          4587 => x"75",
          4588 => x"52",
          4589 => x"70",
          4590 => x"34",
          4591 => x"70",
          4592 => x"3d",
          4593 => x"3d",
          4594 => x"79",
          4595 => x"74",
          4596 => x"56",
          4597 => x"81",
          4598 => x"71",
          4599 => x"16",
          4600 => x"52",
          4601 => x"86",
          4602 => x"2e",
          4603 => x"82",
          4604 => x"86",
          4605 => x"fe",
          4606 => x"76",
          4607 => x"39",
          4608 => x"8a",
          4609 => x"51",
          4610 => x"71",
          4611 => x"33",
          4612 => x"0c",
          4613 => x"04",
          4614 => x"8c",
          4615 => x"80",
          4616 => x"dc",
          4617 => x"3d",
          4618 => x"80",
          4619 => x"33",
          4620 => x"7a",
          4621 => x"38",
          4622 => x"16",
          4623 => x"16",
          4624 => x"17",
          4625 => x"fa",
          4626 => x"8c",
          4627 => x"2e",
          4628 => x"b7",
          4629 => x"dc",
          4630 => x"34",
          4631 => x"70",
          4632 => x"31",
          4633 => x"59",
          4634 => x"77",
          4635 => x"82",
          4636 => x"74",
          4637 => x"81",
          4638 => x"81",
          4639 => x"53",
          4640 => x"16",
          4641 => x"e3",
          4642 => x"81",
          4643 => x"8c",
          4644 => x"3d",
          4645 => x"3d",
          4646 => x"56",
          4647 => x"74",
          4648 => x"2e",
          4649 => x"51",
          4650 => x"82",
          4651 => x"57",
          4652 => x"08",
          4653 => x"54",
          4654 => x"16",
          4655 => x"33",
          4656 => x"3f",
          4657 => x"08",
          4658 => x"38",
          4659 => x"57",
          4660 => x"0c",
          4661 => x"dc",
          4662 => x"0d",
          4663 => x"0d",
          4664 => x"57",
          4665 => x"82",
          4666 => x"58",
          4667 => x"08",
          4668 => x"76",
          4669 => x"83",
          4670 => x"06",
          4671 => x"84",
          4672 => x"78",
          4673 => x"81",
          4674 => x"38",
          4675 => x"82",
          4676 => x"52",
          4677 => x"52",
          4678 => x"3f",
          4679 => x"52",
          4680 => x"51",
          4681 => x"84",
          4682 => x"d2",
          4683 => x"fc",
          4684 => x"8a",
          4685 => x"52",
          4686 => x"51",
          4687 => x"90",
          4688 => x"84",
          4689 => x"fc",
          4690 => x"17",
          4691 => x"a0",
          4692 => x"86",
          4693 => x"08",
          4694 => x"b0",
          4695 => x"55",
          4696 => x"81",
          4697 => x"f8",
          4698 => x"84",
          4699 => x"53",
          4700 => x"17",
          4701 => x"d7",
          4702 => x"dc",
          4703 => x"83",
          4704 => x"77",
          4705 => x"0c",
          4706 => x"04",
          4707 => x"77",
          4708 => x"12",
          4709 => x"55",
          4710 => x"56",
          4711 => x"8d",
          4712 => x"22",
          4713 => x"ac",
          4714 => x"57",
          4715 => x"8c",
          4716 => x"3d",
          4717 => x"3d",
          4718 => x"70",
          4719 => x"57",
          4720 => x"81",
          4721 => x"98",
          4722 => x"81",
          4723 => x"74",
          4724 => x"72",
          4725 => x"f5",
          4726 => x"24",
          4727 => x"81",
          4728 => x"81",
          4729 => x"83",
          4730 => x"38",
          4731 => x"76",
          4732 => x"70",
          4733 => x"16",
          4734 => x"74",
          4735 => x"96",
          4736 => x"dc",
          4737 => x"38",
          4738 => x"06",
          4739 => x"33",
          4740 => x"89",
          4741 => x"08",
          4742 => x"54",
          4743 => x"fc",
          4744 => x"8c",
          4745 => x"fe",
          4746 => x"ff",
          4747 => x"11",
          4748 => x"2b",
          4749 => x"81",
          4750 => x"2a",
          4751 => x"51",
          4752 => x"e2",
          4753 => x"ff",
          4754 => x"da",
          4755 => x"2a",
          4756 => x"05",
          4757 => x"fc",
          4758 => x"8c",
          4759 => x"c6",
          4760 => x"83",
          4761 => x"05",
          4762 => x"f9",
          4763 => x"8c",
          4764 => x"ff",
          4765 => x"ae",
          4766 => x"2a",
          4767 => x"05",
          4768 => x"fc",
          4769 => x"8c",
          4770 => x"38",
          4771 => x"83",
          4772 => x"05",
          4773 => x"f8",
          4774 => x"8c",
          4775 => x"0a",
          4776 => x"39",
          4777 => x"82",
          4778 => x"89",
          4779 => x"f8",
          4780 => x"7c",
          4781 => x"56",
          4782 => x"77",
          4783 => x"38",
          4784 => x"08",
          4785 => x"38",
          4786 => x"72",
          4787 => x"9d",
          4788 => x"24",
          4789 => x"81",
          4790 => x"82",
          4791 => x"83",
          4792 => x"38",
          4793 => x"76",
          4794 => x"70",
          4795 => x"18",
          4796 => x"76",
          4797 => x"9e",
          4798 => x"dc",
          4799 => x"8c",
          4800 => x"d9",
          4801 => x"ff",
          4802 => x"05",
          4803 => x"81",
          4804 => x"54",
          4805 => x"80",
          4806 => x"77",
          4807 => x"f0",
          4808 => x"8f",
          4809 => x"51",
          4810 => x"34",
          4811 => x"17",
          4812 => x"2a",
          4813 => x"05",
          4814 => x"fa",
          4815 => x"8c",
          4816 => x"82",
          4817 => x"81",
          4818 => x"83",
          4819 => x"b4",
          4820 => x"2a",
          4821 => x"8f",
          4822 => x"2a",
          4823 => x"f0",
          4824 => x"06",
          4825 => x"72",
          4826 => x"ec",
          4827 => x"2a",
          4828 => x"05",
          4829 => x"fa",
          4830 => x"8c",
          4831 => x"82",
          4832 => x"80",
          4833 => x"83",
          4834 => x"52",
          4835 => x"fe",
          4836 => x"b4",
          4837 => x"a4",
          4838 => x"76",
          4839 => x"17",
          4840 => x"75",
          4841 => x"3f",
          4842 => x"08",
          4843 => x"dc",
          4844 => x"77",
          4845 => x"77",
          4846 => x"fc",
          4847 => x"b4",
          4848 => x"51",
          4849 => x"c9",
          4850 => x"dc",
          4851 => x"06",
          4852 => x"72",
          4853 => x"3f",
          4854 => x"17",
          4855 => x"8c",
          4856 => x"3d",
          4857 => x"3d",
          4858 => x"7e",
          4859 => x"56",
          4860 => x"75",
          4861 => x"74",
          4862 => x"27",
          4863 => x"80",
          4864 => x"ff",
          4865 => x"75",
          4866 => x"3f",
          4867 => x"08",
          4868 => x"dc",
          4869 => x"38",
          4870 => x"54",
          4871 => x"81",
          4872 => x"39",
          4873 => x"08",
          4874 => x"39",
          4875 => x"51",
          4876 => x"82",
          4877 => x"58",
          4878 => x"08",
          4879 => x"c7",
          4880 => x"dc",
          4881 => x"d2",
          4882 => x"dc",
          4883 => x"cf",
          4884 => x"74",
          4885 => x"fc",
          4886 => x"8c",
          4887 => x"38",
          4888 => x"fe",
          4889 => x"08",
          4890 => x"74",
          4891 => x"38",
          4892 => x"17",
          4893 => x"33",
          4894 => x"73",
          4895 => x"77",
          4896 => x"26",
          4897 => x"80",
          4898 => x"8c",
          4899 => x"3d",
          4900 => x"3d",
          4901 => x"71",
          4902 => x"5b",
          4903 => x"8c",
          4904 => x"77",
          4905 => x"38",
          4906 => x"78",
          4907 => x"81",
          4908 => x"79",
          4909 => x"f9",
          4910 => x"55",
          4911 => x"dc",
          4912 => x"e0",
          4913 => x"dc",
          4914 => x"8c",
          4915 => x"2e",
          4916 => x"98",
          4917 => x"8c",
          4918 => x"82",
          4919 => x"58",
          4920 => x"70",
          4921 => x"80",
          4922 => x"38",
          4923 => x"09",
          4924 => x"e2",
          4925 => x"56",
          4926 => x"76",
          4927 => x"82",
          4928 => x"7a",
          4929 => x"3f",
          4930 => x"8c",
          4931 => x"2e",
          4932 => x"86",
          4933 => x"dc",
          4934 => x"8c",
          4935 => x"70",
          4936 => x"07",
          4937 => x"7c",
          4938 => x"dc",
          4939 => x"51",
          4940 => x"81",
          4941 => x"8c",
          4942 => x"2e",
          4943 => x"17",
          4944 => x"74",
          4945 => x"73",
          4946 => x"27",
          4947 => x"58",
          4948 => x"80",
          4949 => x"56",
          4950 => x"98",
          4951 => x"26",
          4952 => x"56",
          4953 => x"81",
          4954 => x"52",
          4955 => x"c6",
          4956 => x"dc",
          4957 => x"b8",
          4958 => x"82",
          4959 => x"81",
          4960 => x"06",
          4961 => x"8c",
          4962 => x"82",
          4963 => x"09",
          4964 => x"72",
          4965 => x"70",
          4966 => x"51",
          4967 => x"80",
          4968 => x"78",
          4969 => x"06",
          4970 => x"73",
          4971 => x"39",
          4972 => x"52",
          4973 => x"f7",
          4974 => x"dc",
          4975 => x"dc",
          4976 => x"82",
          4977 => x"07",
          4978 => x"55",
          4979 => x"2e",
          4980 => x"80",
          4981 => x"75",
          4982 => x"76",
          4983 => x"3f",
          4984 => x"08",
          4985 => x"38",
          4986 => x"0c",
          4987 => x"fe",
          4988 => x"08",
          4989 => x"74",
          4990 => x"ff",
          4991 => x"0c",
          4992 => x"81",
          4993 => x"84",
          4994 => x"39",
          4995 => x"81",
          4996 => x"8c",
          4997 => x"8c",
          4998 => x"dc",
          4999 => x"39",
          5000 => x"55",
          5001 => x"dc",
          5002 => x"0d",
          5003 => x"0d",
          5004 => x"55",
          5005 => x"82",
          5006 => x"58",
          5007 => x"8c",
          5008 => x"d8",
          5009 => x"74",
          5010 => x"3f",
          5011 => x"08",
          5012 => x"08",
          5013 => x"59",
          5014 => x"77",
          5015 => x"70",
          5016 => x"c8",
          5017 => x"84",
          5018 => x"56",
          5019 => x"58",
          5020 => x"97",
          5021 => x"75",
          5022 => x"52",
          5023 => x"51",
          5024 => x"82",
          5025 => x"80",
          5026 => x"8a",
          5027 => x"32",
          5028 => x"72",
          5029 => x"2a",
          5030 => x"56",
          5031 => x"dc",
          5032 => x"0d",
          5033 => x"0d",
          5034 => x"08",
          5035 => x"74",
          5036 => x"26",
          5037 => x"74",
          5038 => x"72",
          5039 => x"74",
          5040 => x"88",
          5041 => x"73",
          5042 => x"33",
          5043 => x"27",
          5044 => x"16",
          5045 => x"9b",
          5046 => x"2a",
          5047 => x"88",
          5048 => x"58",
          5049 => x"80",
          5050 => x"16",
          5051 => x"0c",
          5052 => x"8a",
          5053 => x"89",
          5054 => x"72",
          5055 => x"38",
          5056 => x"51",
          5057 => x"82",
          5058 => x"54",
          5059 => x"08",
          5060 => x"38",
          5061 => x"8c",
          5062 => x"8b",
          5063 => x"08",
          5064 => x"08",
          5065 => x"82",
          5066 => x"74",
          5067 => x"cb",
          5068 => x"75",
          5069 => x"3f",
          5070 => x"08",
          5071 => x"73",
          5072 => x"98",
          5073 => x"82",
          5074 => x"2e",
          5075 => x"39",
          5076 => x"39",
          5077 => x"13",
          5078 => x"74",
          5079 => x"16",
          5080 => x"18",
          5081 => x"77",
          5082 => x"0c",
          5083 => x"04",
          5084 => x"7a",
          5085 => x"12",
          5086 => x"59",
          5087 => x"80",
          5088 => x"86",
          5089 => x"98",
          5090 => x"14",
          5091 => x"55",
          5092 => x"81",
          5093 => x"83",
          5094 => x"77",
          5095 => x"81",
          5096 => x"0c",
          5097 => x"55",
          5098 => x"76",
          5099 => x"17",
          5100 => x"74",
          5101 => x"9b",
          5102 => x"39",
          5103 => x"ff",
          5104 => x"2a",
          5105 => x"81",
          5106 => x"52",
          5107 => x"e6",
          5108 => x"dc",
          5109 => x"55",
          5110 => x"8c",
          5111 => x"80",
          5112 => x"55",
          5113 => x"08",
          5114 => x"f4",
          5115 => x"08",
          5116 => x"08",
          5117 => x"38",
          5118 => x"77",
          5119 => x"84",
          5120 => x"39",
          5121 => x"52",
          5122 => x"86",
          5123 => x"dc",
          5124 => x"55",
          5125 => x"08",
          5126 => x"c4",
          5127 => x"82",
          5128 => x"81",
          5129 => x"81",
          5130 => x"dc",
          5131 => x"b0",
          5132 => x"dc",
          5133 => x"51",
          5134 => x"82",
          5135 => x"a0",
          5136 => x"15",
          5137 => x"75",
          5138 => x"3f",
          5139 => x"08",
          5140 => x"76",
          5141 => x"77",
          5142 => x"9c",
          5143 => x"55",
          5144 => x"dc",
          5145 => x"0d",
          5146 => x"0d",
          5147 => x"08",
          5148 => x"80",
          5149 => x"fc",
          5150 => x"8c",
          5151 => x"82",
          5152 => x"80",
          5153 => x"8c",
          5154 => x"98",
          5155 => x"78",
          5156 => x"3f",
          5157 => x"08",
          5158 => x"dc",
          5159 => x"38",
          5160 => x"08",
          5161 => x"70",
          5162 => x"58",
          5163 => x"2e",
          5164 => x"83",
          5165 => x"82",
          5166 => x"55",
          5167 => x"81",
          5168 => x"07",
          5169 => x"2e",
          5170 => x"16",
          5171 => x"2e",
          5172 => x"88",
          5173 => x"82",
          5174 => x"56",
          5175 => x"51",
          5176 => x"82",
          5177 => x"54",
          5178 => x"08",
          5179 => x"9b",
          5180 => x"2e",
          5181 => x"83",
          5182 => x"73",
          5183 => x"0c",
          5184 => x"04",
          5185 => x"76",
          5186 => x"54",
          5187 => x"82",
          5188 => x"83",
          5189 => x"76",
          5190 => x"53",
          5191 => x"2e",
          5192 => x"90",
          5193 => x"51",
          5194 => x"82",
          5195 => x"90",
          5196 => x"53",
          5197 => x"dc",
          5198 => x"0d",
          5199 => x"0d",
          5200 => x"83",
          5201 => x"54",
          5202 => x"55",
          5203 => x"3f",
          5204 => x"51",
          5205 => x"2e",
          5206 => x"8b",
          5207 => x"2a",
          5208 => x"51",
          5209 => x"86",
          5210 => x"f7",
          5211 => x"7d",
          5212 => x"75",
          5213 => x"98",
          5214 => x"2e",
          5215 => x"98",
          5216 => x"78",
          5217 => x"3f",
          5218 => x"08",
          5219 => x"dc",
          5220 => x"38",
          5221 => x"70",
          5222 => x"73",
          5223 => x"58",
          5224 => x"8b",
          5225 => x"bf",
          5226 => x"ff",
          5227 => x"53",
          5228 => x"34",
          5229 => x"08",
          5230 => x"e5",
          5231 => x"81",
          5232 => x"2e",
          5233 => x"70",
          5234 => x"57",
          5235 => x"9e",
          5236 => x"2e",
          5237 => x"8c",
          5238 => x"df",
          5239 => x"72",
          5240 => x"81",
          5241 => x"76",
          5242 => x"2e",
          5243 => x"52",
          5244 => x"fc",
          5245 => x"dc",
          5246 => x"8c",
          5247 => x"38",
          5248 => x"fe",
          5249 => x"39",
          5250 => x"16",
          5251 => x"8c",
          5252 => x"3d",
          5253 => x"3d",
          5254 => x"08",
          5255 => x"52",
          5256 => x"c5",
          5257 => x"dc",
          5258 => x"8c",
          5259 => x"38",
          5260 => x"52",
          5261 => x"de",
          5262 => x"dc",
          5263 => x"8c",
          5264 => x"38",
          5265 => x"8c",
          5266 => x"9c",
          5267 => x"ea",
          5268 => x"53",
          5269 => x"9c",
          5270 => x"ea",
          5271 => x"0b",
          5272 => x"74",
          5273 => x"0c",
          5274 => x"04",
          5275 => x"75",
          5276 => x"12",
          5277 => x"53",
          5278 => x"9a",
          5279 => x"dc",
          5280 => x"9c",
          5281 => x"e5",
          5282 => x"0b",
          5283 => x"85",
          5284 => x"fa",
          5285 => x"7a",
          5286 => x"0b",
          5287 => x"98",
          5288 => x"2e",
          5289 => x"80",
          5290 => x"55",
          5291 => x"17",
          5292 => x"33",
          5293 => x"51",
          5294 => x"2e",
          5295 => x"85",
          5296 => x"06",
          5297 => x"e5",
          5298 => x"2e",
          5299 => x"8b",
          5300 => x"70",
          5301 => x"34",
          5302 => x"71",
          5303 => x"05",
          5304 => x"15",
          5305 => x"27",
          5306 => x"15",
          5307 => x"80",
          5308 => x"34",
          5309 => x"52",
          5310 => x"88",
          5311 => x"17",
          5312 => x"52",
          5313 => x"3f",
          5314 => x"08",
          5315 => x"12",
          5316 => x"3f",
          5317 => x"08",
          5318 => x"98",
          5319 => x"da",
          5320 => x"dc",
          5321 => x"23",
          5322 => x"04",
          5323 => x"7f",
          5324 => x"5b",
          5325 => x"33",
          5326 => x"73",
          5327 => x"38",
          5328 => x"80",
          5329 => x"38",
          5330 => x"8c",
          5331 => x"08",
          5332 => x"aa",
          5333 => x"41",
          5334 => x"33",
          5335 => x"73",
          5336 => x"81",
          5337 => x"81",
          5338 => x"dc",
          5339 => x"70",
          5340 => x"07",
          5341 => x"73",
          5342 => x"88",
          5343 => x"70",
          5344 => x"73",
          5345 => x"38",
          5346 => x"ab",
          5347 => x"52",
          5348 => x"91",
          5349 => x"dc",
          5350 => x"98",
          5351 => x"61",
          5352 => x"5a",
          5353 => x"a0",
          5354 => x"e7",
          5355 => x"70",
          5356 => x"79",
          5357 => x"73",
          5358 => x"81",
          5359 => x"38",
          5360 => x"33",
          5361 => x"ae",
          5362 => x"70",
          5363 => x"82",
          5364 => x"51",
          5365 => x"54",
          5366 => x"79",
          5367 => x"74",
          5368 => x"57",
          5369 => x"af",
          5370 => x"70",
          5371 => x"51",
          5372 => x"dc",
          5373 => x"73",
          5374 => x"38",
          5375 => x"82",
          5376 => x"19",
          5377 => x"54",
          5378 => x"82",
          5379 => x"54",
          5380 => x"78",
          5381 => x"81",
          5382 => x"54",
          5383 => x"81",
          5384 => x"af",
          5385 => x"77",
          5386 => x"70",
          5387 => x"25",
          5388 => x"07",
          5389 => x"51",
          5390 => x"2e",
          5391 => x"39",
          5392 => x"80",
          5393 => x"33",
          5394 => x"73",
          5395 => x"81",
          5396 => x"81",
          5397 => x"dc",
          5398 => x"70",
          5399 => x"07",
          5400 => x"73",
          5401 => x"b5",
          5402 => x"2e",
          5403 => x"83",
          5404 => x"76",
          5405 => x"07",
          5406 => x"2e",
          5407 => x"8b",
          5408 => x"77",
          5409 => x"30",
          5410 => x"71",
          5411 => x"53",
          5412 => x"55",
          5413 => x"38",
          5414 => x"5c",
          5415 => x"75",
          5416 => x"73",
          5417 => x"38",
          5418 => x"06",
          5419 => x"11",
          5420 => x"75",
          5421 => x"3f",
          5422 => x"08",
          5423 => x"38",
          5424 => x"33",
          5425 => x"54",
          5426 => x"e6",
          5427 => x"8c",
          5428 => x"2e",
          5429 => x"ff",
          5430 => x"74",
          5431 => x"38",
          5432 => x"75",
          5433 => x"17",
          5434 => x"57",
          5435 => x"a7",
          5436 => x"81",
          5437 => x"e5",
          5438 => x"8c",
          5439 => x"38",
          5440 => x"54",
          5441 => x"89",
          5442 => x"70",
          5443 => x"57",
          5444 => x"54",
          5445 => x"81",
          5446 => x"f7",
          5447 => x"7e",
          5448 => x"2e",
          5449 => x"33",
          5450 => x"e5",
          5451 => x"06",
          5452 => x"7a",
          5453 => x"a0",
          5454 => x"38",
          5455 => x"55",
          5456 => x"84",
          5457 => x"39",
          5458 => x"8b",
          5459 => x"7b",
          5460 => x"7a",
          5461 => x"3f",
          5462 => x"08",
          5463 => x"dc",
          5464 => x"38",
          5465 => x"52",
          5466 => x"aa",
          5467 => x"dc",
          5468 => x"8c",
          5469 => x"c2",
          5470 => x"08",
          5471 => x"55",
          5472 => x"ff",
          5473 => x"15",
          5474 => x"54",
          5475 => x"34",
          5476 => x"70",
          5477 => x"81",
          5478 => x"58",
          5479 => x"8b",
          5480 => x"74",
          5481 => x"3f",
          5482 => x"08",
          5483 => x"38",
          5484 => x"51",
          5485 => x"ff",
          5486 => x"ab",
          5487 => x"55",
          5488 => x"bb",
          5489 => x"2e",
          5490 => x"80",
          5491 => x"85",
          5492 => x"06",
          5493 => x"58",
          5494 => x"80",
          5495 => x"75",
          5496 => x"73",
          5497 => x"b5",
          5498 => x"0b",
          5499 => x"80",
          5500 => x"39",
          5501 => x"54",
          5502 => x"85",
          5503 => x"75",
          5504 => x"81",
          5505 => x"73",
          5506 => x"1b",
          5507 => x"2a",
          5508 => x"51",
          5509 => x"80",
          5510 => x"90",
          5511 => x"ff",
          5512 => x"05",
          5513 => x"f5",
          5514 => x"8c",
          5515 => x"1c",
          5516 => x"39",
          5517 => x"dc",
          5518 => x"0d",
          5519 => x"0d",
          5520 => x"7b",
          5521 => x"73",
          5522 => x"55",
          5523 => x"2e",
          5524 => x"75",
          5525 => x"57",
          5526 => x"26",
          5527 => x"ba",
          5528 => x"70",
          5529 => x"ba",
          5530 => x"06",
          5531 => x"73",
          5532 => x"70",
          5533 => x"51",
          5534 => x"89",
          5535 => x"82",
          5536 => x"ff",
          5537 => x"56",
          5538 => x"2e",
          5539 => x"80",
          5540 => x"dc",
          5541 => x"08",
          5542 => x"76",
          5543 => x"58",
          5544 => x"81",
          5545 => x"ff",
          5546 => x"53",
          5547 => x"26",
          5548 => x"13",
          5549 => x"06",
          5550 => x"9f",
          5551 => x"99",
          5552 => x"e0",
          5553 => x"ff",
          5554 => x"72",
          5555 => x"2a",
          5556 => x"72",
          5557 => x"06",
          5558 => x"ff",
          5559 => x"30",
          5560 => x"70",
          5561 => x"07",
          5562 => x"9f",
          5563 => x"54",
          5564 => x"80",
          5565 => x"81",
          5566 => x"59",
          5567 => x"25",
          5568 => x"8b",
          5569 => x"24",
          5570 => x"76",
          5571 => x"78",
          5572 => x"82",
          5573 => x"51",
          5574 => x"dc",
          5575 => x"0d",
          5576 => x"0d",
          5577 => x"0b",
          5578 => x"ff",
          5579 => x"0c",
          5580 => x"51",
          5581 => x"84",
          5582 => x"dc",
          5583 => x"38",
          5584 => x"51",
          5585 => x"82",
          5586 => x"83",
          5587 => x"54",
          5588 => x"82",
          5589 => x"09",
          5590 => x"e3",
          5591 => x"b4",
          5592 => x"57",
          5593 => x"2e",
          5594 => x"83",
          5595 => x"74",
          5596 => x"70",
          5597 => x"25",
          5598 => x"51",
          5599 => x"38",
          5600 => x"2e",
          5601 => x"b5",
          5602 => x"81",
          5603 => x"80",
          5604 => x"e0",
          5605 => x"8c",
          5606 => x"82",
          5607 => x"80",
          5608 => x"85",
          5609 => x"a0",
          5610 => x"16",
          5611 => x"3f",
          5612 => x"08",
          5613 => x"dc",
          5614 => x"83",
          5615 => x"74",
          5616 => x"0c",
          5617 => x"04",
          5618 => x"61",
          5619 => x"80",
          5620 => x"58",
          5621 => x"0c",
          5622 => x"e1",
          5623 => x"dc",
          5624 => x"56",
          5625 => x"8c",
          5626 => x"86",
          5627 => x"8c",
          5628 => x"29",
          5629 => x"05",
          5630 => x"53",
          5631 => x"80",
          5632 => x"38",
          5633 => x"76",
          5634 => x"74",
          5635 => x"72",
          5636 => x"38",
          5637 => x"51",
          5638 => x"82",
          5639 => x"81",
          5640 => x"81",
          5641 => x"72",
          5642 => x"80",
          5643 => x"38",
          5644 => x"70",
          5645 => x"53",
          5646 => x"86",
          5647 => x"a7",
          5648 => x"34",
          5649 => x"34",
          5650 => x"14",
          5651 => x"b2",
          5652 => x"dc",
          5653 => x"06",
          5654 => x"54",
          5655 => x"72",
          5656 => x"76",
          5657 => x"38",
          5658 => x"70",
          5659 => x"53",
          5660 => x"85",
          5661 => x"70",
          5662 => x"5b",
          5663 => x"82",
          5664 => x"81",
          5665 => x"76",
          5666 => x"81",
          5667 => x"38",
          5668 => x"56",
          5669 => x"83",
          5670 => x"70",
          5671 => x"80",
          5672 => x"83",
          5673 => x"dc",
          5674 => x"8c",
          5675 => x"76",
          5676 => x"05",
          5677 => x"16",
          5678 => x"56",
          5679 => x"d7",
          5680 => x"8d",
          5681 => x"72",
          5682 => x"54",
          5683 => x"57",
          5684 => x"95",
          5685 => x"73",
          5686 => x"3f",
          5687 => x"08",
          5688 => x"57",
          5689 => x"89",
          5690 => x"56",
          5691 => x"d7",
          5692 => x"76",
          5693 => x"f1",
          5694 => x"76",
          5695 => x"e9",
          5696 => x"51",
          5697 => x"82",
          5698 => x"83",
          5699 => x"53",
          5700 => x"2e",
          5701 => x"84",
          5702 => x"ca",
          5703 => x"da",
          5704 => x"dc",
          5705 => x"ff",
          5706 => x"8d",
          5707 => x"14",
          5708 => x"3f",
          5709 => x"08",
          5710 => x"15",
          5711 => x"14",
          5712 => x"34",
          5713 => x"33",
          5714 => x"81",
          5715 => x"54",
          5716 => x"72",
          5717 => x"91",
          5718 => x"ff",
          5719 => x"29",
          5720 => x"33",
          5721 => x"72",
          5722 => x"72",
          5723 => x"38",
          5724 => x"06",
          5725 => x"2e",
          5726 => x"56",
          5727 => x"80",
          5728 => x"da",
          5729 => x"8c",
          5730 => x"82",
          5731 => x"88",
          5732 => x"8f",
          5733 => x"56",
          5734 => x"38",
          5735 => x"51",
          5736 => x"82",
          5737 => x"83",
          5738 => x"55",
          5739 => x"80",
          5740 => x"da",
          5741 => x"8c",
          5742 => x"80",
          5743 => x"da",
          5744 => x"8c",
          5745 => x"ff",
          5746 => x"8d",
          5747 => x"2e",
          5748 => x"88",
          5749 => x"14",
          5750 => x"05",
          5751 => x"75",
          5752 => x"38",
          5753 => x"52",
          5754 => x"51",
          5755 => x"3f",
          5756 => x"08",
          5757 => x"dc",
          5758 => x"82",
          5759 => x"8c",
          5760 => x"ff",
          5761 => x"26",
          5762 => x"57",
          5763 => x"f5",
          5764 => x"82",
          5765 => x"f5",
          5766 => x"81",
          5767 => x"8d",
          5768 => x"2e",
          5769 => x"82",
          5770 => x"16",
          5771 => x"16",
          5772 => x"70",
          5773 => x"7a",
          5774 => x"0c",
          5775 => x"83",
          5776 => x"06",
          5777 => x"de",
          5778 => x"ae",
          5779 => x"dc",
          5780 => x"ff",
          5781 => x"56",
          5782 => x"38",
          5783 => x"38",
          5784 => x"51",
          5785 => x"82",
          5786 => x"a8",
          5787 => x"82",
          5788 => x"39",
          5789 => x"80",
          5790 => x"38",
          5791 => x"15",
          5792 => x"53",
          5793 => x"8d",
          5794 => x"15",
          5795 => x"76",
          5796 => x"51",
          5797 => x"13",
          5798 => x"8d",
          5799 => x"15",
          5800 => x"c5",
          5801 => x"90",
          5802 => x"0b",
          5803 => x"ff",
          5804 => x"15",
          5805 => x"2e",
          5806 => x"81",
          5807 => x"e4",
          5808 => x"b6",
          5809 => x"dc",
          5810 => x"ff",
          5811 => x"81",
          5812 => x"06",
          5813 => x"81",
          5814 => x"51",
          5815 => x"82",
          5816 => x"80",
          5817 => x"8c",
          5818 => x"15",
          5819 => x"14",
          5820 => x"3f",
          5821 => x"08",
          5822 => x"06",
          5823 => x"d4",
          5824 => x"81",
          5825 => x"38",
          5826 => x"d8",
          5827 => x"8c",
          5828 => x"8b",
          5829 => x"2e",
          5830 => x"b3",
          5831 => x"14",
          5832 => x"3f",
          5833 => x"08",
          5834 => x"e4",
          5835 => x"81",
          5836 => x"84",
          5837 => x"d7",
          5838 => x"8c",
          5839 => x"15",
          5840 => x"14",
          5841 => x"3f",
          5842 => x"08",
          5843 => x"76",
          5844 => x"8d",
          5845 => x"05",
          5846 => x"8d",
          5847 => x"86",
          5848 => x"0b",
          5849 => x"80",
          5850 => x"8c",
          5851 => x"3d",
          5852 => x"3d",
          5853 => x"89",
          5854 => x"2e",
          5855 => x"08",
          5856 => x"2e",
          5857 => x"33",
          5858 => x"2e",
          5859 => x"13",
          5860 => x"22",
          5861 => x"76",
          5862 => x"06",
          5863 => x"13",
          5864 => x"c0",
          5865 => x"dc",
          5866 => x"52",
          5867 => x"71",
          5868 => x"55",
          5869 => x"53",
          5870 => x"0c",
          5871 => x"8c",
          5872 => x"3d",
          5873 => x"3d",
          5874 => x"05",
          5875 => x"89",
          5876 => x"52",
          5877 => x"3f",
          5878 => x"0b",
          5879 => x"08",
          5880 => x"82",
          5881 => x"84",
          5882 => x"8c",
          5883 => x"55",
          5884 => x"2e",
          5885 => x"74",
          5886 => x"73",
          5887 => x"38",
          5888 => x"78",
          5889 => x"54",
          5890 => x"92",
          5891 => x"89",
          5892 => x"84",
          5893 => x"b0",
          5894 => x"dc",
          5895 => x"82",
          5896 => x"88",
          5897 => x"eb",
          5898 => x"02",
          5899 => x"e7",
          5900 => x"59",
          5901 => x"80",
          5902 => x"38",
          5903 => x"70",
          5904 => x"d0",
          5905 => x"3d",
          5906 => x"58",
          5907 => x"82",
          5908 => x"55",
          5909 => x"08",
          5910 => x"7a",
          5911 => x"8c",
          5912 => x"56",
          5913 => x"82",
          5914 => x"55",
          5915 => x"08",
          5916 => x"80",
          5917 => x"70",
          5918 => x"57",
          5919 => x"83",
          5920 => x"77",
          5921 => x"73",
          5922 => x"ab",
          5923 => x"2e",
          5924 => x"84",
          5925 => x"06",
          5926 => x"51",
          5927 => x"82",
          5928 => x"55",
          5929 => x"b2",
          5930 => x"06",
          5931 => x"b8",
          5932 => x"2a",
          5933 => x"51",
          5934 => x"2e",
          5935 => x"55",
          5936 => x"77",
          5937 => x"74",
          5938 => x"77",
          5939 => x"81",
          5940 => x"73",
          5941 => x"af",
          5942 => x"7a",
          5943 => x"3f",
          5944 => x"08",
          5945 => x"b2",
          5946 => x"8e",
          5947 => x"ea",
          5948 => x"a0",
          5949 => x"34",
          5950 => x"52",
          5951 => x"bd",
          5952 => x"62",
          5953 => x"d4",
          5954 => x"54",
          5955 => x"15",
          5956 => x"2e",
          5957 => x"7a",
          5958 => x"51",
          5959 => x"75",
          5960 => x"d4",
          5961 => x"be",
          5962 => x"dc",
          5963 => x"8c",
          5964 => x"ca",
          5965 => x"74",
          5966 => x"02",
          5967 => x"70",
          5968 => x"81",
          5969 => x"56",
          5970 => x"86",
          5971 => x"82",
          5972 => x"81",
          5973 => x"06",
          5974 => x"80",
          5975 => x"75",
          5976 => x"73",
          5977 => x"38",
          5978 => x"92",
          5979 => x"7a",
          5980 => x"3f",
          5981 => x"08",
          5982 => x"8c",
          5983 => x"55",
          5984 => x"08",
          5985 => x"77",
          5986 => x"81",
          5987 => x"73",
          5988 => x"38",
          5989 => x"07",
          5990 => x"11",
          5991 => x"0c",
          5992 => x"0c",
          5993 => x"52",
          5994 => x"3f",
          5995 => x"08",
          5996 => x"08",
          5997 => x"63",
          5998 => x"5a",
          5999 => x"82",
          6000 => x"82",
          6001 => x"8c",
          6002 => x"7a",
          6003 => x"17",
          6004 => x"23",
          6005 => x"34",
          6006 => x"1a",
          6007 => x"9c",
          6008 => x"0b",
          6009 => x"77",
          6010 => x"81",
          6011 => x"73",
          6012 => x"8d",
          6013 => x"dc",
          6014 => x"81",
          6015 => x"8c",
          6016 => x"1a",
          6017 => x"22",
          6018 => x"7b",
          6019 => x"a8",
          6020 => x"78",
          6021 => x"3f",
          6022 => x"08",
          6023 => x"dc",
          6024 => x"83",
          6025 => x"82",
          6026 => x"ff",
          6027 => x"06",
          6028 => x"55",
          6029 => x"56",
          6030 => x"76",
          6031 => x"51",
          6032 => x"27",
          6033 => x"70",
          6034 => x"5a",
          6035 => x"76",
          6036 => x"74",
          6037 => x"83",
          6038 => x"73",
          6039 => x"38",
          6040 => x"51",
          6041 => x"82",
          6042 => x"85",
          6043 => x"8e",
          6044 => x"2a",
          6045 => x"08",
          6046 => x"0c",
          6047 => x"79",
          6048 => x"73",
          6049 => x"0c",
          6050 => x"04",
          6051 => x"60",
          6052 => x"40",
          6053 => x"80",
          6054 => x"3d",
          6055 => x"78",
          6056 => x"3f",
          6057 => x"08",
          6058 => x"dc",
          6059 => x"91",
          6060 => x"74",
          6061 => x"38",
          6062 => x"c4",
          6063 => x"33",
          6064 => x"87",
          6065 => x"2e",
          6066 => x"95",
          6067 => x"91",
          6068 => x"56",
          6069 => x"81",
          6070 => x"34",
          6071 => x"a0",
          6072 => x"08",
          6073 => x"31",
          6074 => x"27",
          6075 => x"5c",
          6076 => x"82",
          6077 => x"19",
          6078 => x"ff",
          6079 => x"74",
          6080 => x"7e",
          6081 => x"ff",
          6082 => x"2a",
          6083 => x"79",
          6084 => x"87",
          6085 => x"08",
          6086 => x"98",
          6087 => x"78",
          6088 => x"3f",
          6089 => x"08",
          6090 => x"27",
          6091 => x"74",
          6092 => x"a3",
          6093 => x"1a",
          6094 => x"08",
          6095 => x"d4",
          6096 => x"8c",
          6097 => x"2e",
          6098 => x"82",
          6099 => x"1a",
          6100 => x"59",
          6101 => x"2e",
          6102 => x"77",
          6103 => x"11",
          6104 => x"55",
          6105 => x"85",
          6106 => x"31",
          6107 => x"76",
          6108 => x"81",
          6109 => x"ca",
          6110 => x"8c",
          6111 => x"d7",
          6112 => x"11",
          6113 => x"74",
          6114 => x"38",
          6115 => x"77",
          6116 => x"78",
          6117 => x"84",
          6118 => x"16",
          6119 => x"08",
          6120 => x"2b",
          6121 => x"cf",
          6122 => x"89",
          6123 => x"39",
          6124 => x"0c",
          6125 => x"83",
          6126 => x"80",
          6127 => x"55",
          6128 => x"83",
          6129 => x"9c",
          6130 => x"7e",
          6131 => x"3f",
          6132 => x"08",
          6133 => x"75",
          6134 => x"08",
          6135 => x"1f",
          6136 => x"7c",
          6137 => x"3f",
          6138 => x"7e",
          6139 => x"0c",
          6140 => x"1b",
          6141 => x"1c",
          6142 => x"fd",
          6143 => x"56",
          6144 => x"dc",
          6145 => x"0d",
          6146 => x"0d",
          6147 => x"64",
          6148 => x"58",
          6149 => x"90",
          6150 => x"52",
          6151 => x"d2",
          6152 => x"dc",
          6153 => x"8c",
          6154 => x"38",
          6155 => x"55",
          6156 => x"86",
          6157 => x"83",
          6158 => x"18",
          6159 => x"2a",
          6160 => x"51",
          6161 => x"56",
          6162 => x"83",
          6163 => x"39",
          6164 => x"19",
          6165 => x"83",
          6166 => x"0b",
          6167 => x"81",
          6168 => x"39",
          6169 => x"7c",
          6170 => x"74",
          6171 => x"38",
          6172 => x"7b",
          6173 => x"ec",
          6174 => x"08",
          6175 => x"06",
          6176 => x"81",
          6177 => x"8a",
          6178 => x"05",
          6179 => x"06",
          6180 => x"bf",
          6181 => x"38",
          6182 => x"55",
          6183 => x"7a",
          6184 => x"98",
          6185 => x"77",
          6186 => x"3f",
          6187 => x"08",
          6188 => x"dc",
          6189 => x"82",
          6190 => x"81",
          6191 => x"38",
          6192 => x"ff",
          6193 => x"98",
          6194 => x"18",
          6195 => x"74",
          6196 => x"7e",
          6197 => x"08",
          6198 => x"2e",
          6199 => x"8d",
          6200 => x"ce",
          6201 => x"8c",
          6202 => x"ee",
          6203 => x"08",
          6204 => x"d1",
          6205 => x"8c",
          6206 => x"2e",
          6207 => x"82",
          6208 => x"1b",
          6209 => x"5a",
          6210 => x"2e",
          6211 => x"78",
          6212 => x"11",
          6213 => x"55",
          6214 => x"85",
          6215 => x"31",
          6216 => x"76",
          6217 => x"81",
          6218 => x"c8",
          6219 => x"8c",
          6220 => x"a6",
          6221 => x"11",
          6222 => x"56",
          6223 => x"27",
          6224 => x"80",
          6225 => x"08",
          6226 => x"2b",
          6227 => x"b4",
          6228 => x"b5",
          6229 => x"80",
          6230 => x"34",
          6231 => x"56",
          6232 => x"8c",
          6233 => x"19",
          6234 => x"38",
          6235 => x"b6",
          6236 => x"dc",
          6237 => x"38",
          6238 => x"12",
          6239 => x"9c",
          6240 => x"18",
          6241 => x"06",
          6242 => x"31",
          6243 => x"76",
          6244 => x"7b",
          6245 => x"08",
          6246 => x"cd",
          6247 => x"8c",
          6248 => x"b6",
          6249 => x"7c",
          6250 => x"08",
          6251 => x"1f",
          6252 => x"cb",
          6253 => x"55",
          6254 => x"16",
          6255 => x"31",
          6256 => x"7f",
          6257 => x"94",
          6258 => x"70",
          6259 => x"8c",
          6260 => x"58",
          6261 => x"76",
          6262 => x"75",
          6263 => x"19",
          6264 => x"39",
          6265 => x"80",
          6266 => x"74",
          6267 => x"80",
          6268 => x"8c",
          6269 => x"3d",
          6270 => x"3d",
          6271 => x"3d",
          6272 => x"70",
          6273 => x"ea",
          6274 => x"dc",
          6275 => x"8c",
          6276 => x"fb",
          6277 => x"33",
          6278 => x"70",
          6279 => x"55",
          6280 => x"2e",
          6281 => x"a0",
          6282 => x"78",
          6283 => x"3f",
          6284 => x"08",
          6285 => x"dc",
          6286 => x"38",
          6287 => x"8b",
          6288 => x"07",
          6289 => x"8b",
          6290 => x"16",
          6291 => x"52",
          6292 => x"dd",
          6293 => x"16",
          6294 => x"15",
          6295 => x"3f",
          6296 => x"0a",
          6297 => x"51",
          6298 => x"76",
          6299 => x"51",
          6300 => x"78",
          6301 => x"83",
          6302 => x"51",
          6303 => x"82",
          6304 => x"90",
          6305 => x"bf",
          6306 => x"73",
          6307 => x"76",
          6308 => x"0c",
          6309 => x"04",
          6310 => x"76",
          6311 => x"fe",
          6312 => x"8c",
          6313 => x"82",
          6314 => x"9c",
          6315 => x"fc",
          6316 => x"51",
          6317 => x"82",
          6318 => x"53",
          6319 => x"08",
          6320 => x"8c",
          6321 => x"0c",
          6322 => x"dc",
          6323 => x"0d",
          6324 => x"0d",
          6325 => x"e6",
          6326 => x"52",
          6327 => x"8c",
          6328 => x"8b",
          6329 => x"dc",
          6330 => x"a0",
          6331 => x"71",
          6332 => x"0c",
          6333 => x"04",
          6334 => x"80",
          6335 => x"d0",
          6336 => x"3d",
          6337 => x"3f",
          6338 => x"08",
          6339 => x"dc",
          6340 => x"38",
          6341 => x"52",
          6342 => x"05",
          6343 => x"3f",
          6344 => x"08",
          6345 => x"dc",
          6346 => x"02",
          6347 => x"33",
          6348 => x"55",
          6349 => x"25",
          6350 => x"7a",
          6351 => x"54",
          6352 => x"a2",
          6353 => x"84",
          6354 => x"06",
          6355 => x"73",
          6356 => x"38",
          6357 => x"70",
          6358 => x"a8",
          6359 => x"dc",
          6360 => x"0c",
          6361 => x"8c",
          6362 => x"2e",
          6363 => x"83",
          6364 => x"74",
          6365 => x"0c",
          6366 => x"04",
          6367 => x"6f",
          6368 => x"80",
          6369 => x"53",
          6370 => x"b8",
          6371 => x"3d",
          6372 => x"3f",
          6373 => x"08",
          6374 => x"dc",
          6375 => x"38",
          6376 => x"7c",
          6377 => x"47",
          6378 => x"54",
          6379 => x"81",
          6380 => x"52",
          6381 => x"52",
          6382 => x"3f",
          6383 => x"08",
          6384 => x"dc",
          6385 => x"38",
          6386 => x"51",
          6387 => x"82",
          6388 => x"57",
          6389 => x"08",
          6390 => x"69",
          6391 => x"da",
          6392 => x"8c",
          6393 => x"76",
          6394 => x"d5",
          6395 => x"8c",
          6396 => x"82",
          6397 => x"82",
          6398 => x"52",
          6399 => x"eb",
          6400 => x"dc",
          6401 => x"8c",
          6402 => x"38",
          6403 => x"51",
          6404 => x"73",
          6405 => x"08",
          6406 => x"76",
          6407 => x"d6",
          6408 => x"8c",
          6409 => x"82",
          6410 => x"80",
          6411 => x"76",
          6412 => x"81",
          6413 => x"82",
          6414 => x"39",
          6415 => x"38",
          6416 => x"bc",
          6417 => x"51",
          6418 => x"76",
          6419 => x"11",
          6420 => x"51",
          6421 => x"73",
          6422 => x"38",
          6423 => x"55",
          6424 => x"16",
          6425 => x"56",
          6426 => x"38",
          6427 => x"73",
          6428 => x"90",
          6429 => x"2e",
          6430 => x"16",
          6431 => x"ff",
          6432 => x"ff",
          6433 => x"58",
          6434 => x"74",
          6435 => x"75",
          6436 => x"18",
          6437 => x"58",
          6438 => x"fe",
          6439 => x"7b",
          6440 => x"06",
          6441 => x"18",
          6442 => x"58",
          6443 => x"80",
          6444 => x"a0",
          6445 => x"29",
          6446 => x"05",
          6447 => x"33",
          6448 => x"56",
          6449 => x"2e",
          6450 => x"16",
          6451 => x"33",
          6452 => x"73",
          6453 => x"16",
          6454 => x"26",
          6455 => x"55",
          6456 => x"91",
          6457 => x"54",
          6458 => x"70",
          6459 => x"34",
          6460 => x"ec",
          6461 => x"70",
          6462 => x"34",
          6463 => x"09",
          6464 => x"38",
          6465 => x"39",
          6466 => x"19",
          6467 => x"33",
          6468 => x"05",
          6469 => x"78",
          6470 => x"80",
          6471 => x"82",
          6472 => x"9e",
          6473 => x"f7",
          6474 => x"7d",
          6475 => x"05",
          6476 => x"57",
          6477 => x"3f",
          6478 => x"08",
          6479 => x"dc",
          6480 => x"38",
          6481 => x"53",
          6482 => x"38",
          6483 => x"54",
          6484 => x"92",
          6485 => x"33",
          6486 => x"70",
          6487 => x"54",
          6488 => x"38",
          6489 => x"15",
          6490 => x"70",
          6491 => x"58",
          6492 => x"82",
          6493 => x"8a",
          6494 => x"89",
          6495 => x"53",
          6496 => x"b7",
          6497 => x"ff",
          6498 => x"ff",
          6499 => x"8c",
          6500 => x"15",
          6501 => x"53",
          6502 => x"ff",
          6503 => x"8c",
          6504 => x"26",
          6505 => x"30",
          6506 => x"70",
          6507 => x"77",
          6508 => x"18",
          6509 => x"51",
          6510 => x"88",
          6511 => x"73",
          6512 => x"52",
          6513 => x"ca",
          6514 => x"dc",
          6515 => x"8c",
          6516 => x"2e",
          6517 => x"82",
          6518 => x"ff",
          6519 => x"38",
          6520 => x"08",
          6521 => x"73",
          6522 => x"73",
          6523 => x"9c",
          6524 => x"27",
          6525 => x"75",
          6526 => x"16",
          6527 => x"17",
          6528 => x"33",
          6529 => x"70",
          6530 => x"55",
          6531 => x"80",
          6532 => x"73",
          6533 => x"cc",
          6534 => x"8c",
          6535 => x"82",
          6536 => x"94",
          6537 => x"dc",
          6538 => x"39",
          6539 => x"51",
          6540 => x"82",
          6541 => x"54",
          6542 => x"be",
          6543 => x"27",
          6544 => x"53",
          6545 => x"08",
          6546 => x"73",
          6547 => x"ff",
          6548 => x"15",
          6549 => x"16",
          6550 => x"ff",
          6551 => x"80",
          6552 => x"73",
          6553 => x"c6",
          6554 => x"8c",
          6555 => x"38",
          6556 => x"16",
          6557 => x"80",
          6558 => x"0b",
          6559 => x"81",
          6560 => x"75",
          6561 => x"8c",
          6562 => x"58",
          6563 => x"54",
          6564 => x"74",
          6565 => x"73",
          6566 => x"90",
          6567 => x"c0",
          6568 => x"90",
          6569 => x"83",
          6570 => x"72",
          6571 => x"38",
          6572 => x"08",
          6573 => x"77",
          6574 => x"80",
          6575 => x"8c",
          6576 => x"3d",
          6577 => x"3d",
          6578 => x"89",
          6579 => x"2e",
          6580 => x"80",
          6581 => x"fc",
          6582 => x"3d",
          6583 => x"e1",
          6584 => x"8c",
          6585 => x"82",
          6586 => x"80",
          6587 => x"76",
          6588 => x"75",
          6589 => x"3f",
          6590 => x"08",
          6591 => x"dc",
          6592 => x"38",
          6593 => x"70",
          6594 => x"57",
          6595 => x"a2",
          6596 => x"33",
          6597 => x"70",
          6598 => x"55",
          6599 => x"2e",
          6600 => x"16",
          6601 => x"51",
          6602 => x"82",
          6603 => x"88",
          6604 => x"54",
          6605 => x"84",
          6606 => x"52",
          6607 => x"e5",
          6608 => x"dc",
          6609 => x"84",
          6610 => x"06",
          6611 => x"55",
          6612 => x"80",
          6613 => x"80",
          6614 => x"54",
          6615 => x"dc",
          6616 => x"0d",
          6617 => x"0d",
          6618 => x"fc",
          6619 => x"52",
          6620 => x"3f",
          6621 => x"08",
          6622 => x"8c",
          6623 => x"0c",
          6624 => x"04",
          6625 => x"77",
          6626 => x"fc",
          6627 => x"53",
          6628 => x"de",
          6629 => x"dc",
          6630 => x"8c",
          6631 => x"df",
          6632 => x"38",
          6633 => x"08",
          6634 => x"cd",
          6635 => x"8c",
          6636 => x"80",
          6637 => x"8c",
          6638 => x"73",
          6639 => x"3f",
          6640 => x"08",
          6641 => x"dc",
          6642 => x"09",
          6643 => x"38",
          6644 => x"39",
          6645 => x"08",
          6646 => x"52",
          6647 => x"b3",
          6648 => x"73",
          6649 => x"3f",
          6650 => x"08",
          6651 => x"30",
          6652 => x"9f",
          6653 => x"8c",
          6654 => x"51",
          6655 => x"72",
          6656 => x"0c",
          6657 => x"04",
          6658 => x"65",
          6659 => x"89",
          6660 => x"96",
          6661 => x"df",
          6662 => x"8c",
          6663 => x"82",
          6664 => x"b2",
          6665 => x"75",
          6666 => x"3f",
          6667 => x"08",
          6668 => x"dc",
          6669 => x"02",
          6670 => x"33",
          6671 => x"55",
          6672 => x"25",
          6673 => x"55",
          6674 => x"80",
          6675 => x"76",
          6676 => x"d4",
          6677 => x"82",
          6678 => x"94",
          6679 => x"f0",
          6680 => x"65",
          6681 => x"53",
          6682 => x"05",
          6683 => x"51",
          6684 => x"82",
          6685 => x"5b",
          6686 => x"08",
          6687 => x"7c",
          6688 => x"08",
          6689 => x"fe",
          6690 => x"08",
          6691 => x"55",
          6692 => x"91",
          6693 => x"0c",
          6694 => x"81",
          6695 => x"39",
          6696 => x"c7",
          6697 => x"dc",
          6698 => x"55",
          6699 => x"2e",
          6700 => x"bf",
          6701 => x"5f",
          6702 => x"92",
          6703 => x"51",
          6704 => x"82",
          6705 => x"ff",
          6706 => x"82",
          6707 => x"81",
          6708 => x"82",
          6709 => x"30",
          6710 => x"dc",
          6711 => x"25",
          6712 => x"19",
          6713 => x"5a",
          6714 => x"08",
          6715 => x"38",
          6716 => x"a4",
          6717 => x"8c",
          6718 => x"58",
          6719 => x"77",
          6720 => x"7d",
          6721 => x"bf",
          6722 => x"8c",
          6723 => x"82",
          6724 => x"80",
          6725 => x"70",
          6726 => x"ff",
          6727 => x"56",
          6728 => x"2e",
          6729 => x"9e",
          6730 => x"51",
          6731 => x"3f",
          6732 => x"08",
          6733 => x"06",
          6734 => x"80",
          6735 => x"19",
          6736 => x"54",
          6737 => x"14",
          6738 => x"c5",
          6739 => x"dc",
          6740 => x"06",
          6741 => x"80",
          6742 => x"19",
          6743 => x"54",
          6744 => x"06",
          6745 => x"79",
          6746 => x"78",
          6747 => x"79",
          6748 => x"84",
          6749 => x"07",
          6750 => x"84",
          6751 => x"82",
          6752 => x"92",
          6753 => x"f9",
          6754 => x"8a",
          6755 => x"53",
          6756 => x"e3",
          6757 => x"8c",
          6758 => x"82",
          6759 => x"81",
          6760 => x"17",
          6761 => x"81",
          6762 => x"17",
          6763 => x"2a",
          6764 => x"51",
          6765 => x"55",
          6766 => x"81",
          6767 => x"17",
          6768 => x"8c",
          6769 => x"81",
          6770 => x"9b",
          6771 => x"dc",
          6772 => x"17",
          6773 => x"51",
          6774 => x"82",
          6775 => x"74",
          6776 => x"56",
          6777 => x"98",
          6778 => x"76",
          6779 => x"c6",
          6780 => x"dc",
          6781 => x"09",
          6782 => x"38",
          6783 => x"8c",
          6784 => x"2e",
          6785 => x"85",
          6786 => x"a3",
          6787 => x"38",
          6788 => x"8c",
          6789 => x"15",
          6790 => x"38",
          6791 => x"53",
          6792 => x"08",
          6793 => x"c3",
          6794 => x"8c",
          6795 => x"94",
          6796 => x"18",
          6797 => x"33",
          6798 => x"54",
          6799 => x"34",
          6800 => x"85",
          6801 => x"18",
          6802 => x"74",
          6803 => x"0c",
          6804 => x"04",
          6805 => x"82",
          6806 => x"ff",
          6807 => x"a1",
          6808 => x"e4",
          6809 => x"dc",
          6810 => x"8c",
          6811 => x"f5",
          6812 => x"a1",
          6813 => x"95",
          6814 => x"58",
          6815 => x"82",
          6816 => x"55",
          6817 => x"08",
          6818 => x"02",
          6819 => x"33",
          6820 => x"70",
          6821 => x"55",
          6822 => x"73",
          6823 => x"75",
          6824 => x"80",
          6825 => x"bd",
          6826 => x"d6",
          6827 => x"81",
          6828 => x"87",
          6829 => x"ad",
          6830 => x"78",
          6831 => x"3f",
          6832 => x"08",
          6833 => x"70",
          6834 => x"55",
          6835 => x"2e",
          6836 => x"78",
          6837 => x"dc",
          6838 => x"08",
          6839 => x"38",
          6840 => x"8c",
          6841 => x"76",
          6842 => x"70",
          6843 => x"b5",
          6844 => x"dc",
          6845 => x"8c",
          6846 => x"e9",
          6847 => x"dc",
          6848 => x"51",
          6849 => x"82",
          6850 => x"55",
          6851 => x"08",
          6852 => x"55",
          6853 => x"82",
          6854 => x"84",
          6855 => x"82",
          6856 => x"80",
          6857 => x"51",
          6858 => x"82",
          6859 => x"82",
          6860 => x"30",
          6861 => x"dc",
          6862 => x"25",
          6863 => x"75",
          6864 => x"38",
          6865 => x"8f",
          6866 => x"75",
          6867 => x"c1",
          6868 => x"8c",
          6869 => x"74",
          6870 => x"51",
          6871 => x"3f",
          6872 => x"08",
          6873 => x"8c",
          6874 => x"3d",
          6875 => x"3d",
          6876 => x"99",
          6877 => x"52",
          6878 => x"d8",
          6879 => x"8c",
          6880 => x"82",
          6881 => x"82",
          6882 => x"5e",
          6883 => x"3d",
          6884 => x"cf",
          6885 => x"8c",
          6886 => x"82",
          6887 => x"86",
          6888 => x"82",
          6889 => x"8c",
          6890 => x"2e",
          6891 => x"82",
          6892 => x"80",
          6893 => x"70",
          6894 => x"06",
          6895 => x"54",
          6896 => x"38",
          6897 => x"52",
          6898 => x"52",
          6899 => x"3f",
          6900 => x"08",
          6901 => x"82",
          6902 => x"83",
          6903 => x"82",
          6904 => x"81",
          6905 => x"06",
          6906 => x"54",
          6907 => x"08",
          6908 => x"81",
          6909 => x"81",
          6910 => x"39",
          6911 => x"38",
          6912 => x"08",
          6913 => x"c4",
          6914 => x"8c",
          6915 => x"82",
          6916 => x"81",
          6917 => x"53",
          6918 => x"19",
          6919 => x"8c",
          6920 => x"ae",
          6921 => x"34",
          6922 => x"0b",
          6923 => x"82",
          6924 => x"52",
          6925 => x"51",
          6926 => x"3f",
          6927 => x"b4",
          6928 => x"c9",
          6929 => x"53",
          6930 => x"53",
          6931 => x"51",
          6932 => x"3f",
          6933 => x"0b",
          6934 => x"34",
          6935 => x"80",
          6936 => x"51",
          6937 => x"78",
          6938 => x"83",
          6939 => x"51",
          6940 => x"82",
          6941 => x"54",
          6942 => x"08",
          6943 => x"88",
          6944 => x"64",
          6945 => x"ff",
          6946 => x"75",
          6947 => x"78",
          6948 => x"3f",
          6949 => x"0b",
          6950 => x"78",
          6951 => x"83",
          6952 => x"51",
          6953 => x"3f",
          6954 => x"08",
          6955 => x"80",
          6956 => x"76",
          6957 => x"ae",
          6958 => x"8c",
          6959 => x"3d",
          6960 => x"3d",
          6961 => x"84",
          6962 => x"f1",
          6963 => x"a8",
          6964 => x"05",
          6965 => x"51",
          6966 => x"82",
          6967 => x"55",
          6968 => x"08",
          6969 => x"78",
          6970 => x"08",
          6971 => x"70",
          6972 => x"b8",
          6973 => x"dc",
          6974 => x"8c",
          6975 => x"b9",
          6976 => x"9b",
          6977 => x"a0",
          6978 => x"55",
          6979 => x"38",
          6980 => x"3d",
          6981 => x"3d",
          6982 => x"51",
          6983 => x"3f",
          6984 => x"52",
          6985 => x"52",
          6986 => x"dd",
          6987 => x"08",
          6988 => x"cb",
          6989 => x"8c",
          6990 => x"82",
          6991 => x"95",
          6992 => x"2e",
          6993 => x"88",
          6994 => x"3d",
          6995 => x"38",
          6996 => x"e5",
          6997 => x"dc",
          6998 => x"09",
          6999 => x"b8",
          7000 => x"c9",
          7001 => x"8c",
          7002 => x"82",
          7003 => x"81",
          7004 => x"56",
          7005 => x"3d",
          7006 => x"52",
          7007 => x"ff",
          7008 => x"02",
          7009 => x"8b",
          7010 => x"16",
          7011 => x"2a",
          7012 => x"51",
          7013 => x"89",
          7014 => x"07",
          7015 => x"17",
          7016 => x"81",
          7017 => x"34",
          7018 => x"70",
          7019 => x"81",
          7020 => x"55",
          7021 => x"80",
          7022 => x"64",
          7023 => x"38",
          7024 => x"51",
          7025 => x"82",
          7026 => x"52",
          7027 => x"b7",
          7028 => x"55",
          7029 => x"08",
          7030 => x"dd",
          7031 => x"dc",
          7032 => x"51",
          7033 => x"3f",
          7034 => x"08",
          7035 => x"11",
          7036 => x"82",
          7037 => x"80",
          7038 => x"16",
          7039 => x"ae",
          7040 => x"06",
          7041 => x"53",
          7042 => x"51",
          7043 => x"78",
          7044 => x"83",
          7045 => x"39",
          7046 => x"08",
          7047 => x"51",
          7048 => x"82",
          7049 => x"55",
          7050 => x"08",
          7051 => x"51",
          7052 => x"3f",
          7053 => x"08",
          7054 => x"8c",
          7055 => x"3d",
          7056 => x"3d",
          7057 => x"db",
          7058 => x"84",
          7059 => x"05",
          7060 => x"82",
          7061 => x"d0",
          7062 => x"3d",
          7063 => x"3f",
          7064 => x"08",
          7065 => x"dc",
          7066 => x"38",
          7067 => x"52",
          7068 => x"05",
          7069 => x"3f",
          7070 => x"08",
          7071 => x"dc",
          7072 => x"02",
          7073 => x"33",
          7074 => x"54",
          7075 => x"aa",
          7076 => x"06",
          7077 => x"8b",
          7078 => x"06",
          7079 => x"07",
          7080 => x"56",
          7081 => x"34",
          7082 => x"0b",
          7083 => x"78",
          7084 => x"a9",
          7085 => x"dc",
          7086 => x"82",
          7087 => x"95",
          7088 => x"ef",
          7089 => x"56",
          7090 => x"3d",
          7091 => x"94",
          7092 => x"f4",
          7093 => x"dc",
          7094 => x"8c",
          7095 => x"cb",
          7096 => x"63",
          7097 => x"d4",
          7098 => x"c0",
          7099 => x"dc",
          7100 => x"8c",
          7101 => x"38",
          7102 => x"05",
          7103 => x"06",
          7104 => x"73",
          7105 => x"16",
          7106 => x"22",
          7107 => x"07",
          7108 => x"1f",
          7109 => x"c2",
          7110 => x"81",
          7111 => x"34",
          7112 => x"b3",
          7113 => x"8c",
          7114 => x"74",
          7115 => x"0c",
          7116 => x"04",
          7117 => x"69",
          7118 => x"80",
          7119 => x"d0",
          7120 => x"3d",
          7121 => x"3f",
          7122 => x"08",
          7123 => x"08",
          7124 => x"8c",
          7125 => x"80",
          7126 => x"57",
          7127 => x"81",
          7128 => x"70",
          7129 => x"55",
          7130 => x"80",
          7131 => x"5d",
          7132 => x"52",
          7133 => x"52",
          7134 => x"a9",
          7135 => x"dc",
          7136 => x"8c",
          7137 => x"d1",
          7138 => x"73",
          7139 => x"3f",
          7140 => x"08",
          7141 => x"dc",
          7142 => x"82",
          7143 => x"82",
          7144 => x"65",
          7145 => x"78",
          7146 => x"7b",
          7147 => x"55",
          7148 => x"34",
          7149 => x"8a",
          7150 => x"38",
          7151 => x"1a",
          7152 => x"34",
          7153 => x"9e",
          7154 => x"70",
          7155 => x"51",
          7156 => x"a0",
          7157 => x"8e",
          7158 => x"2e",
          7159 => x"86",
          7160 => x"34",
          7161 => x"30",
          7162 => x"80",
          7163 => x"7a",
          7164 => x"c1",
          7165 => x"2e",
          7166 => x"a0",
          7167 => x"51",
          7168 => x"3f",
          7169 => x"08",
          7170 => x"dc",
          7171 => x"7b",
          7172 => x"55",
          7173 => x"73",
          7174 => x"38",
          7175 => x"73",
          7176 => x"38",
          7177 => x"15",
          7178 => x"ff",
          7179 => x"82",
          7180 => x"7b",
          7181 => x"8c",
          7182 => x"3d",
          7183 => x"3d",
          7184 => x"9c",
          7185 => x"05",
          7186 => x"51",
          7187 => x"82",
          7188 => x"82",
          7189 => x"56",
          7190 => x"dc",
          7191 => x"38",
          7192 => x"52",
          7193 => x"52",
          7194 => x"c0",
          7195 => x"70",
          7196 => x"ff",
          7197 => x"55",
          7198 => x"27",
          7199 => x"78",
          7200 => x"ff",
          7201 => x"05",
          7202 => x"55",
          7203 => x"3f",
          7204 => x"08",
          7205 => x"38",
          7206 => x"70",
          7207 => x"ff",
          7208 => x"82",
          7209 => x"80",
          7210 => x"74",
          7211 => x"07",
          7212 => x"4e",
          7213 => x"82",
          7214 => x"55",
          7215 => x"70",
          7216 => x"06",
          7217 => x"99",
          7218 => x"e0",
          7219 => x"ff",
          7220 => x"54",
          7221 => x"27",
          7222 => x"f9",
          7223 => x"55",
          7224 => x"a3",
          7225 => x"81",
          7226 => x"ff",
          7227 => x"82",
          7228 => x"93",
          7229 => x"75",
          7230 => x"76",
          7231 => x"38",
          7232 => x"77",
          7233 => x"86",
          7234 => x"39",
          7235 => x"27",
          7236 => x"88",
          7237 => x"78",
          7238 => x"5a",
          7239 => x"57",
          7240 => x"81",
          7241 => x"81",
          7242 => x"33",
          7243 => x"06",
          7244 => x"57",
          7245 => x"fe",
          7246 => x"3d",
          7247 => x"55",
          7248 => x"2e",
          7249 => x"76",
          7250 => x"38",
          7251 => x"55",
          7252 => x"33",
          7253 => x"a0",
          7254 => x"06",
          7255 => x"17",
          7256 => x"38",
          7257 => x"43",
          7258 => x"3d",
          7259 => x"ff",
          7260 => x"82",
          7261 => x"54",
          7262 => x"08",
          7263 => x"81",
          7264 => x"ff",
          7265 => x"82",
          7266 => x"54",
          7267 => x"08",
          7268 => x"80",
          7269 => x"54",
          7270 => x"80",
          7271 => x"8c",
          7272 => x"2e",
          7273 => x"80",
          7274 => x"54",
          7275 => x"80",
          7276 => x"52",
          7277 => x"bd",
          7278 => x"8c",
          7279 => x"82",
          7280 => x"b1",
          7281 => x"82",
          7282 => x"52",
          7283 => x"ab",
          7284 => x"54",
          7285 => x"15",
          7286 => x"78",
          7287 => x"ff",
          7288 => x"79",
          7289 => x"83",
          7290 => x"51",
          7291 => x"3f",
          7292 => x"08",
          7293 => x"74",
          7294 => x"0c",
          7295 => x"04",
          7296 => x"60",
          7297 => x"05",
          7298 => x"33",
          7299 => x"05",
          7300 => x"40",
          7301 => x"da",
          7302 => x"dc",
          7303 => x"8c",
          7304 => x"bd",
          7305 => x"33",
          7306 => x"b5",
          7307 => x"2e",
          7308 => x"1a",
          7309 => x"90",
          7310 => x"33",
          7311 => x"70",
          7312 => x"55",
          7313 => x"38",
          7314 => x"97",
          7315 => x"82",
          7316 => x"58",
          7317 => x"7e",
          7318 => x"70",
          7319 => x"55",
          7320 => x"56",
          7321 => x"f5",
          7322 => x"7d",
          7323 => x"70",
          7324 => x"2a",
          7325 => x"08",
          7326 => x"08",
          7327 => x"5d",
          7328 => x"77",
          7329 => x"98",
          7330 => x"26",
          7331 => x"57",
          7332 => x"59",
          7333 => x"52",
          7334 => x"ae",
          7335 => x"15",
          7336 => x"98",
          7337 => x"26",
          7338 => x"55",
          7339 => x"08",
          7340 => x"99",
          7341 => x"dc",
          7342 => x"ff",
          7343 => x"8c",
          7344 => x"38",
          7345 => x"75",
          7346 => x"81",
          7347 => x"93",
          7348 => x"80",
          7349 => x"2e",
          7350 => x"ff",
          7351 => x"58",
          7352 => x"7d",
          7353 => x"38",
          7354 => x"55",
          7355 => x"b4",
          7356 => x"56",
          7357 => x"09",
          7358 => x"38",
          7359 => x"53",
          7360 => x"51",
          7361 => x"3f",
          7362 => x"08",
          7363 => x"dc",
          7364 => x"38",
          7365 => x"ff",
          7366 => x"5c",
          7367 => x"84",
          7368 => x"5c",
          7369 => x"12",
          7370 => x"80",
          7371 => x"78",
          7372 => x"7c",
          7373 => x"90",
          7374 => x"c0",
          7375 => x"90",
          7376 => x"15",
          7377 => x"90",
          7378 => x"54",
          7379 => x"91",
          7380 => x"31",
          7381 => x"84",
          7382 => x"07",
          7383 => x"16",
          7384 => x"73",
          7385 => x"0c",
          7386 => x"04",
          7387 => x"6b",
          7388 => x"05",
          7389 => x"33",
          7390 => x"5a",
          7391 => x"bd",
          7392 => x"80",
          7393 => x"dc",
          7394 => x"f8",
          7395 => x"dc",
          7396 => x"82",
          7397 => x"70",
          7398 => x"74",
          7399 => x"38",
          7400 => x"82",
          7401 => x"81",
          7402 => x"81",
          7403 => x"ff",
          7404 => x"82",
          7405 => x"81",
          7406 => x"81",
          7407 => x"83",
          7408 => x"c0",
          7409 => x"2a",
          7410 => x"51",
          7411 => x"74",
          7412 => x"99",
          7413 => x"53",
          7414 => x"51",
          7415 => x"3f",
          7416 => x"08",
          7417 => x"55",
          7418 => x"92",
          7419 => x"80",
          7420 => x"38",
          7421 => x"06",
          7422 => x"2e",
          7423 => x"48",
          7424 => x"87",
          7425 => x"79",
          7426 => x"78",
          7427 => x"26",
          7428 => x"19",
          7429 => x"74",
          7430 => x"38",
          7431 => x"e4",
          7432 => x"2a",
          7433 => x"70",
          7434 => x"59",
          7435 => x"7a",
          7436 => x"56",
          7437 => x"80",
          7438 => x"51",
          7439 => x"74",
          7440 => x"99",
          7441 => x"53",
          7442 => x"51",
          7443 => x"3f",
          7444 => x"8c",
          7445 => x"ac",
          7446 => x"2a",
          7447 => x"82",
          7448 => x"43",
          7449 => x"83",
          7450 => x"66",
          7451 => x"60",
          7452 => x"90",
          7453 => x"31",
          7454 => x"80",
          7455 => x"8a",
          7456 => x"56",
          7457 => x"26",
          7458 => x"77",
          7459 => x"81",
          7460 => x"74",
          7461 => x"38",
          7462 => x"55",
          7463 => x"83",
          7464 => x"81",
          7465 => x"80",
          7466 => x"38",
          7467 => x"55",
          7468 => x"5e",
          7469 => x"89",
          7470 => x"5a",
          7471 => x"09",
          7472 => x"e1",
          7473 => x"38",
          7474 => x"57",
          7475 => x"fc",
          7476 => x"5a",
          7477 => x"9d",
          7478 => x"26",
          7479 => x"fc",
          7480 => x"10",
          7481 => x"22",
          7482 => x"74",
          7483 => x"38",
          7484 => x"ee",
          7485 => x"66",
          7486 => x"e1",
          7487 => x"dc",
          7488 => x"84",
          7489 => x"89",
          7490 => x"a0",
          7491 => x"82",
          7492 => x"fc",
          7493 => x"56",
          7494 => x"f0",
          7495 => x"80",
          7496 => x"d3",
          7497 => x"38",
          7498 => x"57",
          7499 => x"fc",
          7500 => x"5a",
          7501 => x"9d",
          7502 => x"26",
          7503 => x"fc",
          7504 => x"10",
          7505 => x"22",
          7506 => x"74",
          7507 => x"38",
          7508 => x"ee",
          7509 => x"66",
          7510 => x"81",
          7511 => x"dc",
          7512 => x"05",
          7513 => x"dc",
          7514 => x"26",
          7515 => x"0b",
          7516 => x"08",
          7517 => x"dc",
          7518 => x"11",
          7519 => x"05",
          7520 => x"83",
          7521 => x"2a",
          7522 => x"a0",
          7523 => x"7d",
          7524 => x"69",
          7525 => x"05",
          7526 => x"72",
          7527 => x"5c",
          7528 => x"59",
          7529 => x"2e",
          7530 => x"89",
          7531 => x"60",
          7532 => x"84",
          7533 => x"5d",
          7534 => x"18",
          7535 => x"68",
          7536 => x"74",
          7537 => x"af",
          7538 => x"31",
          7539 => x"53",
          7540 => x"52",
          7541 => x"85",
          7542 => x"dc",
          7543 => x"83",
          7544 => x"06",
          7545 => x"8c",
          7546 => x"ff",
          7547 => x"dd",
          7548 => x"83",
          7549 => x"2a",
          7550 => x"be",
          7551 => x"39",
          7552 => x"09",
          7553 => x"c5",
          7554 => x"f5",
          7555 => x"dc",
          7556 => x"38",
          7557 => x"79",
          7558 => x"80",
          7559 => x"38",
          7560 => x"96",
          7561 => x"06",
          7562 => x"2e",
          7563 => x"5e",
          7564 => x"82",
          7565 => x"9f",
          7566 => x"38",
          7567 => x"38",
          7568 => x"81",
          7569 => x"fc",
          7570 => x"ab",
          7571 => x"7d",
          7572 => x"81",
          7573 => x"7d",
          7574 => x"78",
          7575 => x"74",
          7576 => x"8e",
          7577 => x"9c",
          7578 => x"53",
          7579 => x"51",
          7580 => x"3f",
          7581 => x"fa",
          7582 => x"51",
          7583 => x"3f",
          7584 => x"8b",
          7585 => x"a1",
          7586 => x"8d",
          7587 => x"83",
          7588 => x"52",
          7589 => x"ff",
          7590 => x"81",
          7591 => x"34",
          7592 => x"70",
          7593 => x"2a",
          7594 => x"54",
          7595 => x"1b",
          7596 => x"88",
          7597 => x"74",
          7598 => x"26",
          7599 => x"83",
          7600 => x"52",
          7601 => x"ff",
          7602 => x"8a",
          7603 => x"a0",
          7604 => x"a1",
          7605 => x"0b",
          7606 => x"bf",
          7607 => x"51",
          7608 => x"3f",
          7609 => x"9a",
          7610 => x"a0",
          7611 => x"52",
          7612 => x"ff",
          7613 => x"7d",
          7614 => x"81",
          7615 => x"38",
          7616 => x"0a",
          7617 => x"1b",
          7618 => x"ce",
          7619 => x"a4",
          7620 => x"a0",
          7621 => x"52",
          7622 => x"ff",
          7623 => x"81",
          7624 => x"51",
          7625 => x"3f",
          7626 => x"1b",
          7627 => x"8c",
          7628 => x"0b",
          7629 => x"34",
          7630 => x"c2",
          7631 => x"53",
          7632 => x"52",
          7633 => x"51",
          7634 => x"88",
          7635 => x"a7",
          7636 => x"a0",
          7637 => x"83",
          7638 => x"52",
          7639 => x"ff",
          7640 => x"ff",
          7641 => x"1c",
          7642 => x"a6",
          7643 => x"53",
          7644 => x"52",
          7645 => x"ff",
          7646 => x"82",
          7647 => x"83",
          7648 => x"52",
          7649 => x"b4",
          7650 => x"60",
          7651 => x"7e",
          7652 => x"d7",
          7653 => x"82",
          7654 => x"83",
          7655 => x"83",
          7656 => x"06",
          7657 => x"75",
          7658 => x"05",
          7659 => x"7e",
          7660 => x"b7",
          7661 => x"53",
          7662 => x"51",
          7663 => x"3f",
          7664 => x"a4",
          7665 => x"51",
          7666 => x"3f",
          7667 => x"e4",
          7668 => x"e4",
          7669 => x"9f",
          7670 => x"18",
          7671 => x"1b",
          7672 => x"f6",
          7673 => x"83",
          7674 => x"ff",
          7675 => x"82",
          7676 => x"78",
          7677 => x"c4",
          7678 => x"60",
          7679 => x"7a",
          7680 => x"ff",
          7681 => x"75",
          7682 => x"53",
          7683 => x"51",
          7684 => x"3f",
          7685 => x"52",
          7686 => x"9f",
          7687 => x"56",
          7688 => x"83",
          7689 => x"06",
          7690 => x"52",
          7691 => x"9e",
          7692 => x"52",
          7693 => x"ff",
          7694 => x"f0",
          7695 => x"1b",
          7696 => x"87",
          7697 => x"55",
          7698 => x"83",
          7699 => x"74",
          7700 => x"ff",
          7701 => x"7c",
          7702 => x"74",
          7703 => x"38",
          7704 => x"54",
          7705 => x"52",
          7706 => x"99",
          7707 => x"8c",
          7708 => x"87",
          7709 => x"53",
          7710 => x"08",
          7711 => x"ff",
          7712 => x"76",
          7713 => x"31",
          7714 => x"cd",
          7715 => x"58",
          7716 => x"ff",
          7717 => x"55",
          7718 => x"83",
          7719 => x"61",
          7720 => x"26",
          7721 => x"57",
          7722 => x"53",
          7723 => x"51",
          7724 => x"3f",
          7725 => x"08",
          7726 => x"76",
          7727 => x"31",
          7728 => x"db",
          7729 => x"7d",
          7730 => x"38",
          7731 => x"83",
          7732 => x"8a",
          7733 => x"7d",
          7734 => x"38",
          7735 => x"81",
          7736 => x"80",
          7737 => x"80",
          7738 => x"7a",
          7739 => x"bc",
          7740 => x"d5",
          7741 => x"ff",
          7742 => x"83",
          7743 => x"77",
          7744 => x"0b",
          7745 => x"81",
          7746 => x"34",
          7747 => x"34",
          7748 => x"34",
          7749 => x"56",
          7750 => x"52",
          7751 => x"d8",
          7752 => x"0b",
          7753 => x"82",
          7754 => x"82",
          7755 => x"56",
          7756 => x"34",
          7757 => x"08",
          7758 => x"60",
          7759 => x"1b",
          7760 => x"96",
          7761 => x"83",
          7762 => x"ff",
          7763 => x"81",
          7764 => x"7a",
          7765 => x"ff",
          7766 => x"81",
          7767 => x"dc",
          7768 => x"80",
          7769 => x"7e",
          7770 => x"e3",
          7771 => x"82",
          7772 => x"90",
          7773 => x"8e",
          7774 => x"81",
          7775 => x"82",
          7776 => x"56",
          7777 => x"dc",
          7778 => x"0d",
          7779 => x"0d",
          7780 => x"59",
          7781 => x"ff",
          7782 => x"57",
          7783 => x"b4",
          7784 => x"f8",
          7785 => x"81",
          7786 => x"52",
          7787 => x"dc",
          7788 => x"2e",
          7789 => x"9c",
          7790 => x"33",
          7791 => x"2e",
          7792 => x"76",
          7793 => x"58",
          7794 => x"57",
          7795 => x"09",
          7796 => x"38",
          7797 => x"78",
          7798 => x"38",
          7799 => x"82",
          7800 => x"8d",
          7801 => x"f7",
          7802 => x"02",
          7803 => x"05",
          7804 => x"77",
          7805 => x"81",
          7806 => x"8d",
          7807 => x"e7",
          7808 => x"08",
          7809 => x"24",
          7810 => x"17",
          7811 => x"8c",
          7812 => x"77",
          7813 => x"16",
          7814 => x"25",
          7815 => x"3d",
          7816 => x"75",
          7817 => x"52",
          7818 => x"cb",
          7819 => x"76",
          7820 => x"70",
          7821 => x"2a",
          7822 => x"51",
          7823 => x"84",
          7824 => x"19",
          7825 => x"8b",
          7826 => x"f9",
          7827 => x"84",
          7828 => x"56",
          7829 => x"a7",
          7830 => x"fc",
          7831 => x"53",
          7832 => x"75",
          7833 => x"a1",
          7834 => x"dc",
          7835 => x"84",
          7836 => x"2e",
          7837 => x"87",
          7838 => x"08",
          7839 => x"ff",
          7840 => x"8c",
          7841 => x"3d",
          7842 => x"3d",
          7843 => x"80",
          7844 => x"52",
          7845 => x"9a",
          7846 => x"74",
          7847 => x"0d",
          7848 => x"0d",
          7849 => x"05",
          7850 => x"86",
          7851 => x"54",
          7852 => x"73",
          7853 => x"fe",
          7854 => x"51",
          7855 => x"98",
          7856 => x"f8",
          7857 => x"70",
          7858 => x"56",
          7859 => x"2e",
          7860 => x"8c",
          7861 => x"79",
          7862 => x"33",
          7863 => x"39",
          7864 => x"73",
          7865 => x"81",
          7866 => x"81",
          7867 => x"39",
          7868 => x"90",
          7869 => x"cc",
          7870 => x"52",
          7871 => x"f0",
          7872 => x"dc",
          7873 => x"dc",
          7874 => x"53",
          7875 => x"58",
          7876 => x"3f",
          7877 => x"08",
          7878 => x"16",
          7879 => x"81",
          7880 => x"38",
          7881 => x"81",
          7882 => x"54",
          7883 => x"c2",
          7884 => x"73",
          7885 => x"0c",
          7886 => x"04",
          7887 => x"73",
          7888 => x"26",
          7889 => x"71",
          7890 => x"f1",
          7891 => x"71",
          7892 => x"fd",
          7893 => x"80",
          7894 => x"d4",
          7895 => x"39",
          7896 => x"51",
          7897 => x"81",
          7898 => x"80",
          7899 => x"fe",
          7900 => x"e4",
          7901 => x"9c",
          7902 => x"39",
          7903 => x"51",
          7904 => x"81",
          7905 => x"80",
          7906 => x"fe",
          7907 => x"c8",
          7908 => x"f0",
          7909 => x"39",
          7910 => x"51",
          7911 => x"ff",
          7912 => x"39",
          7913 => x"51",
          7914 => x"ff",
          7915 => x"39",
          7916 => x"51",
          7917 => x"80",
          7918 => x"39",
          7919 => x"51",
          7920 => x"80",
          7921 => x"39",
          7922 => x"51",
          7923 => x"80",
          7924 => x"39",
          7925 => x"51",
          7926 => x"3f",
          7927 => x"04",
          7928 => x"77",
          7929 => x"74",
          7930 => x"8a",
          7931 => x"75",
          7932 => x"51",
          7933 => x"e8",
          7934 => x"fe",
          7935 => x"82",
          7936 => x"52",
          7937 => x"d2",
          7938 => x"8c",
          7939 => x"79",
          7940 => x"82",
          7941 => x"fe",
          7942 => x"87",
          7943 => x"ec",
          7944 => x"02",
          7945 => x"e3",
          7946 => x"57",
          7947 => x"30",
          7948 => x"73",
          7949 => x"59",
          7950 => x"77",
          7951 => x"83",
          7952 => x"74",
          7953 => x"81",
          7954 => x"55",
          7955 => x"81",
          7956 => x"53",
          7957 => x"3d",
          7958 => x"ff",
          7959 => x"82",
          7960 => x"57",
          7961 => x"08",
          7962 => x"8c",
          7963 => x"c0",
          7964 => x"82",
          7965 => x"59",
          7966 => x"05",
          7967 => x"53",
          7968 => x"51",
          7969 => x"82",
          7970 => x"57",
          7971 => x"08",
          7972 => x"55",
          7973 => x"89",
          7974 => x"75",
          7975 => x"d8",
          7976 => x"d8",
          7977 => x"f0",
          7978 => x"70",
          7979 => x"25",
          7980 => x"9f",
          7981 => x"51",
          7982 => x"74",
          7983 => x"38",
          7984 => x"53",
          7985 => x"88",
          7986 => x"51",
          7987 => x"76",
          7988 => x"8c",
          7989 => x"3d",
          7990 => x"3d",
          7991 => x"84",
          7992 => x"33",
          7993 => x"57",
          7994 => x"52",
          7995 => x"af",
          7996 => x"dc",
          7997 => x"75",
          7998 => x"38",
          7999 => x"98",
          8000 => x"60",
          8001 => x"82",
          8002 => x"7e",
          8003 => x"77",
          8004 => x"dc",
          8005 => x"39",
          8006 => x"82",
          8007 => x"89",
          8008 => x"f3",
          8009 => x"61",
          8010 => x"05",
          8011 => x"33",
          8012 => x"68",
          8013 => x"5c",
          8014 => x"7a",
          8015 => x"bc",
          8016 => x"a9",
          8017 => x"c4",
          8018 => x"bd",
          8019 => x"74",
          8020 => x"fc",
          8021 => x"2e",
          8022 => x"a0",
          8023 => x"80",
          8024 => x"18",
          8025 => x"27",
          8026 => x"22",
          8027 => x"c8",
          8028 => x"f9",
          8029 => x"82",
          8030 => x"fe",
          8031 => x"82",
          8032 => x"c3",
          8033 => x"53",
          8034 => x"8e",
          8035 => x"52",
          8036 => x"51",
          8037 => x"3f",
          8038 => x"81",
          8039 => x"ee",
          8040 => x"15",
          8041 => x"74",
          8042 => x"7a",
          8043 => x"72",
          8044 => x"81",
          8045 => x"f4",
          8046 => x"39",
          8047 => x"51",
          8048 => x"3f",
          8049 => x"a0",
          8050 => x"e0",
          8051 => x"39",
          8052 => x"51",
          8053 => x"3f",
          8054 => x"79",
          8055 => x"74",
          8056 => x"55",
          8057 => x"72",
          8058 => x"38",
          8059 => x"53",
          8060 => x"83",
          8061 => x"75",
          8062 => x"81",
          8063 => x"53",
          8064 => x"8b",
          8065 => x"fe",
          8066 => x"73",
          8067 => x"a0",
          8068 => x"98",
          8069 => x"55",
          8070 => x"81",
          8071 => x"ed",
          8072 => x"18",
          8073 => x"58",
          8074 => x"3f",
          8075 => x"08",
          8076 => x"98",
          8077 => x"76",
          8078 => x"81",
          8079 => x"fe",
          8080 => x"82",
          8081 => x"98",
          8082 => x"2c",
          8083 => x"70",
          8084 => x"32",
          8085 => x"72",
          8086 => x"07",
          8087 => x"58",
          8088 => x"57",
          8089 => x"d7",
          8090 => x"2e",
          8091 => x"85",
          8092 => x"8c",
          8093 => x"53",
          8094 => x"fd",
          8095 => x"53",
          8096 => x"dc",
          8097 => x"0d",
          8098 => x"0d",
          8099 => x"33",
          8100 => x"53",
          8101 => x"52",
          8102 => x"d1",
          8103 => x"8c",
          8104 => x"e7",
          8105 => x"82",
          8106 => x"82",
          8107 => x"88",
          8108 => x"82",
          8109 => x"fe",
          8110 => x"74",
          8111 => x"38",
          8112 => x"3f",
          8113 => x"04",
          8114 => x"87",
          8115 => x"08",
          8116 => x"b1",
          8117 => x"fe",
          8118 => x"82",
          8119 => x"fe",
          8120 => x"80",
          8121 => x"ac",
          8122 => x"2a",
          8123 => x"51",
          8124 => x"2e",
          8125 => x"51",
          8126 => x"3f",
          8127 => x"51",
          8128 => x"3f",
          8129 => x"d9",
          8130 => x"82",
          8131 => x"06",
          8132 => x"80",
          8133 => x"81",
          8134 => x"f8",
          8135 => x"dc",
          8136 => x"f0",
          8137 => x"fe",
          8138 => x"72",
          8139 => x"81",
          8140 => x"71",
          8141 => x"38",
          8142 => x"d8",
          8143 => x"82",
          8144 => x"da",
          8145 => x"51",
          8146 => x"3f",
          8147 => x"70",
          8148 => x"52",
          8149 => x"95",
          8150 => x"fe",
          8151 => x"82",
          8152 => x"fe",
          8153 => x"80",
          8154 => x"a8",
          8155 => x"2a",
          8156 => x"51",
          8157 => x"2e",
          8158 => x"51",
          8159 => x"3f",
          8160 => x"51",
          8161 => x"3f",
          8162 => x"d8",
          8163 => x"86",
          8164 => x"06",
          8165 => x"80",
          8166 => x"81",
          8167 => x"f4",
          8168 => x"a8",
          8169 => x"ec",
          8170 => x"fe",
          8171 => x"72",
          8172 => x"81",
          8173 => x"71",
          8174 => x"38",
          8175 => x"d7",
          8176 => x"83",
          8177 => x"d9",
          8178 => x"51",
          8179 => x"3f",
          8180 => x"70",
          8181 => x"52",
          8182 => x"95",
          8183 => x"fe",
          8184 => x"82",
          8185 => x"fe",
          8186 => x"80",
          8187 => x"a4",
          8188 => x"99",
          8189 => x"0d",
          8190 => x"0d",
          8191 => x"05",
          8192 => x"70",
          8193 => x"80",
          8194 => x"fe",
          8195 => x"82",
          8196 => x"54",
          8197 => x"81",
          8198 => x"90",
          8199 => x"f4",
          8200 => x"83",
          8201 => x"dc",
          8202 => x"82",
          8203 => x"07",
          8204 => x"71",
          8205 => x"54",
          8206 => x"c8",
          8207 => x"c8",
          8208 => x"81",
          8209 => x"06",
          8210 => x"a3",
          8211 => x"52",
          8212 => x"b9",
          8213 => x"dc",
          8214 => x"8c",
          8215 => x"dc",
          8216 => x"e9",
          8217 => x"39",
          8218 => x"51",
          8219 => x"82",
          8220 => x"c8",
          8221 => x"c8",
          8222 => x"82",
          8223 => x"06",
          8224 => x"52",
          8225 => x"fa",
          8226 => x"0b",
          8227 => x"0c",
          8228 => x"04",
          8229 => x"80",
          8230 => x"a3",
          8231 => x"5d",
          8232 => x"51",
          8233 => x"3f",
          8234 => x"08",
          8235 => x"59",
          8236 => x"09",
          8237 => x"38",
          8238 => x"52",
          8239 => x"52",
          8240 => x"bf",
          8241 => x"78",
          8242 => x"a0",
          8243 => x"f6",
          8244 => x"dc",
          8245 => x"88",
          8246 => x"a4",
          8247 => x"39",
          8248 => x"5d",
          8249 => x"51",
          8250 => x"3f",
          8251 => x"46",
          8252 => x"52",
          8253 => x"81",
          8254 => x"ff",
          8255 => x"f3",
          8256 => x"8c",
          8257 => x"2b",
          8258 => x"51",
          8259 => x"c2",
          8260 => x"38",
          8261 => x"24",
          8262 => x"bd",
          8263 => x"38",
          8264 => x"90",
          8265 => x"2e",
          8266 => x"78",
          8267 => x"da",
          8268 => x"39",
          8269 => x"2e",
          8270 => x"78",
          8271 => x"85",
          8272 => x"bf",
          8273 => x"38",
          8274 => x"78",
          8275 => x"89",
          8276 => x"80",
          8277 => x"38",
          8278 => x"2e",
          8279 => x"78",
          8280 => x"89",
          8281 => x"b4",
          8282 => x"83",
          8283 => x"38",
          8284 => x"24",
          8285 => x"81",
          8286 => x"fd",
          8287 => x"39",
          8288 => x"2e",
          8289 => x"8a",
          8290 => x"3d",
          8291 => x"53",
          8292 => x"51",
          8293 => x"3f",
          8294 => x"08",
          8295 => x"c4",
          8296 => x"fe",
          8297 => x"ff",
          8298 => x"fe",
          8299 => x"82",
          8300 => x"80",
          8301 => x"38",
          8302 => x"f8",
          8303 => x"84",
          8304 => x"ee",
          8305 => x"8c",
          8306 => x"38",
          8307 => x"08",
          8308 => x"e0",
          8309 => x"b1",
          8310 => x"5c",
          8311 => x"27",
          8312 => x"61",
          8313 => x"70",
          8314 => x"0c",
          8315 => x"f5",
          8316 => x"39",
          8317 => x"80",
          8318 => x"84",
          8319 => x"ed",
          8320 => x"8c",
          8321 => x"2e",
          8322 => x"b4",
          8323 => x"11",
          8324 => x"05",
          8325 => x"ca",
          8326 => x"dc",
          8327 => x"fd",
          8328 => x"3d",
          8329 => x"53",
          8330 => x"51",
          8331 => x"3f",
          8332 => x"08",
          8333 => x"ac",
          8334 => x"f0",
          8335 => x"c9",
          8336 => x"79",
          8337 => x"8c",
          8338 => x"79",
          8339 => x"5b",
          8340 => x"61",
          8341 => x"eb",
          8342 => x"ff",
          8343 => x"ff",
          8344 => x"fe",
          8345 => x"82",
          8346 => x"80",
          8347 => x"38",
          8348 => x"fc",
          8349 => x"84",
          8350 => x"ec",
          8351 => x"8c",
          8352 => x"2e",
          8353 => x"b4",
          8354 => x"11",
          8355 => x"05",
          8356 => x"ce",
          8357 => x"dc",
          8358 => x"fc",
          8359 => x"84",
          8360 => x"e4",
          8361 => x"5a",
          8362 => x"a8",
          8363 => x"33",
          8364 => x"5a",
          8365 => x"2e",
          8366 => x"55",
          8367 => x"33",
          8368 => x"82",
          8369 => x"fe",
          8370 => x"81",
          8371 => x"05",
          8372 => x"39",
          8373 => x"51",
          8374 => x"b4",
          8375 => x"11",
          8376 => x"05",
          8377 => x"fa",
          8378 => x"dc",
          8379 => x"38",
          8380 => x"33",
          8381 => x"2e",
          8382 => x"87",
          8383 => x"80",
          8384 => x"88",
          8385 => x"78",
          8386 => x"38",
          8387 => x"08",
          8388 => x"82",
          8389 => x"59",
          8390 => x"88",
          8391 => x"e8",
          8392 => x"39",
          8393 => x"33",
          8394 => x"2e",
          8395 => x"87",
          8396 => x"9a",
          8397 => x"9e",
          8398 => x"80",
          8399 => x"82",
          8400 => x"44",
          8401 => x"88",
          8402 => x"80",
          8403 => x"3d",
          8404 => x"53",
          8405 => x"51",
          8406 => x"3f",
          8407 => x"08",
          8408 => x"82",
          8409 => x"59",
          8410 => x"89",
          8411 => x"dc",
          8412 => x"cc",
          8413 => x"a1",
          8414 => x"80",
          8415 => x"82",
          8416 => x"43",
          8417 => x"88",
          8418 => x"78",
          8419 => x"38",
          8420 => x"08",
          8421 => x"82",
          8422 => x"59",
          8423 => x"88",
          8424 => x"f4",
          8425 => x"39",
          8426 => x"33",
          8427 => x"2e",
          8428 => x"87",
          8429 => x"88",
          8430 => x"88",
          8431 => x"43",
          8432 => x"f8",
          8433 => x"84",
          8434 => x"ea",
          8435 => x"8c",
          8436 => x"2e",
          8437 => x"62",
          8438 => x"88",
          8439 => x"81",
          8440 => x"32",
          8441 => x"72",
          8442 => x"70",
          8443 => x"51",
          8444 => x"80",
          8445 => x"7a",
          8446 => x"38",
          8447 => x"85",
          8448 => x"e2",
          8449 => x"55",
          8450 => x"53",
          8451 => x"51",
          8452 => x"82",
          8453 => x"fe",
          8454 => x"f9",
          8455 => x"3d",
          8456 => x"53",
          8457 => x"51",
          8458 => x"3f",
          8459 => x"08",
          8460 => x"b0",
          8461 => x"fe",
          8462 => x"ff",
          8463 => x"fe",
          8464 => x"82",
          8465 => x"80",
          8466 => x"63",
          8467 => x"cb",
          8468 => x"34",
          8469 => x"44",
          8470 => x"fc",
          8471 => x"84",
          8472 => x"e8",
          8473 => x"8c",
          8474 => x"38",
          8475 => x"63",
          8476 => x"52",
          8477 => x"51",
          8478 => x"3f",
          8479 => x"79",
          8480 => x"c3",
          8481 => x"79",
          8482 => x"ae",
          8483 => x"38",
          8484 => x"a0",
          8485 => x"fe",
          8486 => x"ff",
          8487 => x"fe",
          8488 => x"82",
          8489 => x"80",
          8490 => x"63",
          8491 => x"cb",
          8492 => x"34",
          8493 => x"44",
          8494 => x"82",
          8495 => x"fe",
          8496 => x"ff",
          8497 => x"3d",
          8498 => x"53",
          8499 => x"51",
          8500 => x"3f",
          8501 => x"08",
          8502 => x"88",
          8503 => x"fe",
          8504 => x"ff",
          8505 => x"fe",
          8506 => x"82",
          8507 => x"80",
          8508 => x"60",
          8509 => x"05",
          8510 => x"82",
          8511 => x"78",
          8512 => x"fe",
          8513 => x"ff",
          8514 => x"fe",
          8515 => x"82",
          8516 => x"df",
          8517 => x"39",
          8518 => x"54",
          8519 => x"d8",
          8520 => x"c9",
          8521 => x"52",
          8522 => x"e6",
          8523 => x"45",
          8524 => x"78",
          8525 => x"ac",
          8526 => x"26",
          8527 => x"82",
          8528 => x"39",
          8529 => x"f0",
          8530 => x"84",
          8531 => x"e9",
          8532 => x"8c",
          8533 => x"2e",
          8534 => x"59",
          8535 => x"22",
          8536 => x"05",
          8537 => x"41",
          8538 => x"82",
          8539 => x"fe",
          8540 => x"ff",
          8541 => x"3d",
          8542 => x"53",
          8543 => x"51",
          8544 => x"3f",
          8545 => x"08",
          8546 => x"d8",
          8547 => x"fe",
          8548 => x"ff",
          8549 => x"fe",
          8550 => x"82",
          8551 => x"80",
          8552 => x"60",
          8553 => x"59",
          8554 => x"41",
          8555 => x"f0",
          8556 => x"84",
          8557 => x"e8",
          8558 => x"8c",
          8559 => x"38",
          8560 => x"60",
          8561 => x"52",
          8562 => x"51",
          8563 => x"3f",
          8564 => x"79",
          8565 => x"ef",
          8566 => x"79",
          8567 => x"ae",
          8568 => x"38",
          8569 => x"9c",
          8570 => x"fe",
          8571 => x"ff",
          8572 => x"fe",
          8573 => x"82",
          8574 => x"80",
          8575 => x"60",
          8576 => x"59",
          8577 => x"41",
          8578 => x"82",
          8579 => x"fe",
          8580 => x"ff",
          8581 => x"3d",
          8582 => x"53",
          8583 => x"51",
          8584 => x"3f",
          8585 => x"08",
          8586 => x"b8",
          8587 => x"82",
          8588 => x"fe",
          8589 => x"63",
          8590 => x"b4",
          8591 => x"11",
          8592 => x"05",
          8593 => x"9a",
          8594 => x"dc",
          8595 => x"f5",
          8596 => x"52",
          8597 => x"51",
          8598 => x"3f",
          8599 => x"2d",
          8600 => x"08",
          8601 => x"fc",
          8602 => x"dc",
          8603 => x"86",
          8604 => x"e2",
          8605 => x"ec",
          8606 => x"c4",
          8607 => x"89",
          8608 => x"b9",
          8609 => x"39",
          8610 => x"51",
          8611 => x"3f",
          8612 => x"a5",
          8613 => x"8c",
          8614 => x"39",
          8615 => x"33",
          8616 => x"2e",
          8617 => x"7d",
          8618 => x"78",
          8619 => x"d3",
          8620 => x"ff",
          8621 => x"fe",
          8622 => x"82",
          8623 => x"5c",
          8624 => x"82",
          8625 => x"7a",
          8626 => x"38",
          8627 => x"8c",
          8628 => x"39",
          8629 => x"b0",
          8630 => x"39",
          8631 => x"56",
          8632 => x"86",
          8633 => x"53",
          8634 => x"52",
          8635 => x"b0",
          8636 => x"e2",
          8637 => x"39",
          8638 => x"52",
          8639 => x"b0",
          8640 => x"e1",
          8641 => x"39",
          8642 => x"86",
          8643 => x"53",
          8644 => x"52",
          8645 => x"b0",
          8646 => x"e1",
          8647 => x"39",
          8648 => x"53",
          8649 => x"52",
          8650 => x"b0",
          8651 => x"e1",
          8652 => x"87",
          8653 => x"8d",
          8654 => x"56",
          8655 => x"54",
          8656 => x"53",
          8657 => x"52",
          8658 => x"b0",
          8659 => x"8a",
          8660 => x"dc",
          8661 => x"dc",
          8662 => x"30",
          8663 => x"80",
          8664 => x"5b",
          8665 => x"7a",
          8666 => x"38",
          8667 => x"7a",
          8668 => x"80",
          8669 => x"81",
          8670 => x"ff",
          8671 => x"7a",
          8672 => x"7d",
          8673 => x"81",
          8674 => x"78",
          8675 => x"ff",
          8676 => x"06",
          8677 => x"82",
          8678 => x"fe",
          8679 => x"f2",
          8680 => x"3d",
          8681 => x"82",
          8682 => x"87",
          8683 => x"70",
          8684 => x"87",
          8685 => x"72",
          8686 => x"a1",
          8687 => x"dc",
          8688 => x"75",
          8689 => x"87",
          8690 => x"73",
          8691 => x"8d",
          8692 => x"8c",
          8693 => x"75",
          8694 => x"94",
          8695 => x"54",
          8696 => x"80",
          8697 => x"fe",
          8698 => x"82",
          8699 => x"90",
          8700 => x"55",
          8701 => x"80",
          8702 => x"fe",
          8703 => x"72",
          8704 => x"08",
          8705 => x"8c",
          8706 => x"87",
          8707 => x"0c",
          8708 => x"0b",
          8709 => x"94",
          8710 => x"0b",
          8711 => x"0c",
          8712 => x"82",
          8713 => x"fe",
          8714 => x"fe",
          8715 => x"82",
          8716 => x"fe",
          8717 => x"82",
          8718 => x"fe",
          8719 => x"81",
          8720 => x"fe",
          8721 => x"81",
          8722 => x"3f",
          8723 => x"80",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"64",
          8762 => x"2f",
          8763 => x"25",
          8764 => x"64",
          8765 => x"2e",
          8766 => x"64",
          8767 => x"6f",
          8768 => x"6f",
          8769 => x"67",
          8770 => x"74",
          8771 => x"00",
          8772 => x"28",
          8773 => x"6d",
          8774 => x"43",
          8775 => x"6e",
          8776 => x"29",
          8777 => x"0a",
          8778 => x"69",
          8779 => x"20",
          8780 => x"6c",
          8781 => x"6e",
          8782 => x"3a",
          8783 => x"20",
          8784 => x"42",
          8785 => x"52",
          8786 => x"20",
          8787 => x"38",
          8788 => x"30",
          8789 => x"2e",
          8790 => x"20",
          8791 => x"44",
          8792 => x"20",
          8793 => x"20",
          8794 => x"38",
          8795 => x"30",
          8796 => x"2e",
          8797 => x"20",
          8798 => x"4e",
          8799 => x"42",
          8800 => x"20",
          8801 => x"38",
          8802 => x"30",
          8803 => x"2e",
          8804 => x"20",
          8805 => x"52",
          8806 => x"20",
          8807 => x"20",
          8808 => x"38",
          8809 => x"30",
          8810 => x"2e",
          8811 => x"20",
          8812 => x"41",
          8813 => x"20",
          8814 => x"20",
          8815 => x"38",
          8816 => x"30",
          8817 => x"2e",
          8818 => x"20",
          8819 => x"44",
          8820 => x"52",
          8821 => x"20",
          8822 => x"76",
          8823 => x"73",
          8824 => x"30",
          8825 => x"2e",
          8826 => x"20",
          8827 => x"49",
          8828 => x"31",
          8829 => x"20",
          8830 => x"6d",
          8831 => x"20",
          8832 => x"30",
          8833 => x"2e",
          8834 => x"20",
          8835 => x"4e",
          8836 => x"43",
          8837 => x"20",
          8838 => x"61",
          8839 => x"6c",
          8840 => x"30",
          8841 => x"2e",
          8842 => x"20",
          8843 => x"49",
          8844 => x"4f",
          8845 => x"42",
          8846 => x"00",
          8847 => x"20",
          8848 => x"42",
          8849 => x"43",
          8850 => x"20",
          8851 => x"4f",
          8852 => x"0a",
          8853 => x"20",
          8854 => x"53",
          8855 => x"00",
          8856 => x"20",
          8857 => x"50",
          8858 => x"00",
          8859 => x"64",
          8860 => x"73",
          8861 => x"3a",
          8862 => x"20",
          8863 => x"50",
          8864 => x"65",
          8865 => x"20",
          8866 => x"74",
          8867 => x"41",
          8868 => x"65",
          8869 => x"3d",
          8870 => x"38",
          8871 => x"00",
          8872 => x"20",
          8873 => x"50",
          8874 => x"65",
          8875 => x"79",
          8876 => x"61",
          8877 => x"41",
          8878 => x"65",
          8879 => x"3d",
          8880 => x"38",
          8881 => x"00",
          8882 => x"20",
          8883 => x"74",
          8884 => x"20",
          8885 => x"72",
          8886 => x"64",
          8887 => x"73",
          8888 => x"20",
          8889 => x"3d",
          8890 => x"38",
          8891 => x"00",
          8892 => x"69",
          8893 => x"0a",
          8894 => x"20",
          8895 => x"50",
          8896 => x"64",
          8897 => x"20",
          8898 => x"20",
          8899 => x"20",
          8900 => x"20",
          8901 => x"3d",
          8902 => x"34",
          8903 => x"00",
          8904 => x"20",
          8905 => x"79",
          8906 => x"6d",
          8907 => x"6f",
          8908 => x"46",
          8909 => x"20",
          8910 => x"20",
          8911 => x"3d",
          8912 => x"2e",
          8913 => x"64",
          8914 => x"0a",
          8915 => x"20",
          8916 => x"44",
          8917 => x"20",
          8918 => x"63",
          8919 => x"72",
          8920 => x"20",
          8921 => x"20",
          8922 => x"3d",
          8923 => x"2e",
          8924 => x"64",
          8925 => x"0a",
          8926 => x"20",
          8927 => x"69",
          8928 => x"6f",
          8929 => x"53",
          8930 => x"4d",
          8931 => x"6f",
          8932 => x"46",
          8933 => x"3d",
          8934 => x"2e",
          8935 => x"64",
          8936 => x"0a",
          8937 => x"6d",
          8938 => x"00",
          8939 => x"65",
          8940 => x"6d",
          8941 => x"6c",
          8942 => x"00",
          8943 => x"56",
          8944 => x"56",
          8945 => x"6e",
          8946 => x"6e",
          8947 => x"77",
          8948 => x"69",
          8949 => x"72",
          8950 => x"78",
          8951 => x"69",
          8952 => x"72",
          8953 => x"69",
          8954 => x"00",
          8955 => x"00",
          8956 => x"30",
          8957 => x"20",
          8958 => x"00",
          8959 => x"61",
          8960 => x"64",
          8961 => x"20",
          8962 => x"65",
          8963 => x"68",
          8964 => x"69",
          8965 => x"72",
          8966 => x"69",
          8967 => x"74",
          8968 => x"4f",
          8969 => x"00",
          8970 => x"61",
          8971 => x"74",
          8972 => x"65",
          8973 => x"72",
          8974 => x"65",
          8975 => x"73",
          8976 => x"79",
          8977 => x"6c",
          8978 => x"64",
          8979 => x"62",
          8980 => x"67",
          8981 => x"00",
          8982 => x"00",
          8983 => x"00",
          8984 => x"00",
          8985 => x"00",
          8986 => x"00",
          8987 => x"00",
          8988 => x"00",
          8989 => x"00",
          8990 => x"00",
          8991 => x"00",
          8992 => x"00",
          8993 => x"00",
          8994 => x"00",
          8995 => x"00",
          8996 => x"00",
          8997 => x"00",
          8998 => x"00",
          8999 => x"00",
          9000 => x"00",
          9001 => x"00",
          9002 => x"00",
          9003 => x"00",
          9004 => x"00",
          9005 => x"00",
          9006 => x"00",
          9007 => x"00",
          9008 => x"00",
          9009 => x"00",
          9010 => x"00",
          9011 => x"00",
          9012 => x"00",
          9013 => x"00",
          9014 => x"00",
          9015 => x"5b",
          9016 => x"5b",
          9017 => x"5b",
          9018 => x"5b",
          9019 => x"5b",
          9020 => x"5b",
          9021 => x"5b",
          9022 => x"5b",
          9023 => x"5b",
          9024 => x"00",
          9025 => x"00",
          9026 => x"44",
          9027 => x"2a",
          9028 => x"3b",
          9029 => x"3f",
          9030 => x"7f",
          9031 => x"41",
          9032 => x"41",
          9033 => x"00",
          9034 => x"fe",
          9035 => x"44",
          9036 => x"2e",
          9037 => x"4f",
          9038 => x"4d",
          9039 => x"20",
          9040 => x"54",
          9041 => x"20",
          9042 => x"4f",
          9043 => x"4d",
          9044 => x"20",
          9045 => x"54",
          9046 => x"20",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"9a",
          9052 => x"41",
          9053 => x"45",
          9054 => x"49",
          9055 => x"92",
          9056 => x"4f",
          9057 => x"99",
          9058 => x"9d",
          9059 => x"49",
          9060 => x"a5",
          9061 => x"a9",
          9062 => x"ad",
          9063 => x"b1",
          9064 => x"b5",
          9065 => x"b9",
          9066 => x"bd",
          9067 => x"c1",
          9068 => x"c5",
          9069 => x"c9",
          9070 => x"cd",
          9071 => x"d1",
          9072 => x"d5",
          9073 => x"d9",
          9074 => x"dd",
          9075 => x"e1",
          9076 => x"e5",
          9077 => x"e9",
          9078 => x"ed",
          9079 => x"f1",
          9080 => x"f5",
          9081 => x"f9",
          9082 => x"fd",
          9083 => x"2e",
          9084 => x"5b",
          9085 => x"22",
          9086 => x"3e",
          9087 => x"00",
          9088 => x"01",
          9089 => x"10",
          9090 => x"00",
          9091 => x"00",
          9092 => x"01",
          9093 => x"04",
          9094 => x"10",
          9095 => x"00",
          9096 => x"69",
          9097 => x"00",
          9098 => x"69",
          9099 => x"6c",
          9100 => x"69",
          9101 => x"00",
          9102 => x"6c",
          9103 => x"00",
          9104 => x"65",
          9105 => x"00",
          9106 => x"63",
          9107 => x"72",
          9108 => x"63",
          9109 => x"00",
          9110 => x"64",
          9111 => x"00",
          9112 => x"64",
          9113 => x"00",
          9114 => x"65",
          9115 => x"65",
          9116 => x"65",
          9117 => x"69",
          9118 => x"69",
          9119 => x"66",
          9120 => x"66",
          9121 => x"61",
          9122 => x"00",
          9123 => x"6d",
          9124 => x"65",
          9125 => x"72",
          9126 => x"65",
          9127 => x"00",
          9128 => x"6e",
          9129 => x"00",
          9130 => x"65",
          9131 => x"00",
          9132 => x"62",
          9133 => x"63",
          9134 => x"62",
          9135 => x"63",
          9136 => x"69",
          9137 => x"00",
          9138 => x"69",
          9139 => x"45",
          9140 => x"72",
          9141 => x"6e",
          9142 => x"6e",
          9143 => x"65",
          9144 => x"72",
          9145 => x"00",
          9146 => x"69",
          9147 => x"6e",
          9148 => x"72",
          9149 => x"79",
          9150 => x"00",
          9151 => x"6f",
          9152 => x"6c",
          9153 => x"6f",
          9154 => x"2e",
          9155 => x"6f",
          9156 => x"74",
          9157 => x"6f",
          9158 => x"2e",
          9159 => x"6e",
          9160 => x"69",
          9161 => x"69",
          9162 => x"61",
          9163 => x"0a",
          9164 => x"63",
          9165 => x"73",
          9166 => x"6e",
          9167 => x"2e",
          9168 => x"69",
          9169 => x"61",
          9170 => x"61",
          9171 => x"65",
          9172 => x"74",
          9173 => x"00",
          9174 => x"69",
          9175 => x"68",
          9176 => x"6c",
          9177 => x"6e",
          9178 => x"69",
          9179 => x"00",
          9180 => x"44",
          9181 => x"20",
          9182 => x"74",
          9183 => x"72",
          9184 => x"63",
          9185 => x"2e",
          9186 => x"72",
          9187 => x"20",
          9188 => x"62",
          9189 => x"69",
          9190 => x"6e",
          9191 => x"69",
          9192 => x"00",
          9193 => x"69",
          9194 => x"6e",
          9195 => x"65",
          9196 => x"6c",
          9197 => x"0a",
          9198 => x"6f",
          9199 => x"6d",
          9200 => x"69",
          9201 => x"20",
          9202 => x"65",
          9203 => x"74",
          9204 => x"66",
          9205 => x"64",
          9206 => x"20",
          9207 => x"6b",
          9208 => x"00",
          9209 => x"6f",
          9210 => x"74",
          9211 => x"6f",
          9212 => x"64",
          9213 => x"00",
          9214 => x"69",
          9215 => x"75",
          9216 => x"6f",
          9217 => x"61",
          9218 => x"6e",
          9219 => x"6e",
          9220 => x"6c",
          9221 => x"0a",
          9222 => x"69",
          9223 => x"69",
          9224 => x"6f",
          9225 => x"64",
          9226 => x"00",
          9227 => x"6e",
          9228 => x"66",
          9229 => x"65",
          9230 => x"6d",
          9231 => x"72",
          9232 => x"00",
          9233 => x"6f",
          9234 => x"61",
          9235 => x"6f",
          9236 => x"20",
          9237 => x"65",
          9238 => x"00",
          9239 => x"61",
          9240 => x"65",
          9241 => x"73",
          9242 => x"63",
          9243 => x"65",
          9244 => x"0a",
          9245 => x"75",
          9246 => x"73",
          9247 => x"00",
          9248 => x"6e",
          9249 => x"77",
          9250 => x"72",
          9251 => x"2e",
          9252 => x"25",
          9253 => x"62",
          9254 => x"73",
          9255 => x"20",
          9256 => x"25",
          9257 => x"62",
          9258 => x"73",
          9259 => x"63",
          9260 => x"00",
          9261 => x"65",
          9262 => x"00",
          9263 => x"30",
          9264 => x"00",
          9265 => x"20",
          9266 => x"30",
          9267 => x"00",
          9268 => x"20",
          9269 => x"20",
          9270 => x"00",
          9271 => x"30",
          9272 => x"00",
          9273 => x"20",
          9274 => x"7c",
          9275 => x"0d",
          9276 => x"4f",
          9277 => x"2a",
          9278 => x"73",
          9279 => x"00",
          9280 => x"37",
          9281 => x"2f",
          9282 => x"30",
          9283 => x"31",
          9284 => x"00",
          9285 => x"5a",
          9286 => x"20",
          9287 => x"20",
          9288 => x"78",
          9289 => x"73",
          9290 => x"20",
          9291 => x"0a",
          9292 => x"50",
          9293 => x"6e",
          9294 => x"72",
          9295 => x"20",
          9296 => x"64",
          9297 => x"0a",
          9298 => x"69",
          9299 => x"20",
          9300 => x"65",
          9301 => x"70",
          9302 => x"00",
          9303 => x"53",
          9304 => x"6e",
          9305 => x"72",
          9306 => x"0a",
          9307 => x"4f",
          9308 => x"20",
          9309 => x"69",
          9310 => x"72",
          9311 => x"74",
          9312 => x"4f",
          9313 => x"20",
          9314 => x"69",
          9315 => x"72",
          9316 => x"74",
          9317 => x"41",
          9318 => x"20",
          9319 => x"69",
          9320 => x"72",
          9321 => x"74",
          9322 => x"41",
          9323 => x"20",
          9324 => x"69",
          9325 => x"72",
          9326 => x"74",
          9327 => x"41",
          9328 => x"20",
          9329 => x"69",
          9330 => x"72",
          9331 => x"74",
          9332 => x"41",
          9333 => x"20",
          9334 => x"69",
          9335 => x"72",
          9336 => x"74",
          9337 => x"65",
          9338 => x"6e",
          9339 => x"70",
          9340 => x"6d",
          9341 => x"2e",
          9342 => x"00",
          9343 => x"6e",
          9344 => x"69",
          9345 => x"74",
          9346 => x"72",
          9347 => x"0a",
          9348 => x"75",
          9349 => x"78",
          9350 => x"62",
          9351 => x"00",
          9352 => x"3a",
          9353 => x"61",
          9354 => x"64",
          9355 => x"20",
          9356 => x"74",
          9357 => x"69",
          9358 => x"73",
          9359 => x"61",
          9360 => x"30",
          9361 => x"6c",
          9362 => x"65",
          9363 => x"69",
          9364 => x"61",
          9365 => x"6c",
          9366 => x"0a",
          9367 => x"20",
          9368 => x"6c",
          9369 => x"69",
          9370 => x"2e",
          9371 => x"00",
          9372 => x"6f",
          9373 => x"6e",
          9374 => x"2e",
          9375 => x"6f",
          9376 => x"72",
          9377 => x"2e",
          9378 => x"00",
          9379 => x"30",
          9380 => x"28",
          9381 => x"78",
          9382 => x"25",
          9383 => x"78",
          9384 => x"38",
          9385 => x"00",
          9386 => x"75",
          9387 => x"4d",
          9388 => x"72",
          9389 => x"00",
          9390 => x"43",
          9391 => x"6c",
          9392 => x"2e",
          9393 => x"30",
          9394 => x"25",
          9395 => x"2d",
          9396 => x"3f",
          9397 => x"00",
          9398 => x"30",
          9399 => x"25",
          9400 => x"2d",
          9401 => x"30",
          9402 => x"25",
          9403 => x"2d",
          9404 => x"78",
          9405 => x"74",
          9406 => x"20",
          9407 => x"65",
          9408 => x"25",
          9409 => x"20",
          9410 => x"0a",
          9411 => x"61",
          9412 => x"6e",
          9413 => x"6f",
          9414 => x"40",
          9415 => x"38",
          9416 => x"2e",
          9417 => x"00",
          9418 => x"61",
          9419 => x"72",
          9420 => x"72",
          9421 => x"20",
          9422 => x"65",
          9423 => x"64",
          9424 => x"00",
          9425 => x"65",
          9426 => x"72",
          9427 => x"67",
          9428 => x"70",
          9429 => x"61",
          9430 => x"6e",
          9431 => x"0a",
          9432 => x"6f",
          9433 => x"72",
          9434 => x"6f",
          9435 => x"67",
          9436 => x"0a",
          9437 => x"50",
          9438 => x"69",
          9439 => x"64",
          9440 => x"73",
          9441 => x"2e",
          9442 => x"00",
          9443 => x"64",
          9444 => x"73",
          9445 => x"00",
          9446 => x"64",
          9447 => x"73",
          9448 => x"61",
          9449 => x"6f",
          9450 => x"6e",
          9451 => x"00",
          9452 => x"75",
          9453 => x"6e",
          9454 => x"2e",
          9455 => x"6e",
          9456 => x"69",
          9457 => x"69",
          9458 => x"72",
          9459 => x"74",
          9460 => x"2e",
          9461 => x"00",
          9462 => x"00",
          9463 => x"00",
          9464 => x"00",
          9465 => x"00",
          9466 => x"01",
          9467 => x"00",
          9468 => x"01",
          9469 => x"81",
          9470 => x"00",
          9471 => x"7f",
          9472 => x"00",
          9473 => x"00",
          9474 => x"00",
          9475 => x"00",
          9476 => x"f5",
          9477 => x"f5",
          9478 => x"f5",
          9479 => x"00",
          9480 => x"01",
          9481 => x"01",
          9482 => x"01",
          9483 => x"00",
          9484 => x"00",
          9485 => x"00",
          9486 => x"00",
          9487 => x"00",
          9488 => x"00",
          9489 => x"00",
          9490 => x"00",
          9491 => x"00",
          9492 => x"00",
          9493 => x"00",
          9494 => x"00",
          9495 => x"00",
          9496 => x"00",
          9497 => x"00",
          9498 => x"00",
          9499 => x"00",
          9500 => x"00",
          9501 => x"00",
          9502 => x"00",
          9503 => x"00",
          9504 => x"00",
          9505 => x"00",
          9506 => x"00",
          9507 => x"00",
          9508 => x"00",
          9509 => x"00",
          9510 => x"00",
          9511 => x"00",
          9512 => x"00",
          9513 => x"00",
          9514 => x"00",
          9515 => x"00",
          9516 => x"00",
          9517 => x"00",
          9518 => x"00",
          9519 => x"00",
          9520 => x"00",
          9521 => x"00",
          9522 => x"00",
          9523 => x"00",
          9524 => x"02",
          9525 => x"00",
          9526 => x"00",
          9527 => x"00",
          9528 => x"04",
          9529 => x"00",
          9530 => x"00",
          9531 => x"00",
          9532 => x"14",
          9533 => x"00",
          9534 => x"00",
          9535 => x"00",
          9536 => x"2b",
          9537 => x"00",
          9538 => x"00",
          9539 => x"00",
          9540 => x"30",
          9541 => x"00",
          9542 => x"00",
          9543 => x"00",
          9544 => x"3c",
          9545 => x"00",
          9546 => x"00",
          9547 => x"00",
          9548 => x"3d",
          9549 => x"00",
          9550 => x"00",
          9551 => x"00",
          9552 => x"3f",
          9553 => x"00",
          9554 => x"00",
          9555 => x"00",
          9556 => x"40",
          9557 => x"00",
          9558 => x"00",
          9559 => x"00",
          9560 => x"41",
          9561 => x"00",
          9562 => x"00",
          9563 => x"00",
          9564 => x"42",
          9565 => x"00",
          9566 => x"00",
          9567 => x"00",
          9568 => x"43",
          9569 => x"00",
          9570 => x"00",
          9571 => x"00",
          9572 => x"50",
          9573 => x"00",
          9574 => x"00",
          9575 => x"00",
          9576 => x"51",
          9577 => x"00",
          9578 => x"00",
          9579 => x"00",
          9580 => x"54",
          9581 => x"00",
          9582 => x"00",
          9583 => x"00",
          9584 => x"55",
          9585 => x"00",
          9586 => x"00",
          9587 => x"00",
          9588 => x"79",
          9589 => x"00",
          9590 => x"00",
          9591 => x"00",
          9592 => x"78",
          9593 => x"00",
          9594 => x"00",
          9595 => x"00",
          9596 => x"82",
          9597 => x"00",
          9598 => x"00",
          9599 => x"00",
          9600 => x"83",
          9601 => x"00",
          9602 => x"00",
          9603 => x"00",
          9604 => x"85",
          9605 => x"00",
          9606 => x"00",
          9607 => x"00",
          9608 => x"87",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"8c",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"8d",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"8e",
          9621 => x"00",
          9622 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e0",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"d0",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cf",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"81",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"9f",
           281 => x"a4",
           282 => x"80",
           283 => x"05",
           284 => x"0b",
           285 => x"04",
           286 => x"9e",
           287 => x"80",
           288 => x"fe",
           289 => x"00",
           290 => x"94",
           291 => x"0d",
           292 => x"08",
           293 => x"52",
           294 => x"05",
           295 => x"de",
           296 => x"70",
           297 => x"85",
           298 => x"0c",
           299 => x"02",
           300 => x"3d",
           301 => x"94",
           302 => x"08",
           303 => x"88",
           304 => x"82",
           305 => x"08",
           306 => x"54",
           307 => x"94",
           308 => x"08",
           309 => x"f9",
           310 => x"0b",
           311 => x"05",
           312 => x"88",
           313 => x"25",
           314 => x"08",
           315 => x"30",
           316 => x"05",
           317 => x"94",
           318 => x"0c",
           319 => x"05",
           320 => x"81",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"0c",
           325 => x"05",
           326 => x"ab",
           327 => x"8c",
           328 => x"94",
           329 => x"0c",
           330 => x"08",
           331 => x"94",
           332 => x"08",
           333 => x"0b",
           334 => x"05",
           335 => x"f0",
           336 => x"08",
           337 => x"80",
           338 => x"8c",
           339 => x"94",
           340 => x"08",
           341 => x"3f",
           342 => x"94",
           343 => x"0c",
           344 => x"fc",
           345 => x"2e",
           346 => x"08",
           347 => x"30",
           348 => x"05",
           349 => x"f8",
           350 => x"88",
           351 => x"3d",
           352 => x"04",
           353 => x"94",
           354 => x"0d",
           355 => x"08",
           356 => x"94",
           357 => x"08",
           358 => x"38",
           359 => x"05",
           360 => x"08",
           361 => x"81",
           362 => x"fc",
           363 => x"08",
           364 => x"80",
           365 => x"94",
           366 => x"08",
           367 => x"8c",
           368 => x"53",
           369 => x"05",
           370 => x"08",
           371 => x"51",
           372 => x"08",
           373 => x"f8",
           374 => x"94",
           375 => x"08",
           376 => x"38",
           377 => x"05",
           378 => x"08",
           379 => x"94",
           380 => x"08",
           381 => x"54",
           382 => x"94",
           383 => x"08",
           384 => x"fd",
           385 => x"0b",
           386 => x"05",
           387 => x"94",
           388 => x"0c",
           389 => x"05",
           390 => x"88",
           391 => x"ac",
           392 => x"fc",
           393 => x"2e",
           394 => x"0b",
           395 => x"05",
           396 => x"38",
           397 => x"05",
           398 => x"08",
           399 => x"94",
           400 => x"08",
           401 => x"fc",
           402 => x"39",
           403 => x"05",
           404 => x"80",
           405 => x"08",
           406 => x"94",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"05",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"05",
           415 => x"08",
           416 => x"94",
           417 => x"08",
           418 => x"08",
           419 => x"94",
           420 => x"08",
           421 => x"08",
           422 => x"ff",
           423 => x"08",
           424 => x"80",
           425 => x"94",
           426 => x"08",
           427 => x"f4",
           428 => x"8d",
           429 => x"f8",
           430 => x"94",
           431 => x"0c",
           432 => x"f4",
           433 => x"0c",
           434 => x"94",
           435 => x"3d",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"c0",
           441 => x"87",
           442 => x"08",
           443 => x"51",
           444 => x"2e",
           445 => x"c0",
           446 => x"51",
           447 => x"87",
           448 => x"08",
           449 => x"06",
           450 => x"38",
           451 => x"8c",
           452 => x"80",
           453 => x"71",
           454 => x"9f",
           455 => x"0b",
           456 => x"33",
           457 => x"3d",
           458 => x"3d",
           459 => x"7d",
           460 => x"80",
           461 => x"0b",
           462 => x"81",
           463 => x"82",
           464 => x"2e",
           465 => x"81",
           466 => x"0b",
           467 => x"8c",
           468 => x"c0",
           469 => x"84",
           470 => x"92",
           471 => x"c0",
           472 => x"70",
           473 => x"81",
           474 => x"53",
           475 => x"a7",
           476 => x"92",
           477 => x"81",
           478 => x"79",
           479 => x"51",
           480 => x"90",
           481 => x"2e",
           482 => x"76",
           483 => x"58",
           484 => x"54",
           485 => x"72",
           486 => x"70",
           487 => x"38",
           488 => x"8c",
           489 => x"ff",
           490 => x"c0",
           491 => x"51",
           492 => x"81",
           493 => x"92",
           494 => x"c0",
           495 => x"70",
           496 => x"51",
           497 => x"80",
           498 => x"80",
           499 => x"70",
           500 => x"81",
           501 => x"87",
           502 => x"08",
           503 => x"2e",
           504 => x"83",
           505 => x"71",
           506 => x"3d",
           507 => x"3d",
           508 => x"11",
           509 => x"71",
           510 => x"88",
           511 => x"84",
           512 => x"fd",
           513 => x"83",
           514 => x"12",
           515 => x"2b",
           516 => x"07",
           517 => x"70",
           518 => x"2b",
           519 => x"07",
           520 => x"53",
           521 => x"52",
           522 => x"04",
           523 => x"79",
           524 => x"9f",
           525 => x"57",
           526 => x"80",
           527 => x"88",
           528 => x"80",
           529 => x"33",
           530 => x"2e",
           531 => x"83",
           532 => x"80",
           533 => x"54",
           534 => x"fe",
           535 => x"88",
           536 => x"08",
           537 => x"3d",
           538 => x"fd",
           539 => x"08",
           540 => x"51",
           541 => x"88",
           542 => x"ff",
           543 => x"39",
           544 => x"82",
           545 => x"06",
           546 => x"2a",
           547 => x"05",
           548 => x"70",
           549 => x"92",
           550 => x"8e",
           551 => x"fe",
           552 => x"08",
           553 => x"55",
           554 => x"55",
           555 => x"89",
           556 => x"fb",
           557 => x"0b",
           558 => x"08",
           559 => x"12",
           560 => x"55",
           561 => x"56",
           562 => x"8d",
           563 => x"33",
           564 => x"94",
           565 => x"57",
           566 => x"0c",
           567 => x"04",
           568 => x"75",
           569 => x"0b",
           570 => x"f4",
           571 => x"51",
           572 => x"83",
           573 => x"06",
           574 => x"14",
           575 => x"3f",
           576 => x"2b",
           577 => x"51",
           578 => x"88",
           579 => x"ff",
           580 => x"88",
           581 => x"0d",
           582 => x"0d",
           583 => x"0b",
           584 => x"55",
           585 => x"23",
           586 => x"53",
           587 => x"88",
           588 => x"08",
           589 => x"38",
           590 => x"39",
           591 => x"73",
           592 => x"83",
           593 => x"06",
           594 => x"14",
           595 => x"8c",
           596 => x"80",
           597 => x"72",
           598 => x"3f",
           599 => x"85",
           600 => x"08",
           601 => x"16",
           602 => x"71",
           603 => x"3d",
           604 => x"3d",
           605 => x"0b",
           606 => x"08",
           607 => x"05",
           608 => x"ff",
           609 => x"57",
           610 => x"2e",
           611 => x"15",
           612 => x"86",
           613 => x"80",
           614 => x"8f",
           615 => x"80",
           616 => x"13",
           617 => x"8c",
           618 => x"72",
           619 => x"0b",
           620 => x"57",
           621 => x"27",
           622 => x"39",
           623 => x"ff",
           624 => x"2a",
           625 => x"a8",
           626 => x"fc",
           627 => x"52",
           628 => x"27",
           629 => x"52",
           630 => x"17",
           631 => x"38",
           632 => x"16",
           633 => x"51",
           634 => x"88",
           635 => x"0c",
           636 => x"80",
           637 => x"0c",
           638 => x"04",
           639 => x"60",
           640 => x"5e",
           641 => x"55",
           642 => x"09",
           643 => x"38",
           644 => x"44",
           645 => x"62",
           646 => x"56",
           647 => x"09",
           648 => x"38",
           649 => x"80",
           650 => x"0c",
           651 => x"51",
           652 => x"26",
           653 => x"51",
           654 => x"88",
           655 => x"7d",
           656 => x"39",
           657 => x"1d",
           658 => x"5a",
           659 => x"a0",
           660 => x"05",
           661 => x"15",
           662 => x"2e",
           663 => x"ef",
           664 => x"59",
           665 => x"08",
           666 => x"81",
           667 => x"ff",
           668 => x"70",
           669 => x"32",
           670 => x"73",
           671 => x"25",
           672 => x"52",
           673 => x"57",
           674 => x"c7",
           675 => x"2e",
           676 => x"83",
           677 => x"77",
           678 => x"07",
           679 => x"2e",
           680 => x"88",
           681 => x"78",
           682 => x"30",
           683 => x"9f",
           684 => x"57",
           685 => x"9b",
           686 => x"8b",
           687 => x"39",
           688 => x"70",
           689 => x"72",
           690 => x"57",
           691 => x"34",
           692 => x"7a",
           693 => x"80",
           694 => x"26",
           695 => x"55",
           696 => x"34",
           697 => x"b1",
           698 => x"80",
           699 => x"54",
           700 => x"85",
           701 => x"06",
           702 => x"1c",
           703 => x"51",
           704 => x"88",
           705 => x"08",
           706 => x"7c",
           707 => x"80",
           708 => x"38",
           709 => x"70",
           710 => x"81",
           711 => x"56",
           712 => x"8b",
           713 => x"08",
           714 => x"5b",
           715 => x"18",
           716 => x"2e",
           717 => x"70",
           718 => x"33",
           719 => x"05",
           720 => x"71",
           721 => x"56",
           722 => x"e2",
           723 => x"75",
           724 => x"38",
           725 => x"9a",
           726 => x"39",
           727 => x"88",
           728 => x"83",
           729 => x"84",
           730 => x"11",
           731 => x"74",
           732 => x"1d",
           733 => x"2a",
           734 => x"51",
           735 => x"89",
           736 => x"92",
           737 => x"8e",
           738 => x"fa",
           739 => x"08",
           740 => x"fd",
           741 => x"88",
           742 => x"0d",
           743 => x"0d",
           744 => x"57",
           745 => x"fe",
           746 => x"76",
           747 => x"3f",
           748 => x"08",
           749 => x"76",
           750 => x"3f",
           751 => x"ff",
           752 => x"82",
           753 => x"d4",
           754 => x"81",
           755 => x"38",
           756 => x"53",
           757 => x"51",
           758 => x"88",
           759 => x"08",
           760 => x"51",
           761 => x"88",
           762 => x"ff",
           763 => x"81",
           764 => x"a9",
           765 => x"80",
           766 => x"52",
           767 => x"aa",
           768 => x"56",
           769 => x"38",
           770 => x"e2",
           771 => x"83",
           772 => x"55",
           773 => x"c6",
           774 => x"81",
           775 => x"0c",
           776 => x"04",
           777 => x"65",
           778 => x"0b",
           779 => x"f4",
           780 => x"3f",
           781 => x"06",
           782 => x"74",
           783 => x"74",
           784 => x"3d",
           785 => x"5a",
           786 => x"88",
           787 => x"06",
           788 => x"2e",
           789 => x"b3",
           790 => x"83",
           791 => x"52",
           792 => x"c6",
           793 => x"ab",
           794 => x"33",
           795 => x"2e",
           796 => x"3d",
           797 => x"f7",
           798 => x"08",
           799 => x"76",
           800 => x"99",
           801 => x"81",
           802 => x"76",
           803 => x"81",
           804 => x"81",
           805 => x"39",
           806 => x"86",
           807 => x"82",
           808 => x"54",
           809 => x"52",
           810 => x"fe",
           811 => x"88",
           812 => x"38",
           813 => x"05",
           814 => x"3f",
           815 => x"ff",
           816 => x"77",
           817 => x"3d",
           818 => x"f6",
           819 => x"08",
           820 => x"05",
           821 => x"29",
           822 => x"ad",
           823 => x"52",
           824 => x"8a",
           825 => x"83",
           826 => x"7a",
           827 => x"0c",
           828 => x"82",
           829 => x"3d",
           830 => x"f5",
           831 => x"08",
           832 => x"95",
           833 => x"51",
           834 => x"88",
           835 => x"ff",
           836 => x"8c",
           837 => x"ef",
           838 => x"e7",
           839 => x"56",
           840 => x"ca",
           841 => x"83",
           842 => x"76",
           843 => x"31",
           844 => x"70",
           845 => x"1d",
           846 => x"71",
           847 => x"5c",
           848 => x"c4",
           849 => x"82",
           850 => x"1b",
           851 => x"e0",
           852 => x"56",
           853 => x"fe",
           854 => x"82",
           855 => x"f6",
           856 => x"38",
           857 => x"39",
           858 => x"80",
           859 => x"38",
           860 => x"76",
           861 => x"81",
           862 => x"95",
           863 => x"51",
           864 => x"88",
           865 => x"0c",
           866 => x"19",
           867 => x"1a",
           868 => x"ff",
           869 => x"1a",
           870 => x"84",
           871 => x"1b",
           872 => x"0b",
           873 => x"78",
           874 => x"9f",
           875 => x"56",
           876 => x"95",
           877 => x"ea",
           878 => x"0b",
           879 => x"08",
           880 => x"74",
           881 => x"df",
           882 => x"81",
           883 => x"3d",
           884 => x"69",
           885 => x"70",
           886 => x"05",
           887 => x"3f",
           888 => x"88",
           889 => x"38",
           890 => x"54",
           891 => x"93",
           892 => x"05",
           893 => x"2a",
           894 => x"51",
           895 => x"80",
           896 => x"83",
           897 => x"75",
           898 => x"3f",
           899 => x"16",
           900 => x"dc",
           901 => x"eb",
           902 => x"9c",
           903 => x"98",
           904 => x"0b",
           905 => x"73",
           906 => x"3d",
           907 => x"3d",
           908 => x"7e",
           909 => x"9f",
           910 => x"5b",
           911 => x"7b",
           912 => x"75",
           913 => x"d1",
           914 => x"33",
           915 => x"84",
           916 => x"2e",
           917 => x"91",
           918 => x"17",
           919 => x"80",
           920 => x"34",
           921 => x"b1",
           922 => x"08",
           923 => x"31",
           924 => x"27",
           925 => x"58",
           926 => x"81",
           927 => x"16",
           928 => x"ff",
           929 => x"74",
           930 => x"82",
           931 => x"05",
           932 => x"06",
           933 => x"06",
           934 => x"9e",
           935 => x"38",
           936 => x"55",
           937 => x"16",
           938 => x"80",
           939 => x"55",
           940 => x"ff",
           941 => x"a4",
           942 => x"16",
           943 => x"f3",
           944 => x"55",
           945 => x"2e",
           946 => x"88",
           947 => x"17",
           948 => x"08",
           949 => x"84",
           950 => x"51",
           951 => x"27",
           952 => x"55",
           953 => x"16",
           954 => x"06",
           955 => x"08",
           956 => x"f0",
           957 => x"08",
           958 => x"98",
           959 => x"98",
           960 => x"75",
           961 => x"16",
           962 => x"78",
           963 => x"e8",
           964 => x"59",
           965 => x"80",
           966 => x"0c",
           967 => x"04",
           968 => x"87",
           969 => x"08",
           970 => x"80",
           971 => x"ea",
           972 => x"08",
           973 => x"c0",
           974 => x"56",
           975 => x"80",
           976 => x"ea",
           977 => x"88",
           978 => x"c0",
           979 => x"87",
           980 => x"08",
           981 => x"80",
           982 => x"ea",
           983 => x"08",
           984 => x"c0",
           985 => x"56",
           986 => x"80",
           987 => x"ea",
           988 => x"88",
           989 => x"c0",
           990 => x"8c",
           991 => x"87",
           992 => x"0c",
           993 => x"0b",
           994 => x"94",
           995 => x"51",
           996 => x"88",
           997 => x"9f",
           998 => x"9b",
           999 => x"ae",
          1000 => x"0b",
          1001 => x"c0",
          1002 => x"55",
          1003 => x"05",
          1004 => x"52",
          1005 => x"f6",
          1006 => x"8d",
          1007 => x"73",
          1008 => x"38",
          1009 => x"e4",
          1010 => x"54",
          1011 => x"54",
          1012 => x"00",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"42",
          1017 => x"54",
          1018 => x"2e",
          1019 => x"00",
          1020 => x"01",
          2048 => x"0b",
          2049 => x"80",
          2050 => x"0b",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"80",
          2058 => x"0b",
          2059 => x"0b",
          2060 => x"93",
          2061 => x"0b",
          2062 => x"0b",
          2063 => x"b3",
          2064 => x"0b",
          2065 => x"0b",
          2066 => x"d3",
          2067 => x"0b",
          2068 => x"0b",
          2069 => x"f3",
          2070 => x"0b",
          2071 => x"0b",
          2072 => x"93",
          2073 => x"0b",
          2074 => x"0b",
          2075 => x"b3",
          2076 => x"0b",
          2077 => x"0b",
          2078 => x"d3",
          2079 => x"0b",
          2080 => x"0b",
          2081 => x"f1",
          2082 => x"0b",
          2083 => x"0b",
          2084 => x"8f",
          2085 => x"0b",
          2086 => x"0b",
          2087 => x"ae",
          2088 => x"0b",
          2089 => x"0b",
          2090 => x"ce",
          2091 => x"0b",
          2092 => x"0b",
          2093 => x"ee",
          2094 => x"0b",
          2095 => x"0b",
          2096 => x"8e",
          2097 => x"0b",
          2098 => x"0b",
          2099 => x"ae",
          2100 => x"0b",
          2101 => x"0b",
          2102 => x"ce",
          2103 => x"0b",
          2104 => x"0b",
          2105 => x"ee",
          2106 => x"0b",
          2107 => x"0b",
          2108 => x"8e",
          2109 => x"0b",
          2110 => x"0b",
          2111 => x"ae",
          2112 => x"0b",
          2113 => x"0b",
          2114 => x"ce",
          2115 => x"0b",
          2116 => x"0b",
          2117 => x"ee",
          2118 => x"0b",
          2119 => x"0b",
          2120 => x"8e",
          2121 => x"0b",
          2122 => x"0b",
          2123 => x"ae",
          2124 => x"0b",
          2125 => x"0b",
          2126 => x"ce",
          2127 => x"0b",
          2128 => x"0b",
          2129 => x"ee",
          2130 => x"0b",
          2131 => x"0b",
          2132 => x"8d",
          2133 => x"0b",
          2134 => x"0b",
          2135 => x"ab",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"00",
          2177 => x"82",
          2178 => x"b8",
          2179 => x"8c",
          2180 => x"80",
          2181 => x"8c",
          2182 => x"c9",
          2183 => x"8c",
          2184 => x"80",
          2185 => x"8c",
          2186 => x"c9",
          2187 => x"8c",
          2188 => x"80",
          2189 => x"8c",
          2190 => x"ca",
          2191 => x"8c",
          2192 => x"80",
          2193 => x"8c",
          2194 => x"d0",
          2195 => x"8c",
          2196 => x"80",
          2197 => x"8c",
          2198 => x"d1",
          2199 => x"8c",
          2200 => x"80",
          2201 => x"8c",
          2202 => x"ca",
          2203 => x"8c",
          2204 => x"80",
          2205 => x"8c",
          2206 => x"d1",
          2207 => x"8c",
          2208 => x"80",
          2209 => x"8c",
          2210 => x"d3",
          2211 => x"8c",
          2212 => x"80",
          2213 => x"8c",
          2214 => x"cf",
          2215 => x"8c",
          2216 => x"80",
          2217 => x"8c",
          2218 => x"ca",
          2219 => x"8c",
          2220 => x"80",
          2221 => x"8c",
          2222 => x"d0",
          2223 => x"8c",
          2224 => x"80",
          2225 => x"8c",
          2226 => x"d0",
          2227 => x"8c",
          2228 => x"80",
          2229 => x"8c",
          2230 => x"ad",
          2231 => x"e8",
          2232 => x"90",
          2233 => x"e8",
          2234 => x"2d",
          2235 => x"08",
          2236 => x"04",
          2237 => x"0c",
          2238 => x"82",
          2239 => x"83",
          2240 => x"82",
          2241 => x"b4",
          2242 => x"8c",
          2243 => x"80",
          2244 => x"8c",
          2245 => x"82",
          2246 => x"e8",
          2247 => x"90",
          2248 => x"e8",
          2249 => x"a5",
          2250 => x"e8",
          2251 => x"90",
          2252 => x"e8",
          2253 => x"96",
          2254 => x"e8",
          2255 => x"90",
          2256 => x"e8",
          2257 => x"8a",
          2258 => x"e8",
          2259 => x"90",
          2260 => x"e8",
          2261 => x"87",
          2262 => x"e8",
          2263 => x"90",
          2264 => x"e8",
          2265 => x"a5",
          2266 => x"e8",
          2267 => x"90",
          2268 => x"e8",
          2269 => x"85",
          2270 => x"e8",
          2271 => x"90",
          2272 => x"e8",
          2273 => x"f8",
          2274 => x"e8",
          2275 => x"90",
          2276 => x"e8",
          2277 => x"c4",
          2278 => x"e8",
          2279 => x"90",
          2280 => x"e8",
          2281 => x"e3",
          2282 => x"e8",
          2283 => x"90",
          2284 => x"e8",
          2285 => x"82",
          2286 => x"e8",
          2287 => x"90",
          2288 => x"e8",
          2289 => x"ec",
          2290 => x"e8",
          2291 => x"90",
          2292 => x"e8",
          2293 => x"d2",
          2294 => x"e8",
          2295 => x"90",
          2296 => x"e8",
          2297 => x"c0",
          2298 => x"e8",
          2299 => x"90",
          2300 => x"e8",
          2301 => x"86",
          2302 => x"e8",
          2303 => x"90",
          2304 => x"e8",
          2305 => x"c0",
          2306 => x"e8",
          2307 => x"90",
          2308 => x"e8",
          2309 => x"c1",
          2310 => x"e8",
          2311 => x"90",
          2312 => x"e8",
          2313 => x"f6",
          2314 => x"e8",
          2315 => x"90",
          2316 => x"e8",
          2317 => x"cf",
          2318 => x"e8",
          2319 => x"90",
          2320 => x"e8",
          2321 => x"fa",
          2322 => x"e8",
          2323 => x"90",
          2324 => x"e8",
          2325 => x"dd",
          2326 => x"e8",
          2327 => x"90",
          2328 => x"e8",
          2329 => x"b2",
          2330 => x"e8",
          2331 => x"90",
          2332 => x"e8",
          2333 => x"bc",
          2334 => x"e8",
          2335 => x"90",
          2336 => x"e8",
          2337 => x"fe",
          2338 => x"e8",
          2339 => x"90",
          2340 => x"e8",
          2341 => x"c4",
          2342 => x"e8",
          2343 => x"90",
          2344 => x"e8",
          2345 => x"ea",
          2346 => x"e8",
          2347 => x"90",
          2348 => x"e8",
          2349 => x"9f",
          2350 => x"e8",
          2351 => x"90",
          2352 => x"e8",
          2353 => x"8b",
          2354 => x"e8",
          2355 => x"90",
          2356 => x"e8",
          2357 => x"ff",
          2358 => x"e8",
          2359 => x"90",
          2360 => x"e8",
          2361 => x"e9",
          2362 => x"e8",
          2363 => x"90",
          2364 => x"e8",
          2365 => x"cd",
          2366 => x"e8",
          2367 => x"90",
          2368 => x"e8",
          2369 => x"2d",
          2370 => x"08",
          2371 => x"04",
          2372 => x"0c",
          2373 => x"82",
          2374 => x"83",
          2375 => x"82",
          2376 => x"b7",
          2377 => x"8c",
          2378 => x"80",
          2379 => x"8c",
          2380 => x"d6",
          2381 => x"8c",
          2382 => x"80",
          2383 => x"8c",
          2384 => x"a4",
          2385 => x"38",
          2386 => x"84",
          2387 => x"0b",
          2388 => x"be",
          2389 => x"51",
          2390 => x"04",
          2391 => x"8c",
          2392 => x"82",
          2393 => x"fd",
          2394 => x"53",
          2395 => x"08",
          2396 => x"52",
          2397 => x"08",
          2398 => x"51",
          2399 => x"82",
          2400 => x"70",
          2401 => x"0c",
          2402 => x"0d",
          2403 => x"0c",
          2404 => x"e8",
          2405 => x"8c",
          2406 => x"3d",
          2407 => x"82",
          2408 => x"8c",
          2409 => x"82",
          2410 => x"88",
          2411 => x"93",
          2412 => x"dc",
          2413 => x"8c",
          2414 => x"85",
          2415 => x"8c",
          2416 => x"82",
          2417 => x"02",
          2418 => x"0c",
          2419 => x"81",
          2420 => x"e8",
          2421 => x"0c",
          2422 => x"8c",
          2423 => x"05",
          2424 => x"e8",
          2425 => x"08",
          2426 => x"08",
          2427 => x"27",
          2428 => x"8c",
          2429 => x"05",
          2430 => x"ae",
          2431 => x"82",
          2432 => x"8c",
          2433 => x"a2",
          2434 => x"e8",
          2435 => x"08",
          2436 => x"e8",
          2437 => x"0c",
          2438 => x"08",
          2439 => x"10",
          2440 => x"08",
          2441 => x"ff",
          2442 => x"8c",
          2443 => x"05",
          2444 => x"80",
          2445 => x"8c",
          2446 => x"05",
          2447 => x"e8",
          2448 => x"08",
          2449 => x"82",
          2450 => x"88",
          2451 => x"8c",
          2452 => x"05",
          2453 => x"8c",
          2454 => x"05",
          2455 => x"e8",
          2456 => x"08",
          2457 => x"08",
          2458 => x"07",
          2459 => x"08",
          2460 => x"82",
          2461 => x"fc",
          2462 => x"2a",
          2463 => x"08",
          2464 => x"82",
          2465 => x"8c",
          2466 => x"2a",
          2467 => x"08",
          2468 => x"ff",
          2469 => x"8c",
          2470 => x"05",
          2471 => x"93",
          2472 => x"e8",
          2473 => x"08",
          2474 => x"e8",
          2475 => x"0c",
          2476 => x"82",
          2477 => x"f8",
          2478 => x"82",
          2479 => x"f4",
          2480 => x"82",
          2481 => x"f4",
          2482 => x"8c",
          2483 => x"3d",
          2484 => x"e8",
          2485 => x"3d",
          2486 => x"79",
          2487 => x"55",
          2488 => x"27",
          2489 => x"75",
          2490 => x"51",
          2491 => x"a9",
          2492 => x"52",
          2493 => x"98",
          2494 => x"81",
          2495 => x"74",
          2496 => x"56",
          2497 => x"52",
          2498 => x"09",
          2499 => x"38",
          2500 => x"dc",
          2501 => x"0d",
          2502 => x"72",
          2503 => x"54",
          2504 => x"84",
          2505 => x"72",
          2506 => x"54",
          2507 => x"84",
          2508 => x"72",
          2509 => x"54",
          2510 => x"84",
          2511 => x"72",
          2512 => x"54",
          2513 => x"84",
          2514 => x"f0",
          2515 => x"8f",
          2516 => x"83",
          2517 => x"38",
          2518 => x"05",
          2519 => x"70",
          2520 => x"0c",
          2521 => x"71",
          2522 => x"38",
          2523 => x"81",
          2524 => x"0d",
          2525 => x"02",
          2526 => x"05",
          2527 => x"53",
          2528 => x"27",
          2529 => x"83",
          2530 => x"80",
          2531 => x"ff",
          2532 => x"ff",
          2533 => x"73",
          2534 => x"05",
          2535 => x"12",
          2536 => x"2e",
          2537 => x"ef",
          2538 => x"8c",
          2539 => x"3d",
          2540 => x"74",
          2541 => x"07",
          2542 => x"2b",
          2543 => x"51",
          2544 => x"a5",
          2545 => x"70",
          2546 => x"0c",
          2547 => x"84",
          2548 => x"72",
          2549 => x"05",
          2550 => x"71",
          2551 => x"53",
          2552 => x"52",
          2553 => x"dd",
          2554 => x"27",
          2555 => x"71",
          2556 => x"53",
          2557 => x"52",
          2558 => x"f2",
          2559 => x"ff",
          2560 => x"3d",
          2561 => x"79",
          2562 => x"83",
          2563 => x"54",
          2564 => x"c3",
          2565 => x"08",
          2566 => x"f7",
          2567 => x"13",
          2568 => x"84",
          2569 => x"06",
          2570 => x"53",
          2571 => x"38",
          2572 => x"74",
          2573 => x"56",
          2574 => x"70",
          2575 => x"fb",
          2576 => x"06",
          2577 => x"82",
          2578 => x"51",
          2579 => x"54",
          2580 => x"dc",
          2581 => x"71",
          2582 => x"53",
          2583 => x"73",
          2584 => x"55",
          2585 => x"38",
          2586 => x"dc",
          2587 => x"0d",
          2588 => x"0d",
          2589 => x"83",
          2590 => x"52",
          2591 => x"71",
          2592 => x"09",
          2593 => x"ff",
          2594 => x"f8",
          2595 => x"80",
          2596 => x"52",
          2597 => x"38",
          2598 => x"08",
          2599 => x"fb",
          2600 => x"06",
          2601 => x"82",
          2602 => x"51",
          2603 => x"70",
          2604 => x"38",
          2605 => x"33",
          2606 => x"2e",
          2607 => x"12",
          2608 => x"52",
          2609 => x"71",
          2610 => x"8c",
          2611 => x"3d",
          2612 => x"3d",
          2613 => x"7c",
          2614 => x"55",
          2615 => x"2e",
          2616 => x"71",
          2617 => x"06",
          2618 => x"2e",
          2619 => x"ff",
          2620 => x"ff",
          2621 => x"71",
          2622 => x"56",
          2623 => x"2e",
          2624 => x"a9",
          2625 => x"2e",
          2626 => x"70",
          2627 => x"51",
          2628 => x"80",
          2629 => x"12",
          2630 => x"15",
          2631 => x"72",
          2632 => x"81",
          2633 => x"71",
          2634 => x"56",
          2635 => x"ff",
          2636 => x"ff",
          2637 => x"31",
          2638 => x"70",
          2639 => x"0c",
          2640 => x"04",
          2641 => x"55",
          2642 => x"88",
          2643 => x"74",
          2644 => x"38",
          2645 => x"52",
          2646 => x"fc",
          2647 => x"80",
          2648 => x"74",
          2649 => x"f7",
          2650 => x"12",
          2651 => x"84",
          2652 => x"06",
          2653 => x"70",
          2654 => x"15",
          2655 => x"55",
          2656 => x"d0",
          2657 => x"76",
          2658 => x"38",
          2659 => x"52",
          2660 => x"80",
          2661 => x"dc",
          2662 => x"0d",
          2663 => x"0d",
          2664 => x"53",
          2665 => x"52",
          2666 => x"82",
          2667 => x"81",
          2668 => x"07",
          2669 => x"52",
          2670 => x"e8",
          2671 => x"8c",
          2672 => x"3d",
          2673 => x"3d",
          2674 => x"08",
          2675 => x"56",
          2676 => x"80",
          2677 => x"33",
          2678 => x"2e",
          2679 => x"86",
          2680 => x"52",
          2681 => x"53",
          2682 => x"13",
          2683 => x"33",
          2684 => x"06",
          2685 => x"70",
          2686 => x"38",
          2687 => x"80",
          2688 => x"74",
          2689 => x"81",
          2690 => x"70",
          2691 => x"81",
          2692 => x"80",
          2693 => x"05",
          2694 => x"76",
          2695 => x"70",
          2696 => x"0c",
          2697 => x"04",
          2698 => x"76",
          2699 => x"80",
          2700 => x"86",
          2701 => x"52",
          2702 => x"99",
          2703 => x"dc",
          2704 => x"80",
          2705 => x"74",
          2706 => x"8c",
          2707 => x"3d",
          2708 => x"3d",
          2709 => x"11",
          2710 => x"52",
          2711 => x"70",
          2712 => x"98",
          2713 => x"33",
          2714 => x"82",
          2715 => x"26",
          2716 => x"84",
          2717 => x"83",
          2718 => x"26",
          2719 => x"85",
          2720 => x"84",
          2721 => x"26",
          2722 => x"86",
          2723 => x"85",
          2724 => x"26",
          2725 => x"88",
          2726 => x"86",
          2727 => x"e7",
          2728 => x"38",
          2729 => x"54",
          2730 => x"87",
          2731 => x"cc",
          2732 => x"87",
          2733 => x"0c",
          2734 => x"c0",
          2735 => x"82",
          2736 => x"c0",
          2737 => x"83",
          2738 => x"c0",
          2739 => x"84",
          2740 => x"c0",
          2741 => x"85",
          2742 => x"c0",
          2743 => x"86",
          2744 => x"c0",
          2745 => x"74",
          2746 => x"a4",
          2747 => x"c0",
          2748 => x"80",
          2749 => x"98",
          2750 => x"52",
          2751 => x"dc",
          2752 => x"0d",
          2753 => x"0d",
          2754 => x"c0",
          2755 => x"81",
          2756 => x"c0",
          2757 => x"5e",
          2758 => x"87",
          2759 => x"08",
          2760 => x"1c",
          2761 => x"98",
          2762 => x"79",
          2763 => x"87",
          2764 => x"08",
          2765 => x"1c",
          2766 => x"98",
          2767 => x"79",
          2768 => x"87",
          2769 => x"08",
          2770 => x"1c",
          2771 => x"98",
          2772 => x"7b",
          2773 => x"87",
          2774 => x"08",
          2775 => x"1c",
          2776 => x"0c",
          2777 => x"ff",
          2778 => x"83",
          2779 => x"58",
          2780 => x"57",
          2781 => x"56",
          2782 => x"55",
          2783 => x"54",
          2784 => x"53",
          2785 => x"ff",
          2786 => x"f1",
          2787 => x"de",
          2788 => x"0d",
          2789 => x"0d",
          2790 => x"33",
          2791 => x"9f",
          2792 => x"52",
          2793 => x"82",
          2794 => x"83",
          2795 => x"fb",
          2796 => x"0b",
          2797 => x"d4",
          2798 => x"ff",
          2799 => x"56",
          2800 => x"84",
          2801 => x"2e",
          2802 => x"c0",
          2803 => x"70",
          2804 => x"2a",
          2805 => x"53",
          2806 => x"80",
          2807 => x"71",
          2808 => x"81",
          2809 => x"70",
          2810 => x"81",
          2811 => x"06",
          2812 => x"80",
          2813 => x"71",
          2814 => x"81",
          2815 => x"70",
          2816 => x"73",
          2817 => x"51",
          2818 => x"80",
          2819 => x"2e",
          2820 => x"c0",
          2821 => x"75",
          2822 => x"82",
          2823 => x"87",
          2824 => x"fb",
          2825 => x"9f",
          2826 => x"0b",
          2827 => x"33",
          2828 => x"06",
          2829 => x"87",
          2830 => x"51",
          2831 => x"86",
          2832 => x"94",
          2833 => x"08",
          2834 => x"70",
          2835 => x"54",
          2836 => x"2e",
          2837 => x"91",
          2838 => x"06",
          2839 => x"d7",
          2840 => x"32",
          2841 => x"51",
          2842 => x"2e",
          2843 => x"93",
          2844 => x"06",
          2845 => x"ff",
          2846 => x"81",
          2847 => x"87",
          2848 => x"52",
          2849 => x"86",
          2850 => x"94",
          2851 => x"72",
          2852 => x"0d",
          2853 => x"0d",
          2854 => x"74",
          2855 => x"ff",
          2856 => x"57",
          2857 => x"80",
          2858 => x"81",
          2859 => x"15",
          2860 => x"87",
          2861 => x"81",
          2862 => x"57",
          2863 => x"c0",
          2864 => x"75",
          2865 => x"38",
          2866 => x"94",
          2867 => x"70",
          2868 => x"81",
          2869 => x"52",
          2870 => x"8c",
          2871 => x"2a",
          2872 => x"51",
          2873 => x"38",
          2874 => x"70",
          2875 => x"51",
          2876 => x"8d",
          2877 => x"2a",
          2878 => x"51",
          2879 => x"be",
          2880 => x"ff",
          2881 => x"c0",
          2882 => x"70",
          2883 => x"38",
          2884 => x"90",
          2885 => x"0c",
          2886 => x"33",
          2887 => x"06",
          2888 => x"70",
          2889 => x"76",
          2890 => x"0c",
          2891 => x"04",
          2892 => x"0b",
          2893 => x"d4",
          2894 => x"ff",
          2895 => x"87",
          2896 => x"51",
          2897 => x"86",
          2898 => x"94",
          2899 => x"08",
          2900 => x"70",
          2901 => x"51",
          2902 => x"2e",
          2903 => x"81",
          2904 => x"87",
          2905 => x"52",
          2906 => x"86",
          2907 => x"94",
          2908 => x"08",
          2909 => x"06",
          2910 => x"0c",
          2911 => x"0d",
          2912 => x"0d",
          2913 => x"87",
          2914 => x"81",
          2915 => x"53",
          2916 => x"84",
          2917 => x"2e",
          2918 => x"c0",
          2919 => x"71",
          2920 => x"2a",
          2921 => x"51",
          2922 => x"52",
          2923 => x"a0",
          2924 => x"ff",
          2925 => x"c0",
          2926 => x"70",
          2927 => x"38",
          2928 => x"90",
          2929 => x"70",
          2930 => x"98",
          2931 => x"51",
          2932 => x"dc",
          2933 => x"0d",
          2934 => x"0d",
          2935 => x"80",
          2936 => x"2a",
          2937 => x"51",
          2938 => x"84",
          2939 => x"c0",
          2940 => x"82",
          2941 => x"87",
          2942 => x"08",
          2943 => x"0c",
          2944 => x"94",
          2945 => x"e0",
          2946 => x"9e",
          2947 => x"87",
          2948 => x"c0",
          2949 => x"82",
          2950 => x"87",
          2951 => x"08",
          2952 => x"0c",
          2953 => x"ac",
          2954 => x"f0",
          2955 => x"9e",
          2956 => x"87",
          2957 => x"c0",
          2958 => x"82",
          2959 => x"87",
          2960 => x"08",
          2961 => x"0c",
          2962 => x"bc",
          2963 => x"80",
          2964 => x"9e",
          2965 => x"88",
          2966 => x"c0",
          2967 => x"82",
          2968 => x"87",
          2969 => x"08",
          2970 => x"88",
          2971 => x"c0",
          2972 => x"82",
          2973 => x"87",
          2974 => x"08",
          2975 => x"0c",
          2976 => x"8c",
          2977 => x"98",
          2978 => x"82",
          2979 => x"80",
          2980 => x"9e",
          2981 => x"84",
          2982 => x"51",
          2983 => x"80",
          2984 => x"81",
          2985 => x"88",
          2986 => x"0b",
          2987 => x"90",
          2988 => x"80",
          2989 => x"52",
          2990 => x"2e",
          2991 => x"52",
          2992 => x"9e",
          2993 => x"87",
          2994 => x"08",
          2995 => x"0a",
          2996 => x"52",
          2997 => x"83",
          2998 => x"71",
          2999 => x"34",
          3000 => x"c0",
          3001 => x"70",
          3002 => x"06",
          3003 => x"70",
          3004 => x"38",
          3005 => x"82",
          3006 => x"80",
          3007 => x"9e",
          3008 => x"a0",
          3009 => x"51",
          3010 => x"80",
          3011 => x"81",
          3012 => x"88",
          3013 => x"0b",
          3014 => x"90",
          3015 => x"80",
          3016 => x"52",
          3017 => x"2e",
          3018 => x"52",
          3019 => x"a2",
          3020 => x"87",
          3021 => x"08",
          3022 => x"80",
          3023 => x"52",
          3024 => x"83",
          3025 => x"71",
          3026 => x"34",
          3027 => x"c0",
          3028 => x"70",
          3029 => x"06",
          3030 => x"70",
          3031 => x"38",
          3032 => x"82",
          3033 => x"80",
          3034 => x"9e",
          3035 => x"81",
          3036 => x"51",
          3037 => x"80",
          3038 => x"81",
          3039 => x"88",
          3040 => x"0b",
          3041 => x"90",
          3042 => x"c0",
          3043 => x"52",
          3044 => x"2e",
          3045 => x"52",
          3046 => x"a6",
          3047 => x"87",
          3048 => x"08",
          3049 => x"06",
          3050 => x"70",
          3051 => x"38",
          3052 => x"82",
          3053 => x"87",
          3054 => x"08",
          3055 => x"06",
          3056 => x"51",
          3057 => x"82",
          3058 => x"80",
          3059 => x"9e",
          3060 => x"84",
          3061 => x"52",
          3062 => x"2e",
          3063 => x"52",
          3064 => x"a9",
          3065 => x"9e",
          3066 => x"83",
          3067 => x"84",
          3068 => x"51",
          3069 => x"aa",
          3070 => x"87",
          3071 => x"08",
          3072 => x"51",
          3073 => x"80",
          3074 => x"81",
          3075 => x"88",
          3076 => x"c0",
          3077 => x"70",
          3078 => x"51",
          3079 => x"ac",
          3080 => x"0d",
          3081 => x"0d",
          3082 => x"51",
          3083 => x"82",
          3084 => x"54",
          3085 => x"88",
          3086 => x"90",
          3087 => x"3f",
          3088 => x"51",
          3089 => x"82",
          3090 => x"54",
          3091 => x"93",
          3092 => x"f8",
          3093 => x"fc",
          3094 => x"52",
          3095 => x"51",
          3096 => x"82",
          3097 => x"54",
          3098 => x"93",
          3099 => x"f0",
          3100 => x"f4",
          3101 => x"52",
          3102 => x"51",
          3103 => x"82",
          3104 => x"54",
          3105 => x"93",
          3106 => x"d8",
          3107 => x"dc",
          3108 => x"52",
          3109 => x"51",
          3110 => x"82",
          3111 => x"54",
          3112 => x"93",
          3113 => x"e0",
          3114 => x"e4",
          3115 => x"52",
          3116 => x"51",
          3117 => x"82",
          3118 => x"54",
          3119 => x"93",
          3120 => x"e8",
          3121 => x"ec",
          3122 => x"52",
          3123 => x"51",
          3124 => x"82",
          3125 => x"54",
          3126 => x"8d",
          3127 => x"a8",
          3128 => x"f3",
          3129 => x"86",
          3130 => x"ab",
          3131 => x"80",
          3132 => x"82",
          3133 => x"52",
          3134 => x"51",
          3135 => x"82",
          3136 => x"54",
          3137 => x"8d",
          3138 => x"aa",
          3139 => x"f4",
          3140 => x"da",
          3141 => x"9d",
          3142 => x"80",
          3143 => x"81",
          3144 => x"87",
          3145 => x"88",
          3146 => x"73",
          3147 => x"38",
          3148 => x"51",
          3149 => x"82",
          3150 => x"54",
          3151 => x"88",
          3152 => x"c8",
          3153 => x"3f",
          3154 => x"33",
          3155 => x"2e",
          3156 => x"f4",
          3157 => x"b2",
          3158 => x"a6",
          3159 => x"80",
          3160 => x"81",
          3161 => x"87",
          3162 => x"f4",
          3163 => x"9a",
          3164 => x"80",
          3165 => x"f4",
          3166 => x"f2",
          3167 => x"84",
          3168 => x"f5",
          3169 => x"e6",
          3170 => x"88",
          3171 => x"f5",
          3172 => x"da",
          3173 => x"f0",
          3174 => x"3f",
          3175 => x"22",
          3176 => x"f8",
          3177 => x"3f",
          3178 => x"08",
          3179 => x"c0",
          3180 => x"e7",
          3181 => x"8c",
          3182 => x"84",
          3183 => x"71",
          3184 => x"82",
          3185 => x"52",
          3186 => x"51",
          3187 => x"82",
          3188 => x"54",
          3189 => x"a8",
          3190 => x"94",
          3191 => x"84",
          3192 => x"51",
          3193 => x"82",
          3194 => x"bd",
          3195 => x"76",
          3196 => x"54",
          3197 => x"08",
          3198 => x"cc",
          3199 => x"3f",
          3200 => x"33",
          3201 => x"2e",
          3202 => x"88",
          3203 => x"bd",
          3204 => x"75",
          3205 => x"3f",
          3206 => x"08",
          3207 => x"29",
          3208 => x"54",
          3209 => x"dc",
          3210 => x"f6",
          3211 => x"be",
          3212 => x"a4",
          3213 => x"3f",
          3214 => x"04",
          3215 => x"02",
          3216 => x"ff",
          3217 => x"84",
          3218 => x"71",
          3219 => x"0b",
          3220 => x"05",
          3221 => x"04",
          3222 => x"51",
          3223 => x"f7",
          3224 => x"39",
          3225 => x"51",
          3226 => x"f7",
          3227 => x"39",
          3228 => x"51",
          3229 => x"f7",
          3230 => x"8e",
          3231 => x"0d",
          3232 => x"80",
          3233 => x"0b",
          3234 => x"84",
          3235 => x"88",
          3236 => x"c0",
          3237 => x"04",
          3238 => x"82",
          3239 => x"89",
          3240 => x"9c",
          3241 => x"ec",
          3242 => x"ec",
          3243 => x"52",
          3244 => x"70",
          3245 => x"26",
          3246 => x"82",
          3247 => x"71",
          3248 => x"8c",
          3249 => x"3d",
          3250 => x"3d",
          3251 => x"84",
          3252 => x"12",
          3253 => x"94",
          3254 => x"16",
          3255 => x"54",
          3256 => x"70",
          3257 => x"38",
          3258 => x"14",
          3259 => x"81",
          3260 => x"76",
          3261 => x"0c",
          3262 => x"75",
          3263 => x"72",
          3264 => x"71",
          3265 => x"70",
          3266 => x"70",
          3267 => x"73",
          3268 => x"74",
          3269 => x"70",
          3270 => x"70",
          3271 => x"8c",
          3272 => x"0c",
          3273 => x"0c",
          3274 => x"0c",
          3275 => x"dc",
          3276 => x"0d",
          3277 => x"0d",
          3278 => x"08",
          3279 => x"56",
          3280 => x"08",
          3281 => x"81",
          3282 => x"84",
          3283 => x"13",
          3284 => x"73",
          3285 => x"06",
          3286 => x"13",
          3287 => x"13",
          3288 => x"13",
          3289 => x"15",
          3290 => x"9f",
          3291 => x"0c",
          3292 => x"08",
          3293 => x"82",
          3294 => x"94",
          3295 => x"82",
          3296 => x"90",
          3297 => x"94",
          3298 => x"73",
          3299 => x"09",
          3300 => x"38",
          3301 => x"70",
          3302 => x"70",
          3303 => x"81",
          3304 => x"84",
          3305 => x"84",
          3306 => x"14",
          3307 => x"08",
          3308 => x"0c",
          3309 => x"0c",
          3310 => x"88",
          3311 => x"88",
          3312 => x"8c",
          3313 => x"82",
          3314 => x"86",
          3315 => x"f9",
          3316 => x"70",
          3317 => x"80",
          3318 => x"38",
          3319 => x"06",
          3320 => x"08",
          3321 => x"08",
          3322 => x"38",
          3323 => x"77",
          3324 => x"38",
          3325 => x"56",
          3326 => x"ff",
          3327 => x"80",
          3328 => x"52",
          3329 => x"3f",
          3330 => x"08",
          3331 => x"08",
          3332 => x"8c",
          3333 => x"80",
          3334 => x"dc",
          3335 => x"30",
          3336 => x"80",
          3337 => x"53",
          3338 => x"54",
          3339 => x"72",
          3340 => x"81",
          3341 => x"38",
          3342 => x"52",
          3343 => x"c8",
          3344 => x"82",
          3345 => x"0c",
          3346 => x"dc",
          3347 => x"0c",
          3348 => x"08",
          3349 => x"82",
          3350 => x"75",
          3351 => x"38",
          3352 => x"53",
          3353 => x"13",
          3354 => x"0c",
          3355 => x"0c",
          3356 => x"0c",
          3357 => x"76",
          3358 => x"53",
          3359 => x"b5",
          3360 => x"82",
          3361 => x"51",
          3362 => x"82",
          3363 => x"54",
          3364 => x"dc",
          3365 => x"0d",
          3366 => x"0d",
          3367 => x"80",
          3368 => x"f0",
          3369 => x"8d",
          3370 => x"0d",
          3371 => x"0d",
          3372 => x"33",
          3373 => x"2e",
          3374 => x"85",
          3375 => x"ed",
          3376 => x"f8",
          3377 => x"80",
          3378 => x"72",
          3379 => x"8c",
          3380 => x"05",
          3381 => x"0c",
          3382 => x"8c",
          3383 => x"71",
          3384 => x"38",
          3385 => x"2d",
          3386 => x"04",
          3387 => x"02",
          3388 => x"82",
          3389 => x"76",
          3390 => x"0c",
          3391 => x"ad",
          3392 => x"8c",
          3393 => x"3d",
          3394 => x"3d",
          3395 => x"73",
          3396 => x"ff",
          3397 => x"71",
          3398 => x"38",
          3399 => x"06",
          3400 => x"54",
          3401 => x"e7",
          3402 => x"0d",
          3403 => x"0d",
          3404 => x"f0",
          3405 => x"8c",
          3406 => x"54",
          3407 => x"81",
          3408 => x"53",
          3409 => x"8e",
          3410 => x"ff",
          3411 => x"14",
          3412 => x"3f",
          3413 => x"82",
          3414 => x"86",
          3415 => x"ec",
          3416 => x"68",
          3417 => x"70",
          3418 => x"33",
          3419 => x"2e",
          3420 => x"75",
          3421 => x"81",
          3422 => x"38",
          3423 => x"70",
          3424 => x"33",
          3425 => x"75",
          3426 => x"81",
          3427 => x"81",
          3428 => x"75",
          3429 => x"81",
          3430 => x"82",
          3431 => x"81",
          3432 => x"56",
          3433 => x"09",
          3434 => x"38",
          3435 => x"71",
          3436 => x"81",
          3437 => x"59",
          3438 => x"9d",
          3439 => x"53",
          3440 => x"95",
          3441 => x"29",
          3442 => x"76",
          3443 => x"79",
          3444 => x"5b",
          3445 => x"e5",
          3446 => x"ec",
          3447 => x"70",
          3448 => x"25",
          3449 => x"32",
          3450 => x"72",
          3451 => x"73",
          3452 => x"58",
          3453 => x"73",
          3454 => x"38",
          3455 => x"79",
          3456 => x"5b",
          3457 => x"75",
          3458 => x"de",
          3459 => x"80",
          3460 => x"89",
          3461 => x"70",
          3462 => x"55",
          3463 => x"cf",
          3464 => x"38",
          3465 => x"24",
          3466 => x"80",
          3467 => x"8e",
          3468 => x"c3",
          3469 => x"73",
          3470 => x"81",
          3471 => x"99",
          3472 => x"c4",
          3473 => x"38",
          3474 => x"73",
          3475 => x"81",
          3476 => x"80",
          3477 => x"38",
          3478 => x"2e",
          3479 => x"f9",
          3480 => x"d8",
          3481 => x"38",
          3482 => x"77",
          3483 => x"08",
          3484 => x"80",
          3485 => x"55",
          3486 => x"8d",
          3487 => x"70",
          3488 => x"51",
          3489 => x"f5",
          3490 => x"2a",
          3491 => x"74",
          3492 => x"53",
          3493 => x"8f",
          3494 => x"fc",
          3495 => x"81",
          3496 => x"80",
          3497 => x"73",
          3498 => x"3f",
          3499 => x"56",
          3500 => x"27",
          3501 => x"a0",
          3502 => x"3f",
          3503 => x"84",
          3504 => x"33",
          3505 => x"93",
          3506 => x"95",
          3507 => x"91",
          3508 => x"8d",
          3509 => x"89",
          3510 => x"fb",
          3511 => x"86",
          3512 => x"2a",
          3513 => x"51",
          3514 => x"2e",
          3515 => x"84",
          3516 => x"86",
          3517 => x"78",
          3518 => x"08",
          3519 => x"32",
          3520 => x"72",
          3521 => x"51",
          3522 => x"74",
          3523 => x"38",
          3524 => x"88",
          3525 => x"7a",
          3526 => x"55",
          3527 => x"3d",
          3528 => x"52",
          3529 => x"e9",
          3530 => x"dc",
          3531 => x"06",
          3532 => x"52",
          3533 => x"3f",
          3534 => x"08",
          3535 => x"27",
          3536 => x"14",
          3537 => x"f8",
          3538 => x"87",
          3539 => x"81",
          3540 => x"b0",
          3541 => x"7d",
          3542 => x"5f",
          3543 => x"75",
          3544 => x"07",
          3545 => x"54",
          3546 => x"26",
          3547 => x"ff",
          3548 => x"84",
          3549 => x"06",
          3550 => x"80",
          3551 => x"96",
          3552 => x"e0",
          3553 => x"73",
          3554 => x"57",
          3555 => x"06",
          3556 => x"54",
          3557 => x"a0",
          3558 => x"2a",
          3559 => x"54",
          3560 => x"38",
          3561 => x"76",
          3562 => x"38",
          3563 => x"fd",
          3564 => x"06",
          3565 => x"38",
          3566 => x"56",
          3567 => x"26",
          3568 => x"3d",
          3569 => x"05",
          3570 => x"ff",
          3571 => x"53",
          3572 => x"d9",
          3573 => x"38",
          3574 => x"56",
          3575 => x"27",
          3576 => x"a0",
          3577 => x"3f",
          3578 => x"3d",
          3579 => x"3d",
          3580 => x"70",
          3581 => x"52",
          3582 => x"73",
          3583 => x"3f",
          3584 => x"04",
          3585 => x"74",
          3586 => x"0c",
          3587 => x"05",
          3588 => x"fa",
          3589 => x"8c",
          3590 => x"80",
          3591 => x"0b",
          3592 => x"0c",
          3593 => x"04",
          3594 => x"82",
          3595 => x"76",
          3596 => x"0c",
          3597 => x"05",
          3598 => x"53",
          3599 => x"72",
          3600 => x"0c",
          3601 => x"04",
          3602 => x"77",
          3603 => x"f4",
          3604 => x"54",
          3605 => x"54",
          3606 => x"80",
          3607 => x"8c",
          3608 => x"71",
          3609 => x"dc",
          3610 => x"06",
          3611 => x"2e",
          3612 => x"72",
          3613 => x"38",
          3614 => x"70",
          3615 => x"25",
          3616 => x"73",
          3617 => x"38",
          3618 => x"86",
          3619 => x"54",
          3620 => x"73",
          3621 => x"ff",
          3622 => x"72",
          3623 => x"74",
          3624 => x"72",
          3625 => x"54",
          3626 => x"81",
          3627 => x"39",
          3628 => x"80",
          3629 => x"51",
          3630 => x"81",
          3631 => x"8c",
          3632 => x"3d",
          3633 => x"3d",
          3634 => x"f4",
          3635 => x"8c",
          3636 => x"53",
          3637 => x"fe",
          3638 => x"82",
          3639 => x"84",
          3640 => x"f8",
          3641 => x"7c",
          3642 => x"70",
          3643 => x"75",
          3644 => x"55",
          3645 => x"2e",
          3646 => x"87",
          3647 => x"76",
          3648 => x"73",
          3649 => x"81",
          3650 => x"81",
          3651 => x"77",
          3652 => x"70",
          3653 => x"58",
          3654 => x"09",
          3655 => x"c2",
          3656 => x"81",
          3657 => x"75",
          3658 => x"55",
          3659 => x"e2",
          3660 => x"90",
          3661 => x"f8",
          3662 => x"8f",
          3663 => x"81",
          3664 => x"75",
          3665 => x"55",
          3666 => x"81",
          3667 => x"27",
          3668 => x"d0",
          3669 => x"55",
          3670 => x"73",
          3671 => x"80",
          3672 => x"14",
          3673 => x"72",
          3674 => x"e0",
          3675 => x"80",
          3676 => x"39",
          3677 => x"55",
          3678 => x"80",
          3679 => x"e0",
          3680 => x"38",
          3681 => x"81",
          3682 => x"53",
          3683 => x"81",
          3684 => x"53",
          3685 => x"8e",
          3686 => x"70",
          3687 => x"55",
          3688 => x"27",
          3689 => x"77",
          3690 => x"74",
          3691 => x"76",
          3692 => x"77",
          3693 => x"70",
          3694 => x"55",
          3695 => x"77",
          3696 => x"38",
          3697 => x"74",
          3698 => x"55",
          3699 => x"dc",
          3700 => x"0d",
          3701 => x"0d",
          3702 => x"56",
          3703 => x"0c",
          3704 => x"70",
          3705 => x"73",
          3706 => x"81",
          3707 => x"81",
          3708 => x"ed",
          3709 => x"2e",
          3710 => x"8e",
          3711 => x"08",
          3712 => x"76",
          3713 => x"56",
          3714 => x"b0",
          3715 => x"06",
          3716 => x"75",
          3717 => x"76",
          3718 => x"70",
          3719 => x"73",
          3720 => x"8b",
          3721 => x"73",
          3722 => x"85",
          3723 => x"82",
          3724 => x"76",
          3725 => x"70",
          3726 => x"ac",
          3727 => x"a0",
          3728 => x"fa",
          3729 => x"53",
          3730 => x"57",
          3731 => x"98",
          3732 => x"39",
          3733 => x"80",
          3734 => x"26",
          3735 => x"86",
          3736 => x"80",
          3737 => x"57",
          3738 => x"74",
          3739 => x"38",
          3740 => x"27",
          3741 => x"14",
          3742 => x"06",
          3743 => x"14",
          3744 => x"06",
          3745 => x"74",
          3746 => x"f9",
          3747 => x"ff",
          3748 => x"89",
          3749 => x"38",
          3750 => x"c5",
          3751 => x"29",
          3752 => x"81",
          3753 => x"76",
          3754 => x"56",
          3755 => x"ba",
          3756 => x"2e",
          3757 => x"30",
          3758 => x"0c",
          3759 => x"82",
          3760 => x"8a",
          3761 => x"fd",
          3762 => x"98",
          3763 => x"2c",
          3764 => x"70",
          3765 => x"10",
          3766 => x"2b",
          3767 => x"54",
          3768 => x"0b",
          3769 => x"12",
          3770 => x"71",
          3771 => x"38",
          3772 => x"11",
          3773 => x"84",
          3774 => x"33",
          3775 => x"52",
          3776 => x"2e",
          3777 => x"83",
          3778 => x"72",
          3779 => x"0c",
          3780 => x"04",
          3781 => x"78",
          3782 => x"9f",
          3783 => x"33",
          3784 => x"71",
          3785 => x"38",
          3786 => x"81",
          3787 => x"f2",
          3788 => x"51",
          3789 => x"72",
          3790 => x"52",
          3791 => x"71",
          3792 => x"52",
          3793 => x"51",
          3794 => x"73",
          3795 => x"3d",
          3796 => x"3d",
          3797 => x"84",
          3798 => x"33",
          3799 => x"bb",
          3800 => x"89",
          3801 => x"84",
          3802 => x"d0",
          3803 => x"51",
          3804 => x"58",
          3805 => x"2e",
          3806 => x"51",
          3807 => x"82",
          3808 => x"70",
          3809 => x"88",
          3810 => x"19",
          3811 => x"56",
          3812 => x"3f",
          3813 => x"08",
          3814 => x"89",
          3815 => x"84",
          3816 => x"d0",
          3817 => x"51",
          3818 => x"80",
          3819 => x"75",
          3820 => x"74",
          3821 => x"3f",
          3822 => x"33",
          3823 => x"74",
          3824 => x"34",
          3825 => x"06",
          3826 => x"27",
          3827 => x"0b",
          3828 => x"34",
          3829 => x"b6",
          3830 => x"a4",
          3831 => x"80",
          3832 => x"82",
          3833 => x"55",
          3834 => x"8c",
          3835 => x"54",
          3836 => x"52",
          3837 => x"c8",
          3838 => x"89",
          3839 => x"8a",
          3840 => x"9e",
          3841 => x"a4",
          3842 => x"cb",
          3843 => x"3d",
          3844 => x"3d",
          3845 => x"80",
          3846 => x"a4",
          3847 => x"d2",
          3848 => x"8c",
          3849 => x"d1",
          3850 => x"a4",
          3851 => x"f8",
          3852 => x"70",
          3853 => x"fa",
          3854 => x"8c",
          3855 => x"2e",
          3856 => x"51",
          3857 => x"82",
          3858 => x"55",
          3859 => x"8c",
          3860 => x"9c",
          3861 => x"dc",
          3862 => x"70",
          3863 => x"80",
          3864 => x"53",
          3865 => x"17",
          3866 => x"52",
          3867 => x"3f",
          3868 => x"09",
          3869 => x"b1",
          3870 => x"0d",
          3871 => x"0d",
          3872 => x"ad",
          3873 => x"5a",
          3874 => x"58",
          3875 => x"89",
          3876 => x"80",
          3877 => x"82",
          3878 => x"81",
          3879 => x"0b",
          3880 => x"08",
          3881 => x"f8",
          3882 => x"70",
          3883 => x"f9",
          3884 => x"8c",
          3885 => x"2e",
          3886 => x"51",
          3887 => x"82",
          3888 => x"81",
          3889 => x"80",
          3890 => x"dc",
          3891 => x"38",
          3892 => x"08",
          3893 => x"17",
          3894 => x"74",
          3895 => x"70",
          3896 => x"07",
          3897 => x"55",
          3898 => x"2e",
          3899 => x"ff",
          3900 => x"89",
          3901 => x"11",
          3902 => x"80",
          3903 => x"82",
          3904 => x"80",
          3905 => x"81",
          3906 => x"ef",
          3907 => x"77",
          3908 => x"06",
          3909 => x"52",
          3910 => x"e6",
          3911 => x"d6",
          3912 => x"3d",
          3913 => x"8c",
          3914 => x"34",
          3915 => x"82",
          3916 => x"a9",
          3917 => x"f6",
          3918 => x"7e",
          3919 => x"72",
          3920 => x"5a",
          3921 => x"2e",
          3922 => x"a2",
          3923 => x"78",
          3924 => x"76",
          3925 => x"81",
          3926 => x"70",
          3927 => x"58",
          3928 => x"2e",
          3929 => x"86",
          3930 => x"26",
          3931 => x"54",
          3932 => x"82",
          3933 => x"70",
          3934 => x"d5",
          3935 => x"8c",
          3936 => x"79",
          3937 => x"51",
          3938 => x"82",
          3939 => x"80",
          3940 => x"15",
          3941 => x"81",
          3942 => x"74",
          3943 => x"38",
          3944 => x"ee",
          3945 => x"81",
          3946 => x"3d",
          3947 => x"f8",
          3948 => x"af",
          3949 => x"dc",
          3950 => x"99",
          3951 => x"78",
          3952 => x"fd",
          3953 => x"8c",
          3954 => x"ff",
          3955 => x"85",
          3956 => x"91",
          3957 => x"70",
          3958 => x"51",
          3959 => x"27",
          3960 => x"80",
          3961 => x"8c",
          3962 => x"3d",
          3963 => x"3d",
          3964 => x"08",
          3965 => x"81",
          3966 => x"5f",
          3967 => x"af",
          3968 => x"89",
          3969 => x"82",
          3970 => x"81",
          3971 => x"89",
          3972 => x"73",
          3973 => x"a8",
          3974 => x"3f",
          3975 => x"08",
          3976 => x"0c",
          3977 => x"08",
          3978 => x"fe",
          3979 => x"82",
          3980 => x"52",
          3981 => x"08",
          3982 => x"3f",
          3983 => x"08",
          3984 => x"38",
          3985 => x"51",
          3986 => x"80",
          3987 => x"89",
          3988 => x"80",
          3989 => x"3d",
          3990 => x"80",
          3991 => x"82",
          3992 => x"56",
          3993 => x"08",
          3994 => x"81",
          3995 => x"38",
          3996 => x"08",
          3997 => x"3f",
          3998 => x"08",
          3999 => x"82",
          4000 => x"25",
          4001 => x"8c",
          4002 => x"05",
          4003 => x"55",
          4004 => x"80",
          4005 => x"ff",
          4006 => x"51",
          4007 => x"74",
          4008 => x"81",
          4009 => x"38",
          4010 => x"0b",
          4011 => x"34",
          4012 => x"dd",
          4013 => x"8c",
          4014 => x"2b",
          4015 => x"51",
          4016 => x"2e",
          4017 => x"81",
          4018 => x"8d",
          4019 => x"98",
          4020 => x"2c",
          4021 => x"33",
          4022 => x"70",
          4023 => x"98",
          4024 => x"84",
          4025 => x"d8",
          4026 => x"15",
          4027 => x"51",
          4028 => x"59",
          4029 => x"58",
          4030 => x"78",
          4031 => x"38",
          4032 => x"b4",
          4033 => x"80",
          4034 => x"ff",
          4035 => x"98",
          4036 => x"80",
          4037 => x"ce",
          4038 => x"74",
          4039 => x"f7",
          4040 => x"8c",
          4041 => x"ff",
          4042 => x"80",
          4043 => x"74",
          4044 => x"34",
          4045 => x"39",
          4046 => x"0a",
          4047 => x"0a",
          4048 => x"2c",
          4049 => x"06",
          4050 => x"73",
          4051 => x"38",
          4052 => x"52",
          4053 => x"ef",
          4054 => x"dc",
          4055 => x"06",
          4056 => x"38",
          4057 => x"56",
          4058 => x"80",
          4059 => x"1c",
          4060 => x"8d",
          4061 => x"98",
          4062 => x"2c",
          4063 => x"33",
          4064 => x"70",
          4065 => x"10",
          4066 => x"2b",
          4067 => x"11",
          4068 => x"51",
          4069 => x"51",
          4070 => x"2e",
          4071 => x"fe",
          4072 => x"f8",
          4073 => x"7d",
          4074 => x"82",
          4075 => x"80",
          4076 => x"fc",
          4077 => x"75",
          4078 => x"34",
          4079 => x"fc",
          4080 => x"3d",
          4081 => x"0c",
          4082 => x"8b",
          4083 => x"38",
          4084 => x"81",
          4085 => x"54",
          4086 => x"82",
          4087 => x"54",
          4088 => x"fd",
          4089 => x"8d",
          4090 => x"73",
          4091 => x"38",
          4092 => x"70",
          4093 => x"55",
          4094 => x"9e",
          4095 => x"54",
          4096 => x"15",
          4097 => x"80",
          4098 => x"ff",
          4099 => x"98",
          4100 => x"88",
          4101 => x"55",
          4102 => x"8d",
          4103 => x"11",
          4104 => x"82",
          4105 => x"73",
          4106 => x"3d",
          4107 => x"82",
          4108 => x"54",
          4109 => x"89",
          4110 => x"54",
          4111 => x"84",
          4112 => x"88",
          4113 => x"80",
          4114 => x"ff",
          4115 => x"98",
          4116 => x"84",
          4117 => x"56",
          4118 => x"25",
          4119 => x"1a",
          4120 => x"54",
          4121 => x"74",
          4122 => x"29",
          4123 => x"05",
          4124 => x"82",
          4125 => x"56",
          4126 => x"75",
          4127 => x"82",
          4128 => x"70",
          4129 => x"98",
          4130 => x"84",
          4131 => x"56",
          4132 => x"25",
          4133 => x"88",
          4134 => x"3f",
          4135 => x"0a",
          4136 => x"0a",
          4137 => x"2c",
          4138 => x"33",
          4139 => x"73",
          4140 => x"38",
          4141 => x"82",
          4142 => x"70",
          4143 => x"55",
          4144 => x"2e",
          4145 => x"82",
          4146 => x"ff",
          4147 => x"82",
          4148 => x"ff",
          4149 => x"82",
          4150 => x"88",
          4151 => x"3f",
          4152 => x"33",
          4153 => x"70",
          4154 => x"8d",
          4155 => x"51",
          4156 => x"74",
          4157 => x"74",
          4158 => x"14",
          4159 => x"73",
          4160 => x"a9",
          4161 => x"80",
          4162 => x"80",
          4163 => x"98",
          4164 => x"84",
          4165 => x"55",
          4166 => x"db",
          4167 => x"e7",
          4168 => x"8d",
          4169 => x"98",
          4170 => x"2c",
          4171 => x"33",
          4172 => x"57",
          4173 => x"fa",
          4174 => x"51",
          4175 => x"74",
          4176 => x"29",
          4177 => x"05",
          4178 => x"82",
          4179 => x"58",
          4180 => x"75",
          4181 => x"fa",
          4182 => x"8d",
          4183 => x"05",
          4184 => x"34",
          4185 => x"c5",
          4186 => x"84",
          4187 => x"f7",
          4188 => x"8c",
          4189 => x"ff",
          4190 => x"98",
          4191 => x"84",
          4192 => x"80",
          4193 => x"38",
          4194 => x"52",
          4195 => x"c2",
          4196 => x"39",
          4197 => x"84",
          4198 => x"8d",
          4199 => x"73",
          4200 => x"8c",
          4201 => x"e6",
          4202 => x"8d",
          4203 => x"05",
          4204 => x"8d",
          4205 => x"81",
          4206 => x"e3",
          4207 => x"88",
          4208 => x"84",
          4209 => x"73",
          4210 => x"e4",
          4211 => x"54",
          4212 => x"84",
          4213 => x"2b",
          4214 => x"75",
          4215 => x"56",
          4216 => x"74",
          4217 => x"74",
          4218 => x"14",
          4219 => x"73",
          4220 => x"b9",
          4221 => x"80",
          4222 => x"80",
          4223 => x"98",
          4224 => x"84",
          4225 => x"55",
          4226 => x"db",
          4227 => x"e5",
          4228 => x"8d",
          4229 => x"98",
          4230 => x"2c",
          4231 => x"33",
          4232 => x"57",
          4233 => x"f9",
          4234 => x"51",
          4235 => x"74",
          4236 => x"29",
          4237 => x"05",
          4238 => x"82",
          4239 => x"58",
          4240 => x"75",
          4241 => x"f8",
          4242 => x"8d",
          4243 => x"81",
          4244 => x"8d",
          4245 => x"56",
          4246 => x"27",
          4247 => x"81",
          4248 => x"82",
          4249 => x"74",
          4250 => x"52",
          4251 => x"3f",
          4252 => x"33",
          4253 => x"06",
          4254 => x"33",
          4255 => x"75",
          4256 => x"38",
          4257 => x"7a",
          4258 => x"89",
          4259 => x"74",
          4260 => x"38",
          4261 => x"d9",
          4262 => x"dc",
          4263 => x"84",
          4264 => x"dc",
          4265 => x"06",
          4266 => x"74",
          4267 => x"c8",
          4268 => x"5b",
          4269 => x"7a",
          4270 => x"88",
          4271 => x"11",
          4272 => x"74",
          4273 => x"38",
          4274 => x"a5",
          4275 => x"dc",
          4276 => x"84",
          4277 => x"dc",
          4278 => x"06",
          4279 => x"74",
          4280 => x"c7",
          4281 => x"1b",
          4282 => x"39",
          4283 => x"74",
          4284 => x"bc",
          4285 => x"ca",
          4286 => x"e2",
          4287 => x"2e",
          4288 => x"93",
          4289 => x"d0",
          4290 => x"80",
          4291 => x"74",
          4292 => x"3f",
          4293 => x"7a",
          4294 => x"88",
          4295 => x"11",
          4296 => x"74",
          4297 => x"38",
          4298 => x"c5",
          4299 => x"dc",
          4300 => x"84",
          4301 => x"dc",
          4302 => x"06",
          4303 => x"74",
          4304 => x"c7",
          4305 => x"1b",
          4306 => x"ff",
          4307 => x"39",
          4308 => x"74",
          4309 => x"d8",
          4310 => x"ca",
          4311 => x"8c",
          4312 => x"8d",
          4313 => x"8c",
          4314 => x"ff",
          4315 => x"53",
          4316 => x"51",
          4317 => x"82",
          4318 => x"82",
          4319 => x"52",
          4320 => x"90",
          4321 => x"39",
          4322 => x"33",
          4323 => x"06",
          4324 => x"33",
          4325 => x"74",
          4326 => x"94",
          4327 => x"54",
          4328 => x"88",
          4329 => x"70",
          4330 => x"e2",
          4331 => x"80",
          4332 => x"88",
          4333 => x"80",
          4334 => x"38",
          4335 => x"ed",
          4336 => x"88",
          4337 => x"54",
          4338 => x"88",
          4339 => x"39",
          4340 => x"8d",
          4341 => x"0b",
          4342 => x"34",
          4343 => x"dc",
          4344 => x"0d",
          4345 => x"0d",
          4346 => x"33",
          4347 => x"70",
          4348 => x"38",
          4349 => x"11",
          4350 => x"82",
          4351 => x"83",
          4352 => x"fc",
          4353 => x"9b",
          4354 => x"84",
          4355 => x"33",
          4356 => x"51",
          4357 => x"80",
          4358 => x"84",
          4359 => x"92",
          4360 => x"51",
          4361 => x"80",
          4362 => x"81",
          4363 => x"72",
          4364 => x"92",
          4365 => x"81",
          4366 => x"0b",
          4367 => x"8c",
          4368 => x"71",
          4369 => x"06",
          4370 => x"80",
          4371 => x"87",
          4372 => x"08",
          4373 => x"38",
          4374 => x"80",
          4375 => x"71",
          4376 => x"c0",
          4377 => x"51",
          4378 => x"87",
          4379 => x"89",
          4380 => x"82",
          4381 => x"33",
          4382 => x"8c",
          4383 => x"3d",
          4384 => x"3d",
          4385 => x"64",
          4386 => x"bf",
          4387 => x"40",
          4388 => x"74",
          4389 => x"cd",
          4390 => x"dc",
          4391 => x"7a",
          4392 => x"81",
          4393 => x"72",
          4394 => x"87",
          4395 => x"11",
          4396 => x"8c",
          4397 => x"92",
          4398 => x"5a",
          4399 => x"58",
          4400 => x"c0",
          4401 => x"76",
          4402 => x"76",
          4403 => x"70",
          4404 => x"81",
          4405 => x"54",
          4406 => x"8e",
          4407 => x"52",
          4408 => x"81",
          4409 => x"81",
          4410 => x"74",
          4411 => x"53",
          4412 => x"83",
          4413 => x"78",
          4414 => x"8f",
          4415 => x"2e",
          4416 => x"c0",
          4417 => x"52",
          4418 => x"87",
          4419 => x"08",
          4420 => x"2e",
          4421 => x"84",
          4422 => x"38",
          4423 => x"87",
          4424 => x"15",
          4425 => x"70",
          4426 => x"52",
          4427 => x"ff",
          4428 => x"39",
          4429 => x"81",
          4430 => x"ff",
          4431 => x"57",
          4432 => x"90",
          4433 => x"80",
          4434 => x"71",
          4435 => x"78",
          4436 => x"38",
          4437 => x"80",
          4438 => x"80",
          4439 => x"81",
          4440 => x"72",
          4441 => x"0c",
          4442 => x"04",
          4443 => x"60",
          4444 => x"8c",
          4445 => x"33",
          4446 => x"5b",
          4447 => x"74",
          4448 => x"e1",
          4449 => x"dc",
          4450 => x"79",
          4451 => x"78",
          4452 => x"06",
          4453 => x"77",
          4454 => x"87",
          4455 => x"11",
          4456 => x"8c",
          4457 => x"92",
          4458 => x"59",
          4459 => x"85",
          4460 => x"98",
          4461 => x"7d",
          4462 => x"0c",
          4463 => x"08",
          4464 => x"70",
          4465 => x"53",
          4466 => x"2e",
          4467 => x"70",
          4468 => x"33",
          4469 => x"18",
          4470 => x"2a",
          4471 => x"51",
          4472 => x"2e",
          4473 => x"c0",
          4474 => x"52",
          4475 => x"87",
          4476 => x"08",
          4477 => x"2e",
          4478 => x"84",
          4479 => x"38",
          4480 => x"87",
          4481 => x"15",
          4482 => x"70",
          4483 => x"52",
          4484 => x"ff",
          4485 => x"39",
          4486 => x"81",
          4487 => x"80",
          4488 => x"52",
          4489 => x"90",
          4490 => x"80",
          4491 => x"71",
          4492 => x"7a",
          4493 => x"38",
          4494 => x"80",
          4495 => x"80",
          4496 => x"81",
          4497 => x"72",
          4498 => x"0c",
          4499 => x"04",
          4500 => x"7a",
          4501 => x"a3",
          4502 => x"88",
          4503 => x"33",
          4504 => x"56",
          4505 => x"3f",
          4506 => x"08",
          4507 => x"83",
          4508 => x"fe",
          4509 => x"87",
          4510 => x"0c",
          4511 => x"76",
          4512 => x"38",
          4513 => x"93",
          4514 => x"2b",
          4515 => x"8c",
          4516 => x"71",
          4517 => x"38",
          4518 => x"71",
          4519 => x"c6",
          4520 => x"39",
          4521 => x"81",
          4522 => x"06",
          4523 => x"71",
          4524 => x"38",
          4525 => x"8c",
          4526 => x"e8",
          4527 => x"98",
          4528 => x"71",
          4529 => x"73",
          4530 => x"92",
          4531 => x"72",
          4532 => x"06",
          4533 => x"f7",
          4534 => x"80",
          4535 => x"88",
          4536 => x"0c",
          4537 => x"80",
          4538 => x"56",
          4539 => x"56",
          4540 => x"82",
          4541 => x"88",
          4542 => x"fe",
          4543 => x"81",
          4544 => x"33",
          4545 => x"07",
          4546 => x"0c",
          4547 => x"3d",
          4548 => x"3d",
          4549 => x"11",
          4550 => x"33",
          4551 => x"71",
          4552 => x"81",
          4553 => x"72",
          4554 => x"75",
          4555 => x"82",
          4556 => x"52",
          4557 => x"54",
          4558 => x"0d",
          4559 => x"0d",
          4560 => x"05",
          4561 => x"52",
          4562 => x"70",
          4563 => x"34",
          4564 => x"51",
          4565 => x"83",
          4566 => x"ff",
          4567 => x"75",
          4568 => x"72",
          4569 => x"54",
          4570 => x"2a",
          4571 => x"70",
          4572 => x"34",
          4573 => x"51",
          4574 => x"81",
          4575 => x"70",
          4576 => x"70",
          4577 => x"3d",
          4578 => x"3d",
          4579 => x"77",
          4580 => x"70",
          4581 => x"38",
          4582 => x"05",
          4583 => x"70",
          4584 => x"34",
          4585 => x"eb",
          4586 => x"0d",
          4587 => x"0d",
          4588 => x"54",
          4589 => x"72",
          4590 => x"54",
          4591 => x"51",
          4592 => x"84",
          4593 => x"fc",
          4594 => x"77",
          4595 => x"53",
          4596 => x"05",
          4597 => x"70",
          4598 => x"33",
          4599 => x"ff",
          4600 => x"52",
          4601 => x"2e",
          4602 => x"80",
          4603 => x"71",
          4604 => x"0c",
          4605 => x"04",
          4606 => x"74",
          4607 => x"89",
          4608 => x"2e",
          4609 => x"11",
          4610 => x"52",
          4611 => x"70",
          4612 => x"dc",
          4613 => x"0d",
          4614 => x"82",
          4615 => x"04",
          4616 => x"8c",
          4617 => x"f7",
          4618 => x"56",
          4619 => x"17",
          4620 => x"74",
          4621 => x"d6",
          4622 => x"b0",
          4623 => x"b4",
          4624 => x"81",
          4625 => x"59",
          4626 => x"82",
          4627 => x"7a",
          4628 => x"06",
          4629 => x"8c",
          4630 => x"17",
          4631 => x"08",
          4632 => x"08",
          4633 => x"08",
          4634 => x"74",
          4635 => x"38",
          4636 => x"55",
          4637 => x"09",
          4638 => x"38",
          4639 => x"18",
          4640 => x"81",
          4641 => x"f9",
          4642 => x"39",
          4643 => x"82",
          4644 => x"8b",
          4645 => x"fa",
          4646 => x"7a",
          4647 => x"57",
          4648 => x"08",
          4649 => x"75",
          4650 => x"3f",
          4651 => x"08",
          4652 => x"dc",
          4653 => x"81",
          4654 => x"b4",
          4655 => x"16",
          4656 => x"be",
          4657 => x"dc",
          4658 => x"85",
          4659 => x"81",
          4660 => x"17",
          4661 => x"8c",
          4662 => x"3d",
          4663 => x"3d",
          4664 => x"52",
          4665 => x"3f",
          4666 => x"08",
          4667 => x"dc",
          4668 => x"38",
          4669 => x"74",
          4670 => x"81",
          4671 => x"38",
          4672 => x"59",
          4673 => x"09",
          4674 => x"e3",
          4675 => x"53",
          4676 => x"08",
          4677 => x"70",
          4678 => x"91",
          4679 => x"d5",
          4680 => x"17",
          4681 => x"3f",
          4682 => x"a4",
          4683 => x"51",
          4684 => x"86",
          4685 => x"f2",
          4686 => x"17",
          4687 => x"3f",
          4688 => x"52",
          4689 => x"51",
          4690 => x"8c",
          4691 => x"84",
          4692 => x"fc",
          4693 => x"17",
          4694 => x"70",
          4695 => x"79",
          4696 => x"52",
          4697 => x"51",
          4698 => x"77",
          4699 => x"80",
          4700 => x"81",
          4701 => x"f9",
          4702 => x"8c",
          4703 => x"2e",
          4704 => x"58",
          4705 => x"dc",
          4706 => x"0d",
          4707 => x"0d",
          4708 => x"98",
          4709 => x"05",
          4710 => x"80",
          4711 => x"27",
          4712 => x"14",
          4713 => x"29",
          4714 => x"05",
          4715 => x"82",
          4716 => x"87",
          4717 => x"f9",
          4718 => x"7a",
          4719 => x"54",
          4720 => x"27",
          4721 => x"76",
          4722 => x"27",
          4723 => x"ff",
          4724 => x"58",
          4725 => x"80",
          4726 => x"82",
          4727 => x"72",
          4728 => x"38",
          4729 => x"72",
          4730 => x"8e",
          4731 => x"39",
          4732 => x"17",
          4733 => x"a4",
          4734 => x"53",
          4735 => x"fd",
          4736 => x"8c",
          4737 => x"9f",
          4738 => x"ff",
          4739 => x"11",
          4740 => x"70",
          4741 => x"18",
          4742 => x"76",
          4743 => x"53",
          4744 => x"82",
          4745 => x"80",
          4746 => x"83",
          4747 => x"b4",
          4748 => x"88",
          4749 => x"79",
          4750 => x"84",
          4751 => x"58",
          4752 => x"80",
          4753 => x"9f",
          4754 => x"80",
          4755 => x"88",
          4756 => x"08",
          4757 => x"51",
          4758 => x"82",
          4759 => x"80",
          4760 => x"10",
          4761 => x"74",
          4762 => x"51",
          4763 => x"82",
          4764 => x"83",
          4765 => x"58",
          4766 => x"87",
          4767 => x"08",
          4768 => x"51",
          4769 => x"82",
          4770 => x"9b",
          4771 => x"2b",
          4772 => x"74",
          4773 => x"51",
          4774 => x"82",
          4775 => x"f0",
          4776 => x"83",
          4777 => x"77",
          4778 => x"0c",
          4779 => x"04",
          4780 => x"7a",
          4781 => x"58",
          4782 => x"81",
          4783 => x"9e",
          4784 => x"17",
          4785 => x"96",
          4786 => x"53",
          4787 => x"81",
          4788 => x"79",
          4789 => x"72",
          4790 => x"38",
          4791 => x"72",
          4792 => x"b8",
          4793 => x"39",
          4794 => x"17",
          4795 => x"a4",
          4796 => x"53",
          4797 => x"fb",
          4798 => x"8c",
          4799 => x"82",
          4800 => x"81",
          4801 => x"83",
          4802 => x"b4",
          4803 => x"78",
          4804 => x"56",
          4805 => x"76",
          4806 => x"38",
          4807 => x"9f",
          4808 => x"33",
          4809 => x"07",
          4810 => x"74",
          4811 => x"83",
          4812 => x"89",
          4813 => x"08",
          4814 => x"51",
          4815 => x"82",
          4816 => x"59",
          4817 => x"08",
          4818 => x"74",
          4819 => x"16",
          4820 => x"84",
          4821 => x"76",
          4822 => x"88",
          4823 => x"81",
          4824 => x"8f",
          4825 => x"53",
          4826 => x"80",
          4827 => x"88",
          4828 => x"08",
          4829 => x"51",
          4830 => x"82",
          4831 => x"59",
          4832 => x"08",
          4833 => x"77",
          4834 => x"06",
          4835 => x"83",
          4836 => x"05",
          4837 => x"f7",
          4838 => x"39",
          4839 => x"a4",
          4840 => x"52",
          4841 => x"ef",
          4842 => x"dc",
          4843 => x"8c",
          4844 => x"38",
          4845 => x"06",
          4846 => x"83",
          4847 => x"18",
          4848 => x"54",
          4849 => x"f6",
          4850 => x"8c",
          4851 => x"0a",
          4852 => x"52",
          4853 => x"83",
          4854 => x"83",
          4855 => x"82",
          4856 => x"8a",
          4857 => x"f8",
          4858 => x"7c",
          4859 => x"59",
          4860 => x"81",
          4861 => x"38",
          4862 => x"08",
          4863 => x"73",
          4864 => x"38",
          4865 => x"52",
          4866 => x"a4",
          4867 => x"dc",
          4868 => x"8c",
          4869 => x"f2",
          4870 => x"82",
          4871 => x"39",
          4872 => x"e6",
          4873 => x"dc",
          4874 => x"de",
          4875 => x"78",
          4876 => x"3f",
          4877 => x"08",
          4878 => x"dc",
          4879 => x"80",
          4880 => x"8c",
          4881 => x"2e",
          4882 => x"8c",
          4883 => x"2e",
          4884 => x"53",
          4885 => x"51",
          4886 => x"82",
          4887 => x"c5",
          4888 => x"08",
          4889 => x"18",
          4890 => x"57",
          4891 => x"90",
          4892 => x"90",
          4893 => x"16",
          4894 => x"54",
          4895 => x"34",
          4896 => x"78",
          4897 => x"38",
          4898 => x"82",
          4899 => x"8a",
          4900 => x"f6",
          4901 => x"7e",
          4902 => x"5b",
          4903 => x"38",
          4904 => x"58",
          4905 => x"88",
          4906 => x"08",
          4907 => x"38",
          4908 => x"39",
          4909 => x"51",
          4910 => x"81",
          4911 => x"8c",
          4912 => x"82",
          4913 => x"8c",
          4914 => x"82",
          4915 => x"ff",
          4916 => x"38",
          4917 => x"82",
          4918 => x"26",
          4919 => x"79",
          4920 => x"08",
          4921 => x"73",
          4922 => x"b9",
          4923 => x"2e",
          4924 => x"80",
          4925 => x"1a",
          4926 => x"08",
          4927 => x"38",
          4928 => x"52",
          4929 => x"af",
          4930 => x"82",
          4931 => x"81",
          4932 => x"06",
          4933 => x"8c",
          4934 => x"82",
          4935 => x"09",
          4936 => x"72",
          4937 => x"70",
          4938 => x"8c",
          4939 => x"51",
          4940 => x"73",
          4941 => x"82",
          4942 => x"80",
          4943 => x"8c",
          4944 => x"81",
          4945 => x"38",
          4946 => x"08",
          4947 => x"73",
          4948 => x"75",
          4949 => x"77",
          4950 => x"56",
          4951 => x"76",
          4952 => x"82",
          4953 => x"26",
          4954 => x"75",
          4955 => x"f8",
          4956 => x"8c",
          4957 => x"2e",
          4958 => x"59",
          4959 => x"08",
          4960 => x"81",
          4961 => x"82",
          4962 => x"59",
          4963 => x"08",
          4964 => x"70",
          4965 => x"25",
          4966 => x"51",
          4967 => x"73",
          4968 => x"75",
          4969 => x"81",
          4970 => x"38",
          4971 => x"f5",
          4972 => x"75",
          4973 => x"f9",
          4974 => x"8c",
          4975 => x"8c",
          4976 => x"70",
          4977 => x"08",
          4978 => x"51",
          4979 => x"80",
          4980 => x"73",
          4981 => x"38",
          4982 => x"52",
          4983 => x"d0",
          4984 => x"dc",
          4985 => x"a5",
          4986 => x"18",
          4987 => x"08",
          4988 => x"18",
          4989 => x"74",
          4990 => x"38",
          4991 => x"18",
          4992 => x"33",
          4993 => x"73",
          4994 => x"97",
          4995 => x"74",
          4996 => x"38",
          4997 => x"55",
          4998 => x"8c",
          4999 => x"85",
          5000 => x"75",
          5001 => x"8c",
          5002 => x"3d",
          5003 => x"3d",
          5004 => x"52",
          5005 => x"3f",
          5006 => x"08",
          5007 => x"82",
          5008 => x"80",
          5009 => x"52",
          5010 => x"c1",
          5011 => x"dc",
          5012 => x"dc",
          5013 => x"0c",
          5014 => x"53",
          5015 => x"15",
          5016 => x"f2",
          5017 => x"56",
          5018 => x"16",
          5019 => x"22",
          5020 => x"27",
          5021 => x"54",
          5022 => x"76",
          5023 => x"33",
          5024 => x"3f",
          5025 => x"08",
          5026 => x"38",
          5027 => x"76",
          5028 => x"70",
          5029 => x"9f",
          5030 => x"56",
          5031 => x"8c",
          5032 => x"3d",
          5033 => x"3d",
          5034 => x"71",
          5035 => x"57",
          5036 => x"0a",
          5037 => x"38",
          5038 => x"53",
          5039 => x"38",
          5040 => x"0c",
          5041 => x"54",
          5042 => x"75",
          5043 => x"73",
          5044 => x"a8",
          5045 => x"73",
          5046 => x"85",
          5047 => x"0b",
          5048 => x"5a",
          5049 => x"27",
          5050 => x"a8",
          5051 => x"18",
          5052 => x"39",
          5053 => x"70",
          5054 => x"58",
          5055 => x"b2",
          5056 => x"76",
          5057 => x"3f",
          5058 => x"08",
          5059 => x"dc",
          5060 => x"bd",
          5061 => x"82",
          5062 => x"27",
          5063 => x"16",
          5064 => x"dc",
          5065 => x"38",
          5066 => x"39",
          5067 => x"55",
          5068 => x"52",
          5069 => x"d5",
          5070 => x"dc",
          5071 => x"0c",
          5072 => x"0c",
          5073 => x"53",
          5074 => x"80",
          5075 => x"85",
          5076 => x"94",
          5077 => x"2a",
          5078 => x"0c",
          5079 => x"06",
          5080 => x"9c",
          5081 => x"58",
          5082 => x"dc",
          5083 => x"0d",
          5084 => x"0d",
          5085 => x"90",
          5086 => x"05",
          5087 => x"f0",
          5088 => x"27",
          5089 => x"0b",
          5090 => x"98",
          5091 => x"84",
          5092 => x"2e",
          5093 => x"76",
          5094 => x"58",
          5095 => x"38",
          5096 => x"15",
          5097 => x"08",
          5098 => x"38",
          5099 => x"88",
          5100 => x"53",
          5101 => x"81",
          5102 => x"c0",
          5103 => x"22",
          5104 => x"89",
          5105 => x"72",
          5106 => x"74",
          5107 => x"f3",
          5108 => x"8c",
          5109 => x"82",
          5110 => x"82",
          5111 => x"27",
          5112 => x"81",
          5113 => x"dc",
          5114 => x"80",
          5115 => x"16",
          5116 => x"dc",
          5117 => x"ca",
          5118 => x"38",
          5119 => x"0c",
          5120 => x"dd",
          5121 => x"08",
          5122 => x"f9",
          5123 => x"8c",
          5124 => x"87",
          5125 => x"dc",
          5126 => x"80",
          5127 => x"55",
          5128 => x"08",
          5129 => x"38",
          5130 => x"8c",
          5131 => x"2e",
          5132 => x"8c",
          5133 => x"75",
          5134 => x"3f",
          5135 => x"08",
          5136 => x"94",
          5137 => x"52",
          5138 => x"c1",
          5139 => x"dc",
          5140 => x"0c",
          5141 => x"0c",
          5142 => x"05",
          5143 => x"80",
          5144 => x"8c",
          5145 => x"3d",
          5146 => x"3d",
          5147 => x"71",
          5148 => x"57",
          5149 => x"51",
          5150 => x"82",
          5151 => x"54",
          5152 => x"08",
          5153 => x"82",
          5154 => x"56",
          5155 => x"52",
          5156 => x"83",
          5157 => x"dc",
          5158 => x"8c",
          5159 => x"d2",
          5160 => x"dc",
          5161 => x"08",
          5162 => x"54",
          5163 => x"e5",
          5164 => x"06",
          5165 => x"58",
          5166 => x"08",
          5167 => x"38",
          5168 => x"75",
          5169 => x"80",
          5170 => x"81",
          5171 => x"7a",
          5172 => x"06",
          5173 => x"39",
          5174 => x"08",
          5175 => x"76",
          5176 => x"3f",
          5177 => x"08",
          5178 => x"dc",
          5179 => x"ff",
          5180 => x"84",
          5181 => x"06",
          5182 => x"54",
          5183 => x"dc",
          5184 => x"0d",
          5185 => x"0d",
          5186 => x"52",
          5187 => x"3f",
          5188 => x"08",
          5189 => x"06",
          5190 => x"51",
          5191 => x"83",
          5192 => x"06",
          5193 => x"14",
          5194 => x"3f",
          5195 => x"08",
          5196 => x"07",
          5197 => x"8c",
          5198 => x"3d",
          5199 => x"3d",
          5200 => x"70",
          5201 => x"06",
          5202 => x"53",
          5203 => x"ed",
          5204 => x"33",
          5205 => x"83",
          5206 => x"06",
          5207 => x"90",
          5208 => x"15",
          5209 => x"3f",
          5210 => x"04",
          5211 => x"7b",
          5212 => x"84",
          5213 => x"58",
          5214 => x"80",
          5215 => x"38",
          5216 => x"52",
          5217 => x"8f",
          5218 => x"dc",
          5219 => x"8c",
          5220 => x"f5",
          5221 => x"08",
          5222 => x"53",
          5223 => x"84",
          5224 => x"39",
          5225 => x"70",
          5226 => x"81",
          5227 => x"51",
          5228 => x"16",
          5229 => x"dc",
          5230 => x"81",
          5231 => x"38",
          5232 => x"ae",
          5233 => x"81",
          5234 => x"54",
          5235 => x"2e",
          5236 => x"8f",
          5237 => x"82",
          5238 => x"76",
          5239 => x"54",
          5240 => x"09",
          5241 => x"38",
          5242 => x"7a",
          5243 => x"80",
          5244 => x"fa",
          5245 => x"8c",
          5246 => x"82",
          5247 => x"89",
          5248 => x"08",
          5249 => x"86",
          5250 => x"98",
          5251 => x"82",
          5252 => x"8b",
          5253 => x"fb",
          5254 => x"70",
          5255 => x"81",
          5256 => x"fc",
          5257 => x"8c",
          5258 => x"82",
          5259 => x"b4",
          5260 => x"08",
          5261 => x"ec",
          5262 => x"8c",
          5263 => x"82",
          5264 => x"a0",
          5265 => x"82",
          5266 => x"52",
          5267 => x"51",
          5268 => x"8b",
          5269 => x"52",
          5270 => x"51",
          5271 => x"81",
          5272 => x"34",
          5273 => x"dc",
          5274 => x"0d",
          5275 => x"0d",
          5276 => x"98",
          5277 => x"70",
          5278 => x"ec",
          5279 => x"8c",
          5280 => x"38",
          5281 => x"53",
          5282 => x"81",
          5283 => x"34",
          5284 => x"04",
          5285 => x"78",
          5286 => x"80",
          5287 => x"34",
          5288 => x"80",
          5289 => x"38",
          5290 => x"18",
          5291 => x"9c",
          5292 => x"70",
          5293 => x"56",
          5294 => x"a0",
          5295 => x"71",
          5296 => x"81",
          5297 => x"81",
          5298 => x"89",
          5299 => x"06",
          5300 => x"73",
          5301 => x"55",
          5302 => x"55",
          5303 => x"81",
          5304 => x"81",
          5305 => x"74",
          5306 => x"75",
          5307 => x"52",
          5308 => x"13",
          5309 => x"08",
          5310 => x"33",
          5311 => x"9c",
          5312 => x"11",
          5313 => x"8a",
          5314 => x"dc",
          5315 => x"96",
          5316 => x"e7",
          5317 => x"dc",
          5318 => x"23",
          5319 => x"e7",
          5320 => x"8c",
          5321 => x"17",
          5322 => x"0d",
          5323 => x"0d",
          5324 => x"5e",
          5325 => x"70",
          5326 => x"55",
          5327 => x"83",
          5328 => x"73",
          5329 => x"91",
          5330 => x"2e",
          5331 => x"1d",
          5332 => x"0c",
          5333 => x"15",
          5334 => x"70",
          5335 => x"56",
          5336 => x"09",
          5337 => x"38",
          5338 => x"80",
          5339 => x"30",
          5340 => x"78",
          5341 => x"54",
          5342 => x"73",
          5343 => x"60",
          5344 => x"54",
          5345 => x"96",
          5346 => x"0b",
          5347 => x"80",
          5348 => x"f6",
          5349 => x"8c",
          5350 => x"85",
          5351 => x"3d",
          5352 => x"5c",
          5353 => x"53",
          5354 => x"51",
          5355 => x"80",
          5356 => x"88",
          5357 => x"5c",
          5358 => x"09",
          5359 => x"d4",
          5360 => x"70",
          5361 => x"71",
          5362 => x"30",
          5363 => x"73",
          5364 => x"51",
          5365 => x"57",
          5366 => x"38",
          5367 => x"75",
          5368 => x"17",
          5369 => x"75",
          5370 => x"30",
          5371 => x"51",
          5372 => x"80",
          5373 => x"38",
          5374 => x"87",
          5375 => x"26",
          5376 => x"77",
          5377 => x"a4",
          5378 => x"27",
          5379 => x"a0",
          5380 => x"39",
          5381 => x"33",
          5382 => x"57",
          5383 => x"27",
          5384 => x"75",
          5385 => x"30",
          5386 => x"32",
          5387 => x"80",
          5388 => x"25",
          5389 => x"56",
          5390 => x"80",
          5391 => x"84",
          5392 => x"58",
          5393 => x"70",
          5394 => x"55",
          5395 => x"09",
          5396 => x"38",
          5397 => x"80",
          5398 => x"30",
          5399 => x"77",
          5400 => x"54",
          5401 => x"81",
          5402 => x"ae",
          5403 => x"06",
          5404 => x"54",
          5405 => x"74",
          5406 => x"80",
          5407 => x"7b",
          5408 => x"30",
          5409 => x"70",
          5410 => x"25",
          5411 => x"07",
          5412 => x"51",
          5413 => x"a7",
          5414 => x"8b",
          5415 => x"39",
          5416 => x"54",
          5417 => x"8c",
          5418 => x"ff",
          5419 => x"ec",
          5420 => x"54",
          5421 => x"e1",
          5422 => x"dc",
          5423 => x"b2",
          5424 => x"70",
          5425 => x"71",
          5426 => x"54",
          5427 => x"82",
          5428 => x"80",
          5429 => x"38",
          5430 => x"76",
          5431 => x"df",
          5432 => x"54",
          5433 => x"81",
          5434 => x"55",
          5435 => x"34",
          5436 => x"52",
          5437 => x"51",
          5438 => x"82",
          5439 => x"bf",
          5440 => x"16",
          5441 => x"26",
          5442 => x"16",
          5443 => x"06",
          5444 => x"17",
          5445 => x"34",
          5446 => x"fd",
          5447 => x"19",
          5448 => x"80",
          5449 => x"79",
          5450 => x"81",
          5451 => x"81",
          5452 => x"85",
          5453 => x"54",
          5454 => x"8f",
          5455 => x"86",
          5456 => x"39",
          5457 => x"f3",
          5458 => x"73",
          5459 => x"80",
          5460 => x"52",
          5461 => x"ce",
          5462 => x"dc",
          5463 => x"8c",
          5464 => x"d7",
          5465 => x"08",
          5466 => x"e6",
          5467 => x"8c",
          5468 => x"82",
          5469 => x"80",
          5470 => x"1b",
          5471 => x"55",
          5472 => x"2e",
          5473 => x"8b",
          5474 => x"06",
          5475 => x"1c",
          5476 => x"33",
          5477 => x"70",
          5478 => x"55",
          5479 => x"38",
          5480 => x"52",
          5481 => x"9f",
          5482 => x"dc",
          5483 => x"8b",
          5484 => x"7a",
          5485 => x"3f",
          5486 => x"75",
          5487 => x"57",
          5488 => x"2e",
          5489 => x"84",
          5490 => x"06",
          5491 => x"75",
          5492 => x"81",
          5493 => x"2a",
          5494 => x"73",
          5495 => x"38",
          5496 => x"54",
          5497 => x"fb",
          5498 => x"80",
          5499 => x"34",
          5500 => x"c1",
          5501 => x"06",
          5502 => x"38",
          5503 => x"39",
          5504 => x"70",
          5505 => x"54",
          5506 => x"86",
          5507 => x"84",
          5508 => x"06",
          5509 => x"73",
          5510 => x"38",
          5511 => x"83",
          5512 => x"b4",
          5513 => x"51",
          5514 => x"82",
          5515 => x"88",
          5516 => x"ea",
          5517 => x"8c",
          5518 => x"3d",
          5519 => x"3d",
          5520 => x"ff",
          5521 => x"71",
          5522 => x"5c",
          5523 => x"80",
          5524 => x"38",
          5525 => x"05",
          5526 => x"a0",
          5527 => x"71",
          5528 => x"38",
          5529 => x"71",
          5530 => x"81",
          5531 => x"38",
          5532 => x"11",
          5533 => x"06",
          5534 => x"70",
          5535 => x"38",
          5536 => x"81",
          5537 => x"05",
          5538 => x"76",
          5539 => x"38",
          5540 => x"fa",
          5541 => x"77",
          5542 => x"57",
          5543 => x"05",
          5544 => x"70",
          5545 => x"33",
          5546 => x"53",
          5547 => x"99",
          5548 => x"e0",
          5549 => x"ff",
          5550 => x"ff",
          5551 => x"70",
          5552 => x"38",
          5553 => x"81",
          5554 => x"51",
          5555 => x"9f",
          5556 => x"72",
          5557 => x"81",
          5558 => x"70",
          5559 => x"72",
          5560 => x"32",
          5561 => x"72",
          5562 => x"73",
          5563 => x"53",
          5564 => x"70",
          5565 => x"38",
          5566 => x"19",
          5567 => x"75",
          5568 => x"38",
          5569 => x"83",
          5570 => x"74",
          5571 => x"59",
          5572 => x"39",
          5573 => x"33",
          5574 => x"8c",
          5575 => x"3d",
          5576 => x"3d",
          5577 => x"80",
          5578 => x"34",
          5579 => x"17",
          5580 => x"75",
          5581 => x"3f",
          5582 => x"8c",
          5583 => x"80",
          5584 => x"16",
          5585 => x"3f",
          5586 => x"08",
          5587 => x"06",
          5588 => x"73",
          5589 => x"2e",
          5590 => x"80",
          5591 => x"0b",
          5592 => x"56",
          5593 => x"e9",
          5594 => x"06",
          5595 => x"57",
          5596 => x"32",
          5597 => x"80",
          5598 => x"51",
          5599 => x"8a",
          5600 => x"e8",
          5601 => x"06",
          5602 => x"53",
          5603 => x"52",
          5604 => x"51",
          5605 => x"82",
          5606 => x"55",
          5607 => x"08",
          5608 => x"38",
          5609 => x"fa",
          5610 => x"86",
          5611 => x"97",
          5612 => x"dc",
          5613 => x"8c",
          5614 => x"2e",
          5615 => x"55",
          5616 => x"dc",
          5617 => x"0d",
          5618 => x"0d",
          5619 => x"05",
          5620 => x"33",
          5621 => x"75",
          5622 => x"fc",
          5623 => x"8c",
          5624 => x"8b",
          5625 => x"82",
          5626 => x"24",
          5627 => x"82",
          5628 => x"84",
          5629 => x"8c",
          5630 => x"55",
          5631 => x"73",
          5632 => x"e6",
          5633 => x"0c",
          5634 => x"06",
          5635 => x"57",
          5636 => x"ae",
          5637 => x"33",
          5638 => x"3f",
          5639 => x"08",
          5640 => x"70",
          5641 => x"55",
          5642 => x"76",
          5643 => x"b8",
          5644 => x"2a",
          5645 => x"51",
          5646 => x"72",
          5647 => x"86",
          5648 => x"74",
          5649 => x"15",
          5650 => x"81",
          5651 => x"d7",
          5652 => x"8c",
          5653 => x"ff",
          5654 => x"06",
          5655 => x"56",
          5656 => x"38",
          5657 => x"8f",
          5658 => x"2a",
          5659 => x"51",
          5660 => x"72",
          5661 => x"80",
          5662 => x"52",
          5663 => x"3f",
          5664 => x"08",
          5665 => x"57",
          5666 => x"09",
          5667 => x"e2",
          5668 => x"74",
          5669 => x"56",
          5670 => x"33",
          5671 => x"72",
          5672 => x"38",
          5673 => x"51",
          5674 => x"82",
          5675 => x"57",
          5676 => x"84",
          5677 => x"ff",
          5678 => x"56",
          5679 => x"25",
          5680 => x"0b",
          5681 => x"56",
          5682 => x"05",
          5683 => x"83",
          5684 => x"2e",
          5685 => x"52",
          5686 => x"c6",
          5687 => x"dc",
          5688 => x"06",
          5689 => x"27",
          5690 => x"16",
          5691 => x"27",
          5692 => x"56",
          5693 => x"84",
          5694 => x"56",
          5695 => x"84",
          5696 => x"14",
          5697 => x"3f",
          5698 => x"08",
          5699 => x"06",
          5700 => x"80",
          5701 => x"06",
          5702 => x"80",
          5703 => x"db",
          5704 => x"8c",
          5705 => x"ff",
          5706 => x"77",
          5707 => x"d8",
          5708 => x"de",
          5709 => x"dc",
          5710 => x"9c",
          5711 => x"c4",
          5712 => x"15",
          5713 => x"14",
          5714 => x"70",
          5715 => x"51",
          5716 => x"56",
          5717 => x"84",
          5718 => x"81",
          5719 => x"71",
          5720 => x"16",
          5721 => x"53",
          5722 => x"23",
          5723 => x"8b",
          5724 => x"73",
          5725 => x"80",
          5726 => x"8d",
          5727 => x"39",
          5728 => x"51",
          5729 => x"82",
          5730 => x"53",
          5731 => x"08",
          5732 => x"72",
          5733 => x"8d",
          5734 => x"ce",
          5735 => x"14",
          5736 => x"3f",
          5737 => x"08",
          5738 => x"06",
          5739 => x"38",
          5740 => x"51",
          5741 => x"82",
          5742 => x"55",
          5743 => x"51",
          5744 => x"82",
          5745 => x"83",
          5746 => x"53",
          5747 => x"80",
          5748 => x"38",
          5749 => x"78",
          5750 => x"2a",
          5751 => x"78",
          5752 => x"86",
          5753 => x"22",
          5754 => x"31",
          5755 => x"ee",
          5756 => x"dc",
          5757 => x"8c",
          5758 => x"2e",
          5759 => x"82",
          5760 => x"80",
          5761 => x"f5",
          5762 => x"83",
          5763 => x"ff",
          5764 => x"38",
          5765 => x"9f",
          5766 => x"38",
          5767 => x"39",
          5768 => x"80",
          5769 => x"38",
          5770 => x"98",
          5771 => x"a0",
          5772 => x"1c",
          5773 => x"0c",
          5774 => x"17",
          5775 => x"76",
          5776 => x"81",
          5777 => x"80",
          5778 => x"d9",
          5779 => x"8c",
          5780 => x"ff",
          5781 => x"8d",
          5782 => x"8e",
          5783 => x"8a",
          5784 => x"14",
          5785 => x"3f",
          5786 => x"08",
          5787 => x"74",
          5788 => x"a2",
          5789 => x"79",
          5790 => x"ee",
          5791 => x"a8",
          5792 => x"15",
          5793 => x"2e",
          5794 => x"10",
          5795 => x"2a",
          5796 => x"05",
          5797 => x"ff",
          5798 => x"53",
          5799 => x"9c",
          5800 => x"81",
          5801 => x"0b",
          5802 => x"ff",
          5803 => x"0c",
          5804 => x"84",
          5805 => x"83",
          5806 => x"06",
          5807 => x"80",
          5808 => x"d8",
          5809 => x"8c",
          5810 => x"ff",
          5811 => x"72",
          5812 => x"81",
          5813 => x"38",
          5814 => x"73",
          5815 => x"3f",
          5816 => x"08",
          5817 => x"82",
          5818 => x"84",
          5819 => x"b2",
          5820 => x"87",
          5821 => x"dc",
          5822 => x"ff",
          5823 => x"82",
          5824 => x"09",
          5825 => x"c8",
          5826 => x"51",
          5827 => x"82",
          5828 => x"84",
          5829 => x"d2",
          5830 => x"06",
          5831 => x"98",
          5832 => x"ee",
          5833 => x"dc",
          5834 => x"85",
          5835 => x"09",
          5836 => x"38",
          5837 => x"51",
          5838 => x"82",
          5839 => x"90",
          5840 => x"a0",
          5841 => x"ca",
          5842 => x"dc",
          5843 => x"0c",
          5844 => x"82",
          5845 => x"81",
          5846 => x"82",
          5847 => x"72",
          5848 => x"80",
          5849 => x"0c",
          5850 => x"82",
          5851 => x"90",
          5852 => x"fb",
          5853 => x"54",
          5854 => x"80",
          5855 => x"73",
          5856 => x"80",
          5857 => x"72",
          5858 => x"80",
          5859 => x"86",
          5860 => x"15",
          5861 => x"71",
          5862 => x"81",
          5863 => x"81",
          5864 => x"d0",
          5865 => x"8c",
          5866 => x"06",
          5867 => x"38",
          5868 => x"54",
          5869 => x"80",
          5870 => x"71",
          5871 => x"82",
          5872 => x"87",
          5873 => x"fa",
          5874 => x"ab",
          5875 => x"58",
          5876 => x"05",
          5877 => x"e6",
          5878 => x"80",
          5879 => x"dc",
          5880 => x"38",
          5881 => x"08",
          5882 => x"8d",
          5883 => x"08",
          5884 => x"80",
          5885 => x"80",
          5886 => x"54",
          5887 => x"84",
          5888 => x"34",
          5889 => x"75",
          5890 => x"2e",
          5891 => x"53",
          5892 => x"53",
          5893 => x"f7",
          5894 => x"8c",
          5895 => x"73",
          5896 => x"0c",
          5897 => x"04",
          5898 => x"67",
          5899 => x"80",
          5900 => x"59",
          5901 => x"78",
          5902 => x"c8",
          5903 => x"06",
          5904 => x"3d",
          5905 => x"99",
          5906 => x"52",
          5907 => x"3f",
          5908 => x"08",
          5909 => x"dc",
          5910 => x"38",
          5911 => x"52",
          5912 => x"52",
          5913 => x"3f",
          5914 => x"08",
          5915 => x"dc",
          5916 => x"02",
          5917 => x"33",
          5918 => x"55",
          5919 => x"25",
          5920 => x"55",
          5921 => x"54",
          5922 => x"81",
          5923 => x"80",
          5924 => x"74",
          5925 => x"81",
          5926 => x"75",
          5927 => x"3f",
          5928 => x"08",
          5929 => x"02",
          5930 => x"91",
          5931 => x"81",
          5932 => x"82",
          5933 => x"06",
          5934 => x"80",
          5935 => x"88",
          5936 => x"39",
          5937 => x"58",
          5938 => x"38",
          5939 => x"70",
          5940 => x"54",
          5941 => x"81",
          5942 => x"52",
          5943 => x"a5",
          5944 => x"dc",
          5945 => x"88",
          5946 => x"62",
          5947 => x"d4",
          5948 => x"54",
          5949 => x"15",
          5950 => x"62",
          5951 => x"e8",
          5952 => x"52",
          5953 => x"51",
          5954 => x"7a",
          5955 => x"83",
          5956 => x"80",
          5957 => x"38",
          5958 => x"08",
          5959 => x"53",
          5960 => x"3d",
          5961 => x"dd",
          5962 => x"8c",
          5963 => x"82",
          5964 => x"82",
          5965 => x"39",
          5966 => x"38",
          5967 => x"33",
          5968 => x"70",
          5969 => x"55",
          5970 => x"2e",
          5971 => x"55",
          5972 => x"77",
          5973 => x"81",
          5974 => x"73",
          5975 => x"38",
          5976 => x"54",
          5977 => x"a0",
          5978 => x"82",
          5979 => x"52",
          5980 => x"a3",
          5981 => x"dc",
          5982 => x"18",
          5983 => x"55",
          5984 => x"dc",
          5985 => x"38",
          5986 => x"70",
          5987 => x"54",
          5988 => x"86",
          5989 => x"c0",
          5990 => x"b0",
          5991 => x"1b",
          5992 => x"1b",
          5993 => x"70",
          5994 => x"d9",
          5995 => x"dc",
          5996 => x"dc",
          5997 => x"0c",
          5998 => x"52",
          5999 => x"3f",
          6000 => x"08",
          6001 => x"08",
          6002 => x"77",
          6003 => x"86",
          6004 => x"1a",
          6005 => x"1a",
          6006 => x"91",
          6007 => x"0b",
          6008 => x"80",
          6009 => x"0c",
          6010 => x"70",
          6011 => x"54",
          6012 => x"81",
          6013 => x"8c",
          6014 => x"2e",
          6015 => x"82",
          6016 => x"94",
          6017 => x"17",
          6018 => x"2b",
          6019 => x"57",
          6020 => x"52",
          6021 => x"9f",
          6022 => x"dc",
          6023 => x"8c",
          6024 => x"26",
          6025 => x"55",
          6026 => x"08",
          6027 => x"81",
          6028 => x"79",
          6029 => x"31",
          6030 => x"70",
          6031 => x"25",
          6032 => x"76",
          6033 => x"81",
          6034 => x"55",
          6035 => x"38",
          6036 => x"0c",
          6037 => x"75",
          6038 => x"54",
          6039 => x"a2",
          6040 => x"7a",
          6041 => x"3f",
          6042 => x"08",
          6043 => x"55",
          6044 => x"89",
          6045 => x"dc",
          6046 => x"1a",
          6047 => x"80",
          6048 => x"54",
          6049 => x"dc",
          6050 => x"0d",
          6051 => x"0d",
          6052 => x"64",
          6053 => x"59",
          6054 => x"90",
          6055 => x"52",
          6056 => x"cf",
          6057 => x"dc",
          6058 => x"8c",
          6059 => x"38",
          6060 => x"55",
          6061 => x"86",
          6062 => x"82",
          6063 => x"19",
          6064 => x"55",
          6065 => x"80",
          6066 => x"38",
          6067 => x"0b",
          6068 => x"82",
          6069 => x"39",
          6070 => x"1a",
          6071 => x"82",
          6072 => x"19",
          6073 => x"08",
          6074 => x"7c",
          6075 => x"74",
          6076 => x"2e",
          6077 => x"94",
          6078 => x"83",
          6079 => x"56",
          6080 => x"38",
          6081 => x"22",
          6082 => x"89",
          6083 => x"55",
          6084 => x"75",
          6085 => x"19",
          6086 => x"39",
          6087 => x"52",
          6088 => x"93",
          6089 => x"dc",
          6090 => x"75",
          6091 => x"38",
          6092 => x"ff",
          6093 => x"98",
          6094 => x"19",
          6095 => x"51",
          6096 => x"82",
          6097 => x"80",
          6098 => x"38",
          6099 => x"08",
          6100 => x"2a",
          6101 => x"80",
          6102 => x"38",
          6103 => x"8a",
          6104 => x"5c",
          6105 => x"27",
          6106 => x"7a",
          6107 => x"54",
          6108 => x"52",
          6109 => x"51",
          6110 => x"82",
          6111 => x"fe",
          6112 => x"83",
          6113 => x"56",
          6114 => x"9f",
          6115 => x"08",
          6116 => x"74",
          6117 => x"38",
          6118 => x"b4",
          6119 => x"16",
          6120 => x"89",
          6121 => x"51",
          6122 => x"77",
          6123 => x"b9",
          6124 => x"1a",
          6125 => x"08",
          6126 => x"84",
          6127 => x"57",
          6128 => x"27",
          6129 => x"56",
          6130 => x"52",
          6131 => x"c7",
          6132 => x"dc",
          6133 => x"38",
          6134 => x"19",
          6135 => x"06",
          6136 => x"52",
          6137 => x"a2",
          6138 => x"31",
          6139 => x"7f",
          6140 => x"94",
          6141 => x"94",
          6142 => x"5c",
          6143 => x"80",
          6144 => x"8c",
          6145 => x"3d",
          6146 => x"3d",
          6147 => x"65",
          6148 => x"5d",
          6149 => x"0c",
          6150 => x"05",
          6151 => x"f6",
          6152 => x"8c",
          6153 => x"82",
          6154 => x"8a",
          6155 => x"33",
          6156 => x"2e",
          6157 => x"56",
          6158 => x"90",
          6159 => x"81",
          6160 => x"06",
          6161 => x"87",
          6162 => x"2e",
          6163 => x"95",
          6164 => x"91",
          6165 => x"56",
          6166 => x"81",
          6167 => x"34",
          6168 => x"8e",
          6169 => x"08",
          6170 => x"56",
          6171 => x"84",
          6172 => x"5c",
          6173 => x"82",
          6174 => x"18",
          6175 => x"ff",
          6176 => x"74",
          6177 => x"7e",
          6178 => x"ff",
          6179 => x"2a",
          6180 => x"7a",
          6181 => x"8c",
          6182 => x"08",
          6183 => x"38",
          6184 => x"39",
          6185 => x"52",
          6186 => x"e7",
          6187 => x"dc",
          6188 => x"8c",
          6189 => x"2e",
          6190 => x"74",
          6191 => x"91",
          6192 => x"2e",
          6193 => x"74",
          6194 => x"88",
          6195 => x"38",
          6196 => x"0c",
          6197 => x"15",
          6198 => x"08",
          6199 => x"06",
          6200 => x"51",
          6201 => x"82",
          6202 => x"fe",
          6203 => x"18",
          6204 => x"51",
          6205 => x"82",
          6206 => x"80",
          6207 => x"38",
          6208 => x"08",
          6209 => x"2a",
          6210 => x"80",
          6211 => x"38",
          6212 => x"8a",
          6213 => x"5b",
          6214 => x"27",
          6215 => x"7b",
          6216 => x"54",
          6217 => x"52",
          6218 => x"51",
          6219 => x"82",
          6220 => x"fe",
          6221 => x"b0",
          6222 => x"31",
          6223 => x"79",
          6224 => x"84",
          6225 => x"16",
          6226 => x"89",
          6227 => x"52",
          6228 => x"cc",
          6229 => x"55",
          6230 => x"16",
          6231 => x"2b",
          6232 => x"39",
          6233 => x"94",
          6234 => x"93",
          6235 => x"cd",
          6236 => x"8c",
          6237 => x"e3",
          6238 => x"b0",
          6239 => x"76",
          6240 => x"94",
          6241 => x"ff",
          6242 => x"71",
          6243 => x"7b",
          6244 => x"38",
          6245 => x"18",
          6246 => x"51",
          6247 => x"82",
          6248 => x"fd",
          6249 => x"53",
          6250 => x"18",
          6251 => x"06",
          6252 => x"51",
          6253 => x"7e",
          6254 => x"83",
          6255 => x"76",
          6256 => x"17",
          6257 => x"1e",
          6258 => x"18",
          6259 => x"0c",
          6260 => x"58",
          6261 => x"74",
          6262 => x"38",
          6263 => x"8c",
          6264 => x"90",
          6265 => x"33",
          6266 => x"55",
          6267 => x"34",
          6268 => x"82",
          6269 => x"90",
          6270 => x"f8",
          6271 => x"8b",
          6272 => x"53",
          6273 => x"f2",
          6274 => x"8c",
          6275 => x"82",
          6276 => x"80",
          6277 => x"16",
          6278 => x"2a",
          6279 => x"51",
          6280 => x"80",
          6281 => x"38",
          6282 => x"52",
          6283 => x"e7",
          6284 => x"dc",
          6285 => x"8c",
          6286 => x"d4",
          6287 => x"08",
          6288 => x"a0",
          6289 => x"73",
          6290 => x"88",
          6291 => x"74",
          6292 => x"51",
          6293 => x"8c",
          6294 => x"9c",
          6295 => x"fb",
          6296 => x"b2",
          6297 => x"15",
          6298 => x"3f",
          6299 => x"15",
          6300 => x"3f",
          6301 => x"0b",
          6302 => x"78",
          6303 => x"3f",
          6304 => x"08",
          6305 => x"81",
          6306 => x"57",
          6307 => x"34",
          6308 => x"dc",
          6309 => x"0d",
          6310 => x"0d",
          6311 => x"54",
          6312 => x"82",
          6313 => x"53",
          6314 => x"08",
          6315 => x"3d",
          6316 => x"73",
          6317 => x"3f",
          6318 => x"08",
          6319 => x"dc",
          6320 => x"82",
          6321 => x"74",
          6322 => x"8c",
          6323 => x"3d",
          6324 => x"3d",
          6325 => x"51",
          6326 => x"8b",
          6327 => x"82",
          6328 => x"24",
          6329 => x"8c",
          6330 => x"8d",
          6331 => x"52",
          6332 => x"dc",
          6333 => x"0d",
          6334 => x"0d",
          6335 => x"3d",
          6336 => x"94",
          6337 => x"c1",
          6338 => x"dc",
          6339 => x"8c",
          6340 => x"e0",
          6341 => x"63",
          6342 => x"d4",
          6343 => x"8d",
          6344 => x"dc",
          6345 => x"8c",
          6346 => x"38",
          6347 => x"05",
          6348 => x"2b",
          6349 => x"80",
          6350 => x"76",
          6351 => x"0c",
          6352 => x"02",
          6353 => x"70",
          6354 => x"81",
          6355 => x"56",
          6356 => x"9e",
          6357 => x"53",
          6358 => x"db",
          6359 => x"8c",
          6360 => x"15",
          6361 => x"82",
          6362 => x"84",
          6363 => x"06",
          6364 => x"55",
          6365 => x"dc",
          6366 => x"0d",
          6367 => x"0d",
          6368 => x"5b",
          6369 => x"80",
          6370 => x"ff",
          6371 => x"9f",
          6372 => x"b5",
          6373 => x"dc",
          6374 => x"8c",
          6375 => x"fc",
          6376 => x"7a",
          6377 => x"08",
          6378 => x"64",
          6379 => x"2e",
          6380 => x"a0",
          6381 => x"70",
          6382 => x"ea",
          6383 => x"dc",
          6384 => x"8c",
          6385 => x"d4",
          6386 => x"7b",
          6387 => x"3f",
          6388 => x"08",
          6389 => x"dc",
          6390 => x"38",
          6391 => x"51",
          6392 => x"82",
          6393 => x"45",
          6394 => x"51",
          6395 => x"82",
          6396 => x"57",
          6397 => x"08",
          6398 => x"80",
          6399 => x"da",
          6400 => x"8c",
          6401 => x"82",
          6402 => x"a4",
          6403 => x"7b",
          6404 => x"3f",
          6405 => x"dc",
          6406 => x"38",
          6407 => x"51",
          6408 => x"82",
          6409 => x"57",
          6410 => x"08",
          6411 => x"38",
          6412 => x"09",
          6413 => x"38",
          6414 => x"e0",
          6415 => x"dc",
          6416 => x"ff",
          6417 => x"74",
          6418 => x"3f",
          6419 => x"78",
          6420 => x"33",
          6421 => x"56",
          6422 => x"91",
          6423 => x"05",
          6424 => x"81",
          6425 => x"56",
          6426 => x"f5",
          6427 => x"54",
          6428 => x"81",
          6429 => x"80",
          6430 => x"78",
          6431 => x"55",
          6432 => x"11",
          6433 => x"18",
          6434 => x"58",
          6435 => x"34",
          6436 => x"ff",
          6437 => x"55",
          6438 => x"34",
          6439 => x"77",
          6440 => x"81",
          6441 => x"ff",
          6442 => x"55",
          6443 => x"34",
          6444 => x"8d",
          6445 => x"84",
          6446 => x"dc",
          6447 => x"70",
          6448 => x"56",
          6449 => x"76",
          6450 => x"81",
          6451 => x"70",
          6452 => x"56",
          6453 => x"82",
          6454 => x"78",
          6455 => x"80",
          6456 => x"27",
          6457 => x"19",
          6458 => x"7a",
          6459 => x"5c",
          6460 => x"55",
          6461 => x"7a",
          6462 => x"5c",
          6463 => x"2e",
          6464 => x"85",
          6465 => x"94",
          6466 => x"81",
          6467 => x"73",
          6468 => x"81",
          6469 => x"7a",
          6470 => x"38",
          6471 => x"76",
          6472 => x"0c",
          6473 => x"04",
          6474 => x"7b",
          6475 => x"fc",
          6476 => x"53",
          6477 => x"bb",
          6478 => x"dc",
          6479 => x"8c",
          6480 => x"fa",
          6481 => x"33",
          6482 => x"f2",
          6483 => x"08",
          6484 => x"27",
          6485 => x"15",
          6486 => x"2a",
          6487 => x"51",
          6488 => x"83",
          6489 => x"94",
          6490 => x"80",
          6491 => x"0c",
          6492 => x"2e",
          6493 => x"79",
          6494 => x"70",
          6495 => x"51",
          6496 => x"2e",
          6497 => x"52",
          6498 => x"fe",
          6499 => x"82",
          6500 => x"ff",
          6501 => x"70",
          6502 => x"fe",
          6503 => x"82",
          6504 => x"73",
          6505 => x"76",
          6506 => x"06",
          6507 => x"0c",
          6508 => x"98",
          6509 => x"58",
          6510 => x"39",
          6511 => x"54",
          6512 => x"73",
          6513 => x"cd",
          6514 => x"8c",
          6515 => x"82",
          6516 => x"81",
          6517 => x"38",
          6518 => x"08",
          6519 => x"9b",
          6520 => x"dc",
          6521 => x"0c",
          6522 => x"0c",
          6523 => x"81",
          6524 => x"76",
          6525 => x"38",
          6526 => x"94",
          6527 => x"94",
          6528 => x"16",
          6529 => x"2a",
          6530 => x"51",
          6531 => x"72",
          6532 => x"38",
          6533 => x"51",
          6534 => x"82",
          6535 => x"54",
          6536 => x"08",
          6537 => x"8c",
          6538 => x"a7",
          6539 => x"74",
          6540 => x"3f",
          6541 => x"08",
          6542 => x"2e",
          6543 => x"74",
          6544 => x"79",
          6545 => x"14",
          6546 => x"38",
          6547 => x"0c",
          6548 => x"94",
          6549 => x"94",
          6550 => x"83",
          6551 => x"72",
          6552 => x"38",
          6553 => x"51",
          6554 => x"82",
          6555 => x"94",
          6556 => x"91",
          6557 => x"53",
          6558 => x"81",
          6559 => x"34",
          6560 => x"39",
          6561 => x"82",
          6562 => x"05",
          6563 => x"08",
          6564 => x"08",
          6565 => x"38",
          6566 => x"0c",
          6567 => x"80",
          6568 => x"72",
          6569 => x"73",
          6570 => x"53",
          6571 => x"8c",
          6572 => x"16",
          6573 => x"38",
          6574 => x"0c",
          6575 => x"82",
          6576 => x"8b",
          6577 => x"f9",
          6578 => x"56",
          6579 => x"80",
          6580 => x"38",
          6581 => x"3d",
          6582 => x"8a",
          6583 => x"51",
          6584 => x"82",
          6585 => x"55",
          6586 => x"08",
          6587 => x"77",
          6588 => x"52",
          6589 => x"b5",
          6590 => x"dc",
          6591 => x"8c",
          6592 => x"c3",
          6593 => x"33",
          6594 => x"55",
          6595 => x"24",
          6596 => x"16",
          6597 => x"2a",
          6598 => x"51",
          6599 => x"80",
          6600 => x"9c",
          6601 => x"77",
          6602 => x"3f",
          6603 => x"08",
          6604 => x"77",
          6605 => x"22",
          6606 => x"74",
          6607 => x"ce",
          6608 => x"8c",
          6609 => x"74",
          6610 => x"81",
          6611 => x"85",
          6612 => x"74",
          6613 => x"38",
          6614 => x"74",
          6615 => x"8c",
          6616 => x"3d",
          6617 => x"3d",
          6618 => x"3d",
          6619 => x"70",
          6620 => x"ff",
          6621 => x"dc",
          6622 => x"82",
          6623 => x"73",
          6624 => x"0d",
          6625 => x"0d",
          6626 => x"3d",
          6627 => x"71",
          6628 => x"e7",
          6629 => x"8c",
          6630 => x"82",
          6631 => x"80",
          6632 => x"93",
          6633 => x"dc",
          6634 => x"51",
          6635 => x"82",
          6636 => x"53",
          6637 => x"82",
          6638 => x"52",
          6639 => x"ac",
          6640 => x"dc",
          6641 => x"8c",
          6642 => x"2e",
          6643 => x"85",
          6644 => x"87",
          6645 => x"dc",
          6646 => x"74",
          6647 => x"d5",
          6648 => x"52",
          6649 => x"89",
          6650 => x"dc",
          6651 => x"70",
          6652 => x"07",
          6653 => x"82",
          6654 => x"06",
          6655 => x"54",
          6656 => x"dc",
          6657 => x"0d",
          6658 => x"0d",
          6659 => x"53",
          6660 => x"53",
          6661 => x"56",
          6662 => x"82",
          6663 => x"55",
          6664 => x"08",
          6665 => x"52",
          6666 => x"81",
          6667 => x"dc",
          6668 => x"8c",
          6669 => x"38",
          6670 => x"05",
          6671 => x"2b",
          6672 => x"80",
          6673 => x"86",
          6674 => x"76",
          6675 => x"38",
          6676 => x"51",
          6677 => x"74",
          6678 => x"0c",
          6679 => x"04",
          6680 => x"63",
          6681 => x"80",
          6682 => x"ec",
          6683 => x"3d",
          6684 => x"3f",
          6685 => x"08",
          6686 => x"dc",
          6687 => x"38",
          6688 => x"73",
          6689 => x"08",
          6690 => x"13",
          6691 => x"58",
          6692 => x"26",
          6693 => x"7c",
          6694 => x"39",
          6695 => x"cc",
          6696 => x"81",
          6697 => x"8c",
          6698 => x"33",
          6699 => x"81",
          6700 => x"06",
          6701 => x"75",
          6702 => x"52",
          6703 => x"05",
          6704 => x"3f",
          6705 => x"08",
          6706 => x"38",
          6707 => x"08",
          6708 => x"38",
          6709 => x"08",
          6710 => x"8c",
          6711 => x"80",
          6712 => x"81",
          6713 => x"59",
          6714 => x"14",
          6715 => x"ca",
          6716 => x"39",
          6717 => x"82",
          6718 => x"57",
          6719 => x"38",
          6720 => x"18",
          6721 => x"ff",
          6722 => x"82",
          6723 => x"5b",
          6724 => x"08",
          6725 => x"7c",
          6726 => x"12",
          6727 => x"52",
          6728 => x"82",
          6729 => x"06",
          6730 => x"14",
          6731 => x"cb",
          6732 => x"dc",
          6733 => x"ff",
          6734 => x"70",
          6735 => x"82",
          6736 => x"51",
          6737 => x"b4",
          6738 => x"bb",
          6739 => x"8c",
          6740 => x"0a",
          6741 => x"70",
          6742 => x"84",
          6743 => x"51",
          6744 => x"ff",
          6745 => x"56",
          6746 => x"38",
          6747 => x"7c",
          6748 => x"0c",
          6749 => x"81",
          6750 => x"74",
          6751 => x"7a",
          6752 => x"0c",
          6753 => x"04",
          6754 => x"79",
          6755 => x"05",
          6756 => x"57",
          6757 => x"82",
          6758 => x"56",
          6759 => x"08",
          6760 => x"91",
          6761 => x"75",
          6762 => x"90",
          6763 => x"81",
          6764 => x"06",
          6765 => x"87",
          6766 => x"2e",
          6767 => x"94",
          6768 => x"73",
          6769 => x"27",
          6770 => x"73",
          6771 => x"8c",
          6772 => x"88",
          6773 => x"76",
          6774 => x"3f",
          6775 => x"08",
          6776 => x"0c",
          6777 => x"39",
          6778 => x"52",
          6779 => x"bf",
          6780 => x"8c",
          6781 => x"2e",
          6782 => x"83",
          6783 => x"82",
          6784 => x"81",
          6785 => x"06",
          6786 => x"56",
          6787 => x"a0",
          6788 => x"82",
          6789 => x"98",
          6790 => x"94",
          6791 => x"08",
          6792 => x"dc",
          6793 => x"51",
          6794 => x"82",
          6795 => x"56",
          6796 => x"8c",
          6797 => x"17",
          6798 => x"07",
          6799 => x"18",
          6800 => x"2e",
          6801 => x"91",
          6802 => x"55",
          6803 => x"dc",
          6804 => x"0d",
          6805 => x"0d",
          6806 => x"3d",
          6807 => x"52",
          6808 => x"da",
          6809 => x"8c",
          6810 => x"82",
          6811 => x"81",
          6812 => x"45",
          6813 => x"52",
          6814 => x"52",
          6815 => x"3f",
          6816 => x"08",
          6817 => x"dc",
          6818 => x"38",
          6819 => x"05",
          6820 => x"2a",
          6821 => x"51",
          6822 => x"55",
          6823 => x"38",
          6824 => x"54",
          6825 => x"81",
          6826 => x"80",
          6827 => x"70",
          6828 => x"54",
          6829 => x"81",
          6830 => x"52",
          6831 => x"c5",
          6832 => x"dc",
          6833 => x"2a",
          6834 => x"51",
          6835 => x"80",
          6836 => x"38",
          6837 => x"8c",
          6838 => x"15",
          6839 => x"86",
          6840 => x"82",
          6841 => x"5c",
          6842 => x"3d",
          6843 => x"c7",
          6844 => x"8c",
          6845 => x"82",
          6846 => x"80",
          6847 => x"8c",
          6848 => x"73",
          6849 => x"3f",
          6850 => x"08",
          6851 => x"dc",
          6852 => x"87",
          6853 => x"39",
          6854 => x"08",
          6855 => x"38",
          6856 => x"08",
          6857 => x"77",
          6858 => x"3f",
          6859 => x"08",
          6860 => x"08",
          6861 => x"8c",
          6862 => x"80",
          6863 => x"55",
          6864 => x"94",
          6865 => x"2e",
          6866 => x"53",
          6867 => x"51",
          6868 => x"82",
          6869 => x"55",
          6870 => x"78",
          6871 => x"fe",
          6872 => x"dc",
          6873 => x"82",
          6874 => x"a0",
          6875 => x"e9",
          6876 => x"53",
          6877 => x"05",
          6878 => x"51",
          6879 => x"82",
          6880 => x"54",
          6881 => x"08",
          6882 => x"78",
          6883 => x"8e",
          6884 => x"58",
          6885 => x"82",
          6886 => x"54",
          6887 => x"08",
          6888 => x"54",
          6889 => x"82",
          6890 => x"84",
          6891 => x"06",
          6892 => x"02",
          6893 => x"33",
          6894 => x"81",
          6895 => x"86",
          6896 => x"f6",
          6897 => x"74",
          6898 => x"70",
          6899 => x"c3",
          6900 => x"dc",
          6901 => x"56",
          6902 => x"08",
          6903 => x"54",
          6904 => x"08",
          6905 => x"81",
          6906 => x"82",
          6907 => x"dc",
          6908 => x"09",
          6909 => x"38",
          6910 => x"b4",
          6911 => x"b0",
          6912 => x"dc",
          6913 => x"51",
          6914 => x"82",
          6915 => x"54",
          6916 => x"08",
          6917 => x"8b",
          6918 => x"b4",
          6919 => x"b7",
          6920 => x"54",
          6921 => x"15",
          6922 => x"90",
          6923 => x"34",
          6924 => x"0a",
          6925 => x"19",
          6926 => x"9f",
          6927 => x"78",
          6928 => x"51",
          6929 => x"a0",
          6930 => x"11",
          6931 => x"05",
          6932 => x"b6",
          6933 => x"ae",
          6934 => x"15",
          6935 => x"78",
          6936 => x"53",
          6937 => x"3f",
          6938 => x"0b",
          6939 => x"77",
          6940 => x"3f",
          6941 => x"08",
          6942 => x"dc",
          6943 => x"82",
          6944 => x"52",
          6945 => x"51",
          6946 => x"3f",
          6947 => x"52",
          6948 => x"aa",
          6949 => x"90",
          6950 => x"34",
          6951 => x"0b",
          6952 => x"78",
          6953 => x"b6",
          6954 => x"dc",
          6955 => x"39",
          6956 => x"52",
          6957 => x"be",
          6958 => x"82",
          6959 => x"99",
          6960 => x"da",
          6961 => x"3d",
          6962 => x"d2",
          6963 => x"53",
          6964 => x"84",
          6965 => x"3d",
          6966 => x"3f",
          6967 => x"08",
          6968 => x"dc",
          6969 => x"38",
          6970 => x"3d",
          6971 => x"3d",
          6972 => x"cc",
          6973 => x"8c",
          6974 => x"82",
          6975 => x"82",
          6976 => x"81",
          6977 => x"81",
          6978 => x"86",
          6979 => x"aa",
          6980 => x"a4",
          6981 => x"a8",
          6982 => x"05",
          6983 => x"ea",
          6984 => x"77",
          6985 => x"70",
          6986 => x"b4",
          6987 => x"3d",
          6988 => x"51",
          6989 => x"82",
          6990 => x"55",
          6991 => x"08",
          6992 => x"6f",
          6993 => x"06",
          6994 => x"a2",
          6995 => x"92",
          6996 => x"81",
          6997 => x"8c",
          6998 => x"2e",
          6999 => x"81",
          7000 => x"51",
          7001 => x"82",
          7002 => x"55",
          7003 => x"08",
          7004 => x"68",
          7005 => x"a8",
          7006 => x"05",
          7007 => x"51",
          7008 => x"3f",
          7009 => x"33",
          7010 => x"8b",
          7011 => x"84",
          7012 => x"06",
          7013 => x"73",
          7014 => x"a0",
          7015 => x"8b",
          7016 => x"54",
          7017 => x"15",
          7018 => x"33",
          7019 => x"70",
          7020 => x"55",
          7021 => x"2e",
          7022 => x"6e",
          7023 => x"df",
          7024 => x"78",
          7025 => x"3f",
          7026 => x"08",
          7027 => x"ff",
          7028 => x"82",
          7029 => x"dc",
          7030 => x"80",
          7031 => x"8c",
          7032 => x"78",
          7033 => x"af",
          7034 => x"dc",
          7035 => x"d4",
          7036 => x"55",
          7037 => x"08",
          7038 => x"81",
          7039 => x"73",
          7040 => x"81",
          7041 => x"63",
          7042 => x"76",
          7043 => x"3f",
          7044 => x"0b",
          7045 => x"87",
          7046 => x"dc",
          7047 => x"77",
          7048 => x"3f",
          7049 => x"08",
          7050 => x"dc",
          7051 => x"78",
          7052 => x"aa",
          7053 => x"dc",
          7054 => x"82",
          7055 => x"a8",
          7056 => x"ed",
          7057 => x"80",
          7058 => x"02",
          7059 => x"df",
          7060 => x"57",
          7061 => x"3d",
          7062 => x"96",
          7063 => x"e9",
          7064 => x"dc",
          7065 => x"8c",
          7066 => x"cf",
          7067 => x"65",
          7068 => x"d4",
          7069 => x"b5",
          7070 => x"dc",
          7071 => x"8c",
          7072 => x"38",
          7073 => x"05",
          7074 => x"06",
          7075 => x"73",
          7076 => x"a7",
          7077 => x"09",
          7078 => x"71",
          7079 => x"06",
          7080 => x"55",
          7081 => x"15",
          7082 => x"81",
          7083 => x"34",
          7084 => x"b4",
          7085 => x"8c",
          7086 => x"74",
          7087 => x"0c",
          7088 => x"04",
          7089 => x"64",
          7090 => x"93",
          7091 => x"52",
          7092 => x"d1",
          7093 => x"8c",
          7094 => x"82",
          7095 => x"80",
          7096 => x"58",
          7097 => x"3d",
          7098 => x"c8",
          7099 => x"8c",
          7100 => x"82",
          7101 => x"b4",
          7102 => x"c7",
          7103 => x"a0",
          7104 => x"55",
          7105 => x"84",
          7106 => x"17",
          7107 => x"2b",
          7108 => x"96",
          7109 => x"b0",
          7110 => x"54",
          7111 => x"15",
          7112 => x"ff",
          7113 => x"82",
          7114 => x"55",
          7115 => x"dc",
          7116 => x"0d",
          7117 => x"0d",
          7118 => x"5a",
          7119 => x"3d",
          7120 => x"99",
          7121 => x"81",
          7122 => x"dc",
          7123 => x"dc",
          7124 => x"82",
          7125 => x"07",
          7126 => x"55",
          7127 => x"2e",
          7128 => x"81",
          7129 => x"55",
          7130 => x"2e",
          7131 => x"7b",
          7132 => x"80",
          7133 => x"70",
          7134 => x"be",
          7135 => x"8c",
          7136 => x"82",
          7137 => x"80",
          7138 => x"52",
          7139 => x"dc",
          7140 => x"dc",
          7141 => x"8c",
          7142 => x"38",
          7143 => x"08",
          7144 => x"08",
          7145 => x"56",
          7146 => x"19",
          7147 => x"59",
          7148 => x"74",
          7149 => x"56",
          7150 => x"ec",
          7151 => x"75",
          7152 => x"74",
          7153 => x"2e",
          7154 => x"16",
          7155 => x"33",
          7156 => x"73",
          7157 => x"38",
          7158 => x"84",
          7159 => x"06",
          7160 => x"7a",
          7161 => x"76",
          7162 => x"07",
          7163 => x"54",
          7164 => x"80",
          7165 => x"80",
          7166 => x"7b",
          7167 => x"53",
          7168 => x"93",
          7169 => x"dc",
          7170 => x"8c",
          7171 => x"38",
          7172 => x"55",
          7173 => x"56",
          7174 => x"8b",
          7175 => x"56",
          7176 => x"83",
          7177 => x"75",
          7178 => x"51",
          7179 => x"3f",
          7180 => x"08",
          7181 => x"82",
          7182 => x"98",
          7183 => x"e6",
          7184 => x"53",
          7185 => x"b8",
          7186 => x"3d",
          7187 => x"3f",
          7188 => x"08",
          7189 => x"08",
          7190 => x"8c",
          7191 => x"98",
          7192 => x"a0",
          7193 => x"70",
          7194 => x"ae",
          7195 => x"6d",
          7196 => x"81",
          7197 => x"57",
          7198 => x"74",
          7199 => x"38",
          7200 => x"81",
          7201 => x"81",
          7202 => x"52",
          7203 => x"89",
          7204 => x"dc",
          7205 => x"a5",
          7206 => x"33",
          7207 => x"54",
          7208 => x"3f",
          7209 => x"08",
          7210 => x"38",
          7211 => x"76",
          7212 => x"05",
          7213 => x"39",
          7214 => x"08",
          7215 => x"15",
          7216 => x"ff",
          7217 => x"73",
          7218 => x"38",
          7219 => x"83",
          7220 => x"56",
          7221 => x"75",
          7222 => x"81",
          7223 => x"33",
          7224 => x"2e",
          7225 => x"52",
          7226 => x"51",
          7227 => x"3f",
          7228 => x"08",
          7229 => x"ff",
          7230 => x"38",
          7231 => x"88",
          7232 => x"8a",
          7233 => x"38",
          7234 => x"ec",
          7235 => x"75",
          7236 => x"74",
          7237 => x"73",
          7238 => x"05",
          7239 => x"17",
          7240 => x"70",
          7241 => x"34",
          7242 => x"70",
          7243 => x"ff",
          7244 => x"55",
          7245 => x"26",
          7246 => x"8b",
          7247 => x"86",
          7248 => x"e5",
          7249 => x"38",
          7250 => x"99",
          7251 => x"05",
          7252 => x"70",
          7253 => x"73",
          7254 => x"81",
          7255 => x"ff",
          7256 => x"ed",
          7257 => x"80",
          7258 => x"91",
          7259 => x"55",
          7260 => x"3f",
          7261 => x"08",
          7262 => x"dc",
          7263 => x"38",
          7264 => x"51",
          7265 => x"3f",
          7266 => x"08",
          7267 => x"dc",
          7268 => x"76",
          7269 => x"67",
          7270 => x"34",
          7271 => x"82",
          7272 => x"84",
          7273 => x"06",
          7274 => x"80",
          7275 => x"2e",
          7276 => x"81",
          7277 => x"ff",
          7278 => x"82",
          7279 => x"54",
          7280 => x"08",
          7281 => x"53",
          7282 => x"08",
          7283 => x"ff",
          7284 => x"67",
          7285 => x"8b",
          7286 => x"53",
          7287 => x"51",
          7288 => x"3f",
          7289 => x"0b",
          7290 => x"79",
          7291 => x"ee",
          7292 => x"dc",
          7293 => x"55",
          7294 => x"dc",
          7295 => x"0d",
          7296 => x"0d",
          7297 => x"88",
          7298 => x"05",
          7299 => x"fc",
          7300 => x"54",
          7301 => x"d2",
          7302 => x"8c",
          7303 => x"82",
          7304 => x"82",
          7305 => x"1a",
          7306 => x"82",
          7307 => x"80",
          7308 => x"8c",
          7309 => x"78",
          7310 => x"1a",
          7311 => x"2a",
          7312 => x"51",
          7313 => x"90",
          7314 => x"82",
          7315 => x"58",
          7316 => x"81",
          7317 => x"39",
          7318 => x"22",
          7319 => x"70",
          7320 => x"56",
          7321 => x"e5",
          7322 => x"14",
          7323 => x"30",
          7324 => x"9f",
          7325 => x"dc",
          7326 => x"19",
          7327 => x"5a",
          7328 => x"81",
          7329 => x"38",
          7330 => x"77",
          7331 => x"82",
          7332 => x"56",
          7333 => x"74",
          7334 => x"ff",
          7335 => x"81",
          7336 => x"55",
          7337 => x"75",
          7338 => x"82",
          7339 => x"dc",
          7340 => x"ff",
          7341 => x"8c",
          7342 => x"2e",
          7343 => x"82",
          7344 => x"8e",
          7345 => x"56",
          7346 => x"09",
          7347 => x"38",
          7348 => x"59",
          7349 => x"77",
          7350 => x"06",
          7351 => x"87",
          7352 => x"39",
          7353 => x"ba",
          7354 => x"55",
          7355 => x"2e",
          7356 => x"15",
          7357 => x"2e",
          7358 => x"83",
          7359 => x"75",
          7360 => x"7e",
          7361 => x"a8",
          7362 => x"dc",
          7363 => x"8c",
          7364 => x"ce",
          7365 => x"16",
          7366 => x"56",
          7367 => x"38",
          7368 => x"19",
          7369 => x"8c",
          7370 => x"7d",
          7371 => x"38",
          7372 => x"0c",
          7373 => x"0c",
          7374 => x"80",
          7375 => x"73",
          7376 => x"98",
          7377 => x"05",
          7378 => x"57",
          7379 => x"26",
          7380 => x"7b",
          7381 => x"0c",
          7382 => x"81",
          7383 => x"84",
          7384 => x"54",
          7385 => x"dc",
          7386 => x"0d",
          7387 => x"0d",
          7388 => x"88",
          7389 => x"05",
          7390 => x"54",
          7391 => x"c5",
          7392 => x"56",
          7393 => x"8c",
          7394 => x"8b",
          7395 => x"8c",
          7396 => x"29",
          7397 => x"05",
          7398 => x"55",
          7399 => x"84",
          7400 => x"34",
          7401 => x"08",
          7402 => x"5f",
          7403 => x"51",
          7404 => x"3f",
          7405 => x"08",
          7406 => x"70",
          7407 => x"57",
          7408 => x"8b",
          7409 => x"82",
          7410 => x"06",
          7411 => x"56",
          7412 => x"38",
          7413 => x"05",
          7414 => x"7e",
          7415 => x"f0",
          7416 => x"dc",
          7417 => x"67",
          7418 => x"2e",
          7419 => x"82",
          7420 => x"8b",
          7421 => x"75",
          7422 => x"80",
          7423 => x"81",
          7424 => x"2e",
          7425 => x"80",
          7426 => x"38",
          7427 => x"0a",
          7428 => x"ff",
          7429 => x"55",
          7430 => x"86",
          7431 => x"8a",
          7432 => x"89",
          7433 => x"2a",
          7434 => x"77",
          7435 => x"59",
          7436 => x"81",
          7437 => x"70",
          7438 => x"07",
          7439 => x"56",
          7440 => x"38",
          7441 => x"05",
          7442 => x"7e",
          7443 => x"80",
          7444 => x"82",
          7445 => x"8a",
          7446 => x"83",
          7447 => x"06",
          7448 => x"08",
          7449 => x"74",
          7450 => x"41",
          7451 => x"56",
          7452 => x"8a",
          7453 => x"61",
          7454 => x"55",
          7455 => x"27",
          7456 => x"93",
          7457 => x"80",
          7458 => x"38",
          7459 => x"70",
          7460 => x"43",
          7461 => x"95",
          7462 => x"06",
          7463 => x"2e",
          7464 => x"77",
          7465 => x"74",
          7466 => x"83",
          7467 => x"06",
          7468 => x"82",
          7469 => x"2e",
          7470 => x"78",
          7471 => x"2e",
          7472 => x"80",
          7473 => x"ae",
          7474 => x"2a",
          7475 => x"81",
          7476 => x"56",
          7477 => x"2e",
          7478 => x"77",
          7479 => x"81",
          7480 => x"79",
          7481 => x"70",
          7482 => x"5a",
          7483 => x"86",
          7484 => x"27",
          7485 => x"52",
          7486 => x"e0",
          7487 => x"8c",
          7488 => x"29",
          7489 => x"70",
          7490 => x"55",
          7491 => x"0b",
          7492 => x"08",
          7493 => x"05",
          7494 => x"ff",
          7495 => x"27",
          7496 => x"88",
          7497 => x"ae",
          7498 => x"2a",
          7499 => x"81",
          7500 => x"56",
          7501 => x"2e",
          7502 => x"77",
          7503 => x"81",
          7504 => x"79",
          7505 => x"70",
          7506 => x"5a",
          7507 => x"86",
          7508 => x"27",
          7509 => x"52",
          7510 => x"e0",
          7511 => x"8c",
          7512 => x"84",
          7513 => x"8c",
          7514 => x"f5",
          7515 => x"81",
          7516 => x"dc",
          7517 => x"8c",
          7518 => x"71",
          7519 => x"83",
          7520 => x"5e",
          7521 => x"89",
          7522 => x"5c",
          7523 => x"1c",
          7524 => x"05",
          7525 => x"ff",
          7526 => x"70",
          7527 => x"31",
          7528 => x"57",
          7529 => x"83",
          7530 => x"06",
          7531 => x"1c",
          7532 => x"5c",
          7533 => x"1d",
          7534 => x"29",
          7535 => x"31",
          7536 => x"55",
          7537 => x"87",
          7538 => x"7c",
          7539 => x"7a",
          7540 => x"31",
          7541 => x"df",
          7542 => x"8c",
          7543 => x"7d",
          7544 => x"81",
          7545 => x"82",
          7546 => x"83",
          7547 => x"80",
          7548 => x"87",
          7549 => x"81",
          7550 => x"fd",
          7551 => x"f8",
          7552 => x"2e",
          7553 => x"80",
          7554 => x"ff",
          7555 => x"8c",
          7556 => x"a0",
          7557 => x"38",
          7558 => x"74",
          7559 => x"86",
          7560 => x"fd",
          7561 => x"81",
          7562 => x"80",
          7563 => x"83",
          7564 => x"39",
          7565 => x"08",
          7566 => x"92",
          7567 => x"b8",
          7568 => x"59",
          7569 => x"27",
          7570 => x"86",
          7571 => x"55",
          7572 => x"09",
          7573 => x"38",
          7574 => x"f5",
          7575 => x"38",
          7576 => x"55",
          7577 => x"86",
          7578 => x"80",
          7579 => x"7a",
          7580 => x"b9",
          7581 => x"81",
          7582 => x"7a",
          7583 => x"8a",
          7584 => x"52",
          7585 => x"ff",
          7586 => x"79",
          7587 => x"7b",
          7588 => x"06",
          7589 => x"51",
          7590 => x"3f",
          7591 => x"1c",
          7592 => x"32",
          7593 => x"96",
          7594 => x"06",
          7595 => x"91",
          7596 => x"a1",
          7597 => x"55",
          7598 => x"ff",
          7599 => x"74",
          7600 => x"06",
          7601 => x"51",
          7602 => x"3f",
          7603 => x"52",
          7604 => x"ff",
          7605 => x"f8",
          7606 => x"34",
          7607 => x"1b",
          7608 => x"d9",
          7609 => x"52",
          7610 => x"ff",
          7611 => x"60",
          7612 => x"51",
          7613 => x"3f",
          7614 => x"09",
          7615 => x"cb",
          7616 => x"b2",
          7617 => x"c3",
          7618 => x"a0",
          7619 => x"52",
          7620 => x"ff",
          7621 => x"82",
          7622 => x"51",
          7623 => x"3f",
          7624 => x"1b",
          7625 => x"95",
          7626 => x"b2",
          7627 => x"a0",
          7628 => x"80",
          7629 => x"1c",
          7630 => x"80",
          7631 => x"93",
          7632 => x"b4",
          7633 => x"1b",
          7634 => x"82",
          7635 => x"52",
          7636 => x"ff",
          7637 => x"7c",
          7638 => x"06",
          7639 => x"51",
          7640 => x"3f",
          7641 => x"a4",
          7642 => x"0b",
          7643 => x"93",
          7644 => x"c8",
          7645 => x"51",
          7646 => x"3f",
          7647 => x"52",
          7648 => x"70",
          7649 => x"9f",
          7650 => x"54",
          7651 => x"52",
          7652 => x"9b",
          7653 => x"56",
          7654 => x"08",
          7655 => x"7d",
          7656 => x"81",
          7657 => x"38",
          7658 => x"86",
          7659 => x"52",
          7660 => x"9b",
          7661 => x"80",
          7662 => x"7a",
          7663 => x"ed",
          7664 => x"85",
          7665 => x"7a",
          7666 => x"8f",
          7667 => x"85",
          7668 => x"83",
          7669 => x"ff",
          7670 => x"ff",
          7671 => x"e8",
          7672 => x"9e",
          7673 => x"52",
          7674 => x"51",
          7675 => x"3f",
          7676 => x"52",
          7677 => x"9e",
          7678 => x"54",
          7679 => x"53",
          7680 => x"51",
          7681 => x"3f",
          7682 => x"16",
          7683 => x"7e",
          7684 => x"d8",
          7685 => x"80",
          7686 => x"ff",
          7687 => x"7f",
          7688 => x"7d",
          7689 => x"81",
          7690 => x"f8",
          7691 => x"ff",
          7692 => x"ff",
          7693 => x"51",
          7694 => x"3f",
          7695 => x"88",
          7696 => x"39",
          7697 => x"f8",
          7698 => x"2e",
          7699 => x"55",
          7700 => x"51",
          7701 => x"3f",
          7702 => x"57",
          7703 => x"83",
          7704 => x"76",
          7705 => x"7a",
          7706 => x"ff",
          7707 => x"82",
          7708 => x"82",
          7709 => x"80",
          7710 => x"dc",
          7711 => x"51",
          7712 => x"3f",
          7713 => x"78",
          7714 => x"74",
          7715 => x"18",
          7716 => x"2e",
          7717 => x"79",
          7718 => x"2e",
          7719 => x"55",
          7720 => x"62",
          7721 => x"74",
          7722 => x"75",
          7723 => x"7e",
          7724 => x"b8",
          7725 => x"dc",
          7726 => x"38",
          7727 => x"78",
          7728 => x"74",
          7729 => x"56",
          7730 => x"93",
          7731 => x"66",
          7732 => x"26",
          7733 => x"56",
          7734 => x"83",
          7735 => x"64",
          7736 => x"77",
          7737 => x"84",
          7738 => x"52",
          7739 => x"9d",
          7740 => x"d4",
          7741 => x"51",
          7742 => x"3f",
          7743 => x"55",
          7744 => x"81",
          7745 => x"34",
          7746 => x"16",
          7747 => x"16",
          7748 => x"16",
          7749 => x"05",
          7750 => x"c1",
          7751 => x"fe",
          7752 => x"fe",
          7753 => x"34",
          7754 => x"08",
          7755 => x"07",
          7756 => x"16",
          7757 => x"dc",
          7758 => x"34",
          7759 => x"c6",
          7760 => x"9c",
          7761 => x"52",
          7762 => x"51",
          7763 => x"3f",
          7764 => x"53",
          7765 => x"51",
          7766 => x"3f",
          7767 => x"8c",
          7768 => x"38",
          7769 => x"52",
          7770 => x"99",
          7771 => x"56",
          7772 => x"08",
          7773 => x"39",
          7774 => x"39",
          7775 => x"39",
          7776 => x"08",
          7777 => x"8c",
          7778 => x"3d",
          7779 => x"3d",
          7780 => x"5b",
          7781 => x"60",
          7782 => x"57",
          7783 => x"25",
          7784 => x"3d",
          7785 => x"55",
          7786 => x"15",
          7787 => x"c9",
          7788 => x"81",
          7789 => x"06",
          7790 => x"3d",
          7791 => x"8d",
          7792 => x"74",
          7793 => x"05",
          7794 => x"17",
          7795 => x"2e",
          7796 => x"c9",
          7797 => x"34",
          7798 => x"83",
          7799 => x"74",
          7800 => x"0c",
          7801 => x"04",
          7802 => x"7b",
          7803 => x"b3",
          7804 => x"57",
          7805 => x"09",
          7806 => x"38",
          7807 => x"51",
          7808 => x"17",
          7809 => x"76",
          7810 => x"88",
          7811 => x"17",
          7812 => x"59",
          7813 => x"81",
          7814 => x"76",
          7815 => x"8b",
          7816 => x"54",
          7817 => x"17",
          7818 => x"51",
          7819 => x"79",
          7820 => x"30",
          7821 => x"9f",
          7822 => x"53",
          7823 => x"75",
          7824 => x"81",
          7825 => x"0c",
          7826 => x"04",
          7827 => x"79",
          7828 => x"56",
          7829 => x"24",
          7830 => x"3d",
          7831 => x"74",
          7832 => x"52",
          7833 => x"cb",
          7834 => x"8c",
          7835 => x"38",
          7836 => x"78",
          7837 => x"06",
          7838 => x"16",
          7839 => x"39",
          7840 => x"82",
          7841 => x"89",
          7842 => x"fd",
          7843 => x"54",
          7844 => x"80",
          7845 => x"ff",
          7846 => x"76",
          7847 => x"3d",
          7848 => x"3d",
          7849 => x"e3",
          7850 => x"53",
          7851 => x"53",
          7852 => x"3f",
          7853 => x"51",
          7854 => x"72",
          7855 => x"3f",
          7856 => x"04",
          7857 => x"7a",
          7858 => x"56",
          7859 => x"80",
          7860 => x"38",
          7861 => x"15",
          7862 => x"16",
          7863 => x"d4",
          7864 => x"54",
          7865 => x"09",
          7866 => x"38",
          7867 => x"f1",
          7868 => x"76",
          7869 => x"89",
          7870 => x"08",
          7871 => x"da",
          7872 => x"8c",
          7873 => x"8c",
          7874 => x"75",
          7875 => x"52",
          7876 => x"be",
          7877 => x"dc",
          7878 => x"84",
          7879 => x"73",
          7880 => x"b2",
          7881 => x"70",
          7882 => x"58",
          7883 => x"27",
          7884 => x"54",
          7885 => x"dc",
          7886 => x"0d",
          7887 => x"0d",
          7888 => x"93",
          7889 => x"38",
          7890 => x"81",
          7891 => x"52",
          7892 => x"81",
          7893 => x"81",
          7894 => x"fd",
          7895 => x"f9",
          7896 => x"e8",
          7897 => x"39",
          7898 => x"51",
          7899 => x"81",
          7900 => x"80",
          7901 => x"fe",
          7902 => x"dd",
          7903 => x"b0",
          7904 => x"39",
          7905 => x"51",
          7906 => x"81",
          7907 => x"80",
          7908 => x"fe",
          7909 => x"c1",
          7910 => x"88",
          7911 => x"81",
          7912 => x"b5",
          7913 => x"b8",
          7914 => x"81",
          7915 => x"a9",
          7916 => x"f8",
          7917 => x"82",
          7918 => x"9d",
          7919 => x"ac",
          7920 => x"82",
          7921 => x"91",
          7922 => x"dc",
          7923 => x"82",
          7924 => x"85",
          7925 => x"80",
          7926 => x"ae",
          7927 => x"0d",
          7928 => x"0d",
          7929 => x"56",
          7930 => x"26",
          7931 => x"52",
          7932 => x"29",
          7933 => x"87",
          7934 => x"51",
          7935 => x"3f",
          7936 => x"08",
          7937 => x"fe",
          7938 => x"82",
          7939 => x"54",
          7940 => x"52",
          7941 => x"51",
          7942 => x"3f",
          7943 => x"04",
          7944 => x"66",
          7945 => x"80",
          7946 => x"5b",
          7947 => x"78",
          7948 => x"07",
          7949 => x"57",
          7950 => x"56",
          7951 => x"26",
          7952 => x"56",
          7953 => x"70",
          7954 => x"51",
          7955 => x"74",
          7956 => x"81",
          7957 => x"8c",
          7958 => x"56",
          7959 => x"3f",
          7960 => x"08",
          7961 => x"dc",
          7962 => x"82",
          7963 => x"87",
          7964 => x"0c",
          7965 => x"08",
          7966 => x"d4",
          7967 => x"80",
          7968 => x"75",
          7969 => x"3f",
          7970 => x"08",
          7971 => x"dc",
          7972 => x"7a",
          7973 => x"2e",
          7974 => x"19",
          7975 => x"59",
          7976 => x"3d",
          7977 => x"cb",
          7978 => x"30",
          7979 => x"80",
          7980 => x"70",
          7981 => x"06",
          7982 => x"56",
          7983 => x"90",
          7984 => x"b4",
          7985 => x"98",
          7986 => x"78",
          7987 => x"3f",
          7988 => x"82",
          7989 => x"96",
          7990 => x"f9",
          7991 => x"02",
          7992 => x"05",
          7993 => x"ff",
          7994 => x"7a",
          7995 => x"fe",
          7996 => x"8c",
          7997 => x"38",
          7998 => x"88",
          7999 => x"2e",
          8000 => x"39",
          8001 => x"54",
          8002 => x"53",
          8003 => x"51",
          8004 => x"8c",
          8005 => x"83",
          8006 => x"76",
          8007 => x"0c",
          8008 => x"04",
          8009 => x"7f",
          8010 => x"8c",
          8011 => x"05",
          8012 => x"15",
          8013 => x"5c",
          8014 => x"5e",
          8015 => x"81",
          8016 => x"f5",
          8017 => x"81",
          8018 => x"ef",
          8019 => x"55",
          8020 => x"80",
          8021 => x"90",
          8022 => x"7b",
          8023 => x"38",
          8024 => x"74",
          8025 => x"7a",
          8026 => x"72",
          8027 => x"81",
          8028 => x"f4",
          8029 => x"39",
          8030 => x"51",
          8031 => x"3f",
          8032 => x"80",
          8033 => x"18",
          8034 => x"27",
          8035 => x"08",
          8036 => x"bc",
          8037 => x"d6",
          8038 => x"82",
          8039 => x"fe",
          8040 => x"84",
          8041 => x"39",
          8042 => x"72",
          8043 => x"38",
          8044 => x"82",
          8045 => x"fe",
          8046 => x"89",
          8047 => x"e4",
          8048 => x"c6",
          8049 => x"55",
          8050 => x"ed",
          8051 => x"80",
          8052 => x"e8",
          8053 => x"b2",
          8054 => x"74",
          8055 => x"38",
          8056 => x"33",
          8057 => x"56",
          8058 => x"83",
          8059 => x"80",
          8060 => x"27",
          8061 => x"53",
          8062 => x"70",
          8063 => x"51",
          8064 => x"2e",
          8065 => x"80",
          8066 => x"38",
          8067 => x"39",
          8068 => x"ed",
          8069 => x"15",
          8070 => x"82",
          8071 => x"fe",
          8072 => x"78",
          8073 => x"5c",
          8074 => x"d5",
          8075 => x"dc",
          8076 => x"70",
          8077 => x"57",
          8078 => x"09",
          8079 => x"38",
          8080 => x"3f",
          8081 => x"08",
          8082 => x"98",
          8083 => x"32",
          8084 => x"9b",
          8085 => x"70",
          8086 => x"75",
          8087 => x"58",
          8088 => x"51",
          8089 => x"24",
          8090 => x"9b",
          8091 => x"06",
          8092 => x"53",
          8093 => x"1e",
          8094 => x"26",
          8095 => x"ff",
          8096 => x"8c",
          8097 => x"3d",
          8098 => x"3d",
          8099 => x"05",
          8100 => x"f0",
          8101 => x"f4",
          8102 => x"f2",
          8103 => x"88",
          8104 => x"fe",
          8105 => x"82",
          8106 => x"82",
          8107 => x"82",
          8108 => x"52",
          8109 => x"51",
          8110 => x"3f",
          8111 => x"85",
          8112 => x"e1",
          8113 => x"0d",
          8114 => x"0d",
          8115 => x"80",
          8116 => x"e7",
          8117 => x"51",
          8118 => x"3f",
          8119 => x"51",
          8120 => x"3f",
          8121 => x"d9",
          8122 => x"81",
          8123 => x"06",
          8124 => x"80",
          8125 => x"81",
          8126 => x"99",
          8127 => x"c8",
          8128 => x"91",
          8129 => x"fe",
          8130 => x"72",
          8131 => x"81",
          8132 => x"71",
          8133 => x"38",
          8134 => x"d8",
          8135 => x"82",
          8136 => x"da",
          8137 => x"51",
          8138 => x"3f",
          8139 => x"70",
          8140 => x"52",
          8141 => x"95",
          8142 => x"fe",
          8143 => x"82",
          8144 => x"fe",
          8145 => x"80",
          8146 => x"c9",
          8147 => x"2a",
          8148 => x"51",
          8149 => x"2e",
          8150 => x"51",
          8151 => x"3f",
          8152 => x"51",
          8153 => x"3f",
          8154 => x"d8",
          8155 => x"85",
          8156 => x"06",
          8157 => x"80",
          8158 => x"81",
          8159 => x"95",
          8160 => x"94",
          8161 => x"8d",
          8162 => x"fe",
          8163 => x"72",
          8164 => x"81",
          8165 => x"71",
          8166 => x"38",
          8167 => x"d7",
          8168 => x"83",
          8169 => x"d9",
          8170 => x"51",
          8171 => x"3f",
          8172 => x"70",
          8173 => x"52",
          8174 => x"95",
          8175 => x"fe",
          8176 => x"82",
          8177 => x"fe",
          8178 => x"80",
          8179 => x"c5",
          8180 => x"2a",
          8181 => x"51",
          8182 => x"2e",
          8183 => x"51",
          8184 => x"3f",
          8185 => x"51",
          8186 => x"3f",
          8187 => x"d7",
          8188 => x"e5",
          8189 => x"3d",
          8190 => x"3d",
          8191 => x"84",
          8192 => x"33",
          8193 => x"56",
          8194 => x"51",
          8195 => x"3f",
          8196 => x"33",
          8197 => x"38",
          8198 => x"84",
          8199 => x"a3",
          8200 => x"b8",
          8201 => x"8c",
          8202 => x"70",
          8203 => x"08",
          8204 => x"82",
          8205 => x"51",
          8206 => x"89",
          8207 => x"89",
          8208 => x"73",
          8209 => x"81",
          8210 => x"82",
          8211 => x"74",
          8212 => x"f2",
          8213 => x"8c",
          8214 => x"2e",
          8215 => x"8c",
          8216 => x"fe",
          8217 => x"8e",
          8218 => x"f4",
          8219 => x"3f",
          8220 => x"89",
          8221 => x"89",
          8222 => x"73",
          8223 => x"81",
          8224 => x"74",
          8225 => x"fe",
          8226 => x"80",
          8227 => x"dc",
          8228 => x"0d",
          8229 => x"0d",
          8230 => x"82",
          8231 => x"5f",
          8232 => x"7c",
          8233 => x"db",
          8234 => x"dc",
          8235 => x"06",
          8236 => x"2e",
          8237 => x"a2",
          8238 => x"a0",
          8239 => x"70",
          8240 => x"ee",
          8241 => x"53",
          8242 => x"8e",
          8243 => x"b5",
          8244 => x"8c",
          8245 => x"2e",
          8246 => x"84",
          8247 => x"bc",
          8248 => x"5f",
          8249 => x"dc",
          8250 => x"9e",
          8251 => x"70",
          8252 => x"f8",
          8253 => x"fe",
          8254 => x"3d",
          8255 => x"51",
          8256 => x"82",
          8257 => x"90",
          8258 => x"2c",
          8259 => x"80",
          8260 => x"b3",
          8261 => x"c2",
          8262 => x"78",
          8263 => x"d5",
          8264 => x"24",
          8265 => x"80",
          8266 => x"38",
          8267 => x"80",
          8268 => x"e9",
          8269 => x"c0",
          8270 => x"38",
          8271 => x"24",
          8272 => x"78",
          8273 => x"92",
          8274 => x"39",
          8275 => x"2e",
          8276 => x"78",
          8277 => x"92",
          8278 => x"c3",
          8279 => x"38",
          8280 => x"2e",
          8281 => x"8a",
          8282 => x"81",
          8283 => x"99",
          8284 => x"83",
          8285 => x"78",
          8286 => x"89",
          8287 => x"9d",
          8288 => x"85",
          8289 => x"38",
          8290 => x"b4",
          8291 => x"11",
          8292 => x"05",
          8293 => x"cb",
          8294 => x"dc",
          8295 => x"fe",
          8296 => x"3d",
          8297 => x"53",
          8298 => x"51",
          8299 => x"3f",
          8300 => x"08",
          8301 => x"ad",
          8302 => x"fe",
          8303 => x"ff",
          8304 => x"fe",
          8305 => x"82",
          8306 => x"86",
          8307 => x"dc",
          8308 => x"84",
          8309 => x"e6",
          8310 => x"63",
          8311 => x"7b",
          8312 => x"38",
          8313 => x"7a",
          8314 => x"5c",
          8315 => x"26",
          8316 => x"e1",
          8317 => x"ff",
          8318 => x"ff",
          8319 => x"fe",
          8320 => x"82",
          8321 => x"80",
          8322 => x"38",
          8323 => x"fc",
          8324 => x"84",
          8325 => x"ed",
          8326 => x"8c",
          8327 => x"2e",
          8328 => x"b4",
          8329 => x"11",
          8330 => x"05",
          8331 => x"b3",
          8332 => x"dc",
          8333 => x"fd",
          8334 => x"84",
          8335 => x"e5",
          8336 => x"5a",
          8337 => x"81",
          8338 => x"59",
          8339 => x"05",
          8340 => x"34",
          8341 => x"42",
          8342 => x"3d",
          8343 => x"53",
          8344 => x"51",
          8345 => x"3f",
          8346 => x"08",
          8347 => x"f5",
          8348 => x"fe",
          8349 => x"ff",
          8350 => x"fe",
          8351 => x"82",
          8352 => x"80",
          8353 => x"38",
          8354 => x"f8",
          8355 => x"84",
          8356 => x"ec",
          8357 => x"8c",
          8358 => x"2e",
          8359 => x"82",
          8360 => x"fe",
          8361 => x"63",
          8362 => x"27",
          8363 => x"70",
          8364 => x"5e",
          8365 => x"7c",
          8366 => x"78",
          8367 => x"79",
          8368 => x"52",
          8369 => x"51",
          8370 => x"3f",
          8371 => x"81",
          8372 => x"d5",
          8373 => x"a4",
          8374 => x"39",
          8375 => x"80",
          8376 => x"84",
          8377 => x"eb",
          8378 => x"8c",
          8379 => x"df",
          8380 => x"a0",
          8381 => x"80",
          8382 => x"82",
          8383 => x"44",
          8384 => x"82",
          8385 => x"59",
          8386 => x"88",
          8387 => x"e0",
          8388 => x"39",
          8389 => x"33",
          8390 => x"2e",
          8391 => x"87",
          8392 => x"ab",
          8393 => x"a3",
          8394 => x"80",
          8395 => x"82",
          8396 => x"44",
          8397 => x"88",
          8398 => x"78",
          8399 => x"38",
          8400 => x"08",
          8401 => x"82",
          8402 => x"fc",
          8403 => x"b4",
          8404 => x"11",
          8405 => x"05",
          8406 => x"87",
          8407 => x"dc",
          8408 => x"38",
          8409 => x"33",
          8410 => x"2e",
          8411 => x"87",
          8412 => x"80",
          8413 => x"88",
          8414 => x"78",
          8415 => x"38",
          8416 => x"08",
          8417 => x"82",
          8418 => x"59",
          8419 => x"88",
          8420 => x"ec",
          8421 => x"39",
          8422 => x"33",
          8423 => x"2e",
          8424 => x"87",
          8425 => x"99",
          8426 => x"9e",
          8427 => x"80",
          8428 => x"82",
          8429 => x"43",
          8430 => x"88",
          8431 => x"05",
          8432 => x"fe",
          8433 => x"ff",
          8434 => x"fe",
          8435 => x"82",
          8436 => x"80",
          8437 => x"80",
          8438 => x"7a",
          8439 => x"38",
          8440 => x"90",
          8441 => x"70",
          8442 => x"2a",
          8443 => x"51",
          8444 => x"78",
          8445 => x"38",
          8446 => x"83",
          8447 => x"82",
          8448 => x"fe",
          8449 => x"a0",
          8450 => x"61",
          8451 => x"63",
          8452 => x"3f",
          8453 => x"51",
          8454 => x"3f",
          8455 => x"b4",
          8456 => x"11",
          8457 => x"05",
          8458 => x"b7",
          8459 => x"dc",
          8460 => x"f9",
          8461 => x"3d",
          8462 => x"53",
          8463 => x"51",
          8464 => x"3f",
          8465 => x"08",
          8466 => x"38",
          8467 => x"80",
          8468 => x"79",
          8469 => x"05",
          8470 => x"fe",
          8471 => x"ff",
          8472 => x"fe",
          8473 => x"82",
          8474 => x"e0",
          8475 => x"39",
          8476 => x"54",
          8477 => x"c4",
          8478 => x"f2",
          8479 => x"52",
          8480 => x"e7",
          8481 => x"45",
          8482 => x"78",
          8483 => x"d5",
          8484 => x"27",
          8485 => x"3d",
          8486 => x"53",
          8487 => x"51",
          8488 => x"3f",
          8489 => x"08",
          8490 => x"38",
          8491 => x"80",
          8492 => x"79",
          8493 => x"05",
          8494 => x"39",
          8495 => x"51",
          8496 => x"3f",
          8497 => x"b4",
          8498 => x"11",
          8499 => x"05",
          8500 => x"81",
          8501 => x"dc",
          8502 => x"f8",
          8503 => x"3d",
          8504 => x"53",
          8505 => x"51",
          8506 => x"3f",
          8507 => x"08",
          8508 => x"38",
          8509 => x"be",
          8510 => x"70",
          8511 => x"23",
          8512 => x"3d",
          8513 => x"53",
          8514 => x"51",
          8515 => x"3f",
          8516 => x"08",
          8517 => x"cd",
          8518 => x"22",
          8519 => x"85",
          8520 => x"e5",
          8521 => x"f8",
          8522 => x"fe",
          8523 => x"79",
          8524 => x"59",
          8525 => x"f7",
          8526 => x"9f",
          8527 => x"60",
          8528 => x"d5",
          8529 => x"fe",
          8530 => x"ff",
          8531 => x"fe",
          8532 => x"82",
          8533 => x"80",
          8534 => x"60",
          8535 => x"05",
          8536 => x"82",
          8537 => x"78",
          8538 => x"39",
          8539 => x"51",
          8540 => x"3f",
          8541 => x"b4",
          8542 => x"11",
          8543 => x"05",
          8544 => x"d1",
          8545 => x"dc",
          8546 => x"f6",
          8547 => x"3d",
          8548 => x"53",
          8549 => x"51",
          8550 => x"3f",
          8551 => x"08",
          8552 => x"38",
          8553 => x"0c",
          8554 => x"05",
          8555 => x"fe",
          8556 => x"ff",
          8557 => x"fe",
          8558 => x"82",
          8559 => x"e4",
          8560 => x"39",
          8561 => x"54",
          8562 => x"e4",
          8563 => x"9e",
          8564 => x"52",
          8565 => x"e4",
          8566 => x"45",
          8567 => x"78",
          8568 => x"81",
          8569 => x"27",
          8570 => x"3d",
          8571 => x"53",
          8572 => x"51",
          8573 => x"3f",
          8574 => x"08",
          8575 => x"38",
          8576 => x"0c",
          8577 => x"05",
          8578 => x"39",
          8579 => x"51",
          8580 => x"3f",
          8581 => x"b4",
          8582 => x"11",
          8583 => x"05",
          8584 => x"bf",
          8585 => x"dc",
          8586 => x"f5",
          8587 => x"52",
          8588 => x"51",
          8589 => x"3f",
          8590 => x"04",
          8591 => x"80",
          8592 => x"84",
          8593 => x"e5",
          8594 => x"8c",
          8595 => x"2e",
          8596 => x"63",
          8597 => x"8c",
          8598 => x"92",
          8599 => x"78",
          8600 => x"dc",
          8601 => x"f4",
          8602 => x"8c",
          8603 => x"82",
          8604 => x"fe",
          8605 => x"f4",
          8606 => x"86",
          8607 => x"dd",
          8608 => x"bd",
          8609 => x"dd",
          8610 => x"e0",
          8611 => x"fa",
          8612 => x"ff",
          8613 => x"d3",
          8614 => x"c9",
          8615 => x"79",
          8616 => x"80",
          8617 => x"38",
          8618 => x"59",
          8619 => x"81",
          8620 => x"3d",
          8621 => x"51",
          8622 => x"3f",
          8623 => x"08",
          8624 => x"7a",
          8625 => x"38",
          8626 => x"89",
          8627 => x"2e",
          8628 => x"cd",
          8629 => x"2e",
          8630 => x"c5",
          8631 => x"f4",
          8632 => x"82",
          8633 => x"80",
          8634 => x"fc",
          8635 => x"ff",
          8636 => x"fe",
          8637 => x"bb",
          8638 => x"9c",
          8639 => x"ff",
          8640 => x"fe",
          8641 => x"ab",
          8642 => x"82",
          8643 => x"80",
          8644 => x"8c",
          8645 => x"ff",
          8646 => x"fe",
          8647 => x"93",
          8648 => x"80",
          8649 => x"98",
          8650 => x"ff",
          8651 => x"fe",
          8652 => x"82",
          8653 => x"82",
          8654 => x"80",
          8655 => x"80",
          8656 => x"80",
          8657 => x"80",
          8658 => x"ff",
          8659 => x"eb",
          8660 => x"8c",
          8661 => x"8c",
          8662 => x"70",
          8663 => x"07",
          8664 => x"5b",
          8665 => x"5a",
          8666 => x"83",
          8667 => x"78",
          8668 => x"78",
          8669 => x"38",
          8670 => x"81",
          8671 => x"59",
          8672 => x"38",
          8673 => x"7d",
          8674 => x"59",
          8675 => x"7e",
          8676 => x"81",
          8677 => x"38",
          8678 => x"51",
          8679 => x"3f",
          8680 => x"fc",
          8681 => x"0b",
          8682 => x"34",
          8683 => x"8c",
          8684 => x"55",
          8685 => x"52",
          8686 => x"bb",
          8687 => x"8c",
          8688 => x"2b",
          8689 => x"53",
          8690 => x"52",
          8691 => x"bb",
          8692 => x"82",
          8693 => x"07",
          8694 => x"c0",
          8695 => x"08",
          8696 => x"84",
          8697 => x"51",
          8698 => x"3f",
          8699 => x"08",
          8700 => x"08",
          8701 => x"84",
          8702 => x"51",
          8703 => x"3f",
          8704 => x"dc",
          8705 => x"0c",
          8706 => x"0b",
          8707 => x"84",
          8708 => x"83",
          8709 => x"94",
          8710 => x"ac",
          8711 => x"f0",
          8712 => x"0b",
          8713 => x"0c",
          8714 => x"3f",
          8715 => x"3f",
          8716 => x"51",
          8717 => x"3f",
          8718 => x"51",
          8719 => x"3f",
          8720 => x"51",
          8721 => x"3f",
          8722 => x"be",
          8723 => x"3f",
          8724 => x"00",
          8725 => x"00",
          8726 => x"00",
          8727 => x"00",
          8728 => x"00",
          8729 => x"00",
          8730 => x"00",
          8731 => x"00",
          8732 => x"00",
          8733 => x"00",
          8734 => x"00",
          8735 => x"00",
          8736 => x"00",
          8737 => x"00",
          8738 => x"00",
          8739 => x"00",
          8740 => x"00",
          8741 => x"00",
          8742 => x"00",
          8743 => x"00",
          8744 => x"00",
          8745 => x"00",
          8746 => x"00",
          8747 => x"00",
          8748 => x"00",
          8749 => x"00",
          8750 => x"00",
          8751 => x"00",
          8752 => x"00",
          8753 => x"00",
          8754 => x"00",
          8755 => x"00",
          8756 => x"00",
          8757 => x"00",
          8758 => x"00",
          8759 => x"00",
          8760 => x"00",
          8761 => x"25",
          8762 => x"64",
          8763 => x"20",
          8764 => x"25",
          8765 => x"64",
          8766 => x"25",
          8767 => x"53",
          8768 => x"43",
          8769 => x"69",
          8770 => x"61",
          8771 => x"6e",
          8772 => x"20",
          8773 => x"6f",
          8774 => x"6f",
          8775 => x"6f",
          8776 => x"67",
          8777 => x"3a",
          8778 => x"76",
          8779 => x"73",
          8780 => x"70",
          8781 => x"65",
          8782 => x"64",
          8783 => x"20",
          8784 => x"57",
          8785 => x"44",
          8786 => x"20",
          8787 => x"30",
          8788 => x"25",
          8789 => x"29",
          8790 => x"20",
          8791 => x"53",
          8792 => x"4d",
          8793 => x"20",
          8794 => x"30",
          8795 => x"25",
          8796 => x"29",
          8797 => x"20",
          8798 => x"49",
          8799 => x"20",
          8800 => x"4d",
          8801 => x"30",
          8802 => x"25",
          8803 => x"29",
          8804 => x"20",
          8805 => x"42",
          8806 => x"20",
          8807 => x"20",
          8808 => x"30",
          8809 => x"25",
          8810 => x"29",
          8811 => x"20",
          8812 => x"52",
          8813 => x"20",
          8814 => x"20",
          8815 => x"30",
          8816 => x"25",
          8817 => x"29",
          8818 => x"20",
          8819 => x"53",
          8820 => x"41",
          8821 => x"20",
          8822 => x"65",
          8823 => x"65",
          8824 => x"25",
          8825 => x"29",
          8826 => x"20",
          8827 => x"54",
          8828 => x"52",
          8829 => x"20",
          8830 => x"69",
          8831 => x"73",
          8832 => x"25",
          8833 => x"29",
          8834 => x"20",
          8835 => x"49",
          8836 => x"20",
          8837 => x"4c",
          8838 => x"68",
          8839 => x"65",
          8840 => x"25",
          8841 => x"29",
          8842 => x"20",
          8843 => x"57",
          8844 => x"42",
          8845 => x"20",
          8846 => x"0a",
          8847 => x"20",
          8848 => x"57",
          8849 => x"32",
          8850 => x"20",
          8851 => x"49",
          8852 => x"4c",
          8853 => x"20",
          8854 => x"50",
          8855 => x"00",
          8856 => x"20",
          8857 => x"53",
          8858 => x"00",
          8859 => x"41",
          8860 => x"65",
          8861 => x"73",
          8862 => x"20",
          8863 => x"43",
          8864 => x"52",
          8865 => x"74",
          8866 => x"63",
          8867 => x"20",
          8868 => x"72",
          8869 => x"20",
          8870 => x"30",
          8871 => x"00",
          8872 => x"20",
          8873 => x"43",
          8874 => x"4d",
          8875 => x"72",
          8876 => x"74",
          8877 => x"20",
          8878 => x"72",
          8879 => x"20",
          8880 => x"30",
          8881 => x"00",
          8882 => x"20",
          8883 => x"53",
          8884 => x"6b",
          8885 => x"61",
          8886 => x"41",
          8887 => x"65",
          8888 => x"20",
          8889 => x"20",
          8890 => x"30",
          8891 => x"00",
          8892 => x"4d",
          8893 => x"3a",
          8894 => x"20",
          8895 => x"5a",
          8896 => x"49",
          8897 => x"20",
          8898 => x"20",
          8899 => x"20",
          8900 => x"20",
          8901 => x"20",
          8902 => x"30",
          8903 => x"00",
          8904 => x"20",
          8905 => x"53",
          8906 => x"65",
          8907 => x"6c",
          8908 => x"20",
          8909 => x"71",
          8910 => x"20",
          8911 => x"20",
          8912 => x"64",
          8913 => x"34",
          8914 => x"7a",
          8915 => x"20",
          8916 => x"53",
          8917 => x"4d",
          8918 => x"6f",
          8919 => x"46",
          8920 => x"20",
          8921 => x"20",
          8922 => x"20",
          8923 => x"64",
          8924 => x"34",
          8925 => x"7a",
          8926 => x"20",
          8927 => x"57",
          8928 => x"62",
          8929 => x"20",
          8930 => x"41",
          8931 => x"6c",
          8932 => x"20",
          8933 => x"71",
          8934 => x"64",
          8935 => x"34",
          8936 => x"7a",
          8937 => x"53",
          8938 => x"6c",
          8939 => x"4d",
          8940 => x"75",
          8941 => x"46",
          8942 => x"00",
          8943 => x"45",
          8944 => x"45",
          8945 => x"69",
          8946 => x"55",
          8947 => x"6f",
          8948 => x"68",
          8949 => x"6f",
          8950 => x"74",
          8951 => x"68",
          8952 => x"6f",
          8953 => x"68",
          8954 => x"00",
          8955 => x"21",
          8956 => x"25",
          8957 => x"20",
          8958 => x"0a",
          8959 => x"46",
          8960 => x"65",
          8961 => x"6f",
          8962 => x"73",
          8963 => x"74",
          8964 => x"68",
          8965 => x"6f",
          8966 => x"66",
          8967 => x"20",
          8968 => x"45",
          8969 => x"0a",
          8970 => x"43",
          8971 => x"6f",
          8972 => x"70",
          8973 => x"63",
          8974 => x"74",
          8975 => x"69",
          8976 => x"72",
          8977 => x"69",
          8978 => x"20",
          8979 => x"61",
          8980 => x"6e",
          8981 => x"00",
          8982 => x"00",
          8983 => x"01",
          8984 => x"00",
          8985 => x"00",
          8986 => x"01",
          8987 => x"00",
          8988 => x"00",
          8989 => x"04",
          8990 => x"00",
          8991 => x"00",
          8992 => x"04",
          8993 => x"00",
          8994 => x"00",
          8995 => x"04",
          8996 => x"00",
          8997 => x"00",
          8998 => x"04",
          8999 => x"00",
          9000 => x"00",
          9001 => x"04",
          9002 => x"00",
          9003 => x"00",
          9004 => x"03",
          9005 => x"00",
          9006 => x"00",
          9007 => x"03",
          9008 => x"00",
          9009 => x"00",
          9010 => x"03",
          9011 => x"00",
          9012 => x"00",
          9013 => x"03",
          9014 => x"00",
          9015 => x"1b",
          9016 => x"1b",
          9017 => x"1b",
          9018 => x"1b",
          9019 => x"1b",
          9020 => x"1b",
          9021 => x"1b",
          9022 => x"1b",
          9023 => x"1b",
          9024 => x"0d",
          9025 => x"08",
          9026 => x"53",
          9027 => x"22",
          9028 => x"3a",
          9029 => x"3e",
          9030 => x"7c",
          9031 => x"46",
          9032 => x"46",
          9033 => x"32",
          9034 => x"eb",
          9035 => x"53",
          9036 => x"35",
          9037 => x"4e",
          9038 => x"41",
          9039 => x"20",
          9040 => x"41",
          9041 => x"20",
          9042 => x"4e",
          9043 => x"41",
          9044 => x"20",
          9045 => x"41",
          9046 => x"20",
          9047 => x"00",
          9048 => x"00",
          9049 => x"00",
          9050 => x"00",
          9051 => x"80",
          9052 => x"8e",
          9053 => x"45",
          9054 => x"49",
          9055 => x"90",
          9056 => x"99",
          9057 => x"59",
          9058 => x"9c",
          9059 => x"41",
          9060 => x"a5",
          9061 => x"a8",
          9062 => x"ac",
          9063 => x"b0",
          9064 => x"b4",
          9065 => x"b8",
          9066 => x"bc",
          9067 => x"c0",
          9068 => x"c4",
          9069 => x"c8",
          9070 => x"cc",
          9071 => x"d0",
          9072 => x"d4",
          9073 => x"d8",
          9074 => x"dc",
          9075 => x"e0",
          9076 => x"e4",
          9077 => x"e8",
          9078 => x"ec",
          9079 => x"f0",
          9080 => x"f4",
          9081 => x"f8",
          9082 => x"fc",
          9083 => x"2b",
          9084 => x"3d",
          9085 => x"5c",
          9086 => x"3c",
          9087 => x"7f",
          9088 => x"00",
          9089 => x"00",
          9090 => x"01",
          9091 => x"00",
          9092 => x"00",
          9093 => x"00",
          9094 => x"00",
          9095 => x"00",
          9096 => x"64",
          9097 => x"74",
          9098 => x"64",
          9099 => x"74",
          9100 => x"66",
          9101 => x"74",
          9102 => x"66",
          9103 => x"64",
          9104 => x"66",
          9105 => x"63",
          9106 => x"6d",
          9107 => x"61",
          9108 => x"6d",
          9109 => x"79",
          9110 => x"6d",
          9111 => x"66",
          9112 => x"6d",
          9113 => x"70",
          9114 => x"6d",
          9115 => x"6d",
          9116 => x"6d",
          9117 => x"68",
          9118 => x"68",
          9119 => x"68",
          9120 => x"68",
          9121 => x"63",
          9122 => x"00",
          9123 => x"6a",
          9124 => x"72",
          9125 => x"61",
          9126 => x"72",
          9127 => x"74",
          9128 => x"69",
          9129 => x"00",
          9130 => x"74",
          9131 => x"00",
          9132 => x"74",
          9133 => x"69",
          9134 => x"6d",
          9135 => x"69",
          9136 => x"6b",
          9137 => x"00",
          9138 => x"44",
          9139 => x"20",
          9140 => x"6f",
          9141 => x"49",
          9142 => x"72",
          9143 => x"20",
          9144 => x"6f",
          9145 => x"00",
          9146 => x"44",
          9147 => x"20",
          9148 => x"20",
          9149 => x"64",
          9150 => x"00",
          9151 => x"4e",
          9152 => x"69",
          9153 => x"66",
          9154 => x"64",
          9155 => x"4e",
          9156 => x"61",
          9157 => x"66",
          9158 => x"64",
          9159 => x"49",
          9160 => x"6c",
          9161 => x"66",
          9162 => x"6e",
          9163 => x"2e",
          9164 => x"41",
          9165 => x"73",
          9166 => x"65",
          9167 => x"64",
          9168 => x"46",
          9169 => x"20",
          9170 => x"65",
          9171 => x"20",
          9172 => x"73",
          9173 => x"0a",
          9174 => x"46",
          9175 => x"20",
          9176 => x"64",
          9177 => x"69",
          9178 => x"6c",
          9179 => x"0a",
          9180 => x"53",
          9181 => x"73",
          9182 => x"69",
          9183 => x"70",
          9184 => x"65",
          9185 => x"64",
          9186 => x"44",
          9187 => x"65",
          9188 => x"6d",
          9189 => x"20",
          9190 => x"69",
          9191 => x"6c",
          9192 => x"0a",
          9193 => x"44",
          9194 => x"20",
          9195 => x"20",
          9196 => x"62",
          9197 => x"2e",
          9198 => x"4e",
          9199 => x"6f",
          9200 => x"74",
          9201 => x"65",
          9202 => x"6c",
          9203 => x"73",
          9204 => x"20",
          9205 => x"6e",
          9206 => x"6e",
          9207 => x"73",
          9208 => x"00",
          9209 => x"46",
          9210 => x"61",
          9211 => x"62",
          9212 => x"65",
          9213 => x"00",
          9214 => x"54",
          9215 => x"6f",
          9216 => x"20",
          9217 => x"72",
          9218 => x"6f",
          9219 => x"61",
          9220 => x"6c",
          9221 => x"2e",
          9222 => x"46",
          9223 => x"20",
          9224 => x"6c",
          9225 => x"65",
          9226 => x"00",
          9227 => x"49",
          9228 => x"66",
          9229 => x"69",
          9230 => x"20",
          9231 => x"6f",
          9232 => x"0a",
          9233 => x"54",
          9234 => x"6d",
          9235 => x"20",
          9236 => x"6e",
          9237 => x"6c",
          9238 => x"0a",
          9239 => x"50",
          9240 => x"6d",
          9241 => x"72",
          9242 => x"6e",
          9243 => x"72",
          9244 => x"2e",
          9245 => x"53",
          9246 => x"65",
          9247 => x"0a",
          9248 => x"55",
          9249 => x"6f",
          9250 => x"65",
          9251 => x"72",
          9252 => x"0a",
          9253 => x"20",
          9254 => x"65",
          9255 => x"73",
          9256 => x"20",
          9257 => x"20",
          9258 => x"65",
          9259 => x"65",
          9260 => x"00",
          9261 => x"72",
          9262 => x"00",
          9263 => x"25",
          9264 => x"00",
          9265 => x"3a",
          9266 => x"25",
          9267 => x"00",
          9268 => x"20",
          9269 => x"20",
          9270 => x"00",
          9271 => x"25",
          9272 => x"00",
          9273 => x"20",
          9274 => x"20",
          9275 => x"7c",
          9276 => x"7a",
          9277 => x"0a",
          9278 => x"25",
          9279 => x"00",
          9280 => x"31",
          9281 => x"34",
          9282 => x"32",
          9283 => x"76",
          9284 => x"31",
          9285 => x"20",
          9286 => x"2c",
          9287 => x"76",
          9288 => x"32",
          9289 => x"25",
          9290 => x"73",
          9291 => x"0a",
          9292 => x"5a",
          9293 => x"49",
          9294 => x"72",
          9295 => x"74",
          9296 => x"6e",
          9297 => x"72",
          9298 => x"54",
          9299 => x"72",
          9300 => x"74",
          9301 => x"75",
          9302 => x"00",
          9303 => x"50",
          9304 => x"69",
          9305 => x"72",
          9306 => x"74",
          9307 => x"49",
          9308 => x"4c",
          9309 => x"20",
          9310 => x"65",
          9311 => x"70",
          9312 => x"49",
          9313 => x"4c",
          9314 => x"20",
          9315 => x"65",
          9316 => x"70",
          9317 => x"55",
          9318 => x"30",
          9319 => x"20",
          9320 => x"65",
          9321 => x"70",
          9322 => x"55",
          9323 => x"30",
          9324 => x"20",
          9325 => x"65",
          9326 => x"70",
          9327 => x"55",
          9328 => x"31",
          9329 => x"20",
          9330 => x"65",
          9331 => x"70",
          9332 => x"55",
          9333 => x"31",
          9334 => x"20",
          9335 => x"65",
          9336 => x"70",
          9337 => x"53",
          9338 => x"69",
          9339 => x"75",
          9340 => x"69",
          9341 => x"2e",
          9342 => x"00",
          9343 => x"45",
          9344 => x"6c",
          9345 => x"20",
          9346 => x"65",
          9347 => x"2e",
          9348 => x"61",
          9349 => x"65",
          9350 => x"2e",
          9351 => x"00",
          9352 => x"30",
          9353 => x"46",
          9354 => x"65",
          9355 => x"6f",
          9356 => x"69",
          9357 => x"6c",
          9358 => x"20",
          9359 => x"63",
          9360 => x"20",
          9361 => x"70",
          9362 => x"73",
          9363 => x"6e",
          9364 => x"6d",
          9365 => x"61",
          9366 => x"2e",
          9367 => x"2a",
          9368 => x"43",
          9369 => x"72",
          9370 => x"2e",
          9371 => x"00",
          9372 => x"43",
          9373 => x"69",
          9374 => x"2e",
          9375 => x"43",
          9376 => x"61",
          9377 => x"67",
          9378 => x"00",
          9379 => x"25",
          9380 => x"78",
          9381 => x"38",
          9382 => x"3e",
          9383 => x"6c",
          9384 => x"30",
          9385 => x"0a",
          9386 => x"44",
          9387 => x"20",
          9388 => x"6f",
          9389 => x"00",
          9390 => x"0a",
          9391 => x"70",
          9392 => x"65",
          9393 => x"25",
          9394 => x"20",
          9395 => x"58",
          9396 => x"3f",
          9397 => x"00",
          9398 => x"25",
          9399 => x"20",
          9400 => x"58",
          9401 => x"25",
          9402 => x"20",
          9403 => x"58",
          9404 => x"45",
          9405 => x"75",
          9406 => x"67",
          9407 => x"64",
          9408 => x"20",
          9409 => x"78",
          9410 => x"2e",
          9411 => x"43",
          9412 => x"69",
          9413 => x"63",
          9414 => x"20",
          9415 => x"30",
          9416 => x"2e",
          9417 => x"00",
          9418 => x"43",
          9419 => x"20",
          9420 => x"75",
          9421 => x"64",
          9422 => x"64",
          9423 => x"25",
          9424 => x"0a",
          9425 => x"52",
          9426 => x"61",
          9427 => x"6e",
          9428 => x"70",
          9429 => x"63",
          9430 => x"6f",
          9431 => x"2e",
          9432 => x"43",
          9433 => x"20",
          9434 => x"6f",
          9435 => x"6e",
          9436 => x"2e",
          9437 => x"5a",
          9438 => x"62",
          9439 => x"25",
          9440 => x"25",
          9441 => x"73",
          9442 => x"00",
          9443 => x"25",
          9444 => x"25",
          9445 => x"73",
          9446 => x"25",
          9447 => x"25",
          9448 => x"42",
          9449 => x"63",
          9450 => x"61",
          9451 => x"0a",
          9452 => x"52",
          9453 => x"69",
          9454 => x"2e",
          9455 => x"45",
          9456 => x"6c",
          9457 => x"20",
          9458 => x"65",
          9459 => x"70",
          9460 => x"2e",
          9461 => x"00",
          9462 => x"00",
          9463 => x"00",
          9464 => x"00",
          9465 => x"00",
          9466 => x"00",
          9467 => x"00",
          9468 => x"00",
          9469 => x"00",
          9470 => x"01",
          9471 => x"01",
          9472 => x"00",
          9473 => x"00",
          9474 => x"00",
          9475 => x"00",
          9476 => x"05",
          9477 => x"05",
          9478 => x"05",
          9479 => x"00",
          9480 => x"01",
          9481 => x"01",
          9482 => x"01",
          9483 => x"01",
          9484 => x"00",
          9485 => x"00",
          9486 => x"00",
          9487 => x"00",
          9488 => x"00",
          9489 => x"00",
          9490 => x"00",
          9491 => x"00",
          9492 => x"00",
          9493 => x"00",
          9494 => x"00",
          9495 => x"00",
          9496 => x"00",
          9497 => x"00",
          9498 => x"00",
          9499 => x"00",
          9500 => x"00",
          9501 => x"00",
          9502 => x"00",
          9503 => x"00",
          9504 => x"00",
          9505 => x"00",
          9506 => x"00",
          9507 => x"00",
          9508 => x"00",
          9509 => x"00",
          9510 => x"00",
          9511 => x"00",
          9512 => x"00",
          9513 => x"00",
          9514 => x"00",
          9515 => x"00",
          9516 => x"01",
          9517 => x"00",
          9518 => x"01",
          9519 => x"00",
          9520 => x"02",
          9521 => x"01",
          9522 => x"00",
          9523 => x"00",
          9524 => x"01",
          9525 => x"00",
          9526 => x"00",
          9527 => x"00",
          9528 => x"01",
          9529 => x"00",
          9530 => x"00",
          9531 => x"00",
          9532 => x"01",
          9533 => x"00",
          9534 => x"00",
          9535 => x"00",
          9536 => x"01",
          9537 => x"00",
          9538 => x"00",
          9539 => x"00",
          9540 => x"01",
          9541 => x"00",
          9542 => x"00",
          9543 => x"00",
          9544 => x"01",
          9545 => x"00",
          9546 => x"00",
          9547 => x"00",
          9548 => x"01",
          9549 => x"00",
          9550 => x"00",
          9551 => x"00",
          9552 => x"01",
          9553 => x"00",
          9554 => x"00",
          9555 => x"00",
          9556 => x"01",
          9557 => x"00",
          9558 => x"00",
          9559 => x"00",
          9560 => x"01",
          9561 => x"00",
          9562 => x"00",
          9563 => x"00",
          9564 => x"01",
          9565 => x"00",
          9566 => x"00",
          9567 => x"00",
          9568 => x"01",
          9569 => x"00",
          9570 => x"00",
          9571 => x"00",
          9572 => x"01",
          9573 => x"00",
          9574 => x"00",
          9575 => x"00",
          9576 => x"01",
          9577 => x"00",
          9578 => x"00",
          9579 => x"00",
          9580 => x"01",
          9581 => x"00",
          9582 => x"00",
          9583 => x"00",
          9584 => x"01",
          9585 => x"00",
          9586 => x"00",
          9587 => x"00",
          9588 => x"01",
          9589 => x"00",
          9590 => x"00",
          9591 => x"00",
          9592 => x"01",
          9593 => x"00",
          9594 => x"00",
          9595 => x"00",
          9596 => x"01",
          9597 => x"00",
          9598 => x"00",
          9599 => x"00",
          9600 => x"01",
          9601 => x"00",
          9602 => x"00",
          9603 => x"00",
          9604 => x"01",
          9605 => x"00",
          9606 => x"00",
          9607 => x"00",
          9608 => x"01",
          9609 => x"00",
          9610 => x"00",
          9611 => x"00",
          9612 => x"01",
          9613 => x"00",
          9614 => x"00",
          9615 => x"00",
          9616 => x"01",
          9617 => x"00",
          9618 => x"00",
          9619 => x"00",
          9620 => x"01",
          9621 => x"00",
          9622 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
