-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use pkgs.config_pkg.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_BIT_BRAM_32BIT_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e9040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"88738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cb2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8a",
           179 => x"fd2d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"80040088",
           281 => x"e2040000",
           282 => x"009fac70",
           283 => x"9fdc278b",
           284 => x"38807170",
           285 => x"8405530c",
           286 => x"88eb0488",
           287 => x"e2519e99",
           288 => x"04940802",
           289 => x"940cfd3d",
           290 => x"0d805394",
           291 => x"088c0508",
           292 => x"52940888",
           293 => x"05085182",
           294 => x"de3f8808",
           295 => x"70880c54",
           296 => x"853d0d94",
           297 => x"0c049408",
           298 => x"02940cfd",
           299 => x"3d0d8153",
           300 => x"94088c05",
           301 => x"08529408",
           302 => x"88050851",
           303 => x"82b93f88",
           304 => x"0870880c",
           305 => x"54853d0d",
           306 => x"940c0494",
           307 => x"0802940c",
           308 => x"f93d0d80",
           309 => x"0b9408fc",
           310 => x"050c9408",
           311 => x"88050880",
           312 => x"25ab3894",
           313 => x"08880508",
           314 => x"30940888",
           315 => x"050c800b",
           316 => x"9408f405",
           317 => x"0c9408fc",
           318 => x"05088838",
           319 => x"810b9408",
           320 => x"f4050c94",
           321 => x"08f40508",
           322 => x"9408fc05",
           323 => x"0c94088c",
           324 => x"05088025",
           325 => x"ab389408",
           326 => x"8c050830",
           327 => x"94088c05",
           328 => x"0c800b94",
           329 => x"08f0050c",
           330 => x"9408fc05",
           331 => x"08883881",
           332 => x"0b9408f0",
           333 => x"050c9408",
           334 => x"f0050894",
           335 => x"08fc050c",
           336 => x"80539408",
           337 => x"8c050852",
           338 => x"94088805",
           339 => x"085181a7",
           340 => x"3f880870",
           341 => x"9408f805",
           342 => x"0c549408",
           343 => x"fc050880",
           344 => x"2e8c3894",
           345 => x"08f80508",
           346 => x"309408f8",
           347 => x"050c9408",
           348 => x"f8050870",
           349 => x"880c5489",
           350 => x"3d0d940c",
           351 => x"04940802",
           352 => x"940cfb3d",
           353 => x"0d800b94",
           354 => x"08fc050c",
           355 => x"94088805",
           356 => x"08802593",
           357 => x"38940888",
           358 => x"05083094",
           359 => x"0888050c",
           360 => x"810b9408",
           361 => x"fc050c94",
           362 => x"088c0508",
           363 => x"80258c38",
           364 => x"94088c05",
           365 => x"08309408",
           366 => x"8c050c81",
           367 => x"5394088c",
           368 => x"05085294",
           369 => x"08880508",
           370 => x"51ad3f88",
           371 => x"08709408",
           372 => x"f8050c54",
           373 => x"9408fc05",
           374 => x"08802e8c",
           375 => x"389408f8",
           376 => x"05083094",
           377 => x"08f8050c",
           378 => x"9408f805",
           379 => x"0870880c",
           380 => x"54873d0d",
           381 => x"940c0494",
           382 => x"0802940c",
           383 => x"fd3d0d81",
           384 => x"0b9408fc",
           385 => x"050c800b",
           386 => x"9408f805",
           387 => x"0c94088c",
           388 => x"05089408",
           389 => x"88050827",
           390 => x"ac389408",
           391 => x"fc050880",
           392 => x"2ea33880",
           393 => x"0b94088c",
           394 => x"05082499",
           395 => x"3894088c",
           396 => x"05081094",
           397 => x"088c050c",
           398 => x"9408fc05",
           399 => x"08109408",
           400 => x"fc050cc9",
           401 => x"399408fc",
           402 => x"0508802e",
           403 => x"80c93894",
           404 => x"088c0508",
           405 => x"94088805",
           406 => x"0826a138",
           407 => x"94088805",
           408 => x"0894088c",
           409 => x"05083194",
           410 => x"0888050c",
           411 => x"9408f805",
           412 => x"089408fc",
           413 => x"05080794",
           414 => x"08f8050c",
           415 => x"9408fc05",
           416 => x"08812a94",
           417 => x"08fc050c",
           418 => x"94088c05",
           419 => x"08812a94",
           420 => x"088c050c",
           421 => x"ffaf3994",
           422 => x"08900508",
           423 => x"802e8f38",
           424 => x"94088805",
           425 => x"08709408",
           426 => x"f4050c51",
           427 => x"8d399408",
           428 => x"f8050870",
           429 => x"9408f405",
           430 => x"0c519408",
           431 => x"f4050888",
           432 => x"0c853d0d",
           433 => x"940c04ff",
           434 => x"3d0d8188",
           435 => x"0b87c092",
           436 => x"8c0c810b",
           437 => x"87c0928c",
           438 => x"0c850b87",
           439 => x"c0988c0c",
           440 => x"87c0928c",
           441 => x"08708206",
           442 => x"51517080",
           443 => x"2e8a3887",
           444 => x"c0988c08",
           445 => x"5170e938",
           446 => x"87c0928c",
           447 => x"08fc8080",
           448 => x"06527193",
           449 => x"3887c098",
           450 => x"8c085170",
           451 => x"802e8838",
           452 => x"710b0b0b",
           453 => x"9fa8340b",
           454 => x"0b0b9fa8",
           455 => x"33880c83",
           456 => x"3d0d04fa",
           457 => x"3d0d787b",
           458 => x"7d565856",
           459 => x"800b0b0b",
           460 => x"0b9fa833",
           461 => x"81065255",
           462 => x"82527075",
           463 => x"2e098106",
           464 => x"819e3885",
           465 => x"0b87c098",
           466 => x"8c0c7987",
           467 => x"c092800c",
           468 => x"840b87c0",
           469 => x"928c0c87",
           470 => x"c0928c08",
           471 => x"70852a70",
           472 => x"81065152",
           473 => x"5370802e",
           474 => x"a73887c0",
           475 => x"92840870",
           476 => x"81ff0676",
           477 => x"79275253",
           478 => x"5173802e",
           479 => x"90387080",
           480 => x"2e8b3871",
           481 => x"76708105",
           482 => x"5834ff14",
           483 => x"54811555",
           484 => x"72a20651",
           485 => x"70802e8b",
           486 => x"3887c098",
           487 => x"8c085170",
           488 => x"ffb53887",
           489 => x"c0988c08",
           490 => x"51709538",
           491 => x"810b87c0",
           492 => x"928c0c87",
           493 => x"c0928c08",
           494 => x"70820651",
           495 => x"5170f438",
           496 => x"8073fc80",
           497 => x"80065252",
           498 => x"70722e09",
           499 => x"81068f38",
           500 => x"87c0988c",
           501 => x"08517072",
           502 => x"2e098106",
           503 => x"83388152",
           504 => x"71880c88",
           505 => x"3d0d04fe",
           506 => x"3d0d7481",
           507 => x"11337133",
           508 => x"71882b07",
           509 => x"880c5351",
           510 => x"843d0d04",
           511 => x"fd3d0d75",
           512 => x"83113382",
           513 => x"12337190",
           514 => x"2b71882b",
           515 => x"07811433",
           516 => x"70720788",
           517 => x"2b753371",
           518 => x"07880c52",
           519 => x"53545654",
           520 => x"52853d0d",
           521 => x"04f93d0d",
           522 => x"790b0b0b",
           523 => x"9fac0857",
           524 => x"57817727",
           525 => x"80ed3876",
           526 => x"88170827",
           527 => x"80e53875",
           528 => x"33557482",
           529 => x"2e893874",
           530 => x"832eae38",
           531 => x"80d53974",
           532 => x"54761083",
           533 => x"fe065376",
           534 => x"882a8c17",
           535 => x"08055288",
           536 => x"3d705255",
           537 => x"fdbd3f88",
           538 => x"08b93874",
           539 => x"51fef83f",
           540 => x"880883ff",
           541 => x"ff0655ad",
           542 => x"39845476",
           543 => x"822b83fc",
           544 => x"06537687",
           545 => x"2a8c1708",
           546 => x"0552883d",
           547 => x"705255fd",
           548 => x"923f8808",
           549 => x"8e387451",
           550 => x"fee23f88",
           551 => x"08f00a06",
           552 => x"55833981",
           553 => x"5574880c",
           554 => x"893d0d04",
           555 => x"fb3d0d0b",
           556 => x"0b0b9fac",
           557 => x"08fe1988",
           558 => x"1208fe05",
           559 => x"55565480",
           560 => x"56747327",
           561 => x"8d388214",
           562 => x"33757129",
           563 => x"94160805",
           564 => x"57537588",
           565 => x"0c873d0d",
           566 => x"04fd3d0d",
           567 => x"7554800b",
           568 => x"0b0b0b9f",
           569 => x"ac087033",
           570 => x"51535371",
           571 => x"832e0981",
           572 => x"068c3894",
           573 => x"1451fdef",
           574 => x"3f880890",
           575 => x"2b539a14",
           576 => x"51fde43f",
           577 => x"880883ff",
           578 => x"ff067307",
           579 => x"880c853d",
           580 => x"0d04fc3d",
           581 => x"0d760b0b",
           582 => x"0b9fac08",
           583 => x"55558075",
           584 => x"23881508",
           585 => x"5372812e",
           586 => x"88388814",
           587 => x"08732685",
           588 => x"388152b0",
           589 => x"39729038",
           590 => x"73335271",
           591 => x"832e0981",
           592 => x"06853890",
           593 => x"14085372",
           594 => x"8c160c72",
           595 => x"802e8b38",
           596 => x"7251fed8",
           597 => x"3f880852",
           598 => x"85399014",
           599 => x"08527190",
           600 => x"160c8052",
           601 => x"71880c86",
           602 => x"3d0d04fa",
           603 => x"3d0d780b",
           604 => x"0b0b9fac",
           605 => x"08712281",
           606 => x"057083ff",
           607 => x"ff065754",
           608 => x"57557380",
           609 => x"2e883890",
           610 => x"15085372",
           611 => x"86388352",
           612 => x"80dc3973",
           613 => x"8f065271",
           614 => x"80cf3881",
           615 => x"1390160c",
           616 => x"8c150853",
           617 => x"728f3883",
           618 => x"0b841722",
           619 => x"57527376",
           620 => x"27bc38b5",
           621 => x"39821633",
           622 => x"ff057484",
           623 => x"2a065271",
           624 => x"a8387251",
           625 => x"fcdf3f81",
           626 => x"52718808",
           627 => x"27a03883",
           628 => x"52880888",
           629 => x"17082796",
           630 => x"3888088c",
           631 => x"160c8808",
           632 => x"51fdc93f",
           633 => x"88089016",
           634 => x"0c737523",
           635 => x"80527188",
           636 => x"0c883d0d",
           637 => x"04f23d0d",
           638 => x"60626458",
           639 => x"5e5c7533",
           640 => x"5574a02e",
           641 => x"09810688",
           642 => x"38811670",
           643 => x"4456ef39",
           644 => x"62703356",
           645 => x"5674af2e",
           646 => x"09810684",
           647 => x"38811643",
           648 => x"800b881d",
           649 => x"0c627033",
           650 => x"5155749f",
           651 => x"268f387b",
           652 => x"51fddf3f",
           653 => x"88085680",
           654 => x"7d3482d3",
           655 => x"39933d84",
           656 => x"1d087058",
           657 => x"5a5f8a55",
           658 => x"a0767081",
           659 => x"055834ff",
           660 => x"155574ff",
           661 => x"2e098106",
           662 => x"ef388070",
           663 => x"595b887f",
           664 => x"085f5a7a",
           665 => x"811c7081",
           666 => x"ff066013",
           667 => x"703370af",
           668 => x"327030a0",
           669 => x"73277180",
           670 => x"25075151",
           671 => x"525b535d",
           672 => x"57557480",
           673 => x"c73876ae",
           674 => x"2e098106",
           675 => x"83388155",
           676 => x"777a2775",
           677 => x"07557480",
           678 => x"2e9f3879",
           679 => x"88327030",
           680 => x"78ae3270",
           681 => x"30707307",
           682 => x"9f2a5351",
           683 => x"57515675",
           684 => x"9b388858",
           685 => x"8b5affab",
           686 => x"39778119",
           687 => x"7081ff06",
           688 => x"721c535a",
           689 => x"57557675",
           690 => x"34ff9839",
           691 => x"7a1e7f0c",
           692 => x"805576a0",
           693 => x"26833881",
           694 => x"55748b1a",
           695 => x"347b51fc",
           696 => x"b13f8808",
           697 => x"80ef38a0",
           698 => x"547b2270",
           699 => x"852b83e0",
           700 => x"06545590",
           701 => x"1c08527c",
           702 => x"51f8a83f",
           703 => x"88085788",
           704 => x"0880fb38",
           705 => x"7c335574",
           706 => x"802e80ee",
           707 => x"388b1d33",
           708 => x"70832a70",
           709 => x"81065156",
           710 => x"5674b238",
           711 => x"8b7d841e",
           712 => x"08880859",
           713 => x"5b5b58ff",
           714 => x"185877ff",
           715 => x"2e9a3879",
           716 => x"7081055b",
           717 => x"33797081",
           718 => x"055b3371",
           719 => x"71315256",
           720 => x"5675802e",
           721 => x"e2388639",
           722 => x"75802e92",
           723 => x"387b51fc",
           724 => x"9a3fff8e",
           725 => x"39880856",
           726 => x"8808b438",
           727 => x"83397656",
           728 => x"841c088b",
           729 => x"11335155",
           730 => x"74a5388b",
           731 => x"1d337084",
           732 => x"2a708106",
           733 => x"51565674",
           734 => x"89388356",
           735 => x"92398156",
           736 => x"8e397c51",
           737 => x"fad33f88",
           738 => x"08881d0c",
           739 => x"fdaf3975",
           740 => x"880c903d",
           741 => x"0d04f93d",
           742 => x"0d797b59",
           743 => x"57825483",
           744 => x"fe537752",
           745 => x"7651f6fb",
           746 => x"3f835688",
           747 => x"0880e738",
           748 => x"7651f8b3",
           749 => x"3f880883",
           750 => x"ffff0655",
           751 => x"82567482",
           752 => x"d4d52e09",
           753 => x"810680ce",
           754 => x"387554b6",
           755 => x"53775276",
           756 => x"51f6d03f",
           757 => x"88085688",
           758 => x"08943876",
           759 => x"51f8883f",
           760 => x"880883ff",
           761 => x"ff065574",
           762 => x"8182c62e",
           763 => x"a9388254",
           764 => x"80d25377",
           765 => x"527651f6",
           766 => x"aa3f8808",
           767 => x"56880894",
           768 => x"387651f7",
           769 => x"e23f8808",
           770 => x"83ffff06",
           771 => x"55748182",
           772 => x"c62e8338",
           773 => x"81567588",
           774 => x"0c893d0d",
           775 => x"04ed3d0d",
           776 => x"6559800b",
           777 => x"0b0b0b9f",
           778 => x"ac0cf59b",
           779 => x"3f880881",
           780 => x"06558256",
           781 => x"7482f238",
           782 => x"7475538d",
           783 => x"3d705357",
           784 => x"5afed33f",
           785 => x"880881ff",
           786 => x"06577681",
           787 => x"2e098106",
           788 => x"b3389054",
           789 => x"83be5374",
           790 => x"527551f5",
           791 => x"c63f8808",
           792 => x"ab388d3d",
           793 => x"33557480",
           794 => x"2eac3895",
           795 => x"3de40551",
           796 => x"f78a3f88",
           797 => x"08880853",
           798 => x"76525afe",
           799 => x"993f8808",
           800 => x"81ff0657",
           801 => x"76832e09",
           802 => x"81068638",
           803 => x"81568299",
           804 => x"3976802e",
           805 => x"86388656",
           806 => x"828f39a4",
           807 => x"548d5379",
           808 => x"527551f4",
           809 => x"fe3f8156",
           810 => x"880881fd",
           811 => x"38953de5",
           812 => x"0551f6b3",
           813 => x"3f880883",
           814 => x"ffff0658",
           815 => x"778c3895",
           816 => x"3df30551",
           817 => x"f6b63f88",
           818 => x"085802af",
           819 => x"05337871",
           820 => x"29028805",
           821 => x"ad057054",
           822 => x"52595bf6",
           823 => x"8a3f8808",
           824 => x"83ffff06",
           825 => x"7a058c1a",
           826 => x"0c8c3d33",
           827 => x"821a3495",
           828 => x"3de00551",
           829 => x"f5f13f88",
           830 => x"08841a23",
           831 => x"953de205",
           832 => x"51f5e43f",
           833 => x"880883ff",
           834 => x"ff065675",
           835 => x"8c38953d",
           836 => x"ef0551f5",
           837 => x"e73f8808",
           838 => x"567a51f5",
           839 => x"ca3f8808",
           840 => x"83ffff06",
           841 => x"76713179",
           842 => x"31841b22",
           843 => x"70842a82",
           844 => x"1d335672",
           845 => x"71315559",
           846 => x"5c5155ee",
           847 => x"c43f8808",
           848 => x"82057088",
           849 => x"1b0c8808",
           850 => x"e08a0556",
           851 => x"567483df",
           852 => x"fe268338",
           853 => x"825783ff",
           854 => x"f6762785",
           855 => x"38835789",
           856 => x"39865676",
           857 => x"802e80c1",
           858 => x"38767934",
           859 => x"76832e09",
           860 => x"81069038",
           861 => x"953dfb05",
           862 => x"51f5813f",
           863 => x"8808901a",
           864 => x"0c88398c",
           865 => x"19081890",
           866 => x"1a0c7983",
           867 => x"ffff068c",
           868 => x"1a081971",
           869 => x"842a0594",
           870 => x"1b0c5580",
           871 => x"0b811a34",
           872 => x"780b0b0b",
           873 => x"9fac0c80",
           874 => x"5675880c",
           875 => x"953d0d04",
           876 => x"ea3d0d0b",
           877 => x"0b0b9fac",
           878 => x"08558554",
           879 => x"74802e80",
           880 => x"df38800b",
           881 => x"81163498",
           882 => x"3de01145",
           883 => x"6954893d",
           884 => x"705457ec",
           885 => x"0551f89d",
           886 => x"3f880854",
           887 => x"880880c0",
           888 => x"38883d33",
           889 => x"5473802e",
           890 => x"933802a7",
           891 => x"05337084",
           892 => x"2a708106",
           893 => x"51555773",
           894 => x"802e8538",
           895 => x"8354a139",
           896 => x"7551f5d5",
           897 => x"3f8808a0",
           898 => x"160c983d",
           899 => x"dc0551f3",
           900 => x"eb3f8808",
           901 => x"9c160c73",
           902 => x"98160c81",
           903 => x"0b811634",
           904 => x"73880c98",
           905 => x"3d0d04f6",
           906 => x"3d0d7d7f",
           907 => x"7e0b0b0b",
           908 => x"9fac0859",
           909 => x"5b5c5880",
           910 => x"7b0c8557",
           911 => x"75802e81",
           912 => x"d1388116",
           913 => x"33810655",
           914 => x"84577480",
           915 => x"2e81c338",
           916 => x"91397481",
           917 => x"17348639",
           918 => x"800b8117",
           919 => x"34815781",
           920 => x"b1399c16",
           921 => x"08981708",
           922 => x"31557478",
           923 => x"27833874",
           924 => x"5877802e",
           925 => x"819a3898",
           926 => x"16087083",
           927 => x"ff065657",
           928 => x"7480c738",
           929 => x"821633ff",
           930 => x"0577892a",
           931 => x"067081ff",
           932 => x"065b5579",
           933 => x"9e387687",
           934 => x"38a01608",
           935 => x"558b39a4",
           936 => x"160851f3",
           937 => x"803f8808",
           938 => x"55817527",
           939 => x"ffaa3874",
           940 => x"a4170ca4",
           941 => x"160851f3",
           942 => x"f33f8808",
           943 => x"55880880",
           944 => x"2eff8f38",
           945 => x"88081aa8",
           946 => x"170c9816",
           947 => x"0883ff06",
           948 => x"84807131",
           949 => x"51557775",
           950 => x"27833877",
           951 => x"55745498",
           952 => x"160883ff",
           953 => x"0653a816",
           954 => x"08527851",
           955 => x"f0b53f88",
           956 => x"08fee538",
           957 => x"98160815",
           958 => x"98170c77",
           959 => x"75317b08",
           960 => x"167c0c58",
           961 => x"78802efe",
           962 => x"e8387419",
           963 => x"59fee239",
           964 => x"80577688",
           965 => x"0c8c3d0d",
           966 => x"04fb3d0d",
           967 => x"9b9086e4",
           968 => x"0b87c094",
           969 => x"8c0c9b90",
           970 => x"86e40b87",
           971 => x"c0949c0c",
           972 => x"8c80830b",
           973 => x"87c09484",
           974 => x"0c8c8083",
           975 => x"0b87c094",
           976 => x"940c9fb0",
           977 => x"51f9d63f",
           978 => x"8808b838",
           979 => x"9f9851fc",
           980 => x"df3f8808",
           981 => x"ae38a080",
           982 => x"0b880887",
           983 => x"c098880c",
           984 => x"55873dfc",
           985 => x"05538480",
           986 => x"527451fd",
           987 => x"ba3f8808",
           988 => x"8d387554",
           989 => x"73802e86",
           990 => x"38731555",
           991 => x"e439a080",
           992 => x"54730480",
           993 => x"54fb3900",
           994 => x"00ffffff",
           995 => x"ff00ffff",
           996 => x"ffff00ff",
           997 => x"ffffff00",
           998 => x"424f4f54",
           999 => x"54494e59",
          1000 => x"2e524f4d",
          1001 => x"00000000",
          1002 => x"01000000",
          2048 => x"0b0b0b84",
          2049 => x"800b0b0b",
          2050 => x"0b89fd04",
          2051 => x"ffffffff",
          2052 => x"ffffffff",
          2053 => x"ffffffff",
          2054 => x"ffffffff",
          2055 => x"ffffffff",
          2056 => x"0b0b0b84",
          2057 => x"80040b0b",
          2058 => x"0b848404",
          2059 => x"0b0b0b84",
          2060 => x"93040b0b",
          2061 => x"0b84a204",
          2062 => x"0b0b0b84",
          2063 => x"b1040b0b",
          2064 => x"0b84c004",
          2065 => x"0b0b0b84",
          2066 => x"cf040b0b",
          2067 => x"0b84de04",
          2068 => x"0b0b0b84",
          2069 => x"ed040b0b",
          2070 => x"0b84fc04",
          2071 => x"0b0b0b85",
          2072 => x"8b040b0b",
          2073 => x"0b859a04",
          2074 => x"0b0b0b85",
          2075 => x"a9040b0b",
          2076 => x"0b85b804",
          2077 => x"0b0b0b85",
          2078 => x"c7040b0b",
          2079 => x"0b85d604",
          2080 => x"0b0b0b85",
          2081 => x"e5040b0b",
          2082 => x"0b85f404",
          2083 => x"0b0b0b86",
          2084 => x"83040b0b",
          2085 => x"0b869304",
          2086 => x"0b0b0b86",
          2087 => x"a3040b0b",
          2088 => x"0b86b304",
          2089 => x"0b0b0b86",
          2090 => x"c3040b0b",
          2091 => x"0b86d304",
          2092 => x"0b0b0b86",
          2093 => x"e3040b0b",
          2094 => x"0b86f304",
          2095 => x"0b0b0b87",
          2096 => x"83040b0b",
          2097 => x"0b879304",
          2098 => x"0b0b0b87",
          2099 => x"a3040b0b",
          2100 => x"0b87b304",
          2101 => x"0b0b0b87",
          2102 => x"c3040b0b",
          2103 => x"0b87d304",
          2104 => x"0b0b0b87",
          2105 => x"e3040b0b",
          2106 => x"0b87f304",
          2107 => x"0b0b0b88",
          2108 => x"83040b0b",
          2109 => x"0b889304",
          2110 => x"0b0b0b88",
          2111 => x"a3040b0b",
          2112 => x"0b88b304",
          2113 => x"0b0b0b88",
          2114 => x"c3040b0b",
          2115 => x"0b88d304",
          2116 => x"0b0b0b88",
          2117 => x"e3040b0b",
          2118 => x"0b88f304",
          2119 => x"0b0b0b89",
          2120 => x"83040b0b",
          2121 => x"0b899304",
          2122 => x"0b0b0b89",
          2123 => x"a2040b0b",
          2124 => x"0b89b104",
          2125 => x"0b0b0b89",
          2126 => x"c0040b0b",
          2127 => x"0b89cf04",
          2128 => x"0b0b0b89",
          2129 => x"de040b0b",
          2130 => x"0b89ed04",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"00000000",
          2137 => x"00000000",
          2138 => x"00000000",
          2139 => x"00000000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"00000000",
          2145 => x"00000000",
          2146 => x"00000000",
          2147 => x"00000000",
          2148 => x"00000000",
          2149 => x"00000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"00000000",
          2153 => x"00000000",
          2154 => x"00000000",
          2155 => x"00000000",
          2156 => x"00000000",
          2157 => x"00000000",
          2158 => x"00000000",
          2159 => x"00000000",
          2160 => x"00000000",
          2161 => x"00000000",
          2162 => x"00000000",
          2163 => x"00000000",
          2164 => x"00000000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"00000000",
          2169 => x"00000000",
          2170 => x"00000000",
          2171 => x"00000000",
          2172 => x"00000000",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"00848004",
          2177 => x"81d3b80c",
          2178 => x"94e72d81",
          2179 => x"d3b80883",
          2180 => x"80900481",
          2181 => x"d3b80c9f",
          2182 => x"a72d81d3",
          2183 => x"b8088380",
          2184 => x"900481d3",
          2185 => x"b80c9fec",
          2186 => x"2d81d3b8",
          2187 => x"08838090",
          2188 => x"0481d3b8",
          2189 => x"0ca08a2d",
          2190 => x"81d3b808",
          2191 => x"83809004",
          2192 => x"81d3b80c",
          2193 => x"a6de2d81",
          2194 => x"d3b80883",
          2195 => x"80900481",
          2196 => x"d3b80ca7",
          2197 => x"f22d81d3",
          2198 => x"b8088380",
          2199 => x"900481d3",
          2200 => x"b80ca0ab",
          2201 => x"2d81d3b8",
          2202 => x"08838090",
          2203 => x"0481d3b8",
          2204 => x"0ca88f2d",
          2205 => x"81d3b808",
          2206 => x"83809004",
          2207 => x"81d3b80c",
          2208 => x"aaa52d81",
          2209 => x"d3b80883",
          2210 => x"80900481",
          2211 => x"d3b80ca6",
          2212 => x"842d81d3",
          2213 => x"b8088380",
          2214 => x"900481d3",
          2215 => x"b80ca69a",
          2216 => x"2d81d3b8",
          2217 => x"08838090",
          2218 => x"0481d3b8",
          2219 => x"0ca6be2d",
          2220 => x"81d3b808",
          2221 => x"83809004",
          2222 => x"81d3b80c",
          2223 => x"96e72d81",
          2224 => x"d3b80883",
          2225 => x"80900481",
          2226 => x"d3b80c97",
          2227 => x"b52d81d3",
          2228 => x"b8088380",
          2229 => x"900481d3",
          2230 => x"b80c8fbf",
          2231 => x"2d81d3b8",
          2232 => x"08838090",
          2233 => x"0481d3b8",
          2234 => x"0c90f72d",
          2235 => x"81d3b808",
          2236 => x"83809004",
          2237 => x"81d3b80c",
          2238 => x"92d12d81",
          2239 => x"d3b80883",
          2240 => x"80900481",
          2241 => x"d3b80c80",
          2242 => x"ded92d81",
          2243 => x"d3b80883",
          2244 => x"80900481",
          2245 => x"d3b80c80",
          2246 => x"edd02d81",
          2247 => x"d3b80883",
          2248 => x"80900481",
          2249 => x"d3b80c80",
          2250 => x"e3df2d81",
          2251 => x"d3b80883",
          2252 => x"80900481",
          2253 => x"d3b80c80",
          2254 => x"e7c62d81",
          2255 => x"d3b80883",
          2256 => x"80900481",
          2257 => x"d3b80c80",
          2258 => x"f2f92d81",
          2259 => x"d3b80883",
          2260 => x"80900481",
          2261 => x"d3b80c80",
          2262 => x"fced2d81",
          2263 => x"d3b80883",
          2264 => x"80900481",
          2265 => x"d3b80c80",
          2266 => x"ec812d81",
          2267 => x"d3b80883",
          2268 => x"80900481",
          2269 => x"d3b80c80",
          2270 => x"f7a42d81",
          2271 => x"d3b80883",
          2272 => x"80900481",
          2273 => x"d3b80c80",
          2274 => x"f8c82d81",
          2275 => x"d3b80883",
          2276 => x"80900481",
          2277 => x"d3b80c80",
          2278 => x"f8f12d81",
          2279 => x"d3b80883",
          2280 => x"80900481",
          2281 => x"d3b80c81",
          2282 => x"82812d81",
          2283 => x"d3b80883",
          2284 => x"80900481",
          2285 => x"d3b80c80",
          2286 => x"fef92d81",
          2287 => x"d3b80883",
          2288 => x"80900481",
          2289 => x"d3b80c81",
          2290 => x"84da2d81",
          2291 => x"d3b80883",
          2292 => x"80900481",
          2293 => x"d3b80c80",
          2294 => x"f9e72d81",
          2295 => x"d3b80883",
          2296 => x"80900481",
          2297 => x"d3b80c81",
          2298 => x"87de2d81",
          2299 => x"d3b80883",
          2300 => x"80900481",
          2301 => x"d3b80c81",
          2302 => x"88e42d81",
          2303 => x"d3b80883",
          2304 => x"80900481",
          2305 => x"d3b80c80",
          2306 => x"eeb02d81",
          2307 => x"d3b80883",
          2308 => x"80900481",
          2309 => x"d3b80c80",
          2310 => x"ee892d81",
          2311 => x"d3b80883",
          2312 => x"80900481",
          2313 => x"d3b80c80",
          2314 => x"efb32d81",
          2315 => x"d3b80883",
          2316 => x"80900481",
          2317 => x"d3b80c80",
          2318 => x"fac12d81",
          2319 => x"d3b80883",
          2320 => x"80900481",
          2321 => x"d3b80c81",
          2322 => x"89dd2d81",
          2323 => x"d3b80883",
          2324 => x"80900481",
          2325 => x"d3b80c81",
          2326 => x"8be82d81",
          2327 => x"d3b80883",
          2328 => x"80900481",
          2329 => x"d3b80c81",
          2330 => x"8fd52d81",
          2331 => x"d3b80883",
          2332 => x"80900481",
          2333 => x"d3b80c80",
          2334 => x"ddea2d81",
          2335 => x"d3b80883",
          2336 => x"80900481",
          2337 => x"d3b80c81",
          2338 => x"92c62d81",
          2339 => x"d3b80883",
          2340 => x"80900481",
          2341 => x"d3b80cad",
          2342 => x"e52d81d3",
          2343 => x"b8088380",
          2344 => x"900481d3",
          2345 => x"b80cafbe",
          2346 => x"2d81d3b8",
          2347 => x"08838090",
          2348 => x"0481d3b8",
          2349 => x"0cb1982d",
          2350 => x"81d3b808",
          2351 => x"83809004",
          2352 => x"81d3b80c",
          2353 => x"8fe82d81",
          2354 => x"d3b80883",
          2355 => x"80900481",
          2356 => x"d3b80c90",
          2357 => x"cd2d81d3",
          2358 => x"b8088380",
          2359 => x"900481d3",
          2360 => x"b80c93da",
          2361 => x"2d81d3b8",
          2362 => x"08838090",
          2363 => x"0481d3b8",
          2364 => x"0c819fc4",
          2365 => x"2d81d3b8",
          2366 => x"08838090",
          2367 => x"0481d3ac",
          2368 => x"7081f6b0",
          2369 => x"278e3880",
          2370 => x"71708405",
          2371 => x"530c0b0b",
          2372 => x"0b8a8004",
          2373 => x"84805181",
          2374 => x"afc1043c",
          2375 => x"0481d3b8",
          2376 => x"080281d3",
          2377 => x"b80cfd3d",
          2378 => x"0d805381",
          2379 => x"d3b8088c",
          2380 => x"05085281",
          2381 => x"d3b80888",
          2382 => x"05085180",
          2383 => x"c53f81d3",
          2384 => x"ac087081",
          2385 => x"d3ac0c54",
          2386 => x"853d0d81",
          2387 => x"d3b80c04",
          2388 => x"81d3b808",
          2389 => x"0281d3b8",
          2390 => x"0cfd3d0d",
          2391 => x"815381d3",
          2392 => x"b8088c05",
          2393 => x"085281d3",
          2394 => x"b8088805",
          2395 => x"0851933f",
          2396 => x"81d3ac08",
          2397 => x"7081d3ac",
          2398 => x"0c54853d",
          2399 => x"0d81d3b8",
          2400 => x"0c0481d3",
          2401 => x"b8080281",
          2402 => x"d3b80cfd",
          2403 => x"3d0d810b",
          2404 => x"81d3b808",
          2405 => x"fc050c80",
          2406 => x"0b81d3b8",
          2407 => x"08f8050c",
          2408 => x"81d3b808",
          2409 => x"8c050881",
          2410 => x"d3b80888",
          2411 => x"050827b9",
          2412 => x"3881d3b8",
          2413 => x"08fc0508",
          2414 => x"802eae38",
          2415 => x"800b81d3",
          2416 => x"b8088c05",
          2417 => x"0824a238",
          2418 => x"81d3b808",
          2419 => x"8c050810",
          2420 => x"81d3b808",
          2421 => x"8c050c81",
          2422 => x"d3b808fc",
          2423 => x"05081081",
          2424 => x"d3b808fc",
          2425 => x"050cffb8",
          2426 => x"3981d3b8",
          2427 => x"08fc0508",
          2428 => x"802e80e1",
          2429 => x"3881d3b8",
          2430 => x"088c0508",
          2431 => x"81d3b808",
          2432 => x"88050826",
          2433 => x"ad3881d3",
          2434 => x"b8088805",
          2435 => x"0881d3b8",
          2436 => x"088c0508",
          2437 => x"3181d3b8",
          2438 => x"0888050c",
          2439 => x"81d3b808",
          2440 => x"f8050881",
          2441 => x"d3b808fc",
          2442 => x"05080781",
          2443 => x"d3b808f8",
          2444 => x"050c81d3",
          2445 => x"b808fc05",
          2446 => x"08812a81",
          2447 => x"d3b808fc",
          2448 => x"050c81d3",
          2449 => x"b8088c05",
          2450 => x"08812a81",
          2451 => x"d3b8088c",
          2452 => x"050cff95",
          2453 => x"3981d3b8",
          2454 => x"08900508",
          2455 => x"802e9338",
          2456 => x"81d3b808",
          2457 => x"88050870",
          2458 => x"81d3b808",
          2459 => x"f4050c51",
          2460 => x"913981d3",
          2461 => x"b808f805",
          2462 => x"087081d3",
          2463 => x"b808f405",
          2464 => x"0c5181d3",
          2465 => x"b808f405",
          2466 => x"0881d3ac",
          2467 => x"0c853d0d",
          2468 => x"81d3b80c",
          2469 => x"04fc3d0d",
          2470 => x"76797102",
          2471 => x"8c059f05",
          2472 => x"33575553",
          2473 => x"55837227",
          2474 => x"8a387483",
          2475 => x"06517080",
          2476 => x"2ea438ff",
          2477 => x"125271ff",
          2478 => x"2e933873",
          2479 => x"73708105",
          2480 => x"5534ff12",
          2481 => x"5271ff2e",
          2482 => x"098106ef",
          2483 => x"387481d3",
          2484 => x"ac0c863d",
          2485 => x"0d047474",
          2486 => x"882b7507",
          2487 => x"7071902b",
          2488 => x"07515451",
          2489 => x"8f7227a5",
          2490 => x"38727170",
          2491 => x"8405530c",
          2492 => x"72717084",
          2493 => x"05530c72",
          2494 => x"71708405",
          2495 => x"530c7271",
          2496 => x"70840553",
          2497 => x"0cf01252",
          2498 => x"718f26dd",
          2499 => x"38837227",
          2500 => x"90387271",
          2501 => x"70840553",
          2502 => x"0cfc1252",
          2503 => x"718326f2",
          2504 => x"387053ff",
          2505 => x"8e39fb3d",
          2506 => x"0d777970",
          2507 => x"72078306",
          2508 => x"53545270",
          2509 => x"93387173",
          2510 => x"73085456",
          2511 => x"54717308",
          2512 => x"2e80c638",
          2513 => x"73755452",
          2514 => x"71337081",
          2515 => x"ff065254",
          2516 => x"70802e9d",
          2517 => x"38723355",
          2518 => x"70752e09",
          2519 => x"81069538",
          2520 => x"81128114",
          2521 => x"71337081",
          2522 => x"ff065456",
          2523 => x"545270e5",
          2524 => x"38723355",
          2525 => x"7381ff06",
          2526 => x"7581ff06",
          2527 => x"71713181",
          2528 => x"d3ac0c52",
          2529 => x"52873d0d",
          2530 => x"04710970",
          2531 => x"f7fbfdff",
          2532 => x"140670f8",
          2533 => x"84828180",
          2534 => x"06515151",
          2535 => x"70973884",
          2536 => x"14841671",
          2537 => x"08545654",
          2538 => x"7175082e",
          2539 => x"dc387375",
          2540 => x"5452ff94",
          2541 => x"39800b81",
          2542 => x"d3ac0c87",
          2543 => x"3d0d04fe",
          2544 => x"3d0d8070",
          2545 => x"54527188",
          2546 => x"2b52879b",
          2547 => x"3f81d3ac",
          2548 => x"0881ff06",
          2549 => x"72078114",
          2550 => x"54528373",
          2551 => x"25e83871",
          2552 => x"81d3ac0c",
          2553 => x"843d0d04",
          2554 => x"fc3d0d76",
          2555 => x"70087053",
          2556 => x"55557380",
          2557 => x"2e80cd38",
          2558 => x"73335170",
          2559 => x"a02e0981",
          2560 => x"068c3881",
          2561 => x"14703352",
          2562 => x"5470a02e",
          2563 => x"f6387352",
          2564 => x"84398112",
          2565 => x"52807233",
          2566 => x"525370a0",
          2567 => x"2e833881",
          2568 => x"53703070",
          2569 => x"9f2a7406",
          2570 => x"515170e6",
          2571 => x"38713351",
          2572 => x"70a02e09",
          2573 => x"81068838",
          2574 => x"80727081",
          2575 => x"05543471",
          2576 => x"750c7351",
          2577 => x"7081d3ac",
          2578 => x"0c863d0d",
          2579 => x"04fc3d0d",
          2580 => x"76537208",
          2581 => x"802e9138",
          2582 => x"863dfc05",
          2583 => x"52725199",
          2584 => x"c43f81d3",
          2585 => x"ac088538",
          2586 => x"80538339",
          2587 => x"74537281",
          2588 => x"d3ac0c86",
          2589 => x"3d0d04f5",
          2590 => x"3d0d7d82",
          2591 => x"1133ff05",
          2592 => x"5b5c815b",
          2593 => x"798b2681",
          2594 => x"bf38831c",
          2595 => x"33ff055a",
          2596 => x"825b799e",
          2597 => x"2681b138",
          2598 => x"841c335a",
          2599 => x"835b7997",
          2600 => x"2681a538",
          2601 => x"851c335a",
          2602 => x"845b79bb",
          2603 => x"26819938",
          2604 => x"861c335a",
          2605 => x"855b79bb",
          2606 => x"26818d38",
          2607 => x"881c225a",
          2608 => x"865b7987",
          2609 => x"e7268180",
          2610 => x"388a1c22",
          2611 => x"5a875b79",
          2612 => x"87e72680",
          2613 => x"f3388a1c",
          2614 => x"2259881c",
          2615 => x"2258861c",
          2616 => x"3357851c",
          2617 => x"3356841c",
          2618 => x"3355831c",
          2619 => x"3354821c",
          2620 => x"33537b22",
          2621 => x"5281b68c",
          2622 => x"5194893f",
          2623 => x"87c0989c",
          2624 => x"5b817b0c",
          2625 => x"7b2287c0",
          2626 => x"98bc0c82",
          2627 => x"1c3387c0",
          2628 => x"98b80c83",
          2629 => x"1c3387c0",
          2630 => x"98b40c84",
          2631 => x"1c3387c0",
          2632 => x"98b00c85",
          2633 => x"1c3387c0",
          2634 => x"98ac0c86",
          2635 => x"1c3387c0",
          2636 => x"98a80c88",
          2637 => x"1c2287c0",
          2638 => x"98a40c8a",
          2639 => x"1c2287c0",
          2640 => x"98a00c80",
          2641 => x"7b0c805b",
          2642 => x"7a81d3ac",
          2643 => x"0c8d3d0d",
          2644 => x"04f53d0d",
          2645 => x"7d5a87c0",
          2646 => x"989c5c81",
          2647 => x"7c0c87c0",
          2648 => x"98bc085b",
          2649 => x"7a7a2387",
          2650 => x"c098b808",
          2651 => x"5b7a821b",
          2652 => x"3487c098",
          2653 => x"b4085b7a",
          2654 => x"831b3487",
          2655 => x"c098b008",
          2656 => x"5b7a841b",
          2657 => x"3487c098",
          2658 => x"ac085b7a",
          2659 => x"851b3487",
          2660 => x"c098a808",
          2661 => x"5b7a861b",
          2662 => x"3487c098",
          2663 => x"a4085b7a",
          2664 => x"881b2387",
          2665 => x"c098a008",
          2666 => x"5b7a8a1b",
          2667 => x"23807c0c",
          2668 => x"8a1a2259",
          2669 => x"881a2258",
          2670 => x"861a3357",
          2671 => x"851a3356",
          2672 => x"841a3355",
          2673 => x"831a3354",
          2674 => x"821a3353",
          2675 => x"79225281",
          2676 => x"b68c5192",
          2677 => x"af3f8d3d",
          2678 => x"0d04803d",
          2679 => x"0d028b05",
          2680 => x"33703070",
          2681 => x"9f2a5151",
          2682 => x"51700b0b",
          2683 => x"81cba434",
          2684 => x"823d0d04",
          2685 => x"fd3d0d75",
          2686 => x"0b0b81cb",
          2687 => x"a4335454",
          2688 => x"87c09484",
          2689 => x"5172802e",
          2690 => x"863887c0",
          2691 => x"94945170",
          2692 => x"0870962a",
          2693 => x"70810651",
          2694 => x"52527080",
          2695 => x"2e8c3871",
          2696 => x"912a7081",
          2697 => x"06515170",
          2698 => x"d7387196",
          2699 => x"2a813270",
          2700 => x"81065151",
          2701 => x"70802e8d",
          2702 => x"3871932a",
          2703 => x"70810651",
          2704 => x"5170ffbc",
          2705 => x"380b0b81",
          2706 => x"cba43351",
          2707 => x"87c09480",
          2708 => x"5270802e",
          2709 => x"863887c0",
          2710 => x"94905273",
          2711 => x"720c7381",
          2712 => x"d3ac0c85",
          2713 => x"3d0d04fd",
          2714 => x"3d0d0297",
          2715 => x"05330b0b",
          2716 => x"81cba433",
          2717 => x"545487c0",
          2718 => x"94845172",
          2719 => x"802e8638",
          2720 => x"87c09494",
          2721 => x"51700870",
          2722 => x"962a7081",
          2723 => x"06515252",
          2724 => x"70802e8c",
          2725 => x"3871912a",
          2726 => x"70810651",
          2727 => x"5170d738",
          2728 => x"71962a81",
          2729 => x"32708106",
          2730 => x"51517080",
          2731 => x"2e8d3871",
          2732 => x"932a7081",
          2733 => x"06515170",
          2734 => x"ffbc380b",
          2735 => x"0b81cba4",
          2736 => x"335187c0",
          2737 => x"94805270",
          2738 => x"802e8638",
          2739 => x"87c09490",
          2740 => x"5273720c",
          2741 => x"853d0d04",
          2742 => x"fb3d0d77",
          2743 => x"54807433",
          2744 => x"52567076",
          2745 => x"2e80f738",
          2746 => x"73708105",
          2747 => x"55330b0b",
          2748 => x"81cba433",
          2749 => x"545587c0",
          2750 => x"94845172",
          2751 => x"802e8638",
          2752 => x"87c09494",
          2753 => x"51700870",
          2754 => x"962a7081",
          2755 => x"06515252",
          2756 => x"70802e8c",
          2757 => x"3871912a",
          2758 => x"70810651",
          2759 => x"5170d738",
          2760 => x"71962a81",
          2761 => x"32708106",
          2762 => x"51517080",
          2763 => x"2e8d3871",
          2764 => x"932a7081",
          2765 => x"06515170",
          2766 => x"ffbc380b",
          2767 => x"0b81cba4",
          2768 => x"335187c0",
          2769 => x"94805270",
          2770 => x"802e8638",
          2771 => x"87c09490",
          2772 => x"5274720c",
          2773 => x"81167433",
          2774 => x"525670ff",
          2775 => x"8b387581",
          2776 => x"d3ac0c87",
          2777 => x"3d0d04ff",
          2778 => x"3d0d0b0b",
          2779 => x"81cba433",
          2780 => x"5287c094",
          2781 => x"84517180",
          2782 => x"2e863887",
          2783 => x"c0949451",
          2784 => x"70087082",
          2785 => x"2a708106",
          2786 => x"51515170",
          2787 => x"802ee238",
          2788 => x"0b0b81cb",
          2789 => x"a4335187",
          2790 => x"c0948052",
          2791 => x"70802e86",
          2792 => x"3887c094",
          2793 => x"90527108",
          2794 => x"7081ff06",
          2795 => x"81d3ac0c",
          2796 => x"51833d0d",
          2797 => x"04ff3d0d",
          2798 => x"0b0b81cb",
          2799 => x"a4335187",
          2800 => x"c0948452",
          2801 => x"70802e86",
          2802 => x"3887c094",
          2803 => x"94527108",
          2804 => x"70822a70",
          2805 => x"81065151",
          2806 => x"51ff5270",
          2807 => x"802ea238",
          2808 => x"0b0b81cb",
          2809 => x"a4335187",
          2810 => x"c0948052",
          2811 => x"70802e86",
          2812 => x"3887c094",
          2813 => x"90527108",
          2814 => x"70982b70",
          2815 => x"982c5153",
          2816 => x"517181d3",
          2817 => x"ac0c833d",
          2818 => x"0d04fd3d",
          2819 => x"0d87c09e",
          2820 => x"80700870",
          2821 => x"9c2a8a06",
          2822 => x"51525370",
          2823 => x"802e839f",
          2824 => x"3881cba8",
          2825 => x"0b87c09e",
          2826 => x"9c08710c",
          2827 => x"841187c0",
          2828 => x"9ea00871",
          2829 => x"0c528811",
          2830 => x"87c09e8c",
          2831 => x"08710c52",
          2832 => x"8c1187c0",
          2833 => x"9e900871",
          2834 => x"0c529011",
          2835 => x"87c09e94",
          2836 => x"08710c52",
          2837 => x"941187c0",
          2838 => x"9e980871",
          2839 => x"0c529811",
          2840 => x"87c09ea4",
          2841 => x"08710c52",
          2842 => x"9c1187c0",
          2843 => x"9ea80871",
          2844 => x"0c52a011",
          2845 => x"87c09eac",
          2846 => x"08710c52",
          2847 => x"73085252",
          2848 => x"70a41323",
          2849 => x"a81287c0",
          2850 => x"9e840871",
          2851 => x"0c51810b",
          2852 => x"ac1334ad",
          2853 => x"1252800b",
          2854 => x"87c09e88",
          2855 => x"0870a080",
          2856 => x"06515253",
          2857 => x"70802e83",
          2858 => x"38815372",
          2859 => x"7234800b",
          2860 => x"87c09e88",
          2861 => x"08708180",
          2862 => x"80065152",
          2863 => x"5270802e",
          2864 => x"83388152",
          2865 => x"7181cbd6",
          2866 => x"34800b87",
          2867 => x"c09e8808",
          2868 => x"7080c080",
          2869 => x"06515252",
          2870 => x"70802e83",
          2871 => x"38815271",
          2872 => x"81cbd734",
          2873 => x"800b87c0",
          2874 => x"9e880870",
          2875 => x"90800651",
          2876 => x"52527080",
          2877 => x"2e833881",
          2878 => x"527181cb",
          2879 => x"d834800b",
          2880 => x"87c09e88",
          2881 => x"08708880",
          2882 => x"06515252",
          2883 => x"70802e83",
          2884 => x"38815271",
          2885 => x"81cbd934",
          2886 => x"800b87c0",
          2887 => x"9e880870",
          2888 => x"84800651",
          2889 => x"52527080",
          2890 => x"2e833881",
          2891 => x"527181cb",
          2892 => x"da34800b",
          2893 => x"87c09e88",
          2894 => x"08708280",
          2895 => x"06515252",
          2896 => x"70802e83",
          2897 => x"38815271",
          2898 => x"81cbdb34",
          2899 => x"800b87c0",
          2900 => x"9e880870",
          2901 => x"81800651",
          2902 => x"52527080",
          2903 => x"2e833881",
          2904 => x"527181cb",
          2905 => x"dc3481cb",
          2906 => x"dd5287c0",
          2907 => x"9e887008",
          2908 => x"7080e006",
          2909 => x"70862c51",
          2910 => x"51525370",
          2911 => x"72708105",
          2912 => x"54347154",
          2913 => x"80730870",
          2914 => x"90065152",
          2915 => x"5270802e",
          2916 => x"83388152",
          2917 => x"71743480",
          2918 => x"0b87c09e",
          2919 => x"88087088",
          2920 => x"06515252",
          2921 => x"70802e83",
          2922 => x"38815271",
          2923 => x"81cbdf34",
          2924 => x"87c09e88",
          2925 => x"08708706",
          2926 => x"51517081",
          2927 => x"cbe03485",
          2928 => x"3d0d04fc",
          2929 => x"3d0d81b6",
          2930 => x"a45184be",
          2931 => x"3f81cbd4",
          2932 => x"33547380",
          2933 => x"2e883881",
          2934 => x"b6b85184",
          2935 => x"ad3f81b6",
          2936 => x"cc5184a6",
          2937 => x"3f81cbd5",
          2938 => x"70335555",
          2939 => x"73802e91",
          2940 => x"38d71508",
          2941 => x"5381cba8",
          2942 => x"085281b6",
          2943 => x"e4518a84",
          2944 => x"3f81cbd6",
          2945 => x"70335555",
          2946 => x"73802e90",
          2947 => x"38de1508",
          2948 => x"53da1508",
          2949 => x"5281b78c",
          2950 => x"5189e93f",
          2951 => x"81cbd770",
          2952 => x"33555573",
          2953 => x"8a388115",
          2954 => x"33547380",
          2955 => x"2e933881",
          2956 => x"cbbc7008",
          2957 => x"54fc1108",
          2958 => x"535481b7",
          2959 => x"b05189c4",
          2960 => x"3f81cbd9",
          2961 => x"33547380",
          2962 => x"2e883881",
          2963 => x"b7d45183",
          2964 => x"b93f81cb",
          2965 => x"da335473",
          2966 => x"802e8838",
          2967 => x"81b7e051",
          2968 => x"83a83f81",
          2969 => x"cbdb3354",
          2970 => x"73802e88",
          2971 => x"3881b7ec",
          2972 => x"5183973f",
          2973 => x"81cbdc70",
          2974 => x"33555573",
          2975 => x"802e8c38",
          2976 => x"81153352",
          2977 => x"81b7f851",
          2978 => x"88fa3f81",
          2979 => x"cbde3354",
          2980 => x"73802e88",
          2981 => x"3881b898",
          2982 => x"5182ef3f",
          2983 => x"81cbdf70",
          2984 => x"33555573",
          2985 => x"802e8c38",
          2986 => x"81153352",
          2987 => x"81b8b451",
          2988 => x"88d23f81",
          2989 => x"b8d05182",
          2990 => x"d13f81cb",
          2991 => x"c0707070",
          2992 => x"84055208",
          2993 => x"5481b8dc",
          2994 => x"53555588",
          2995 => x"b73f7308",
          2996 => x"5281b984",
          2997 => x"5188ad3f",
          2998 => x"88150852",
          2999 => x"81b9ac51",
          3000 => x"88a23f8c",
          3001 => x"15225281",
          3002 => x"b9d45188",
          3003 => x"973f9015",
          3004 => x"085281b9",
          3005 => x"fc51888c",
          3006 => x"3f863d0d",
          3007 => x"04ff3d0d",
          3008 => x"028e0533",
          3009 => x"52718526",
          3010 => x"bb387110",
          3011 => x"100b0b81",
          3012 => x"b0a80552",
          3013 => x"71080481",
          3014 => x"baa451f7",
          3015 => x"bb3fac39",
          3016 => x"81baac51",
          3017 => x"f7b23fa3",
          3018 => x"3981bab4",
          3019 => x"51f7a93f",
          3020 => x"9a3981ba",
          3021 => x"bc51f7a0",
          3022 => x"3f913981",
          3023 => x"bac051f7",
          3024 => x"973f8839",
          3025 => x"81bac851",
          3026 => x"f78e3f83",
          3027 => x"3d0d0471",
          3028 => x"88800c04",
          3029 => x"800b87c0",
          3030 => x"96840c04",
          3031 => x"ff3d0d87",
          3032 => x"c0968470",
          3033 => x"08525280",
          3034 => x"720c7074",
          3035 => x"077081cb",
          3036 => x"e40c720c",
          3037 => x"833d0d04",
          3038 => x"ff3d0d87",
          3039 => x"c0968470",
          3040 => x"0881cbe4",
          3041 => x"0c528072",
          3042 => x"0c730970",
          3043 => x"81cbe408",
          3044 => x"067081cb",
          3045 => x"e40c730c",
          3046 => x"51833d0d",
          3047 => x"0481cbe4",
          3048 => x"0887c096",
          3049 => x"840c04fe",
          3050 => x"3d0d0293",
          3051 => x"05335372",
          3052 => x"8a2e0981",
          3053 => x"0685388d",
          3054 => x"51ed3f81",
          3055 => x"d3c40880",
          3056 => x"2e953881",
          3057 => x"d3c40852",
          3058 => x"72723481",
          3059 => x"d3c40881",
          3060 => x"0581d3c4",
          3061 => x"0c923981",
          3062 => x"d3bc0880",
          3063 => x"2e8a3872",
          3064 => x"5181d3bc",
          3065 => x"0852712d",
          3066 => x"843d0d04",
          3067 => x"fe3d0d02",
          3068 => x"97053381",
          3069 => x"d3bc0876",
          3070 => x"81d3bc0c",
          3071 => x"5451ffa7",
          3072 => x"3f7281d3",
          3073 => x"bc0c843d",
          3074 => x"0d04fe3d",
          3075 => x"0d747033",
          3076 => x"53537180",
          3077 => x"2e913872",
          3078 => x"70810554",
          3079 => x"3351ff87",
          3080 => x"3f723352",
          3081 => x"71f13884",
          3082 => x"3d0d04fd",
          3083 => x"3d0d7681",
          3084 => x"d3bc0877",
          3085 => x"81d3bc0c",
          3086 => x"71335455",
          3087 => x"5371802e",
          3088 => x"91387270",
          3089 => x"81055433",
          3090 => x"51fedc3f",
          3091 => x"72335271",
          3092 => x"f1387381",
          3093 => x"d3bc0c85",
          3094 => x"3d0d04ec",
          3095 => x"3d0d6668",
          3096 => x"5d597870",
          3097 => x"81055a33",
          3098 => x"5675802e",
          3099 => x"85923875",
          3100 => x"a52e8838",
          3101 => x"7551feaf",
          3102 => x"3fe83980",
          3103 => x"707a7081",
          3104 => x"055c3358",
          3105 => x"5e5a75b0",
          3106 => x"2e098106",
          3107 => x"8c388179",
          3108 => x"7081055b",
          3109 => x"33575d92",
          3110 => x"3975ad2e",
          3111 => x"0981068a",
          3112 => x"38827970",
          3113 => x"81055b33",
          3114 => x"575d75aa",
          3115 => x"2e098106",
          3116 => x"92387b84",
          3117 => x"1d71087b",
          3118 => x"7081055d",
          3119 => x"33595c5d",
          3120 => x"539f39d0",
          3121 => x"16537289",
          3122 => x"26973879",
          3123 => x"8a2916d0",
          3124 => x"05797081",
          3125 => x"055b33d0",
          3126 => x"1155575a",
          3127 => x"897327eb",
          3128 => x"387580ec",
          3129 => x"32703070",
          3130 => x"72078025",
          3131 => x"7880cc32",
          3132 => x"70307072",
          3133 => x"07802573",
          3134 => x"07535952",
          3135 => x"52545473",
          3136 => x"802e8c38",
          3137 => x"7c840779",
          3138 => x"7081055b",
          3139 => x"33575d75",
          3140 => x"802e83ec",
          3141 => x"38755580",
          3142 => x"e0762789",
          3143 => x"38e01670",
          3144 => x"81ff0656",
          3145 => x"53ffbe15",
          3146 => x"53729626",
          3147 => x"81983872",
          3148 => x"101081b0",
          3149 => x"c0055372",
          3150 => x"08047b84",
          3151 => x"1d710857",
          3152 => x"5d538075",
          3153 => x"33545472",
          3154 => x"742e8d38",
          3155 => x"81147016",
          3156 => x"70335154",
          3157 => x"5472f538",
          3158 => x"7c812a70",
          3159 => x"81065153",
          3160 => x"72a33873",
          3161 => x"81155553",
          3162 => x"727a2799",
          3163 => x"387c812a",
          3164 => x"810656a0",
          3165 => x"51fcb03f",
          3166 => x"758b3873",
          3167 => x"81155553",
          3168 => x"797326ef",
          3169 => x"387451fd",
          3170 => x"813f7381",
          3171 => x"15555372",
          3172 => x"7a27fdce",
          3173 => x"38a051fc",
          3174 => x"8e3f7381",
          3175 => x"15555379",
          3176 => x"7326f238",
          3177 => x"fdbc397b",
          3178 => x"841d8312",
          3179 => x"33535d53",
          3180 => x"fbf53ffd",
          3181 => x"ad39825b",
          3182 => x"9539885b",
          3183 => x"91398a5b",
          3184 => x"8d39905b",
          3185 => x"89397551",
          3186 => x"fbdd3ffd",
          3187 => x"95397c82",
          3188 => x"2a708106",
          3189 => x"51537280",
          3190 => x"2e8b387b",
          3191 => x"841d7108",
          3192 => x"595d539c",
          3193 => x"397480c4",
          3194 => x"2e098106",
          3195 => x"8b387b84",
          3196 => x"1d710859",
          3197 => x"5d538939",
          3198 => x"7b841d71",
          3199 => x"08595d53",
          3200 => x"7480c432",
          3201 => x"70307072",
          3202 => x"07802570",
          3203 => x"807b2406",
          3204 => x"51525553",
          3205 => x"72802e88",
          3206 => x"3876307d",
          3207 => x"90075e57",
          3208 => x"80587a52",
          3209 => x"7651e6a8",
          3210 => x"3f81d3ac",
          3211 => x"0881ff06",
          3212 => x"7b537752",
          3213 => x"55e5e63f",
          3214 => x"81d3ac08",
          3215 => x"57897527",
          3216 => x"993874a7",
          3217 => x"167081ff",
          3218 => x"06575454",
          3219 => x"7580f82e",
          3220 => x"89388714",
          3221 => x"7081ff06",
          3222 => x"5653963d",
          3223 => x"7805e005",
          3224 => x"b0165454",
          3225 => x"72743481",
          3226 => x"18773070",
          3227 => x"79079f2a",
          3228 => x"709f7427",
          3229 => x"06515154",
          3230 => x"5872ffa6",
          3231 => x"387c842a",
          3232 => x"70810651",
          3233 => x"5372802e",
          3234 => x"8e38963d",
          3235 => x"7805e005",
          3236 => x"53ad7334",
          3237 => x"81185877",
          3238 => x"7d810654",
          3239 => x"54b05572",
          3240 => x"8338a055",
          3241 => x"7c812a70",
          3242 => x"81065153",
          3243 => x"72a33873",
          3244 => x"81155553",
          3245 => x"727a2799",
          3246 => x"387c812a",
          3247 => x"81065674",
          3248 => x"51f9e43f",
          3249 => x"758b3873",
          3250 => x"81155553",
          3251 => x"797326ef",
          3252 => x"38ff1897",
          3253 => x"3de00511",
          3254 => x"70335354",
          3255 => x"58f9c83f",
          3256 => x"77ef3873",
          3257 => x"81155553",
          3258 => x"727a27fa",
          3259 => x"f538a051",
          3260 => x"f9b53f73",
          3261 => x"81155553",
          3262 => x"797326f2",
          3263 => x"38fae339",
          3264 => x"963d0d04",
          3265 => x"fd3d0d86",
          3266 => x"3d707084",
          3267 => x"05520855",
          3268 => x"527351fa",
          3269 => x"c63f853d",
          3270 => x"0d04fe3d",
          3271 => x"0d7481d3",
          3272 => x"c40c853d",
          3273 => x"88055275",
          3274 => x"51fab03f",
          3275 => x"81d3c408",
          3276 => x"53807334",
          3277 => x"800b81d3",
          3278 => x"c40c843d",
          3279 => x"0d04fd3d",
          3280 => x"0d81d3bc",
          3281 => x"087681d3",
          3282 => x"bc0c873d",
          3283 => x"88055377",
          3284 => x"5253fa87",
          3285 => x"3f7281d3",
          3286 => x"bc0c853d",
          3287 => x"0d04fa3d",
          3288 => x"0d787a57",
          3289 => x"57805381",
          3290 => x"d3c00873",
          3291 => x"2e80fa38",
          3292 => x"86397353",
          3293 => x"80f33980",
          3294 => x"5581d3c0",
          3295 => x"0852712d",
          3296 => x"81d3ac08",
          3297 => x"81ff0654",
          3298 => x"73802ee6",
          3299 => x"38738d2e",
          3300 => x"80ca3873",
          3301 => x"88327030",
          3302 => x"76307078",
          3303 => x"079f2a72",
          3304 => x"80250652",
          3305 => x"54515372",
          3306 => x"802e8e38",
          3307 => x"ff157481",
          3308 => x"ff065255",
          3309 => x"f7f13fc1",
          3310 => x"399f7425",
          3311 => x"ffbb38ff",
          3312 => x"16527472",
          3313 => x"25ffb238",
          3314 => x"76155273",
          3315 => x"72348115",
          3316 => x"7481ff06",
          3317 => x"5255f7cf",
          3318 => x"3fff9e39",
          3319 => x"74175280",
          3320 => x"72348a51",
          3321 => x"f7c13f81",
          3322 => x"537281d3",
          3323 => x"ac0c883d",
          3324 => x"0d04fe3d",
          3325 => x"0d81d3c0",
          3326 => x"087581d3",
          3327 => x"c00c7753",
          3328 => x"765253fe",
          3329 => x"d93f7281",
          3330 => x"d3c00c84",
          3331 => x"3d0d04f8",
          3332 => x"3d0d7a7c",
          3333 => x"5a558070",
          3334 => x"7a0c7508",
          3335 => x"70335654",
          3336 => x"5873a02e",
          3337 => x"09810692",
          3338 => x"38740881",
          3339 => x"05750c74",
          3340 => x"08703355",
          3341 => x"5373a02e",
          3342 => x"f03873ad",
          3343 => x"2e098106",
          3344 => x"8e388175",
          3345 => x"0811760c",
          3346 => x"75087033",
          3347 => x"56545873",
          3348 => x"b02e0981",
          3349 => x"0680d338",
          3350 => x"74088105",
          3351 => x"750c7408",
          3352 => x"70335553",
          3353 => x"7380e22e",
          3354 => x"9a387380",
          3355 => x"f82e0981",
          3356 => x"06a13890",
          3357 => x"0b811476",
          3358 => x"0c750870",
          3359 => x"33565457",
          3360 => x"80c13982",
          3361 => x"75088105",
          3362 => x"760c7508",
          3363 => x"70335654",
          3364 => x"57b13981",
          3365 => x"56a07427",
          3366 => x"818238d0",
          3367 => x"14538056",
          3368 => x"88578973",
          3369 => x"279d3880",
          3370 => x"f339d014",
          3371 => x"53805672",
          3372 => x"892680e8",
          3373 => x"388b3980",
          3374 => x"5680e139",
          3375 => x"805680dc",
          3376 => x"398a5780",
          3377 => x"56a07427",
          3378 => x"80c53880",
          3379 => x"e0742789",
          3380 => x"38e01470",
          3381 => x"81ff0655",
          3382 => x"53d01470",
          3383 => x"81ff0655",
          3384 => x"53907427",
          3385 => x"8e38f914",
          3386 => x"7081ff06",
          3387 => x"55538974",
          3388 => x"27c53873",
          3389 => x"7727c538",
          3390 => x"76762914",
          3391 => x"75088105",
          3392 => x"760c7508",
          3393 => x"70335654",
          3394 => x"5673a026",
          3395 => x"ffbd3877",
          3396 => x"802e8438",
          3397 => x"75305675",
          3398 => x"790c8156",
          3399 => x"7581d3ac",
          3400 => x"0c8a3d0d",
          3401 => x"04f83d0d",
          3402 => x"7a7c5a55",
          3403 => x"80707a0c",
          3404 => x"75087033",
          3405 => x"56545873",
          3406 => x"a02e0981",
          3407 => x"06923874",
          3408 => x"08810575",
          3409 => x"0c740870",
          3410 => x"33555373",
          3411 => x"a02ef038",
          3412 => x"73ad2e09",
          3413 => x"81068e38",
          3414 => x"81750811",
          3415 => x"760c7508",
          3416 => x"70335654",
          3417 => x"5873b02e",
          3418 => x"09810680",
          3419 => x"d3387408",
          3420 => x"8105750c",
          3421 => x"74087033",
          3422 => x"55537380",
          3423 => x"e22e9a38",
          3424 => x"7380f82e",
          3425 => x"098106a1",
          3426 => x"38900b81",
          3427 => x"14760c75",
          3428 => x"08703356",
          3429 => x"545780c1",
          3430 => x"39827508",
          3431 => x"8105760c",
          3432 => x"75087033",
          3433 => x"565457b1",
          3434 => x"398156a0",
          3435 => x"74278182",
          3436 => x"38d01453",
          3437 => x"80568857",
          3438 => x"8973279d",
          3439 => x"3880f339",
          3440 => x"d0145380",
          3441 => x"56728926",
          3442 => x"80e8388b",
          3443 => x"39805680",
          3444 => x"e1398056",
          3445 => x"80dc398a",
          3446 => x"578056a0",
          3447 => x"742780c5",
          3448 => x"3880e074",
          3449 => x"278938e0",
          3450 => x"147081ff",
          3451 => x"065553d0",
          3452 => x"147081ff",
          3453 => x"06555390",
          3454 => x"74278e38",
          3455 => x"f9147081",
          3456 => x"ff065553",
          3457 => x"897427c5",
          3458 => x"38737727",
          3459 => x"c5387676",
          3460 => x"29147508",
          3461 => x"8105760c",
          3462 => x"75087033",
          3463 => x"56545673",
          3464 => x"a026ffbd",
          3465 => x"3877802e",
          3466 => x"84387530",
          3467 => x"5675790c",
          3468 => x"81567581",
          3469 => x"d3ac0c8a",
          3470 => x"3d0d04ff",
          3471 => x"3d0d028f",
          3472 => x"05335181",
          3473 => x"52707226",
          3474 => x"873881cb",
          3475 => x"e8113352",
          3476 => x"7181d3ac",
          3477 => x"0c833d0d",
          3478 => x"04fd3d0d",
          3479 => x"02970533",
          3480 => x"0284059b",
          3481 => x"05335553",
          3482 => x"83517281",
          3483 => x"2680ed38",
          3484 => x"72902987",
          3485 => x"c0928c05",
          3486 => x"51885273",
          3487 => x"802e8438",
          3488 => x"81885271",
          3489 => x"710c7290",
          3490 => x"2987c092",
          3491 => x"8c055181",
          3492 => x"710c850b",
          3493 => x"87c0988c",
          3494 => x"0c705287",
          3495 => x"c0988c54",
          3496 => x"71087082",
          3497 => x"06515170",
          3498 => x"802e8738",
          3499 => x"73085170",
          3500 => x"ef387290",
          3501 => x"2987c092",
          3502 => x"8c057008",
          3503 => x"fc808006",
          3504 => x"53517192",
          3505 => x"3887c098",
          3506 => x"8c085170",
          3507 => x"802e8738",
          3508 => x"7181cbe8",
          3509 => x"143481cb",
          3510 => x"e8133351",
          3511 => x"7081d3ac",
          3512 => x"0c853d0d",
          3513 => x"04f23d0d",
          3514 => x"61636502",
          3515 => x"8c0580c3",
          3516 => x"05335641",
          3517 => x"5d588373",
          3518 => x"525bfebf",
          3519 => x"3f81d3ac",
          3520 => x"0881067b",
          3521 => x"55527181",
          3522 => x"ac388070",
          3523 => x"585d87c0",
          3524 => x"988c7384",
          3525 => x"2b87c092",
          3526 => x"8c1187c0",
          3527 => x"92841272",
          3528 => x"425c575b",
          3529 => x"5685760c",
          3530 => x"87c09280",
          3531 => x"1a7c710c",
          3532 => x"5284750c",
          3533 => x"74087085",
          3534 => x"2a708106",
          3535 => x"51535471",
          3536 => x"802e8e38",
          3537 => x"78085271",
          3538 => x"78708105",
          3539 => x"5a348117",
          3540 => x"5773a206",
          3541 => x"5271802e",
          3542 => x"87387508",
          3543 => x"5271d538",
          3544 => x"75085271",
          3545 => x"802e8738",
          3546 => x"7684802e",
          3547 => x"99388175",
          3548 => x"0c87c092",
          3549 => x"8c1e5372",
          3550 => x"08708206",
          3551 => x"515271f7",
          3552 => x"38ff1b5b",
          3553 => x"8d398480",
          3554 => x"1c811e70",
          3555 => x"81ff065f",
          3556 => x"535c7a80",
          3557 => x"2e903873",
          3558 => x"fc808006",
          3559 => x"52718738",
          3560 => x"7e7d26ff",
          3561 => x"803873fc",
          3562 => x"80800652",
          3563 => x"71802e83",
          3564 => x"38815271",
          3565 => x"547381d3",
          3566 => x"ac0c903d",
          3567 => x"0d04f33d",
          3568 => x"0d606264",
          3569 => x"028c05bf",
          3570 => x"05335640",
          3571 => x"5c578373",
          3572 => x"525afce7",
          3573 => x"3f81d3ac",
          3574 => x"0881067a",
          3575 => x"55527181",
          3576 => x"ae38805c",
          3577 => x"87c0988c",
          3578 => x"73842b87",
          3579 => x"c0928c11",
          3580 => x"87c09284",
          3581 => x"1272415b",
          3582 => x"575a5685",
          3583 => x"760c87c0",
          3584 => x"9280197b",
          3585 => x"710c5282",
          3586 => x"750c8053",
          3587 => x"74087084",
          3588 => x"2a708106",
          3589 => x"51535471",
          3590 => x"802e8c38",
          3591 => x"76708105",
          3592 => x"5833780c",
          3593 => x"81135373",
          3594 => x"812a7081",
          3595 => x"06515271",
          3596 => x"802e8738",
          3597 => x"75085271",
          3598 => x"d3387508",
          3599 => x"5271802e",
          3600 => x"87387284",
          3601 => x"802e9938",
          3602 => x"81750c87",
          3603 => x"c0928c1d",
          3604 => x"53720870",
          3605 => x"82065152",
          3606 => x"71f738ff",
          3607 => x"1a5a8d39",
          3608 => x"811c7081",
          3609 => x"ff068480",
          3610 => x"1d5d5d52",
          3611 => x"79802e90",
          3612 => x"3873fc80",
          3613 => x"80065271",
          3614 => x"87387d7c",
          3615 => x"26fefc38",
          3616 => x"73fc8080",
          3617 => x"06527180",
          3618 => x"2e833881",
          3619 => x"52715473",
          3620 => x"81d3ac0c",
          3621 => x"8f3d0d04",
          3622 => x"f73d0d7d",
          3623 => x"028405af",
          3624 => x"05330288",
          3625 => x"05b30533",
          3626 => x"71545556",
          3627 => x"56fb8c3f",
          3628 => x"81d3ac08",
          3629 => x"81065283",
          3630 => x"5471bc38",
          3631 => x"81547274",
          3632 => x"2ea23872",
          3633 => x"74248838",
          3634 => x"72802e8a",
          3635 => x"38a73972",
          3636 => x"832e9a38",
          3637 => x"a0397490",
          3638 => x"2987c092",
          3639 => x"8c057008",
          3640 => x"51529439",
          3641 => x"88800a76",
          3642 => x"0c80548b",
          3643 => x"39818076",
          3644 => x"0c805483",
          3645 => x"39845473",
          3646 => x"81d3ac0c",
          3647 => x"8b3d0d04",
          3648 => x"ff3d0d73",
          3649 => x"70338112",
          3650 => x"3370882b",
          3651 => x"720781d3",
          3652 => x"ac0c5252",
          3653 => x"52833d0d",
          3654 => x"04fd3d0d",
          3655 => x"75831133",
          3656 => x"82123371",
          3657 => x"902b7188",
          3658 => x"2b078114",
          3659 => x"33710774",
          3660 => x"3371882b",
          3661 => x"0781d3ac",
          3662 => x"0c515456",
          3663 => x"5452853d",
          3664 => x"0d04ff3d",
          3665 => x"0d730284",
          3666 => x"05920522",
          3667 => x"52527072",
          3668 => x"70810554",
          3669 => x"3470882a",
          3670 => x"51707234",
          3671 => x"833d0d04",
          3672 => x"ff3d0d73",
          3673 => x"75525270",
          3674 => x"72708105",
          3675 => x"54347088",
          3676 => x"2a517072",
          3677 => x"70810554",
          3678 => x"3470882a",
          3679 => x"51707270",
          3680 => x"81055434",
          3681 => x"70882a51",
          3682 => x"70723483",
          3683 => x"3d0d04fe",
          3684 => x"3d0d7675",
          3685 => x"77545451",
          3686 => x"70802e93",
          3687 => x"38717081",
          3688 => x"05533373",
          3689 => x"70810555",
          3690 => x"34ff1151",
          3691 => x"70ef3884",
          3692 => x"3d0d04fe",
          3693 => x"3d0d7577",
          3694 => x"76545253",
          3695 => x"72727081",
          3696 => x"055434ff",
          3697 => x"115170f4",
          3698 => x"38843d0d",
          3699 => x"04fc3d0d",
          3700 => x"78777956",
          3701 => x"56537470",
          3702 => x"81055633",
          3703 => x"74708105",
          3704 => x"56337171",
          3705 => x"31ff1656",
          3706 => x"52525272",
          3707 => x"802e8638",
          3708 => x"71802ee2",
          3709 => x"387181d3",
          3710 => x"ac0c863d",
          3711 => x"0d04fe3d",
          3712 => x"0d747671",
          3713 => x"33535452",
          3714 => x"70802e99",
          3715 => x"3870732e",
          3716 => x"94388112",
          3717 => x"70335252",
          3718 => x"70802e89",
          3719 => x"3870732e",
          3720 => x"098106ee",
          3721 => x"38713381",
          3722 => x"d3ac0c84",
          3723 => x"3d0d0480",
          3724 => x"0b81d3ac",
          3725 => x"0c04800b",
          3726 => x"81d3ac0c",
          3727 => x"04f93d0d",
          3728 => x"7956800b",
          3729 => x"83173356",
          3730 => x"5874782e",
          3731 => x"80d73881",
          3732 => x"54b01608",
          3733 => x"53b41670",
          3734 => x"53811733",
          3735 => x"5257fade",
          3736 => x"3f81d3ac",
          3737 => x"08782e09",
          3738 => x"8106b838",
          3739 => x"81d3ac08",
          3740 => x"831734b0",
          3741 => x"1608a417",
          3742 => x"08315574",
          3743 => x"9c170827",
          3744 => x"a4388216",
          3745 => x"33557482",
          3746 => x"2e098106",
          3747 => x"98388154",
          3748 => x"b016089c",
          3749 => x"17080553",
          3750 => x"76528116",
          3751 => x"3351fa9e",
          3752 => x"3f833981",
          3753 => x"587781d3",
          3754 => x"ac0c893d",
          3755 => x"0d04fa3d",
          3756 => x"0d787a56",
          3757 => x"578056b0",
          3758 => x"1708752e",
          3759 => x"af387651",
          3760 => x"fefb3f81",
          3761 => x"d3ac0856",
          3762 => x"81d3ac08",
          3763 => x"9f388154",
          3764 => x"7453b417",
          3765 => x"52811733",
          3766 => x"51f88a3f",
          3767 => x"81d3ac08",
          3768 => x"802e8538",
          3769 => x"ff558156",
          3770 => x"74b0180c",
          3771 => x"7581d3ac",
          3772 => x"0c883d0d",
          3773 => x"04f83d0d",
          3774 => x"7a705257",
          3775 => x"febf3f81",
          3776 => x"d3ac0858",
          3777 => x"81d3ac08",
          3778 => x"81913876",
          3779 => x"33557483",
          3780 => x"2e098106",
          3781 => x"80f03884",
          3782 => x"17335978",
          3783 => x"812e0981",
          3784 => x"0680e338",
          3785 => x"84805381",
          3786 => x"d3ac0852",
          3787 => x"b4177052",
          3788 => x"56fd803f",
          3789 => x"82d4d552",
          3790 => x"84b21751",
          3791 => x"fc843f84",
          3792 => x"8b85a4d2",
          3793 => x"527551fc",
          3794 => x"973f868a",
          3795 => x"85e4f252",
          3796 => x"84981751",
          3797 => x"fc8a3f90",
          3798 => x"17085284",
          3799 => x"9c1751fb",
          3800 => x"ff3f8c17",
          3801 => x"085284a0",
          3802 => x"1751fbf4",
          3803 => x"3fa01708",
          3804 => x"810570b0",
          3805 => x"190c7955",
          3806 => x"53755281",
          3807 => x"173351f8",
          3808 => x"bd3f7784",
          3809 => x"18348053",
          3810 => x"80528117",
          3811 => x"3351fa88",
          3812 => x"3f81d3ac",
          3813 => x"08802e83",
          3814 => x"38815877",
          3815 => x"81d3ac0c",
          3816 => x"8a3d0d04",
          3817 => x"fb3d0d77",
          3818 => x"fe1a9812",
          3819 => x"08fe0555",
          3820 => x"56548056",
          3821 => x"7473278d",
          3822 => x"388a1422",
          3823 => x"707629ac",
          3824 => x"16080557",
          3825 => x"537581d3",
          3826 => x"ac0c873d",
          3827 => x"0d04f93d",
          3828 => x"0d7a7a70",
          3829 => x"08565455",
          3830 => x"81752788",
          3831 => x"38981408",
          3832 => x"75268638",
          3833 => x"815681d9",
          3834 => x"39ff7433",
          3835 => x"54567282",
          3836 => x"2e80f538",
          3837 => x"72822489",
          3838 => x"3872812e",
          3839 => x"8d3881bf",
          3840 => x"3972832e",
          3841 => x"818e3881",
          3842 => x"b6397481",
          3843 => x"2a157089",
          3844 => x"2aa41608",
          3845 => x"05537452",
          3846 => x"57fd933f",
          3847 => x"81d3ac08",
          3848 => x"819f3876",
          3849 => x"83ff0614",
          3850 => x"b4113381",
          3851 => x"1970892a",
          3852 => x"a4180805",
          3853 => x"55765459",
          3854 => x"5953fcf2",
          3855 => x"3f81d3ac",
          3856 => x"0880fe38",
          3857 => x"7683ff06",
          3858 => x"14b41133",
          3859 => x"70882b7a",
          3860 => x"07778106",
          3861 => x"71842a5a",
          3862 => x"525a5153",
          3863 => x"7280e238",
          3864 => x"779fff06",
          3865 => x"5680da39",
          3866 => x"74882aa4",
          3867 => x"15080552",
          3868 => x"7351fcba",
          3869 => x"3f81d3ac",
          3870 => x"0880c638",
          3871 => x"741583ff",
          3872 => x"067405b4",
          3873 => x"0551f8f8",
          3874 => x"3f81d3ac",
          3875 => x"0883ffff",
          3876 => x"0656ae39",
          3877 => x"74872aa4",
          3878 => x"15080552",
          3879 => x"7351fc8e",
          3880 => x"3f81d3ac",
          3881 => x"089b3874",
          3882 => x"822b83fc",
          3883 => x"067405b4",
          3884 => x"0551f8e5",
          3885 => x"3f81d3ac",
          3886 => x"08f00a06",
          3887 => x"56833981",
          3888 => x"567581d3",
          3889 => x"ac0c893d",
          3890 => x"0d04f73d",
          3891 => x"0d7b7d7f",
          3892 => x"58555582",
          3893 => x"57817427",
          3894 => x"82af3873",
          3895 => x"98160827",
          3896 => x"82a73874",
          3897 => x"33537277",
          3898 => x"2e81a838",
          3899 => x"72772489",
          3900 => x"3872812e",
          3901 => x"8d388291",
          3902 => x"3972832e",
          3903 => x"81c93882",
          3904 => x"88397381",
          3905 => x"2a147089",
          3906 => x"2aa41708",
          3907 => x"05537552",
          3908 => x"59fb9b3f",
          3909 => x"81d3ac08",
          3910 => x"5781d3ac",
          3911 => x"0881ea38",
          3912 => x"7883ff06",
          3913 => x"15b41181",
          3914 => x"1b768106",
          3915 => x"565b5158",
          3916 => x"75577280",
          3917 => x"2e8f3875",
          3918 => x"842b9ff0",
          3919 => x"0678338f",
          3920 => x"06710758",
          3921 => x"53767834",
          3922 => x"810b8316",
          3923 => x"3478892a",
          3924 => x"a4160805",
          3925 => x"527451fa",
          3926 => x"d53f81d3",
          3927 => x"ac085781",
          3928 => x"d3ac0881",
          3929 => x"a4387883",
          3930 => x"ff0615b4",
          3931 => x"11758106",
          3932 => x"78842a57",
          3933 => x"55515872",
          3934 => x"8f387588",
          3935 => x"2a783357",
          3936 => x"8f067681",
          3937 => x"f0060754",
          3938 => x"73783481",
          3939 => x"0b831634",
          3940 => x"80f73973",
          3941 => x"882aa416",
          3942 => x"08055274",
          3943 => x"51fa8f3f",
          3944 => x"81d3ac08",
          3945 => x"5781d3ac",
          3946 => x"0880de38",
          3947 => x"7583ffff",
          3948 => x"06527314",
          3949 => x"83ff0675",
          3950 => x"05b40551",
          3951 => x"f7843f81",
          3952 => x"0b831634",
          3953 => x"80c33973",
          3954 => x"872aa416",
          3955 => x"08055274",
          3956 => x"51f9db3f",
          3957 => x"81d3ac08",
          3958 => x"5781d3ac",
          3959 => x"08ab3875",
          3960 => x"f00a0674",
          3961 => x"822b83fc",
          3962 => x"067611b4",
          3963 => x"05705451",
          3964 => x"5456f6a5",
          3965 => x"3f81d3ac",
          3966 => x"088f0a06",
          3967 => x"76075272",
          3968 => x"51f6dd3f",
          3969 => x"810b8316",
          3970 => x"347681d3",
          3971 => x"ac0c8b3d",
          3972 => x"0d04f93d",
          3973 => x"0d797b7d",
          3974 => x"72085858",
          3975 => x"55578174",
          3976 => x"27883898",
          3977 => x"15087426",
          3978 => x"86388256",
          3979 => x"818e3975",
          3980 => x"802eaa38",
          3981 => x"ff537552",
          3982 => x"7451fd8e",
          3983 => x"3f81d3ac",
          3984 => x"085681d3",
          3985 => x"ac0880f4",
          3986 => x"38933982",
          3987 => x"5680ed39",
          3988 => x"815680e8",
          3989 => x"3981d3ac",
          3990 => x"085680e0",
          3991 => x"39735276",
          3992 => x"51faeb3f",
          3993 => x"81d3ac08",
          3994 => x"5681d3ac",
          3995 => x"08802e80",
          3996 => x"c93881d3",
          3997 => x"ac08812e",
          3998 => x"d23881d3",
          3999 => x"ac08ff2e",
          4000 => x"cf388053",
          4001 => x"73527451",
          4002 => x"fcc03f81",
          4003 => x"d3ac08c5",
          4004 => x"38981508",
          4005 => x"fe055490",
          4006 => x"15087427",
          4007 => x"93389015",
          4008 => x"08810590",
          4009 => x"160c8415",
          4010 => x"33810754",
          4011 => x"73841634",
          4012 => x"75549815",
          4013 => x"087626ff",
          4014 => x"a4388056",
          4015 => x"7581d3ac",
          4016 => x"0c893d0d",
          4017 => x"04f53d0d",
          4018 => x"7d7f7108",
          4019 => x"5b5c5c7a",
          4020 => x"95388c19",
          4021 => x"08587780",
          4022 => x"2e883898",
          4023 => x"19087826",
          4024 => x"b7388158",
          4025 => x"b3397a52",
          4026 => x"7b51f9e2",
          4027 => x"3f815574",
          4028 => x"81d3ac08",
          4029 => x"2782e938",
          4030 => x"81d3ac08",
          4031 => x"5581d3ac",
          4032 => x"08ff2e82",
          4033 => x"db3881d3",
          4034 => x"ac085598",
          4035 => x"190881d3",
          4036 => x"ac082682",
          4037 => x"cb387a58",
          4038 => x"80559019",
          4039 => x"08752e82",
          4040 => x"bf388057",
          4041 => x"777b2e09",
          4042 => x"810680db",
          4043 => x"38811b57",
          4044 => x"98190877",
          4045 => x"26833882",
          4046 => x"5776527b",
          4047 => x"51f98f3f",
          4048 => x"81d3ac08",
          4049 => x"56805a81",
          4050 => x"d3ac0881",
          4051 => x"2e098106",
          4052 => x"863881d3",
          4053 => x"ac085a75",
          4054 => x"ff327030",
          4055 => x"70720780",
          4056 => x"25707d07",
          4057 => x"79535152",
          4058 => x"56547381",
          4059 => x"f3387580",
          4060 => x"2e95388c",
          4061 => x"19085681",
          4062 => x"76278a38",
          4063 => x"75981a08",
          4064 => x"27833875",
          4065 => x"58805776",
          4066 => x"80de3877",
          4067 => x"57811757",
          4068 => x"98190877",
          4069 => x"26893882",
          4070 => x"57767826",
          4071 => x"81b63876",
          4072 => x"527b51f8",
          4073 => x"a93f81d3",
          4074 => x"ac085681",
          4075 => x"d3ac0880",
          4076 => x"2eb63880",
          4077 => x"5a81d3ac",
          4078 => x"08812e09",
          4079 => x"81068638",
          4080 => x"81d3ac08",
          4081 => x"5a75ff32",
          4082 => x"70307072",
          4083 => x"07802570",
          4084 => x"7d075152",
          4085 => x"56547380",
          4086 => x"ff387678",
          4087 => x"2e098106",
          4088 => x"ffab3880",
          4089 => x"5580f939",
          4090 => x"ff537652",
          4091 => x"7851f9da",
          4092 => x"3f81d3ac",
          4093 => x"0881d3ac",
          4094 => x"08307081",
          4095 => x"d3ac0807",
          4096 => x"80257d30",
          4097 => x"707f079f",
          4098 => x"2a720652",
          4099 => x"57515656",
          4100 => x"74802e8f",
          4101 => x"3876537a",
          4102 => x"527851f9",
          4103 => x"ad3f81d3",
          4104 => x"ac085675",
          4105 => x"a638768c",
          4106 => x"1a0c9819",
          4107 => x"08fe0554",
          4108 => x"90190874",
          4109 => x"26893890",
          4110 => x"1908ff05",
          4111 => x"901a0c84",
          4112 => x"19338107",
          4113 => x"5473841a",
          4114 => x"349439ff",
          4115 => x"5775812e",
          4116 => x"8d388939",
          4117 => x"80558939",
          4118 => x"75558539",
          4119 => x"81577655",
          4120 => x"7481d3ac",
          4121 => x"0c8d3d0d",
          4122 => x"04f73d0d",
          4123 => x"7b705257",
          4124 => x"f3cb3f81",
          4125 => x"5581d3ac",
          4126 => x"0880db38",
          4127 => x"7c527651",
          4128 => x"f6a23f81",
          4129 => x"d3ac0881",
          4130 => x"d3ac08b0",
          4131 => x"190c5a84",
          4132 => x"80538052",
          4133 => x"b4177052",
          4134 => x"55f2983f",
          4135 => x"74598158",
          4136 => x"80568439",
          4137 => x"7716568a",
          4138 => x"17225575",
          4139 => x"75279738",
          4140 => x"7754751a",
          4141 => x"53785281",
          4142 => x"173351ee",
          4143 => x"813f81d3",
          4144 => x"ac08802e",
          4145 => x"df38800b",
          4146 => x"8a182256",
          4147 => x"5874762e",
          4148 => x"83388158",
          4149 => x"77557481",
          4150 => x"d3ac0c8b",
          4151 => x"3d0d04f8",
          4152 => x"3d0d7a7c",
          4153 => x"71085856",
          4154 => x"5774f080",
          4155 => x"0a268a38",
          4156 => x"749f0653",
          4157 => x"72802e86",
          4158 => x"38825881",
          4159 => x"ae397490",
          4160 => x"180c8817",
          4161 => x"085473aa",
          4162 => x"38753353",
          4163 => x"82732785",
          4164 => x"38a81608",
          4165 => x"54739b38",
          4166 => x"74852a53",
          4167 => x"820b8817",
          4168 => x"225a5872",
          4169 => x"79278183",
          4170 => x"38a81608",
          4171 => x"98180c80",
          4172 => x"d1398a16",
          4173 => x"2270892b",
          4174 => x"54587275",
          4175 => x"26b63873",
          4176 => x"527651f5",
          4177 => x"893f81d3",
          4178 => x"ac085481",
          4179 => x"d3ac08ff",
          4180 => x"2ebf3881",
          4181 => x"0b81d3ac",
          4182 => x"08278b38",
          4183 => x"98160881",
          4184 => x"d3ac0826",
          4185 => x"86388258",
          4186 => x"80c13974",
          4187 => x"73315574",
          4188 => x"7327cc38",
          4189 => x"73527551",
          4190 => x"f4aa3f81",
          4191 => x"d3ac0898",
          4192 => x"180c7394",
          4193 => x"180c8258",
          4194 => x"98170880",
          4195 => x"2e9d3885",
          4196 => x"39815897",
          4197 => x"3974892a",
          4198 => x"98180805",
          4199 => x"98180c74",
          4200 => x"83ff0616",
          4201 => x"b4059c18",
          4202 => x"0c805877",
          4203 => x"81d3ac0c",
          4204 => x"8a3d0d04",
          4205 => x"f93d0d79",
          4206 => x"7b710890",
          4207 => x"1308a005",
          4208 => x"59595955",
          4209 => x"f0800a76",
          4210 => x"27863880",
          4211 => x"0b98160c",
          4212 => x"84539815",
          4213 => x"08802e81",
          4214 => x"da387583",
          4215 => x"ff065473",
          4216 => x"81c13898",
          4217 => x"15088105",
          4218 => x"98160c94",
          4219 => x"15089838",
          4220 => x"75852a88",
          4221 => x"18225953",
          4222 => x"77732681",
          4223 => x"a6387398",
          4224 => x"160c8453",
          4225 => x"81ad398a",
          4226 => x"1722ff11",
          4227 => x"77892a06",
          4228 => x"51537281",
          4229 => x"8e389415",
          4230 => x"08527451",
          4231 => x"f3b03f81",
          4232 => x"d3ac0854",
          4233 => x"8253810b",
          4234 => x"81d3ac08",
          4235 => x"27818438",
          4236 => x"815381d3",
          4237 => x"ac08ff2e",
          4238 => x"80f93898",
          4239 => x"170881d3",
          4240 => x"ac082680",
          4241 => x"cc38778a",
          4242 => x"38779816",
          4243 => x"0c845380",
          4244 => x"e2399415",
          4245 => x"08527451",
          4246 => x"f8eb3f81",
          4247 => x"d3ac0854",
          4248 => x"875381d3",
          4249 => x"ac08802e",
          4250 => x"80c93882",
          4251 => x"5381d3ac",
          4252 => x"08812ebf",
          4253 => x"38815381",
          4254 => x"d3ac08ff",
          4255 => x"2eb53881",
          4256 => x"d3ac0852",
          4257 => x"7651fbe1",
          4258 => x"3f815381",
          4259 => x"d3ac08a3",
          4260 => x"38739416",
          4261 => x"0c735276",
          4262 => x"51f2893f",
          4263 => x"81d3ac08",
          4264 => x"98160c75",
          4265 => x"90160c75",
          4266 => x"83ff0617",
          4267 => x"b4059c16",
          4268 => x"0c805372",
          4269 => x"81d3ac0c",
          4270 => x"893d0d04",
          4271 => x"f83d0d7a",
          4272 => x"7c71085a",
          4273 => x"5a568052",
          4274 => x"7551fc93",
          4275 => x"3f81d3ac",
          4276 => x"085481d3",
          4277 => x"ac0880e1",
          4278 => x"3881d3ac",
          4279 => x"08579816",
          4280 => x"08527751",
          4281 => x"efc83f81",
          4282 => x"d3ac0854",
          4283 => x"81d3ac08",
          4284 => x"80c73881",
          4285 => x"d3ac089c",
          4286 => x"17087033",
          4287 => x"51545572",
          4288 => x"81e52e09",
          4289 => x"81068338",
          4290 => x"81557230",
          4291 => x"70802576",
          4292 => x"07515372",
          4293 => x"802e8b38",
          4294 => x"81175776",
          4295 => x"792e9a38",
          4296 => x"83398057",
          4297 => x"81527551",
          4298 => x"fd8a3f81",
          4299 => x"d3ac0854",
          4300 => x"81d3ac08",
          4301 => x"802effa6",
          4302 => x"3873842e",
          4303 => x"09810683",
          4304 => x"38875473",
          4305 => x"81d3ac0c",
          4306 => x"8a3d0d04",
          4307 => x"fd3d0d76",
          4308 => x"9a115254",
          4309 => x"ebaa3f81",
          4310 => x"d3ac0883",
          4311 => x"ffff0676",
          4312 => x"70335153",
          4313 => x"5371832e",
          4314 => x"09810690",
          4315 => x"38941451",
          4316 => x"eb8e3f81",
          4317 => x"d3ac0890",
          4318 => x"2b730753",
          4319 => x"7281d3ac",
          4320 => x"0c853d0d",
          4321 => x"04fc3d0d",
          4322 => x"77797083",
          4323 => x"ffff0654",
          4324 => x"9a125355",
          4325 => x"55ebab3f",
          4326 => x"76703351",
          4327 => x"5372832e",
          4328 => x"0981068b",
          4329 => x"3873902a",
          4330 => x"52941551",
          4331 => x"eb943f86",
          4332 => x"3d0d04f7",
          4333 => x"3d0d7b7d",
          4334 => x"5b568476",
          4335 => x"085a5898",
          4336 => x"1608802e",
          4337 => x"81863898",
          4338 => x"16085278",
          4339 => x"51eddf3f",
          4340 => x"81d3ac08",
          4341 => x"5881d3ac",
          4342 => x"0880f138",
          4343 => x"9c160870",
          4344 => x"33565374",
          4345 => x"86388458",
          4346 => x"80e2399c",
          4347 => x"16088b11",
          4348 => x"3370bf06",
          4349 => x"7081ff06",
          4350 => x"5a515153",
          4351 => x"72861734",
          4352 => x"7481e532",
          4353 => x"703076ae",
          4354 => x"32703070",
          4355 => x"73069f2a",
          4356 => x"53515551",
          4357 => x"5473802e",
          4358 => x"9b38768f",
          4359 => x"2e963880",
          4360 => x"77df0654",
          4361 => x"5472882e",
          4362 => x"09810683",
          4363 => x"38815473",
          4364 => x"7a2e9938",
          4365 => x"80527551",
          4366 => x"fafa3f81",
          4367 => x"d3ac0858",
          4368 => x"81d3ac08",
          4369 => x"87389816",
          4370 => x"08fefc38",
          4371 => x"77802e86",
          4372 => x"38800b98",
          4373 => x"170c7781",
          4374 => x"d3ac0c8b",
          4375 => x"3d0d04f8",
          4376 => x"3d0d7a70",
          4377 => x"08595680",
          4378 => x"527551f8",
          4379 => x"f23f81d3",
          4380 => x"ac085481",
          4381 => x"d3ac0880",
          4382 => x"ef388639",
          4383 => x"845780e6",
          4384 => x"39981608",
          4385 => x"527751ec",
          4386 => x"a53f81d3",
          4387 => x"ac085781",
          4388 => x"d3ac0880",
          4389 => x"d1389c16",
          4390 => x"08703351",
          4391 => x"5473802e",
          4392 => x"db389c16",
          4393 => x"088b1133",
          4394 => x"bf065555",
          4395 => x"73861734",
          4396 => x"8b153370",
          4397 => x"832a7081",
          4398 => x"06515559",
          4399 => x"7393388b",
          4400 => x"53a01652",
          4401 => x"7451ea85",
          4402 => x"3f81d3ac",
          4403 => x"08802e96",
          4404 => x"38805275",
          4405 => x"51f9dd3f",
          4406 => x"81d3ac08",
          4407 => x"5781d3ac",
          4408 => x"08802eff",
          4409 => x"9c387654",
          4410 => x"7381d3ac",
          4411 => x"0c8a3d0d",
          4412 => x"04fb3d0d",
          4413 => x"77700857",
          4414 => x"54815273",
          4415 => x"51fbbd3f",
          4416 => x"81d3ac08",
          4417 => x"5581d3ac",
          4418 => x"08b43898",
          4419 => x"14085275",
          4420 => x"51eb9b3f",
          4421 => x"81d3ac08",
          4422 => x"5581d3ac",
          4423 => x"08a038a0",
          4424 => x"5381d3ac",
          4425 => x"08529c14",
          4426 => x"0851e987",
          4427 => x"3f8b53a0",
          4428 => x"14529c14",
          4429 => x"0851e8d7",
          4430 => x"3f810b83",
          4431 => x"17347481",
          4432 => x"d3ac0c87",
          4433 => x"3d0d04fc",
          4434 => x"3d0d7670",
          4435 => x"08981208",
          4436 => x"54705356",
          4437 => x"53ead73f",
          4438 => x"81d3ac08",
          4439 => x"5481d3ac",
          4440 => x"088d389c",
          4441 => x"130853e5",
          4442 => x"7334810b",
          4443 => x"83163473",
          4444 => x"81d3ac0c",
          4445 => x"863d0d04",
          4446 => x"fa3d0d78",
          4447 => x"7a575780",
          4448 => x"0b891734",
          4449 => x"98170880",
          4450 => x"2e818938",
          4451 => x"80705555",
          4452 => x"9c170814",
          4453 => x"70338116",
          4454 => x"56545272",
          4455 => x"a02ead38",
          4456 => x"72852e09",
          4457 => x"81068438",
          4458 => x"81e55373",
          4459 => x"892e0981",
          4460 => x"068e3875",
          4461 => x"15880552",
          4462 => x"ae0b8113",
          4463 => x"34811555",
          4464 => x"75158805",
          4465 => x"52728113",
          4466 => x"34811555",
          4467 => x"8a7427c0",
          4468 => x"38751588",
          4469 => x"0552800b",
          4470 => x"8113349c",
          4471 => x"1708528b",
          4472 => x"12338817",
          4473 => x"349c1708",
          4474 => x"9c0551e6",
          4475 => x"ac3f81d3",
          4476 => x"ac08760c",
          4477 => x"9c170896",
          4478 => x"0551e684",
          4479 => x"3f81d3ac",
          4480 => x"08861723",
          4481 => x"9c170898",
          4482 => x"0551e5f4",
          4483 => x"3f81d3ac",
          4484 => x"08841723",
          4485 => x"883d0d04",
          4486 => x"f53d0d7e",
          4487 => x"70087fa0",
          4488 => x"055d5a5c",
          4489 => x"8b53a052",
          4490 => x"7a51e787",
          4491 => x"3f807058",
          4492 => x"58887933",
          4493 => x"555a73ae",
          4494 => x"2e098106",
          4495 => x"80df3878",
          4496 => x"17703381",
          4497 => x"1971ae32",
          4498 => x"7030709f",
          4499 => x"2a738226",
          4500 => x"07515153",
          4501 => x"59575473",
          4502 => x"8c387a18",
          4503 => x"54757434",
          4504 => x"811858db",
          4505 => x"3975af32",
          4506 => x"70307780",
          4507 => x"dc327030",
          4508 => x"7073069f",
          4509 => x"2a535156",
          4510 => x"51557480",
          4511 => x"2e893886",
          4512 => x"5475a026",
          4513 => x"82e43876",
          4514 => x"197c0ca4",
          4515 => x"54a07627",
          4516 => x"8338a054",
          4517 => x"738b1c34",
          4518 => x"805482ce",
          4519 => x"39781770",
          4520 => x"33811959",
          4521 => x"5754a076",
          4522 => x"27828c38",
          4523 => x"75af3270",
          4524 => x"307780dc",
          4525 => x"32703072",
          4526 => x"80257180",
          4527 => x"25075351",
          4528 => x"56515574",
          4529 => x"802eb538",
          4530 => x"84398117",
          4531 => x"5780771a",
          4532 => x"70335155",
          4533 => x"5a73af2e",
          4534 => x"09810683",
          4535 => x"38815a80",
          4536 => x"771a7033",
          4537 => x"51555573",
          4538 => x"80dc2e09",
          4539 => x"81068338",
          4540 => x"81557975",
          4541 => x"075473d2",
          4542 => x"3881bc39",
          4543 => x"75ae3270",
          4544 => x"30708025",
          4545 => x"7a7d2707",
          4546 => x"51515473",
          4547 => x"802ea238",
          4548 => x"798b3270",
          4549 => x"3077ae32",
          4550 => x"70307280",
          4551 => x"25719f2a",
          4552 => x"07535156",
          4553 => x"51557481",
          4554 => x"b1388858",
          4555 => x"8b5afeed",
          4556 => x"3975982b",
          4557 => x"54738025",
          4558 => x"8c387580",
          4559 => x"ff0681bb",
          4560 => x"dc113357",
          4561 => x"547551e5",
          4562 => x"e63f81d3",
          4563 => x"ac08802e",
          4564 => x"b9387817",
          4565 => x"70338119",
          4566 => x"71545956",
          4567 => x"54e5d73f",
          4568 => x"81d3ac08",
          4569 => x"802e8938",
          4570 => x"ff1a5473",
          4571 => x"78268638",
          4572 => x"865480f6",
          4573 => x"397a1854",
          4574 => x"75743481",
          4575 => x"187b1155",
          4576 => x"58747434",
          4577 => x"811858fe",
          4578 => x"94397552",
          4579 => x"81bad451",
          4580 => x"e4ec3f81",
          4581 => x"d3ac0880",
          4582 => x"c538ff9f",
          4583 => x"16547399",
          4584 => x"268938e0",
          4585 => x"167081ff",
          4586 => x"0657547a",
          4587 => x"18547574",
          4588 => x"34811858",
          4589 => x"fde73976",
          4590 => x"197c0c86",
          4591 => x"5477802e",
          4592 => x"a9387a33",
          4593 => x"547381e5",
          4594 => x"2e098106",
          4595 => x"8438857b",
          4596 => x"348454a0",
          4597 => x"76278d38",
          4598 => x"89398654",
          4599 => x"8d398654",
          4600 => x"89398054",
          4601 => x"738b1c34",
          4602 => x"80547381",
          4603 => x"d3ac0c8d",
          4604 => x"3d0d04fa",
          4605 => x"3d0d7870",
          4606 => x"08585680",
          4607 => x"7a703351",
          4608 => x"545572af",
          4609 => x"2e833881",
          4610 => x"55807a70",
          4611 => x"33515454",
          4612 => x"7280dc2e",
          4613 => x"83388154",
          4614 => x"74740653",
          4615 => x"72802e8c",
          4616 => x"38941708",
          4617 => x"88170cb3",
          4618 => x"39811a5a",
          4619 => x"807a7033",
          4620 => x"51545572",
          4621 => x"af2e0981",
          4622 => x"06833881",
          4623 => x"55807a70",
          4624 => x"33515454",
          4625 => x"7280dc2e",
          4626 => x"09810683",
          4627 => x"38815474",
          4628 => x"74075372",
          4629 => x"d438800b",
          4630 => x"88170c79",
          4631 => x"70335153",
          4632 => x"729f269b",
          4633 => x"38ff800b",
          4634 => x"ab173480",
          4635 => x"527551f0",
          4636 => x"ee3f81d3",
          4637 => x"ac085581",
          4638 => x"aa398555",
          4639 => x"81a53989",
          4640 => x"3d840552",
          4641 => x"7551fb90",
          4642 => x"3f81d3ac",
          4643 => x"085581d3",
          4644 => x"ac08818f",
          4645 => x"387551f7",
          4646 => x"c63f81d3",
          4647 => x"ac08ab17",
          4648 => x"33555581",
          4649 => x"d3ac0880",
          4650 => x"2e80c238",
          4651 => x"81d3ac08",
          4652 => x"842e0981",
          4653 => x"0680ec38",
          4654 => x"73852a70",
          4655 => x"81065153",
          4656 => x"72802e9a",
          4657 => x"3873822a",
          4658 => x"70810651",
          4659 => x"5372802e",
          4660 => x"ffad38ff",
          4661 => x"800bab17",
          4662 => x"34805580",
          4663 => x"c6397382",
          4664 => x"2a708106",
          4665 => x"515372bb",
          4666 => x"388555b7",
          4667 => x"3973822a",
          4668 => x"70810651",
          4669 => x"5372ac38",
          4670 => x"86163370",
          4671 => x"842a7081",
          4672 => x"06515454",
          4673 => x"72802efe",
          4674 => x"f1389016",
          4675 => x"0883ff06",
          4676 => x"17b40552",
          4677 => x"7651f4b4",
          4678 => x"3f81d3ac",
          4679 => x"0888170c",
          4680 => x"fedd3974",
          4681 => x"81d3ac0c",
          4682 => x"883d0d04",
          4683 => x"f63d0d7c",
          4684 => x"59ff7908",
          4685 => x"70725459",
          4686 => x"565a7480",
          4687 => x"2e81d038",
          4688 => x"76708105",
          4689 => x"583370ba",
          4690 => x"32703072",
          4691 => x"a026719f",
          4692 => x"2a065151",
          4693 => x"525370e8",
          4694 => x"3872ba2e",
          4695 => x"09810681",
          4696 => x"a9387433",
          4697 => x"d0115252",
          4698 => x"70892692",
          4699 => x"38821572",
          4700 => x"81ff06d0",
          4701 => x"11515951",
          4702 => x"70772e80",
          4703 => x"ff38800b",
          4704 => x"81bbcc5c",
          4705 => x"58771010",
          4706 => x"1b70087a",
          4707 => x"08575751",
          4708 => x"75708105",
          4709 => x"57337570",
          4710 => x"81055733",
          4711 => x"ff9f1253",
          4712 => x"54547099",
          4713 => x"268938e0",
          4714 => x"147081ff",
          4715 => x"065551ff",
          4716 => x"9f135170",
          4717 => x"99268938",
          4718 => x"e0137081",
          4719 => x"ff065451",
          4720 => x"73307474",
          4721 => x"32703070",
          4722 => x"72078025",
          4723 => x"739f2a06",
          4724 => x"53555351",
          4725 => x"70ffb938",
          4726 => x"73307578",
          4727 => x"32703070",
          4728 => x"72079f2a",
          4729 => x"739f2a07",
          4730 => x"53555351",
          4731 => x"70802e8c",
          4732 => x"38811858",
          4733 => x"837825ff",
          4734 => x"8c388b39",
          4735 => x"77832486",
          4736 => x"3877777a",
          4737 => x"0c5a7951",
          4738 => x"863981d3",
          4739 => x"dc335170",
          4740 => x"81d3ac0c",
          4741 => x"8c3d0d04",
          4742 => x"fb3d0d77",
          4743 => x"56800b83",
          4744 => x"1734ff0b",
          4745 => x"b0170c78",
          4746 => x"527551e1",
          4747 => x"813f8455",
          4748 => x"81d3ac08",
          4749 => x"81843884",
          4750 => x"b21651dd",
          4751 => x"c33f81d3",
          4752 => x"ac0883ff",
          4753 => x"ff065483",
          4754 => x"557382d4",
          4755 => x"d52e0981",
          4756 => x"0680e738",
          4757 => x"800bb417",
          4758 => x"33555573",
          4759 => x"81e92e09",
          4760 => x"81068338",
          4761 => x"81557381",
          4762 => x"eb327030",
          4763 => x"70802577",
          4764 => x"07515154",
          4765 => x"738e38b4",
          4766 => x"16335473",
          4767 => x"81e82e09",
          4768 => x"8106b538",
          4769 => x"835381ba",
          4770 => x"e45280ea",
          4771 => x"1651debd",
          4772 => x"3f81d3ac",
          4773 => x"085581d3",
          4774 => x"ac08802e",
          4775 => x"9d388553",
          4776 => x"81bae852",
          4777 => x"81861651",
          4778 => x"dea33f81",
          4779 => x"d3ac0855",
          4780 => x"81d3ac08",
          4781 => x"802e8338",
          4782 => x"82557481",
          4783 => x"d3ac0c87",
          4784 => x"3d0d04f3",
          4785 => x"3d0d6002",
          4786 => x"840580c7",
          4787 => x"05335854",
          4788 => x"80740c7f",
          4789 => x"51fcd53f",
          4790 => x"81d3ac08",
          4791 => x"588b5680",
          4792 => x"0b81d3ac",
          4793 => x"0824879e",
          4794 => x"3881d3ac",
          4795 => x"08101081",
          4796 => x"d3c80570",
          4797 => x"0856538c",
          4798 => x"5674802e",
          4799 => x"87883874",
          4800 => x"740c7681",
          4801 => x"fe067533",
          4802 => x"54577280",
          4803 => x"2eaf3881",
          4804 => x"153351d6",
          4805 => x"a63f81d3",
          4806 => x"ac0881ff",
          4807 => x"06708106",
          4808 => x"54547299",
          4809 => x"3876802e",
          4810 => x"8f387382",
          4811 => x"2a708106",
          4812 => x"51538a56",
          4813 => x"7286cf38",
          4814 => x"805686ca",
          4815 => x"39807534",
          4816 => x"77811634",
          4817 => x"81528115",
          4818 => x"3351d68d",
          4819 => x"3f81d3ac",
          4820 => x"0881ff06",
          4821 => x"70810654",
          4822 => x"54835672",
          4823 => x"86a83876",
          4824 => x"802e8f38",
          4825 => x"73822a70",
          4826 => x"81065153",
          4827 => x"8a567286",
          4828 => x"95388070",
          4829 => x"5375525a",
          4830 => x"fd9e3f81",
          4831 => x"d3ac0881",
          4832 => x"ff065776",
          4833 => x"822e0981",
          4834 => x"0680e438",
          4835 => x"79547390",
          4836 => x"2915903d",
          4837 => x"75101005",
          4838 => x"f00583f6",
          4839 => x"12335559",
          4840 => x"56805772",
          4841 => x"772e8d38",
          4842 => x"83fa1651",
          4843 => x"daeb3f81",
          4844 => x"d3ac0857",
          4845 => x"76780c81",
          4846 => x"14548374",
          4847 => x"27d03880",
          4848 => x"548f3d74",
          4849 => x"101005f0",
          4850 => x"11085b53",
          4851 => x"83577980",
          4852 => x"2e903879",
          4853 => x"527451fc",
          4854 => x"bf3f81d3",
          4855 => x"ac0881ff",
          4856 => x"06578177",
          4857 => x"27893881",
          4858 => x"14548374",
          4859 => x"27d33881",
          4860 => x"5676842e",
          4861 => x"8590388d",
          4862 => x"56768126",
          4863 => x"858838bf",
          4864 => x"1551d9fc",
          4865 => x"3f81d3ac",
          4866 => x"0883ffff",
          4867 => x"06538d56",
          4868 => x"7284802e",
          4869 => x"09810684",
          4870 => x"ed3880ca",
          4871 => x"1551d9e0",
          4872 => x"3f81d3ac",
          4873 => x"0883ffff",
          4874 => x"0654738d",
          4875 => x"3880d815",
          4876 => x"51d9e63f",
          4877 => x"81d3ac08",
          4878 => x"54739c16",
          4879 => x"0c80c415",
          4880 => x"33821634",
          4881 => x"80c41533",
          4882 => x"ff05538d",
          4883 => x"56728126",
          4884 => x"84b43882",
          4885 => x"15337471",
          4886 => x"2980c117",
          4887 => x"33525553",
          4888 => x"728a1623",
          4889 => x"7283ffff",
          4890 => x"06537280",
          4891 => x"2e8b38ff",
          4892 => x"13730653",
          4893 => x"72802e86",
          4894 => x"388d5684",
          4895 => x"893980c5",
          4896 => x"1551d8fc",
          4897 => x"3f81d3ac",
          4898 => x"08881623",
          4899 => x"81d3ac08",
          4900 => x"83ffff06",
          4901 => x"8f06538d",
          4902 => x"567283ea",
          4903 => x"3880c715",
          4904 => x"51d8dd3f",
          4905 => x"81d3ac08",
          4906 => x"83ffff06",
          4907 => x"53728d38",
          4908 => x"80d41551",
          4909 => x"d8e33f81",
          4910 => x"d3ac0853",
          4911 => x"80c21551",
          4912 => x"d8be3f81",
          4913 => x"d3ac0883",
          4914 => x"ffff0659",
          4915 => x"8d567880",
          4916 => x"2e83b338",
          4917 => x"88152274",
          4918 => x"1a71842a",
          4919 => x"0559568d",
          4920 => x"56777326",
          4921 => x"83a0388a",
          4922 => x"15225272",
          4923 => x"783151ff",
          4924 => x"b0ab3f81",
          4925 => x"d3ac0853",
          4926 => x"8d5681d3",
          4927 => x"ac08802e",
          4928 => x"83843880",
          4929 => x"5781d3ac",
          4930 => x"0880ffff",
          4931 => x"fff52683",
          4932 => x"38835772",
          4933 => x"83fff526",
          4934 => x"83388257",
          4935 => x"729ff526",
          4936 => x"83388157",
          4937 => x"8d567680",
          4938 => x"2e82db38",
          4939 => x"82139816",
          4940 => x"0c79a016",
          4941 => x"0c7919a4",
          4942 => x"160c771a",
          4943 => x"ac160c76",
          4944 => x"832e0981",
          4945 => x"06b73880",
          4946 => x"de1551d7",
          4947 => x"b33f81d3",
          4948 => x"ac0883ff",
          4949 => x"ff06538d",
          4950 => x"567282aa",
          4951 => x"38881522",
          4952 => x"538d5672",
          4953 => x"82a03880",
          4954 => x"e01551d7",
          4955 => x"ac3f81d3",
          4956 => x"ac08a816",
          4957 => x"0c981508",
          4958 => x"822b53b6",
          4959 => x"39881522",
          4960 => x"538d5672",
          4961 => x"802e81fe",
          4962 => x"38a41508",
          4963 => x"14a8160c",
          4964 => x"76822e09",
          4965 => x"81068838",
          4966 => x"98150810",
          4967 => x"53943998",
          4968 => x"15081098",
          4969 => x"16080570",
          4970 => x"812a9817",
          4971 => x"08810605",
          4972 => x"515383ff",
          4973 => x"13892a53",
          4974 => x"8d56729c",
          4975 => x"16082681",
          4976 => x"c538ff0b",
          4977 => x"90160cff",
          4978 => x"0b8c160c",
          4979 => x"ff800b84",
          4980 => x"16347683",
          4981 => x"2e098106",
          4982 => x"81923880",
          4983 => x"e41551d6",
          4984 => x"9f3f81d3",
          4985 => x"ac0883ff",
          4986 => x"ff065372",
          4987 => x"812e0981",
          4988 => x"0680f938",
          4989 => x"811a5274",
          4990 => x"51d9b33f",
          4991 => x"81d3ac08",
          4992 => x"80ea3881",
          4993 => x"d3ac0884",
          4994 => x"163484b2",
          4995 => x"1551d5f0",
          4996 => x"3f81d3ac",
          4997 => x"0883ffff",
          4998 => x"06537282",
          4999 => x"d4d52e09",
          5000 => x"810680c8",
          5001 => x"38b41551",
          5002 => x"d5ef3f81",
          5003 => x"d3ac0884",
          5004 => x"8b85a4d2",
          5005 => x"2e098106",
          5006 => x"b3388498",
          5007 => x"1551d5d9",
          5008 => x"3f81d3ac",
          5009 => x"08868a85",
          5010 => x"e4f22e09",
          5011 => x"81069d38",
          5012 => x"849c1551",
          5013 => x"d5c33f81",
          5014 => x"d3ac0890",
          5015 => x"160c84a0",
          5016 => x"1551d5b5",
          5017 => x"3f81d3ac",
          5018 => x"088c160c",
          5019 => x"76753481",
          5020 => x"d3d82281",
          5021 => x"05537281",
          5022 => x"d3d82372",
          5023 => x"86162380",
          5024 => x"0b94160c",
          5025 => x"80567581",
          5026 => x"d3ac0c8f",
          5027 => x"3d0d04fb",
          5028 => x"3d0d7754",
          5029 => x"89557380",
          5030 => x"2eb53873",
          5031 => x"08802eaf",
          5032 => x"38730870",
          5033 => x"33535371",
          5034 => x"802ea438",
          5035 => x"84142286",
          5036 => x"14225752",
          5037 => x"71762e09",
          5038 => x"81069438",
          5039 => x"81133351",
          5040 => x"cef93f81",
          5041 => x"d3ac0881",
          5042 => x"06527183",
          5043 => x"38715580",
          5044 => x"5374732e",
          5045 => x"09810684",
          5046 => x"38730853",
          5047 => x"7873710c",
          5048 => x"527481d3",
          5049 => x"ac0c873d",
          5050 => x"0d04fa3d",
          5051 => x"0d02ab05",
          5052 => x"337a5889",
          5053 => x"3dfc0552",
          5054 => x"56f4b13f",
          5055 => x"81d3ac08",
          5056 => x"558b5480",
          5057 => x"0b81d3ac",
          5058 => x"082480c4",
          5059 => x"3881d3ac",
          5060 => x"08101081",
          5061 => x"d3c80570",
          5062 => x"08515473",
          5063 => x"802e8438",
          5064 => x"80743478",
          5065 => x"802e8638",
          5066 => x"78548074",
          5067 => x"34741010",
          5068 => x"81d3c805",
          5069 => x"79710c54",
          5070 => x"75547580",
          5071 => x"2e923880",
          5072 => x"53893d70",
          5073 => x"53840551",
          5074 => x"f6f93f81",
          5075 => x"d3ac0854",
          5076 => x"7381d3ac",
          5077 => x"0c883d0d",
          5078 => x"04eb3d0d",
          5079 => x"67028405",
          5080 => x"80e70533",
          5081 => x"58588955",
          5082 => x"77802e84",
          5083 => x"e93876bf",
          5084 => x"06705498",
          5085 => x"3dd00553",
          5086 => x"993d8405",
          5087 => x"5257f6c3",
          5088 => x"3f81d3ac",
          5089 => x"085681d3",
          5090 => x"ac0884c5",
          5091 => x"387a5c68",
          5092 => x"52973dd4",
          5093 => x"0551f0db",
          5094 => x"3f81d3ac",
          5095 => x"085681d3",
          5096 => x"ac089238",
          5097 => x"0280d705",
          5098 => x"3370982b",
          5099 => x"56597480",
          5100 => x"25833886",
          5101 => x"56769c06",
          5102 => x"5574802e",
          5103 => x"81c33875",
          5104 => x"802e9c38",
          5105 => x"75842e09",
          5106 => x"81068e38",
          5107 => x"973dd405",
          5108 => x"51ea9e3f",
          5109 => x"81d3ac08",
          5110 => x"56768807",
          5111 => x"57a03902",
          5112 => x"b2053391",
          5113 => x"06557480",
          5114 => x"2e853887",
          5115 => x"56903976",
          5116 => x"822a7081",
          5117 => x"06515574",
          5118 => x"802e8338",
          5119 => x"88567583",
          5120 => x"d0387683",
          5121 => x"2a708106",
          5122 => x"51557480",
          5123 => x"2e81a738",
          5124 => x"62527a51",
          5125 => x"e6b63f81",
          5126 => x"d3ac0859",
          5127 => x"8288b20a",
          5128 => x"52628e05",
          5129 => x"51d2b93f",
          5130 => x"6255a00b",
          5131 => x"8b163475",
          5132 => x"5362527a",
          5133 => x"51e6ce3f",
          5134 => x"7552629c",
          5135 => x"0551d2a0",
          5136 => x"3f7a5581",
          5137 => x"0b831634",
          5138 => x"78802e80",
          5139 => x"e9387ab0",
          5140 => x"11087755",
          5141 => x"7a54993d",
          5142 => x"d4055351",
          5143 => x"55dbb33f",
          5144 => x"81d3ac08",
          5145 => x"5681d3ac",
          5146 => x"0882e638",
          5147 => x"74527a51",
          5148 => x"d4bc3f81",
          5149 => x"d3ac087b",
          5150 => x"ff1b8c12",
          5151 => x"0c5656b6",
          5152 => x"397582cd",
          5153 => x"3802b205",
          5154 => x"3370842a",
          5155 => x"70810651",
          5156 => x"56597480",
          5157 => x"2e853884",
          5158 => x"569c3976",
          5159 => x"812a7081",
          5160 => x"06515574",
          5161 => x"802e8f38",
          5162 => x"02b20533",
          5163 => x"81065574",
          5164 => x"802e8338",
          5165 => x"87567582",
          5166 => x"98387683",
          5167 => x"2a708106",
          5168 => x"51557480",
          5169 => x"2e863876",
          5170 => x"80c00757",
          5171 => x"7ab01108",
          5172 => x"a01a0c63",
          5173 => x"a41a0c55",
          5174 => x"7581f638",
          5175 => x"62527451",
          5176 => x"e4ea3f81",
          5177 => x"d3ac0888",
          5178 => x"190c629c",
          5179 => x"0551d0a9",
          5180 => x"3f81d3ac",
          5181 => x"088c190c",
          5182 => x"74780c86",
          5183 => x"15228419",
          5184 => x"23769019",
          5185 => x"34759119",
          5186 => x"34759c19",
          5187 => x"0c759419",
          5188 => x"0c848053",
          5189 => x"7552a818",
          5190 => x"51d1983f",
          5191 => x"76852a70",
          5192 => x"81065155",
          5193 => x"74802e81",
          5194 => x"a3388c18",
          5195 => x"08802e81",
          5196 => x"9b388c18",
          5197 => x"0894190c",
          5198 => x"7a8a1122",
          5199 => x"70892b88",
          5200 => x"1b088c1c",
          5201 => x"085d5a5c",
          5202 => x"5155a539",
          5203 => x"76527751",
          5204 => x"d4fc3f81",
          5205 => x"d3ac0857",
          5206 => x"81d3ac08",
          5207 => x"81268338",
          5208 => x"825676ff",
          5209 => x"2e098106",
          5210 => x"83388156",
          5211 => x"787a3159",
          5212 => x"75307077",
          5213 => x"07802570",
          5214 => x"7b7d2606",
          5215 => x"51515574",
          5216 => x"cb387698",
          5217 => x"190c7580",
          5218 => x"c8387883",
          5219 => x"ff065574",
          5220 => x"802eb938",
          5221 => x"76527a51",
          5222 => x"d48a3f81",
          5223 => x"d3ac0885",
          5224 => x"388256a8",
          5225 => x"3978892a",
          5226 => x"81d3ac08",
          5227 => x"05709c1a",
          5228 => x"0c558154",
          5229 => x"7453a818",
          5230 => x"527a8111",
          5231 => x"335255ca",
          5232 => x"a43f81d3",
          5233 => x"ac08802e",
          5234 => x"83388156",
          5235 => x"75802e84",
          5236 => x"3880780c",
          5237 => x"75557481",
          5238 => x"d3ac0c97",
          5239 => x"3d0d04f3",
          5240 => x"3d0d7f62",
          5241 => x"64635f5f",
          5242 => x"5a57807d",
          5243 => x"0c8f3dfc",
          5244 => x"05527651",
          5245 => x"f9993f81",
          5246 => x"d3ac0855",
          5247 => x"81d3ac08",
          5248 => x"8a389117",
          5249 => x"33557480",
          5250 => x"2e863874",
          5251 => x"5683ae39",
          5252 => x"90173381",
          5253 => x"06558756",
          5254 => x"74802e83",
          5255 => x"a038bd39",
          5256 => x"820b9118",
          5257 => x"34825683",
          5258 => x"9439810b",
          5259 => x"91183481",
          5260 => x"56838a39",
          5261 => x"820b9118",
          5262 => x"34825683",
          5263 => x"8039810b",
          5264 => x"91183481",
          5265 => x"5682f639",
          5266 => x"810b9118",
          5267 => x"34815682",
          5268 => x"ec39810b",
          5269 => x"91183481",
          5270 => x"5682e239",
          5271 => x"8c170894",
          5272 => x"18083155",
          5273 => x"74792783",
          5274 => x"38745978",
          5275 => x"802e82cb",
          5276 => x"38941708",
          5277 => x"7083ff06",
          5278 => x"56567482",
          5279 => x"83387d8a",
          5280 => x"1122ff05",
          5281 => x"77892a06",
          5282 => x"5c557aa8",
          5283 => x"38758738",
          5284 => x"88170855",
          5285 => x"8f399817",
          5286 => x"08527651",
          5287 => x"d2b03f81",
          5288 => x"d3ac0855",
          5289 => x"817527fe",
          5290 => x"f73874ff",
          5291 => x"2efefb38",
          5292 => x"7498180c",
          5293 => x"98170852",
          5294 => x"7d51d1e8",
          5295 => x"3f81d3ac",
          5296 => x"08802efe",
          5297 => x"ef3881d3",
          5298 => x"ac081b79",
          5299 => x"892a5b58",
          5300 => x"79802e80",
          5301 => x"d738791b",
          5302 => x"7e8a1122",
          5303 => x"51565674",
          5304 => x"76278538",
          5305 => x"747b315a",
          5306 => x"79547753",
          5307 => x"7b527d81",
          5308 => x"11335255",
          5309 => x"c7ef3f81",
          5310 => x"d3ac08fe",
          5311 => x"c1389017",
          5312 => x"3370982b",
          5313 => x"56567480",
          5314 => x"259b389c",
          5315 => x"17087831",
          5316 => x"55747a27",
          5317 => x"90388480",
          5318 => x"53a81752",
          5319 => x"74848029",
          5320 => x"1c51cceb",
          5321 => x"3f79892b",
          5322 => x"5680f939",
          5323 => x"9c170878",
          5324 => x"2e80c938",
          5325 => x"90173370",
          5326 => x"982b5656",
          5327 => x"748025a5",
          5328 => x"3881549c",
          5329 => x"170853a8",
          5330 => x"17527d81",
          5331 => x"11335255",
          5332 => x"c8ec3f81",
          5333 => x"d3ac08fd",
          5334 => x"ef389017",
          5335 => x"3380ff06",
          5336 => x"55749018",
          5337 => x"34815477",
          5338 => x"53a81752",
          5339 => x"7d811133",
          5340 => x"5255c6f1",
          5341 => x"3f81d3ac",
          5342 => x"08fdd738",
          5343 => x"779c180c",
          5344 => x"94170883",
          5345 => x"ff068480",
          5346 => x"71315755",
          5347 => x"78762783",
          5348 => x"38785675",
          5349 => x"53941708",
          5350 => x"83ff0617",
          5351 => x"a805527b",
          5352 => x"51cbec3f",
          5353 => x"7876317d",
          5354 => x"08177e0c",
          5355 => x"761d9419",
          5356 => x"0818941a",
          5357 => x"0c5d5978",
          5358 => x"fdb73880",
          5359 => x"567581d3",
          5360 => x"ac0c8f3d",
          5361 => x"0d04f33d",
          5362 => x"0d7f6264",
          5363 => x"635f5f5a",
          5364 => x"57807d0c",
          5365 => x"8f3dfc05",
          5366 => x"527651f5",
          5367 => x"b23f81d3",
          5368 => x"ac085581",
          5369 => x"d3ac088a",
          5370 => x"38911733",
          5371 => x"5574802e",
          5372 => x"86387456",
          5373 => x"84823990",
          5374 => x"17337081",
          5375 => x"2a708106",
          5376 => x"51565687",
          5377 => x"5674802e",
          5378 => x"83ee38bd",
          5379 => x"39820b91",
          5380 => x"18348256",
          5381 => x"83e23981",
          5382 => x"0b911834",
          5383 => x"815683d8",
          5384 => x"39810b91",
          5385 => x"18348156",
          5386 => x"83ce3982",
          5387 => x"0b911834",
          5388 => x"825683c4",
          5389 => x"39810b91",
          5390 => x"18348156",
          5391 => x"83ba3981",
          5392 => x"0b911834",
          5393 => x"815683b0",
          5394 => x"39941708",
          5395 => x"19557494",
          5396 => x"18082786",
          5397 => x"38941708",
          5398 => x"09597880",
          5399 => x"2e838c38",
          5400 => x"94170870",
          5401 => x"83ff0656",
          5402 => x"567482a8",
          5403 => x"387d8a11",
          5404 => x"22ff0577",
          5405 => x"892a065c",
          5406 => x"557a80c6",
          5407 => x"38759638",
          5408 => x"88170855",
          5409 => x"74a3387a",
          5410 => x"527651d4",
          5411 => x"b83f81d3",
          5412 => x"ac08558f",
          5413 => x"39981708",
          5414 => x"527651d4",
          5415 => x"a83f81d3",
          5416 => x"ac085574",
          5417 => x"802e82c3",
          5418 => x"3874812e",
          5419 => x"fedf3874",
          5420 => x"ff2efee3",
          5421 => x"38749818",
          5422 => x"0c881708",
          5423 => x"85387488",
          5424 => x"180c9017",
          5425 => x"3370982b",
          5426 => x"56587480",
          5427 => x"25a53881",
          5428 => x"549c1708",
          5429 => x"53a81752",
          5430 => x"7d811133",
          5431 => x"5255c5de",
          5432 => x"3f81d3ac",
          5433 => x"08feba38",
          5434 => x"90173380",
          5435 => x"ff065574",
          5436 => x"90183498",
          5437 => x"1708527d",
          5438 => x"51cda93f",
          5439 => x"81d3ac08",
          5440 => x"802efea7",
          5441 => x"3881d3ac",
          5442 => x"081b7989",
          5443 => x"2a5b5879",
          5444 => x"802e80d5",
          5445 => x"38791b7e",
          5446 => x"8a112251",
          5447 => x"56567476",
          5448 => x"27853874",
          5449 => x"7b315a79",
          5450 => x"5477537b",
          5451 => x"527d8111",
          5452 => x"335255c5",
          5453 => x"893f81d3",
          5454 => x"ac08fdf9",
          5455 => x"389c1708",
          5456 => x"78315574",
          5457 => x"7a279b38",
          5458 => x"84805374",
          5459 => x"8480291c",
          5460 => x"52a81751",
          5461 => x"c8b93f90",
          5462 => x"173380ff",
          5463 => x"06557490",
          5464 => x"18347989",
          5465 => x"2b5680db",
          5466 => x"399c1708",
          5467 => x"782ea138",
          5468 => x"9417088c",
          5469 => x"18082798",
          5470 => x"38815477",
          5471 => x"53a81752",
          5472 => x"7d811133",
          5473 => x"5255c2dd",
          5474 => x"3f81d3ac",
          5475 => x"08fdb038",
          5476 => x"779c180c",
          5477 => x"94170883",
          5478 => x"ff068480",
          5479 => x"71315755",
          5480 => x"78762783",
          5481 => x"38785675",
          5482 => x"537b5294",
          5483 => x"170883ff",
          5484 => x"0617a805",
          5485 => x"51c7d83f",
          5486 => x"901733ff",
          5487 => x"80075574",
          5488 => x"90183478",
          5489 => x"76317d08",
          5490 => x"177e0c76",
          5491 => x"1d941908",
          5492 => x"1870941b",
          5493 => x"0c8c1a08",
          5494 => x"58585d59",
          5495 => x"74762783",
          5496 => x"38755574",
          5497 => x"8c180c78",
          5498 => x"fcf63890",
          5499 => x"173380c0",
          5500 => x"07557490",
          5501 => x"18348056",
          5502 => x"7581d3ac",
          5503 => x"0c8f3d0d",
          5504 => x"04f73d0d",
          5505 => x"7b8c3dfc",
          5506 => x"05537052",
          5507 => x"58f1803f",
          5508 => x"81d3ac08",
          5509 => x"5781d3ac",
          5510 => x"0881aa38",
          5511 => x"90183370",
          5512 => x"862a7081",
          5513 => x"06515656",
          5514 => x"74802e81",
          5515 => x"98387598",
          5516 => x"2b557480",
          5517 => x"25a73881",
          5518 => x"549c1808",
          5519 => x"53a81852",
          5520 => x"79811133",
          5521 => x"5255c2f6",
          5522 => x"3f815581",
          5523 => x"d3ac0880",
          5524 => x"f6389018",
          5525 => x"3380ff06",
          5526 => x"55749019",
          5527 => x"34a01808",
          5528 => x"527951c8",
          5529 => x"c93f81d3",
          5530 => x"ac085781",
          5531 => x"d3ac0880",
          5532 => x"d438a418",
          5533 => x"088b1133",
          5534 => x"a0075656",
          5535 => x"748b1734",
          5536 => x"88180853",
          5537 => x"75527708",
          5538 => x"51d9fa3f",
          5539 => x"8c180852",
          5540 => x"9c1651c5",
          5541 => x"cb3f8288",
          5542 => x"b20a5296",
          5543 => x"1651c5c0",
          5544 => x"3f765292",
          5545 => x"1651c59a",
          5546 => x"3f795581",
          5547 => x"0b831634",
          5548 => x"7951c8c1",
          5549 => x"3f81d3ac",
          5550 => x"08901933",
          5551 => x"81bf0656",
          5552 => x"57749019",
          5553 => x"34765574",
          5554 => x"81d3ac0c",
          5555 => x"8b3d0d04",
          5556 => x"fc3d0d76",
          5557 => x"705254fe",
          5558 => x"a83f81d3",
          5559 => x"ac085381",
          5560 => x"d3ac089c",
          5561 => x"38863dfc",
          5562 => x"05527351",
          5563 => x"efa13f81",
          5564 => x"d3ac0853",
          5565 => x"81d3ac08",
          5566 => x"873881d3",
          5567 => x"ac08740c",
          5568 => x"7281d3ac",
          5569 => x"0c863d0d",
          5570 => x"04fe3d0d",
          5571 => x"853d51e4",
          5572 => x"9b3f8b53",
          5573 => x"800b81d3",
          5574 => x"ac08248b",
          5575 => x"3881d3ac",
          5576 => x"0881d3dc",
          5577 => x"34805372",
          5578 => x"81d3ac0c",
          5579 => x"843d0d04",
          5580 => x"ef3d0d80",
          5581 => x"53933dd0",
          5582 => x"0552943d",
          5583 => x"51e7843f",
          5584 => x"81d3ac08",
          5585 => x"5581d3ac",
          5586 => x"0880df38",
          5587 => x"76586352",
          5588 => x"933dd405",
          5589 => x"51e19c3f",
          5590 => x"81d3ac08",
          5591 => x"5581d3ac",
          5592 => x"08be3802",
          5593 => x"80c70533",
          5594 => x"70982b55",
          5595 => x"56738025",
          5596 => x"8938767a",
          5597 => x"94120c54",
          5598 => x"a73902a2",
          5599 => x"05337084",
          5600 => x"2a708106",
          5601 => x"51555673",
          5602 => x"802e9338",
          5603 => x"767f5370",
          5604 => x"5254d7b8",
          5605 => x"3f81d3ac",
          5606 => x"0894150c",
          5607 => x"83398555",
          5608 => x"74842e09",
          5609 => x"81068338",
          5610 => x"85557481",
          5611 => x"d3ac0c93",
          5612 => x"3d0d04e1",
          5613 => x"3d0da33d",
          5614 => x"08a33d08",
          5615 => x"5b5c807a",
          5616 => x"348053a1",
          5617 => x"3dffb805",
          5618 => x"52a23d51",
          5619 => x"e5f53f81",
          5620 => x"d3ac0857",
          5621 => x"81d3ac08",
          5622 => x"8393387e",
          5623 => x"467b7f94",
          5624 => x"11084a55",
          5625 => x"68565974",
          5626 => x"802e81f9",
          5627 => x"38963d70",
          5628 => x"943d405e",
          5629 => x"5ba0527a",
          5630 => x"51d1e43f",
          5631 => x"81d3ac08",
          5632 => x"5781d3ac",
          5633 => x"0881de38",
          5634 => x"6b527e51",
          5635 => x"c5a03f81",
          5636 => x"d3ac0857",
          5637 => x"81d3ac08",
          5638 => x"81cb386c",
          5639 => x"527e51d6",
          5640 => x"ab3f81d3",
          5641 => x"ac084876",
          5642 => x"527a51d1",
          5643 => x"b23f81d3",
          5644 => x"ac085781",
          5645 => x"d3ac0881",
          5646 => x"ac387c54",
          5647 => x"80527351",
          5648 => x"d6f13f81",
          5649 => x"d3ac0857",
          5650 => x"81d3ac08",
          5651 => x"a4386c52",
          5652 => x"7e51d5f8",
          5653 => x"3f81d3ac",
          5654 => x"08752e95",
          5655 => x"38765273",
          5656 => x"51d2d13f",
          5657 => x"81d3ac08",
          5658 => x"5781d3ac",
          5659 => x"08802ecc",
          5660 => x"3876842e",
          5661 => x"09810683",
          5662 => x"38825776",
          5663 => x"81ef38a1",
          5664 => x"3dffbc11",
          5665 => x"53d40551",
          5666 => x"d9ee3f76",
          5667 => x"933d7079",
          5668 => x"12811133",
          5669 => x"51525755",
          5670 => x"5673802e",
          5671 => x"8e388116",
          5672 => x"70168111",
          5673 => x"33515556",
          5674 => x"73f43881",
          5675 => x"16547874",
          5676 => x"27853891",
          5677 => x"57af3975",
          5678 => x"802e9938",
          5679 => x"7d58ff19",
          5680 => x"a33d0811",
          5681 => x"ff18701b",
          5682 => x"57585659",
          5683 => x"81143375",
          5684 => x"3475eb38",
          5685 => x"ff19a33d",
          5686 => x"08115559",
          5687 => x"af743467",
          5688 => x"5574fe91",
          5689 => x"38768185",
          5690 => x"38787c2e",
          5691 => x"0981068c",
          5692 => x"38ff19a3",
          5693 => x"3d081155",
          5694 => x"59af7434",
          5695 => x"807081d3",
          5696 => x"dc337010",
          5697 => x"1081bbcc",
          5698 => x"05700870",
          5699 => x"33525257",
          5700 => x"57575873",
          5701 => x"782e8d38",
          5702 => x"81167016",
          5703 => x"70335155",
          5704 => x"5673f538",
          5705 => x"82165473",
          5706 => x"7926a538",
          5707 => x"80587776",
          5708 => x"27943877",
          5709 => x"15547333",
          5710 => x"7a708105",
          5711 => x"5c348118",
          5712 => x"58757826",
          5713 => x"ee38ba7a",
          5714 => x"7081055c",
          5715 => x"34811858",
          5716 => x"77833891",
          5717 => x"57769638",
          5718 => x"a23d0819",
          5719 => x"811a5a54",
          5720 => x"73337a70",
          5721 => x"81055c34",
          5722 => x"7b7926ec",
          5723 => x"38807a34",
          5724 => x"7681d3ac",
          5725 => x"0ca13d0d",
          5726 => x"04f43d0d",
          5727 => x"7e60903d",
          5728 => x"fc055471",
          5729 => x"535957ea",
          5730 => x"863f81d3",
          5731 => x"ac085a81",
          5732 => x"d3ac088a",
          5733 => x"38911733",
          5734 => x"5a79802e",
          5735 => x"86387955",
          5736 => x"83f9398c",
          5737 => x"17087827",
          5738 => x"94389017",
          5739 => x"3370812a",
          5740 => x"70810651",
          5741 => x"56567485",
          5742 => x"388c1708",
          5743 => x"58941708",
          5744 => x"56807094",
          5745 => x"190c5b77",
          5746 => x"7b2e82b3",
          5747 => x"387c8a11",
          5748 => x"2270892b",
          5749 => x"5b515575",
          5750 => x"7b2eb638",
          5751 => x"7852ff18",
          5752 => x"51ff96b9",
          5753 => x"3f81d3ac",
          5754 => x"08ff177a",
          5755 => x"54705357",
          5756 => x"55ff96a9",
          5757 => x"3f81d3ac",
          5758 => x"08752695",
          5759 => x"38783076",
          5760 => x"0694180c",
          5761 => x"77941808",
          5762 => x"31981808",
          5763 => x"575880c9",
          5764 => x"39881708",
          5765 => x"5675be38",
          5766 => x"75527651",
          5767 => x"c9a73f81",
          5768 => x"d3ac0856",
          5769 => x"81d3ac08",
          5770 => x"812e0981",
          5771 => x"068b3882",
          5772 => x"0b911834",
          5773 => x"825582e3",
          5774 => x"3981d3ac",
          5775 => x"08ff2e09",
          5776 => x"81068b38",
          5777 => x"810b9118",
          5778 => x"34815582",
          5779 => x"ce3981d3",
          5780 => x"ac088818",
          5781 => x"0c759818",
          5782 => x"0c75802e",
          5783 => x"81a13878",
          5784 => x"782780ea",
          5785 => x"38777931",
          5786 => x"9418081a",
          5787 => x"94190c90",
          5788 => x"18337081",
          5789 => x"2a708106",
          5790 => x"51575d58",
          5791 => x"74802e9a",
          5792 => x"38755276",
          5793 => x"51c8be3f",
          5794 => x"81d3ac08",
          5795 => x"5681d3ac",
          5796 => x"08943881",
          5797 => x"d3ac0858",
          5798 => x"b5397552",
          5799 => x"7651c2ae",
          5800 => x"3f81d3ac",
          5801 => x"085675ff",
          5802 => x"2e81e138",
          5803 => x"8176278a",
          5804 => x"387c5598",
          5805 => x"15087626",
          5806 => x"8b38820b",
          5807 => x"91183482",
          5808 => x"5581d839",
          5809 => x"7598180c",
          5810 => x"777926ff",
          5811 => x"98389417",
          5812 => x"08189418",
          5813 => x"0c7783ff",
          5814 => x"06557480",
          5815 => x"2ea13875",
          5816 => x"527c51c1",
          5817 => x"bf3f81d3",
          5818 => x"ac088b38",
          5819 => x"820b9118",
          5820 => x"34825581",
          5821 => x"a6397789",
          5822 => x"2a81d3ac",
          5823 => x"08055b8c",
          5824 => x"17089418",
          5825 => x"08279238",
          5826 => x"9417088c",
          5827 => x"180c9017",
          5828 => x"3380c007",
          5829 => x"55749018",
          5830 => x"34941708",
          5831 => x"83ff0655",
          5832 => x"74802e80",
          5833 => x"f4389c17",
          5834 => x"087b2e80",
          5835 => x"ec389017",
          5836 => x"3370982b",
          5837 => x"565c7480",
          5838 => x"25b03881",
          5839 => x"549c1708",
          5840 => x"53a81752",
          5841 => x"7c811133",
          5842 => x"5255ffb8",
          5843 => x"f13f81d3",
          5844 => x"ac08802e",
          5845 => x"8a38810b",
          5846 => x"91183481",
          5847 => x"55bd3990",
          5848 => x"173380ff",
          5849 => x"06557490",
          5850 => x"18348154",
          5851 => x"7a53a817",
          5852 => x"527c8111",
          5853 => x"335255ff",
          5854 => x"b6eb3f81",
          5855 => x"d3ac0880",
          5856 => x"2e933881",
          5857 => x"0b911834",
          5858 => x"81559039",
          5859 => x"810b9118",
          5860 => x"34815587",
          5861 => x"397a9c18",
          5862 => x"0c795574",
          5863 => x"81d3ac0c",
          5864 => x"8e3d0d04",
          5865 => x"f93d0d79",
          5866 => x"56895475",
          5867 => x"802e818f",
          5868 => x"38805389",
          5869 => x"3dfc0552",
          5870 => x"8a3d8405",
          5871 => x"51de843f",
          5872 => x"81d3ac08",
          5873 => x"5581d3ac",
          5874 => x"0880ef38",
          5875 => x"77760c7a",
          5876 => x"527551d8",
          5877 => x"9e3f81d3",
          5878 => x"ac085581",
          5879 => x"d3ac0880",
          5880 => x"ca38ab16",
          5881 => x"3370982b",
          5882 => x"55578074",
          5883 => x"24a63886",
          5884 => x"16337084",
          5885 => x"2a708106",
          5886 => x"51555773",
          5887 => x"802e9338",
          5888 => x"9c160852",
          5889 => x"7751cec4",
          5890 => x"3f81d3ac",
          5891 => x"0888170c",
          5892 => x"83398555",
          5893 => x"74953877",
          5894 => x"54861422",
          5895 => x"84172374",
          5896 => x"527551c9",
          5897 => x"ba3f81d3",
          5898 => x"ac085574",
          5899 => x"842e0981",
          5900 => x"06833885",
          5901 => x"5574802e",
          5902 => x"84388076",
          5903 => x"0c745473",
          5904 => x"81d3ac0c",
          5905 => x"893d0d04",
          5906 => x"fc3d0d76",
          5907 => x"873dfc05",
          5908 => x"53705254",
          5909 => x"e4b93f81",
          5910 => x"d3ac0853",
          5911 => x"81d3ac08",
          5912 => x"873881d3",
          5913 => x"ac08740c",
          5914 => x"7281d3ac",
          5915 => x"0c863d0d",
          5916 => x"04fb3d0d",
          5917 => x"7779893d",
          5918 => x"fc055471",
          5919 => x"535654e4",
          5920 => x"8e3f81d3",
          5921 => x"ac085381",
          5922 => x"d3ac0880",
          5923 => x"d1387492",
          5924 => x"3881d3ac",
          5925 => x"08527351",
          5926 => x"c8c53f81",
          5927 => x"d3ac0853",
          5928 => x"bd398052",
          5929 => x"7351ce8b",
          5930 => x"3f81d3ac",
          5931 => x"085381d3",
          5932 => x"ac08842e",
          5933 => x"09810683",
          5934 => x"38805372",
          5935 => x"a1387452",
          5936 => x"7351d1b4",
          5937 => x"3f725273",
          5938 => x"51c9e93f",
          5939 => x"81d3ac08",
          5940 => x"5381d3ac",
          5941 => x"08842e09",
          5942 => x"81068338",
          5943 => x"80537281",
          5944 => x"d3ac0c87",
          5945 => x"3d0d04ef",
          5946 => x"3d0d6456",
          5947 => x"8053883d",
          5948 => x"7053953d",
          5949 => x"5254dbcb",
          5950 => x"3f81d3ac",
          5951 => x"085581d3",
          5952 => x"ac08b538",
          5953 => x"63527351",
          5954 => x"d5e93f81",
          5955 => x"d3ac0855",
          5956 => x"81d3ac08",
          5957 => x"a3380280",
          5958 => x"c7053370",
          5959 => x"982b5557",
          5960 => x"73802585",
          5961 => x"38865590",
          5962 => x"3975802e",
          5963 => x"8b387552",
          5964 => x"933dd405",
          5965 => x"51d0c13f",
          5966 => x"7481d3ac",
          5967 => x"0c933d0d",
          5968 => x"04f23d0d",
          5969 => x"6163555a",
          5970 => x"8053903d",
          5971 => x"ec055291",
          5972 => x"3d51daef",
          5973 => x"3f81d3ac",
          5974 => x"085981d3",
          5975 => x"ac088284",
          5976 => x"387a740c",
          5977 => x"73089811",
          5978 => x"08fe0555",
          5979 => x"55901508",
          5980 => x"74269338",
          5981 => x"9015087a",
          5982 => x"0c81e939",
          5983 => x"815981cf",
          5984 => x"39825981",
          5985 => x"ca39807b",
          5986 => x"70335656",
          5987 => x"5773812e",
          5988 => x"09810680",
          5989 => x"c0388275",
          5990 => x"5d567552",
          5991 => x"903df005",
          5992 => x"51ffbcaa",
          5993 => x"3f81d3ac",
          5994 => x"08ff2ed0",
          5995 => x"3881d3ac",
          5996 => x"08812ecd",
          5997 => x"3881d3ac",
          5998 => x"08307081",
          5999 => x"d3ac0807",
          6000 => x"80257805",
          6001 => x"81187d53",
          6002 => x"58585498",
          6003 => x"14087626",
          6004 => x"c93880fb",
          6005 => x"397a9811",
          6006 => x"08a41208",
          6007 => x"5a575480",
          6008 => x"55749838",
          6009 => x"77528118",
          6010 => x"7b5258ff",
          6011 => x"b9c03f81",
          6012 => x"d3ac0859",
          6013 => x"81d3ac08",
          6014 => x"80d5387a",
          6015 => x"70335154",
          6016 => x"73822e09",
          6017 => x"8106a038",
          6018 => x"7a15b405",
          6019 => x"51ffb5f0",
          6020 => x"3f81d3ac",
          6021 => x"0883ffff",
          6022 => x"06703070",
          6023 => x"80251982",
          6024 => x"18585951",
          6025 => x"549d397a",
          6026 => x"15b40551",
          6027 => x"ffb5ea3f",
          6028 => x"81d3ac08",
          6029 => x"f00a0670",
          6030 => x"30708025",
          6031 => x"19841858",
          6032 => x"59515474",
          6033 => x"83ff06ff",
          6034 => x"17575575",
          6035 => x"ff933876",
          6036 => x"7a0c7a77",
          6037 => x"90120c54",
          6038 => x"7a841133",
          6039 => x"81075555",
          6040 => x"73841634",
          6041 => x"7881d3ac",
          6042 => x"0c903d0d",
          6043 => x"04f83d0d",
          6044 => x"7a8b3dfc",
          6045 => x"05537052",
          6046 => x"58e0943f",
          6047 => x"81d3ac08",
          6048 => x"5781d3ac",
          6049 => x"088a3891",
          6050 => x"18335776",
          6051 => x"802e8638",
          6052 => x"765681dc",
          6053 => x"39901833",
          6054 => x"70812a70",
          6055 => x"81065156",
          6056 => x"56875674",
          6057 => x"802e81c8",
          6058 => x"38941808",
          6059 => x"8c190827",
          6060 => x"81bc3894",
          6061 => x"18089a38",
          6062 => x"80538818",
          6063 => x"08527751",
          6064 => x"ffbecf3f",
          6065 => x"81d3ac08",
          6066 => x"57800b88",
          6067 => x"190c80ca",
          6068 => x"39981808",
          6069 => x"527751ff",
          6070 => x"b9f43f81",
          6071 => x"d3ac0881",
          6072 => x"d3ac08ff",
          6073 => x"32703070",
          6074 => x"72078025",
          6075 => x"52575856",
          6076 => x"81d3ac08",
          6077 => x"812e0981",
          6078 => x"06833882",
          6079 => x"57769b38",
          6080 => x"78557598",
          6081 => x"16082792",
          6082 => x"38981808",
          6083 => x"53755277",
          6084 => x"51ffbdfe",
          6085 => x"3f81d3ac",
          6086 => x"08579418",
          6087 => x"088c190c",
          6088 => x"90183380",
          6089 => x"c0075574",
          6090 => x"90193476",
          6091 => x"b9387498",
          6092 => x"2b557480",
          6093 => x"25ab3881",
          6094 => x"549c1808",
          6095 => x"53a81852",
          6096 => x"78811133",
          6097 => x"5255ffb0",
          6098 => x"f53f81d3",
          6099 => x"ac08802e",
          6100 => x"85388157",
          6101 => x"8c399018",
          6102 => x"3380ff06",
          6103 => x"55749019",
          6104 => x"3476802e",
          6105 => x"89387691",
          6106 => x"19347656",
          6107 => x"83397656",
          6108 => x"7581d3ac",
          6109 => x"0c8a3d0d",
          6110 => x"04e33d0d",
          6111 => x"81baf051",
          6112 => x"ff96d53f",
          6113 => x"82539f3d",
          6114 => x"ffa40552",
          6115 => x"a03d51d6",
          6116 => x"b23f81d3",
          6117 => x"ac085681",
          6118 => x"d3ac0882",
          6119 => x"d33881ba",
          6120 => x"f451ff96",
          6121 => x"b33f7744",
          6122 => x"6f529f3d",
          6123 => x"d40551d0",
          6124 => x"c23f81d3",
          6125 => x"ac0881ba",
          6126 => x"f85256ff",
          6127 => x"969a3f75",
          6128 => x"82ae3802",
          6129 => x"80f70533",
          6130 => x"70852a70",
          6131 => x"81065155",
          6132 => x"5573802e",
          6133 => x"83388656",
          6134 => x"75829538",
          6135 => x"81bafc51",
          6136 => x"ff95f53f",
          6137 => x"0280f705",
          6138 => x"3370982b",
          6139 => x"55557380",
          6140 => x"25853886",
          6141 => x"56903902",
          6142 => x"80d20533",
          6143 => x"81065473",
          6144 => x"802e8338",
          6145 => x"87567581",
          6146 => x"e7386a52",
          6147 => x"7751c6bc",
          6148 => x"3f81d3ac",
          6149 => x"08028405",
          6150 => x"80d20533",
          6151 => x"70842a70",
          6152 => x"81065156",
          6153 => x"56577380",
          6154 => x"2e80e538",
          6155 => x"81bb8051",
          6156 => x"ff95a53f",
          6157 => x"87785556",
          6158 => x"94140877",
          6159 => x"2e80d138",
          6160 => x"81bb8451",
          6161 => x"ff95913f",
          6162 => x"7759765b",
          6163 => x"81bb8851",
          6164 => x"ff95853f",
          6165 => x"8052893d",
          6166 => x"705254c1",
          6167 => x"823f81d3",
          6168 => x"ac085681",
          6169 => x"d3ac0881",
          6170 => x"873881d3",
          6171 => x"ac085273",
          6172 => x"51c6c03f",
          6173 => x"81d3ac08",
          6174 => x"5681d3ac",
          6175 => x"08833887",
          6176 => x"56758432",
          6177 => x"70307072",
          6178 => x"079f2c78",
          6179 => x"06585654",
          6180 => x"7580dd38",
          6181 => x"81bb8c51",
          6182 => x"ff94bd3f",
          6183 => x"9f3dd405",
          6184 => x"51c9a43f",
          6185 => x"81d3ac08",
          6186 => x"81d3ac08",
          6187 => x"307081d3",
          6188 => x"ac080780",
          6189 => x"25793070",
          6190 => x"7b079f2a",
          6191 => x"72065257",
          6192 => x"51565674",
          6193 => x"802e9b38",
          6194 => x"81bb9051",
          6195 => x"ff94893f",
          6196 => x"80537652",
          6197 => x"9f3dd405",
          6198 => x"51ffbab6",
          6199 => x"3f81d3ac",
          6200 => x"0856758c",
          6201 => x"387751ff",
          6202 => x"b48b3f81",
          6203 => x"d3ac0856",
          6204 => x"81bb9451",
          6205 => x"ff93e13f",
          6206 => x"7581d3ac",
          6207 => x"0c9f3d0d",
          6208 => x"04ea3d0d",
          6209 => x"8253983d",
          6210 => x"c0055299",
          6211 => x"3d51d3b3",
          6212 => x"3f81d3ac",
          6213 => x"085581d3",
          6214 => x"ac0882b5",
          6215 => x"38775d68",
          6216 => x"52983dd4",
          6217 => x"0551cdcb",
          6218 => x"3f81d3ac",
          6219 => x"085581d3",
          6220 => x"ac088338",
          6221 => x"88557484",
          6222 => x"2e098106",
          6223 => x"82933802",
          6224 => x"80db0533",
          6225 => x"70852a70",
          6226 => x"81065155",
          6227 => x"5673802e",
          6228 => x"83388655",
          6229 => x"74842e09",
          6230 => x"810681f5",
          6231 => x"38775980",
          6232 => x"52983dc4",
          6233 => x"0551ffba",
          6234 => x"dc3f81d3",
          6235 => x"ac085680",
          6236 => x"5581d3ac",
          6237 => x"08752e09",
          6238 => x"81068338",
          6239 => x"87557581",
          6240 => x"2e098106",
          6241 => x"83388255",
          6242 => x"75ff2e09",
          6243 => x"81068338",
          6244 => x"81558288",
          6245 => x"b20a5774",
          6246 => x"81aa3875",
          6247 => x"527751ff",
          6248 => x"bdc73f81",
          6249 => x"d3ac0855",
          6250 => x"81d3ac08",
          6251 => x"8196388b",
          6252 => x"53a052b4",
          6253 => x"1851ffaf",
          6254 => x"fa3f7754",
          6255 => x"ae0bb415",
          6256 => x"34775490",
          6257 => x"0bbf1534",
          6258 => x"765280ca",
          6259 => x"1851ffaf",
          6260 => x"8f3f7553",
          6261 => x"b4185277",
          6262 => x"51c3aa3f",
          6263 => x"a053b418",
          6264 => x"5280d418",
          6265 => x"51ffafa7",
          6266 => x"3f7754ae",
          6267 => x"0b80d515",
          6268 => x"347e5380",
          6269 => x"d4185277",
          6270 => x"51c38a3f",
          6271 => x"7754810b",
          6272 => x"83153498",
          6273 => x"3dd40551",
          6274 => x"c5e73f81",
          6275 => x"d3ac0855",
          6276 => x"81d3ac08",
          6277 => x"af387652",
          6278 => x"63960551",
          6279 => x"ffaec13f",
          6280 => x"75536352",
          6281 => x"7751c2dd",
          6282 => x"3f635490",
          6283 => x"0b8b1534",
          6284 => x"7754810b",
          6285 => x"83153477",
          6286 => x"51ffb1b9",
          6287 => x"3f81d3ac",
          6288 => x"08558e39",
          6289 => x"80537552",
          6290 => x"983dc405",
          6291 => x"51ffb7c2",
          6292 => x"3f7481d3",
          6293 => x"ac0c983d",
          6294 => x"0d04db3d",
          6295 => x"0da83d84",
          6296 => x"0551cdc8",
          6297 => x"3f8253a7",
          6298 => x"3dff8405",
          6299 => x"52a83d51",
          6300 => x"d0d13f81",
          6301 => x"d3ac0855",
          6302 => x"81d3ac08",
          6303 => x"82d73877",
          6304 => x"4ca83d08",
          6305 => x"52a73dd4",
          6306 => x"0551cae7",
          6307 => x"3f81d3ac",
          6308 => x"085581d3",
          6309 => x"ac0882bd",
          6310 => x"38028197",
          6311 => x"053381a0",
          6312 => x"06547380",
          6313 => x"2e833886",
          6314 => x"557482a9",
          6315 => x"38a053a3",
          6316 => x"3d0852a7",
          6317 => x"3dff8805",
          6318 => x"51ffadd3",
          6319 => x"3fac53a7",
          6320 => x"3dd40552",
          6321 => x"913d7052",
          6322 => x"54ffadc3",
          6323 => x"3fa93d08",
          6324 => x"527351ca",
          6325 => x"9e3f81d3",
          6326 => x"ac085581",
          6327 => x"d3ac0894",
          6328 => x"38626e2e",
          6329 => x"0981068a",
          6330 => x"38845564",
          6331 => x"a13d082e",
          6332 => x"83388855",
          6333 => x"74842e09",
          6334 => x"810681b8",
          6335 => x"38a73dff",
          6336 => x"a80551c3",
          6337 => x"ec3f81d3",
          6338 => x"ac085581",
          6339 => x"d3ac0881",
          6340 => x"c4386756",
          6341 => x"9353a73d",
          6342 => x"ff950552",
          6343 => x"8d1651ff",
          6344 => x"aced3f02",
          6345 => x"ab05338b",
          6346 => x"17348b16",
          6347 => x"3370842a",
          6348 => x"70810651",
          6349 => x"55577389",
          6350 => x"3876a007",
          6351 => x"54738b17",
          6352 => x"34775481",
          6353 => x"0b831534",
          6354 => x"8b163370",
          6355 => x"842a7081",
          6356 => x"06515557",
          6357 => x"73802e80",
          6358 => x"db386d63",
          6359 => x"2e80d538",
          6360 => x"75527751",
          6361 => x"ffbfe53f",
          6362 => x"81d3ac08",
          6363 => x"527751ff",
          6364 => x"b0b23f82",
          6365 => x"5581d3ac",
          6366 => x"08802eb8",
          6367 => x"3881d3ac",
          6368 => x"08527751",
          6369 => x"ffaea73f",
          6370 => x"81d3ac08",
          6371 => x"80d41957",
          6372 => x"5581d3ac",
          6373 => x"08bf3881",
          6374 => x"16335473",
          6375 => x"ae2e0981",
          6376 => x"06923862",
          6377 => x"53755277",
          6378 => x"51ffbfd9",
          6379 => x"3f775481",
          6380 => x"0b831534",
          6381 => x"749f38a7",
          6382 => x"3dd40551",
          6383 => x"c3893f81",
          6384 => x"d3ac0855",
          6385 => x"81d3ac08",
          6386 => x"8c387751",
          6387 => x"ffaea63f",
          6388 => x"81d3ac08",
          6389 => x"557481d3",
          6390 => x"ac0ca73d",
          6391 => x"0d04ed3d",
          6392 => x"0d0280db",
          6393 => x"05330284",
          6394 => x"0580df05",
          6395 => x"33575782",
          6396 => x"53953dd0",
          6397 => x"0552963d",
          6398 => x"51cdc83f",
          6399 => x"81d3ac08",
          6400 => x"5581d3ac",
          6401 => x"0880d438",
          6402 => x"785a6552",
          6403 => x"953dd405",
          6404 => x"51c7e03f",
          6405 => x"81d3ac08",
          6406 => x"5581d3ac",
          6407 => x"08bd3802",
          6408 => x"80cf0533",
          6409 => x"81a00654",
          6410 => x"73802e83",
          6411 => x"38865574",
          6412 => x"aa3875a7",
          6413 => x"06617109",
          6414 => x"8b123371",
          6415 => x"067a7406",
          6416 => x"07515755",
          6417 => x"56748b15",
          6418 => x"34785481",
          6419 => x"0b831534",
          6420 => x"7851ffad",
          6421 => x"a03f81d3",
          6422 => x"ac085574",
          6423 => x"81d3ac0c",
          6424 => x"953d0d04",
          6425 => x"ee3d0d65",
          6426 => x"56825394",
          6427 => x"3dd00552",
          6428 => x"953d51cc",
          6429 => x"ce3f81d3",
          6430 => x"ac085581",
          6431 => x"d3ac0880",
          6432 => x"d3387759",
          6433 => x"6452943d",
          6434 => x"d40551c6",
          6435 => x"e63f81d3",
          6436 => x"ac085581",
          6437 => x"d3ac08bc",
          6438 => x"380280cb",
          6439 => x"053381a0",
          6440 => x"06547380",
          6441 => x"2e833886",
          6442 => x"5574a938",
          6443 => x"86162284",
          6444 => x"17227090",
          6445 => x"2b720754",
          6446 => x"57547f96",
          6447 => x"0551ffa9",
          6448 => x"9f3f7754",
          6449 => x"810b8315",
          6450 => x"347751ff",
          6451 => x"aca73f81",
          6452 => x"d3ac0855",
          6453 => x"7481d3ac",
          6454 => x"0c943d0d",
          6455 => x"04ea3d0d",
          6456 => x"696b5c59",
          6457 => x"8053983d",
          6458 => x"d0055299",
          6459 => x"3d51cbd3",
          6460 => x"3f81d3ac",
          6461 => x"0881d3ac",
          6462 => x"08307081",
          6463 => x"d3ac0807",
          6464 => x"80257b30",
          6465 => x"707d079f",
          6466 => x"2a720652",
          6467 => x"57515656",
          6468 => x"74802e80",
          6469 => x"f6387b5d",
          6470 => x"805f8052",
          6471 => x"8d3d7052",
          6472 => x"54ffb7bb",
          6473 => x"3f81d3ac",
          6474 => x"085681d3",
          6475 => x"ac0880ce",
          6476 => x"38815273",
          6477 => x"51ffbcfb",
          6478 => x"3f81d3ac",
          6479 => x"085681d3",
          6480 => x"ac08bb38",
          6481 => x"81d3ac08",
          6482 => x"81d3ac08",
          6483 => x"655c5858",
          6484 => x"79178118",
          6485 => x"7a1a5658",
          6486 => x"55743374",
          6487 => x"34811858",
          6488 => x"8a7727ec",
          6489 => x"38771954",
          6490 => x"80743477",
          6491 => x"802e8f38",
          6492 => x"ff187911",
          6493 => x"70335155",
          6494 => x"5873a02e",
          6495 => x"e8387584",
          6496 => x"2e098106",
          6497 => x"86388079",
          6498 => x"34805675",
          6499 => x"30707707",
          6500 => x"80257c30",
          6501 => x"707e079f",
          6502 => x"2a720652",
          6503 => x"56515574",
          6504 => x"802ebc38",
          6505 => x"7ba01108",
          6506 => x"5351ffaa",
          6507 => x"813f81d3",
          6508 => x"ac085681",
          6509 => x"d3ac08a7",
          6510 => x"387b7033",
          6511 => x"515480c3",
          6512 => x"5873832e",
          6513 => x"8b3880e4",
          6514 => x"5873842e",
          6515 => x"8338a758",
          6516 => x"7b18b405",
          6517 => x"51ffa6c1",
          6518 => x"3f81d3ac",
          6519 => x"087b0c75",
          6520 => x"81d3ac0c",
          6521 => x"983d0d04",
          6522 => x"e83d0d82",
          6523 => x"539a3dff",
          6524 => x"b805529b",
          6525 => x"3d51c9cb",
          6526 => x"3f81d3ac",
          6527 => x"085581d3",
          6528 => x"ac0883c8",
          6529 => x"388b53a0",
          6530 => x"529a3dff",
          6531 => x"bc0551ff",
          6532 => x"a7a13f80",
          6533 => x"6b707133",
          6534 => x"52575557",
          6535 => x"9f742781",
          6536 => x"b5387433",
          6537 => x"6b81054c",
          6538 => x"7081ff06",
          6539 => x"5256ffa7",
          6540 => x"fe3f81d3",
          6541 => x"ac08802e",
          6542 => x"a2386a70",
          6543 => x"33705351",
          6544 => x"54ffa7f2",
          6545 => x"3f81d3ac",
          6546 => x"08802e8d",
          6547 => x"3875882b",
          6548 => x"74076b81",
          6549 => x"054c5683",
          6550 => x"398056ff",
          6551 => x"9f165473",
          6552 => x"99268a38",
          6553 => x"e0167083",
          6554 => x"ffff0657",
          6555 => x"5480ff76",
          6556 => x"27873881",
          6557 => x"badc1633",
          6558 => x"5675802e",
          6559 => x"a3387552",
          6560 => x"81bcdc51",
          6561 => x"ffa6f73f",
          6562 => x"81d3ac08",
          6563 => x"933881ff",
          6564 => x"76278838",
          6565 => x"76892688",
          6566 => x"388b398a",
          6567 => x"77278638",
          6568 => x"865582a8",
          6569 => x"3981ff76",
          6570 => x"2793389a",
          6571 => x"3d7705ff",
          6572 => x"bc057688",
          6573 => x"2a555573",
          6574 => x"75348117",
          6575 => x"579a3d77",
          6576 => x"05ffbc05",
          6577 => x"54757434",
          6578 => x"81176b70",
          6579 => x"33565657",
          6580 => x"739f26fe",
          6581 => x"cd38893d",
          6582 => x"33548655",
          6583 => x"7381e52e",
          6584 => x"81ea3876",
          6585 => x"802ea838",
          6586 => x"029f0570",
          6587 => x"78127033",
          6588 => x"51525654",
          6589 => x"73a02e09",
          6590 => x"81069438",
          6591 => x"ff175776",
          6592 => x"802e8c38",
          6593 => x"76157033",
          6594 => x"515473a0",
          6595 => x"2eee3877",
          6596 => x"5f804180",
          6597 => x"528f3d70",
          6598 => x"5255ffb3",
          6599 => x"c23f81d3",
          6600 => x"ac085481",
          6601 => x"d3ac0881",
          6602 => x"a1388152",
          6603 => x"7451ffb9",
          6604 => x"823f81d3",
          6605 => x"ac085481",
          6606 => x"d3ac08b0",
          6607 => x"3876802e",
          6608 => x"91388b53",
          6609 => x"9a3dffbc",
          6610 => x"05526551",
          6611 => x"ffa4c03f",
          6612 => x"86396554",
          6613 => x"e5743477",
          6614 => x"54810b83",
          6615 => x"15347751",
          6616 => x"ffa7923f",
          6617 => x"81d3ac08",
          6618 => x"5480df39",
          6619 => x"81d3ac08",
          6620 => x"842e0981",
          6621 => x"0680d338",
          6622 => x"80547674",
          6623 => x"2e80cb38",
          6624 => x"81529a3d",
          6625 => x"d40551ff",
          6626 => x"b6b23f81",
          6627 => x"d3ac0854",
          6628 => x"81d3ac08",
          6629 => x"b538a053",
          6630 => x"81d3ac08",
          6631 => x"526551ff",
          6632 => x"a4913f65",
          6633 => x"54880b8b",
          6634 => x"15348b53",
          6635 => x"9a3dffbc",
          6636 => x"05526551",
          6637 => x"ffa3d83f",
          6638 => x"7754810b",
          6639 => x"83153477",
          6640 => x"51ffa6b1",
          6641 => x"3f81d3ac",
          6642 => x"08547355",
          6643 => x"7481d3ac",
          6644 => x"0c9a3d0d",
          6645 => x"04f13d0d",
          6646 => x"61630288",
          6647 => x"0580cf05",
          6648 => x"33943dfc",
          6649 => x"05557254",
          6650 => x"5e5c58cd",
          6651 => x"a23f81d3",
          6652 => x"ac085781",
          6653 => x"d3ac088a",
          6654 => x"38911833",
          6655 => x"5776802e",
          6656 => x"86387654",
          6657 => x"82b7397a",
          6658 => x"802e9538",
          6659 => x"8c180890",
          6660 => x"38901833",
          6661 => x"70812a70",
          6662 => x"81065155",
          6663 => x"55739038",
          6664 => x"87548299",
          6665 => x"39825781",
          6666 => x"89398157",
          6667 => x"8184397f",
          6668 => x"8a112270",
          6669 => x"892b7055",
          6670 => x"7d545851",
          6671 => x"54fef9dd",
          6672 => x"3fff167b",
          6673 => x"06703070",
          6674 => x"72079f2a",
          6675 => x"81d3ac08",
          6676 => x"05628c11",
          6677 => x"085d5240",
          6678 => x"5555805f",
          6679 => x"81792788",
          6680 => x"38981408",
          6681 => x"79268338",
          6682 => x"82597879",
          6683 => x"565d805a",
          6684 => x"74527751",
          6685 => x"ffa6d73f",
          6686 => x"81d3ac08",
          6687 => x"81166156",
          6688 => x"56569814",
          6689 => x"08752683",
          6690 => x"38825575",
          6691 => x"812eff95",
          6692 => x"3875ff2e",
          6693 => x"ff943875",
          6694 => x"8b38811a",
          6695 => x"5a797e2e",
          6696 => x"91388539",
          6697 => x"745d805a",
          6698 => x"74792e09",
          6699 => x"8106c138",
          6700 => x"87577681",
          6701 => x"86387b80",
          6702 => x"2eb9387c",
          6703 => x"7e57557d",
          6704 => x"802eb338",
          6705 => x"81155475",
          6706 => x"812e0981",
          6707 => x"068338ff",
          6708 => x"54735374",
          6709 => x"527f51ff",
          6710 => x"a7f03f81",
          6711 => x"d3ac0857",
          6712 => x"81d3ac08",
          6713 => x"91387481",
          6714 => x"16ff1858",
          6715 => x"565f75d4",
          6716 => x"388439ff",
          6717 => x"1d5f7680",
          6718 => x"c2387f7f",
          6719 => x"8c120c54",
          6720 => x"7b802eb7",
          6721 => x"387c8819",
          6722 => x"0c7a8c19",
          6723 => x"0c901833",
          6724 => x"80c00754",
          6725 => x"73901934",
          6726 => x"7f981108",
          6727 => x"fe055555",
          6728 => x"90150874",
          6729 => x"26953890",
          6730 => x"15087e31",
          6731 => x"90160c7f",
          6732 => x"84113381",
          6733 => x"07555573",
          6734 => x"84163476",
          6735 => x"547381d3",
          6736 => x"ac0c913d",
          6737 => x"0d04ea3d",
          6738 => x"0d6a0284",
          6739 => x"0580e705",
          6740 => x"339b3d53",
          6741 => x"5e58ffbf",
          6742 => x"d33f81d3",
          6743 => x"ac08568b",
          6744 => x"57800b81",
          6745 => x"d3ac0824",
          6746 => x"8cd13881",
          6747 => x"d3ac0810",
          6748 => x"1081d3c8",
          6749 => x"05557408",
          6750 => x"802e8738",
          6751 => x"74085580",
          6752 => x"75347581",
          6753 => x"ff065a81",
          6754 => x"527951ff",
          6755 => x"99cb3f81",
          6756 => x"d3ac0881",
          6757 => x"ff067081",
          6758 => x"06565683",
          6759 => x"57748c9b",
          6760 => x"3875822a",
          6761 => x"70810651",
          6762 => x"558a5774",
          6763 => x"8c8d3898",
          6764 => x"3dfc0553",
          6765 => x"83527951",
          6766 => x"ff9ddd3f",
          6767 => x"81d3ac08",
          6768 => x"98386680",
          6769 => x"2e933866",
          6770 => x"82808026",
          6771 => x"8c3866ff",
          6772 => x"05670655",
          6773 => x"74802e83",
          6774 => x"38814784",
          6775 => x"805e7780",
          6776 => x"2e86387d",
          6777 => x"78269238",
          6778 => x"7781800a",
          6779 => x"268b38ff",
          6780 => x"18780655",
          6781 => x"74802e86",
          6782 => x"3893578b",
          6783 => x"be397d52",
          6784 => x"7751fef6",
          6785 => x"983f81d3",
          6786 => x"ac086c7f",
          6787 => x"546e5340",
          6788 => x"58fef689",
          6789 => x"3f81d3ac",
          6790 => x"087e81d3",
          6791 => x"ac082960",
          6792 => x"30706207",
          6793 => x"802581d3",
          6794 => x"ac083070",
          6795 => x"81d3ac08",
          6796 => x"07802572",
          6797 => x"07525951",
          6798 => x"58464191",
          6799 => x"57758afb",
          6800 => x"38983df8",
          6801 => x"05538152",
          6802 => x"7951ff9c",
          6803 => x"cb3f8157",
          6804 => x"81d3ac08",
          6805 => x"8ae5387c",
          6806 => x"832a7081",
          6807 => x"06515580",
          6808 => x"4474642e",
          6809 => x"09810683",
          6810 => x"38bf448e",
          6811 => x"57636626",
          6812 => x"8ac93865",
          6813 => x"6431468e",
          6814 => x"5780ff66",
          6815 => x"278abc38",
          6816 => x"93577781",
          6817 => x"80268ab3",
          6818 => x"387c812a",
          6819 => x"70810651",
          6820 => x"5574802e",
          6821 => x"95387c87",
          6822 => x"06557482",
          6823 => x"2e88387c",
          6824 => x"81065574",
          6825 => x"85388342",
          6826 => x"8f397c81",
          6827 => x"06559357",
          6828 => x"82427480",
          6829 => x"2e8a8438",
          6830 => x"77596183",
          6831 => x"2e098106",
          6832 => x"80f13877",
          6833 => x"b4386591",
          6834 => x"2a785c57",
          6835 => x"810b81bd",
          6836 => x"80707122",
          6837 => x"52585659",
          6838 => x"74802e9d",
          6839 => x"38747726",
          6840 => x"9838811b",
          6841 => x"79107110",
          6842 => x"18702251",
          6843 => x"575a5b74",
          6844 => x"802e8638",
          6845 => x"767527ea",
          6846 => x"38785265",
          6847 => x"51fef49d",
          6848 => x"3f81d3ac",
          6849 => x"0881d3ac",
          6850 => x"0810101f",
          6851 => x"7f548705",
          6852 => x"5256fef4",
          6853 => x"883f81d3",
          6854 => x"ac085ca0",
          6855 => x"5b800bfc",
          6856 => x"808a1756",
          6857 => x"43fdfff0",
          6858 => x"0a752781",
          6859 => x"8b388e57",
          6860 => x"89893977",
          6861 => x"b438658c",
          6862 => x"2a785c57",
          6863 => x"810b81bc",
          6864 => x"f0707122",
          6865 => x"52585659",
          6866 => x"74802e9d",
          6867 => x"38747726",
          6868 => x"9838811b",
          6869 => x"79107110",
          6870 => x"18702251",
          6871 => x"575a5b74",
          6872 => x"802e8638",
          6873 => x"767527ea",
          6874 => x"38785265",
          6875 => x"51fef3ad",
          6876 => x"3f81d3ac",
          6877 => x"08108405",
          6878 => x"5781d3ac",
          6879 => x"089ff526",
          6880 => x"9238810b",
          6881 => x"81d3ac08",
          6882 => x"83291170",
          6883 => x"722a8305",
          6884 => x"5158427d",
          6885 => x"52761eff",
          6886 => x"0551fef3",
          6887 => x"803f81d3",
          6888 => x"ac085c81",
          6889 => x"7e535b81",
          6890 => x"808051fe",
          6891 => x"f2ef3f81",
          6892 => x"d3ac0883",
          6893 => x"ffff0643",
          6894 => x"631b7c11",
          6895 => x"64056811",
          6896 => x"ff056930",
          6897 => x"70720673",
          6898 => x"31525859",
          6899 => x"57406183",
          6900 => x"2e098106",
          6901 => x"8938761b",
          6902 => x"6018415b",
          6903 => x"8439761c",
          6904 => x"5c789029",
          6905 => x"16706531",
          6906 => x"51557466",
          6907 => x"2687be38",
          6908 => x"657b317c",
          6909 => x"31795370",
          6910 => x"64315256",
          6911 => x"fef29e3f",
          6912 => x"81d3ac08",
          6913 => x"5661832e",
          6914 => x"0981069b",
          6915 => x"3881d3ac",
          6916 => x"0883fff5",
          6917 => x"26913877",
          6918 => x"89387881",
          6919 => x"2a5877fd",
          6920 => x"97388e57",
          6921 => x"87953961",
          6922 => x"822e0981",
          6923 => x"0680d338",
          6924 => x"83fff576",
          6925 => x"27b43877",
          6926 => x"8f387819",
          6927 => x"557480c0",
          6928 => x"26863874",
          6929 => x"58fcf139",
          6930 => x"7c812a81",
          6931 => x"06557480",
          6932 => x"2e863883",
          6933 => x"42fce139",
          6934 => x"778b3878",
          6935 => x"19588180",
          6936 => x"7827fcd4",
          6937 => x"388e5786",
          6938 => x"d239759f",
          6939 => x"f5269338",
          6940 => x"778b3878",
          6941 => x"19588180",
          6942 => x"7827fcbc",
          6943 => x"388e5786",
          6944 => x"ba398055",
          6945 => x"61812e09",
          6946 => x"81068338",
          6947 => x"6155759f",
          6948 => x"f5267506",
          6949 => x"558e5774",
          6950 => x"86a1387d",
          6951 => x"5380527e",
          6952 => x"51ff9a8f",
          6953 => x"3f8b5381",
          6954 => x"bb98527e",
          6955 => x"51ff99df",
          6956 => x"3f7d528b",
          6957 => x"1f51ff99",
          6958 => x"893f787f",
          6959 => x"8d05347a",
          6960 => x"83ffff06",
          6961 => x"528e1f51",
          6962 => x"ff98f73f",
          6963 => x"817f9005",
          6964 => x"34618332",
          6965 => x"70307096",
          6966 => x"2a848006",
          6967 => x"54515591",
          6968 => x"1f51ff98",
          6969 => x"dd3f6583",
          6970 => x"ffff2690",
          6971 => x"380280d6",
          6972 => x"05225293",
          6973 => x"1f51ff98",
          6974 => x"c93f8a39",
          6975 => x"6552a01f",
          6976 => x"51ff98dc",
          6977 => x"3ff87f95",
          6978 => x"0534bf52",
          6979 => x"981f51ff",
          6980 => x"98b03f81",
          6981 => x"ff529a1f",
          6982 => x"51ff98a6",
          6983 => x"3f63529c",
          6984 => x"1f51ff98",
          6985 => x"bb3f6183",
          6986 => x"2e098106",
          6987 => x"80cf3882",
          6988 => x"88b20a52",
          6989 => x"80c31f51",
          6990 => x"ff98a53f",
          6991 => x"7b52a41f",
          6992 => x"51ff989c",
          6993 => x"3f8252ac",
          6994 => x"1f51ff98",
          6995 => x"933f8152",
          6996 => x"b01f51ff",
          6997 => x"97ec3f86",
          6998 => x"52b21f51",
          6999 => x"ff97e33f",
          7000 => x"ff807f80",
          7001 => x"c00534a9",
          7002 => x"7f80c205",
          7003 => x"34935381",
          7004 => x"bba45280",
          7005 => x"c71f51ff",
          7006 => x"98953fb2",
          7007 => x"398288b2",
          7008 => x"0a52a71f",
          7009 => x"51ff97d8",
          7010 => x"3f7b83ff",
          7011 => x"ff065296",
          7012 => x"1f51ff97",
          7013 => x"ad3fff80",
          7014 => x"7fa40534",
          7015 => x"a97fa605",
          7016 => x"34935381",
          7017 => x"bbb852ab",
          7018 => x"1f51ff97",
          7019 => x"e23f82d4",
          7020 => x"d55283fe",
          7021 => x"1f51ff97",
          7022 => x"893f8154",
          7023 => x"63537e52",
          7024 => x"7951ff93",
          7025 => x"f93f8157",
          7026 => x"81d3ac08",
          7027 => x"83ed3861",
          7028 => x"832e0981",
          7029 => x"0680f038",
          7030 => x"81546386",
          7031 => x"05537e52",
          7032 => x"7951ff93",
          7033 => x"d93f7d53",
          7034 => x"80527e51",
          7035 => x"ff97c43f",
          7036 => x"848b85a4",
          7037 => x"d2527e51",
          7038 => x"ff96e53f",
          7039 => x"868a85e4",
          7040 => x"f25283e4",
          7041 => x"1f51ff96",
          7042 => x"d73fff16",
          7043 => x"5283e81f",
          7044 => x"51ff96cc",
          7045 => x"3f825283",
          7046 => x"ec1f51ff",
          7047 => x"96c23f82",
          7048 => x"d4d55283",
          7049 => x"fe1f51ff",
          7050 => x"96983f81",
          7051 => x"54638705",
          7052 => x"537e5279",
          7053 => x"51ff9386",
          7054 => x"3f815463",
          7055 => x"8105537e",
          7056 => x"527951ff",
          7057 => x"92f83f64",
          7058 => x"5380527e",
          7059 => x"51ff96e3",
          7060 => x"3f7f5680",
          7061 => x"5b61832e",
          7062 => x"0981069e",
          7063 => x"38f8527e",
          7064 => x"51ff95fc",
          7065 => x"3fff5284",
          7066 => x"1f51ff95",
          7067 => x"f33ff00a",
          7068 => x"52881f51",
          7069 => x"ff95e93f",
          7070 => x"953987ff",
          7071 => x"fff85561",
          7072 => x"812e8338",
          7073 => x"f8557452",
          7074 => x"7e51ff95",
          7075 => x"d33f7b55",
          7076 => x"60577461",
          7077 => x"26833874",
          7078 => x"57765475",
          7079 => x"537e5279",
          7080 => x"51ff929a",
          7081 => x"3f81d3ac",
          7082 => x"08828638",
          7083 => x"7d538052",
          7084 => x"7e51ff95",
          7085 => x"fe3f7616",
          7086 => x"75783156",
          7087 => x"5674d138",
          7088 => x"811b5b7a",
          7089 => x"802eff8d",
          7090 => x"38785561",
          7091 => x"832e8338",
          7092 => x"62556057",
          7093 => x"74612683",
          7094 => x"38745776",
          7095 => x"5475537e",
          7096 => x"527951ff",
          7097 => x"91d83f81",
          7098 => x"d3ac0881",
          7099 => x"c8387616",
          7100 => x"75783156",
          7101 => x"5674db38",
          7102 => x"8c576183",
          7103 => x"2e933886",
          7104 => x"576583ff",
          7105 => x"ff268a38",
          7106 => x"84576182",
          7107 => x"2e833881",
          7108 => x"577c832a",
          7109 => x"81065877",
          7110 => x"80ff387d",
          7111 => x"5377527e",
          7112 => x"51ff958f",
          7113 => x"3f82d4d5",
          7114 => x"5283fe1f",
          7115 => x"51ff9492",
          7116 => x"3f83be1f",
          7117 => x"56777634",
          7118 => x"810b8117",
          7119 => x"34810b82",
          7120 => x"17347783",
          7121 => x"17347684",
          7122 => x"17346366",
          7123 => x"055780fd",
          7124 => x"c1527651",
          7125 => x"feebc63f",
          7126 => x"fe0b8517",
          7127 => x"3481d3ac",
          7128 => x"08822abf",
          7129 => x"07557486",
          7130 => x"173481d3",
          7131 => x"ac088717",
          7132 => x"34635283",
          7133 => x"c61f51ff",
          7134 => x"93e63f65",
          7135 => x"5283ca1f",
          7136 => x"51ff93dc",
          7137 => x"3f815477",
          7138 => x"537e5279",
          7139 => x"51ff90ae",
          7140 => x"3f815781",
          7141 => x"d3ac08a3",
          7142 => x"38805380",
          7143 => x"527951ff",
          7144 => x"91f63f81",
          7145 => x"5781d3ac",
          7146 => x"0891388d",
          7147 => x"398e578b",
          7148 => x"39815787",
          7149 => x"39815783",
          7150 => x"39805776",
          7151 => x"81d3ac0c",
          7152 => x"983d0d04",
          7153 => x"ff3d0d73",
          7154 => x"52719326",
          7155 => x"81e23871",
          7156 => x"101081b1",
          7157 => x"9c055271",
          7158 => x"080481c1",
          7159 => x"dc51ff80",
          7160 => x"a93f81d4",
          7161 => x"3981c1e8",
          7162 => x"51ff809e",
          7163 => x"3f81c939",
          7164 => x"81c1fc51",
          7165 => x"ff80933f",
          7166 => x"81be3981",
          7167 => x"c29051ff",
          7168 => x"80883f81",
          7169 => x"b33981c2",
          7170 => x"a051feff",
          7171 => x"fd3f81a8",
          7172 => x"3981c2b0",
          7173 => x"51fefff2",
          7174 => x"3f819d39",
          7175 => x"81c2c451",
          7176 => x"feffe73f",
          7177 => x"81923981",
          7178 => x"c2d451fe",
          7179 => x"ffdc3f81",
          7180 => x"873981c2",
          7181 => x"ec51feff",
          7182 => x"d13f80fc",
          7183 => x"3981c384",
          7184 => x"51feffc6",
          7185 => x"3f80f139",
          7186 => x"81c39c51",
          7187 => x"feffbb3f",
          7188 => x"80e63981",
          7189 => x"c3b851fe",
          7190 => x"ffb03f80",
          7191 => x"db3981c3",
          7192 => x"cc51feff",
          7193 => x"a53f80d0",
          7194 => x"3981c3f8",
          7195 => x"51feff9a",
          7196 => x"3f80c539",
          7197 => x"81c48c51",
          7198 => x"feff8f3f",
          7199 => x"bb3981c4",
          7200 => x"ac51feff",
          7201 => x"853fb139",
          7202 => x"81c4c051",
          7203 => x"fefefb3f",
          7204 => x"a73981c4",
          7205 => x"d851fefe",
          7206 => x"f13f9d39",
          7207 => x"81c4f051",
          7208 => x"fefee73f",
          7209 => x"933981c5",
          7210 => x"8851fefe",
          7211 => x"dd3f8939",
          7212 => x"81c59451",
          7213 => x"fefed33f",
          7214 => x"833d0d04",
          7215 => x"fb3d0d77",
          7216 => x"79565674",
          7217 => x"87e72693",
          7218 => x"38745275",
          7219 => x"87e82951",
          7220 => x"fee8ca3f",
          7221 => x"81d3ac08",
          7222 => x"559a3987",
          7223 => x"e8527451",
          7224 => x"fee8ba3f",
          7225 => x"81d3ac08",
          7226 => x"527551fe",
          7227 => x"e8af3f81",
          7228 => x"d3ac0855",
          7229 => x"74547953",
          7230 => x"755281c5",
          7231 => x"a451ff84",
          7232 => x"833f873d",
          7233 => x"0d04feec",
          7234 => x"3d0d8197",
          7235 => x"3d088199",
          7236 => x"3d080288",
          7237 => x"0584e305",
          7238 => x"33717330",
          7239 => x"70750780",
          7240 => x"2587ff75",
          7241 => x"27075459",
          7242 => x"5a5c5758",
          7243 => x"93557581",
          7244 => x"87388153",
          7245 => x"77528196",
          7246 => x"3dfbd805",
          7247 => x"51ffbc99",
          7248 => x"3f81d3ac",
          7249 => x"085881d3",
          7250 => x"ac08bb38",
          7251 => x"81d3ac08",
          7252 => x"87c09888",
          7253 => x"0c81d3ac",
          7254 => x"08598196",
          7255 => x"3dfbd411",
          7256 => x"55558480",
          7257 => x"537652fb",
          7258 => x"d81551c0",
          7259 => x"f23f81d3",
          7260 => x"ac085881",
          7261 => x"d3ac088e",
          7262 => x"387a802e",
          7263 => x"89387a19",
          7264 => x"7b185859",
          7265 => x"d5398196",
          7266 => x"3dfbd805",
          7267 => x"51cac13f",
          7268 => x"77307079",
          7269 => x"0780257b",
          7270 => x"30709f2a",
          7271 => x"72065157",
          7272 => x"51567480",
          7273 => x"2e903881",
          7274 => x"c5c85387",
          7275 => x"c0988808",
          7276 => x"527851fe",
          7277 => x"873f7755",
          7278 => x"7481d3ac",
          7279 => x"0c81963d",
          7280 => x"0d04f83d",
          7281 => x"0d02b705",
          7282 => x"3357ff7d",
          7283 => x"57598053",
          7284 => x"7b527a51",
          7285 => x"feb03f81",
          7286 => x"d3ac08a4",
          7287 => x"3876802e",
          7288 => x"88387681",
          7289 => x"2e983898",
          7290 => x"39615560",
          7291 => x"5481d3ac",
          7292 => x"537f527e",
          7293 => x"51752d81",
          7294 => x"d3ac0859",
          7295 => x"83397504",
          7296 => x"7881d3ac",
          7297 => x"0c8a3d0d",
          7298 => x"04fb3d0d",
          7299 => x"029f0533",
          7300 => x"81c5d053",
          7301 => x"81c5d852",
          7302 => x"56ff81e8",
          7303 => x"3f81cbcc",
          7304 => x"70225255",
          7305 => x"fef9d63f",
          7306 => x"81c5e454",
          7307 => x"81c5f053",
          7308 => x"81153352",
          7309 => x"81c5f851",
          7310 => x"ff81c93f",
          7311 => x"75802e85",
          7312 => x"38fef6ff",
          7313 => x"3f873d0d",
          7314 => x"04fe3d0d",
          7315 => x"87c09680",
          7316 => x"0853fef9",
          7317 => x"ff3f8151",
          7318 => x"feeeff3f",
          7319 => x"81c69451",
          7320 => x"fef0f53f",
          7321 => x"8051feee",
          7322 => x"f13f7281",
          7323 => x"2a708106",
          7324 => x"51527180",
          7325 => x"2e953881",
          7326 => x"51feeede",
          7327 => x"3f81c6b0",
          7328 => x"51fef0d4",
          7329 => x"3f8051fe",
          7330 => x"eed03f72",
          7331 => x"822a7081",
          7332 => x"06515271",
          7333 => x"802e9538",
          7334 => x"8151feee",
          7335 => x"bd3f81c6",
          7336 => x"c451fef0",
          7337 => x"b33f8051",
          7338 => x"feeeaf3f",
          7339 => x"72832a70",
          7340 => x"81065152",
          7341 => x"71802e95",
          7342 => x"388151fe",
          7343 => x"ee9c3f81",
          7344 => x"c6d451fe",
          7345 => x"f0923f80",
          7346 => x"51feee8e",
          7347 => x"3f72842a",
          7348 => x"70810651",
          7349 => x"5271802e",
          7350 => x"95388151",
          7351 => x"feedfb3f",
          7352 => x"81c6e851",
          7353 => x"feeff13f",
          7354 => x"8051feed",
          7355 => x"ed3f7285",
          7356 => x"2a708106",
          7357 => x"51527180",
          7358 => x"2e953881",
          7359 => x"51feedda",
          7360 => x"3f81c6fc",
          7361 => x"51feefd0",
          7362 => x"3f8051fe",
          7363 => x"edcc3f72",
          7364 => x"862a7081",
          7365 => x"06515271",
          7366 => x"802e9538",
          7367 => x"8151feed",
          7368 => x"b93f81c7",
          7369 => x"9051feef",
          7370 => x"af3f8051",
          7371 => x"feedab3f",
          7372 => x"72872a70",
          7373 => x"81065152",
          7374 => x"71802e95",
          7375 => x"388151fe",
          7376 => x"ed983f81",
          7377 => x"c7a451fe",
          7378 => x"ef8e3f80",
          7379 => x"51feed8a",
          7380 => x"3f72882a",
          7381 => x"70810651",
          7382 => x"5271802e",
          7383 => x"95388151",
          7384 => x"feecf73f",
          7385 => x"81c7b851",
          7386 => x"feeeed3f",
          7387 => x"8051feec",
          7388 => x"e93ffef8",
          7389 => x"a83f843d",
          7390 => x"0d04fa3d",
          7391 => x"0d787008",
          7392 => x"70555657",
          7393 => x"74802e80",
          7394 => x"ed388e39",
          7395 => x"74770c85",
          7396 => x"14335380",
          7397 => x"e1398115",
          7398 => x"55807533",
          7399 => x"545472a0",
          7400 => x"2e833881",
          7401 => x"54723070",
          7402 => x"9f2a7506",
          7403 => x"515372e6",
          7404 => x"38743353",
          7405 => x"72a02e09",
          7406 => x"81068838",
          7407 => x"80757081",
          7408 => x"05573480",
          7409 => x"56759029",
          7410 => x"81cbec05",
          7411 => x"77085370",
          7412 => x"085254fe",
          7413 => x"e6d03f81",
          7414 => x"d3ac088b",
          7415 => x"38841433",
          7416 => x"5372812e",
          7417 => x"ffa63881",
          7418 => x"167081ff",
          7419 => x"065753bb",
          7420 => x"7627d238",
          7421 => x"ff537281",
          7422 => x"d3ac0c88",
          7423 => x"3d0d04ce",
          7424 => x"3d0d8070",
          7425 => x"81f6ac72",
          7426 => x"710c5d5e",
          7427 => x"5c8c5a81",
          7428 => x"527b51ff",
          7429 => x"84c33f81",
          7430 => x"d3ac0881",
          7431 => x"ff065978",
          7432 => x"7c2e0981",
          7433 => x"069f3881",
          7434 => x"c7f85296",
          7435 => x"3d705259",
          7436 => x"fefde73f",
          7437 => x"7b537852",
          7438 => x"eab01b51",
          7439 => x"ffb5ab3f",
          7440 => x"81d3ac08",
          7441 => x"5a79802e",
          7442 => x"8b3881c7",
          7443 => x"fc51fefd",
          7444 => x"b33f8539",
          7445 => x"81705e5c",
          7446 => x"81c8b451",
          7447 => x"fef7ab3f",
          7448 => x"963d7043",
          7449 => x"5980f870",
          7450 => x"545a8052",
          7451 => x"7851fee4",
          7452 => x"a43f7952",
          7453 => x"6151fefd",
          7454 => x"e53fb43d",
          7455 => x"fef80551",
          7456 => x"fdf83f81",
          7457 => x"d3ac0890",
          7458 => x"2b70902c",
          7459 => x"51597881",
          7460 => x"872685af",
          7461 => x"38781010",
          7462 => x"81b1ec05",
          7463 => x"59780804",
          7464 => x"b43dfef4",
          7465 => x"1153fef8",
          7466 => x"0551fefe",
          7467 => x"e23f81d3",
          7468 => x"ac088c38",
          7469 => x"81c8b851",
          7470 => x"fefcc93f",
          7471 => x"ff9a39b4",
          7472 => x"3dfef011",
          7473 => x"53fef805",
          7474 => x"51fefec3",
          7475 => x"3f81d3ac",
          7476 => x"08802e88",
          7477 => x"38816025",
          7478 => x"83388040",
          7479 => x"02bf0533",
          7480 => x"520280c3",
          7481 => x"053351ff",
          7482 => x"82ef3f81",
          7483 => x"d3ac0881",
          7484 => x"ff065978",
          7485 => x"8e3881c8",
          7486 => x"c851fef6",
          7487 => x"8d3f815d",
          7488 => x"fed63981",
          7489 => x"c8d851fe",
          7490 => x"f6803ffe",
          7491 => x"cb39b43d",
          7492 => x"fef41153",
          7493 => x"fef80551",
          7494 => x"fefdf43f",
          7495 => x"81d3ac08",
          7496 => x"802efeb4",
          7497 => x"38805380",
          7498 => x"520280c3",
          7499 => x"053351ff",
          7500 => x"86e63f81",
          7501 => x"d3ac0852",
          7502 => x"81c8f051",
          7503 => x"fefbc53f",
          7504 => x"fe9639b4",
          7505 => x"3dfef411",
          7506 => x"53fef805",
          7507 => x"51fefdbf",
          7508 => x"3f81d3ac",
          7509 => x"08802e87",
          7510 => x"38608926",
          7511 => x"fdfa38b4",
          7512 => x"3dfef011",
          7513 => x"53fef805",
          7514 => x"51fefda3",
          7515 => x"3f81d3ac",
          7516 => x"08863881",
          7517 => x"d3ac0840",
          7518 => x"605381c8",
          7519 => x"f852963d",
          7520 => x"705259fe",
          7521 => x"fb943f02",
          7522 => x"bf053353",
          7523 => x"78526084",
          7524 => x"b42981e0",
          7525 => x"dc0551ff",
          7526 => x"b2d03f81",
          7527 => x"d3ac0880",
          7528 => x"2e8c3881",
          7529 => x"d3ac0851",
          7530 => x"f49a3ffd",
          7531 => x"ab3981c8",
          7532 => x"c851fef4",
          7533 => x"d53f815c",
          7534 => x"fd9e39b4",
          7535 => x"3dfef805",
          7536 => x"51fee4a4",
          7537 => x"3f81d3ac",
          7538 => x"08b53dfe",
          7539 => x"f805525b",
          7540 => x"fee4fa3f",
          7541 => x"815381d3",
          7542 => x"ac08527a",
          7543 => x"51f6a73f",
          7544 => x"81d3ac08",
          7545 => x"802efcf0",
          7546 => x"3881d3ac",
          7547 => x"0851f3d4",
          7548 => x"3ffce539",
          7549 => x"b43dfef8",
          7550 => x"0551fee3",
          7551 => x"eb3f81d3",
          7552 => x"ac08b53d",
          7553 => x"fef80552",
          7554 => x"5bfee4c1",
          7555 => x"3f81d3ac",
          7556 => x"08b53dfe",
          7557 => x"f805525a",
          7558 => x"fee4b23f",
          7559 => x"81d3ac08",
          7560 => x"b53dfef8",
          7561 => x"055259fe",
          7562 => x"e4a33f81",
          7563 => x"cba85881",
          7564 => x"d3e05780",
          7565 => x"56805581",
          7566 => x"d3ac0881",
          7567 => x"ff065478",
          7568 => x"5379527a",
          7569 => x"51f6fb3f",
          7570 => x"81d3ac08",
          7571 => x"802efc88",
          7572 => x"3881d3ac",
          7573 => x"0851f2ec",
          7574 => x"3ffbfd39",
          7575 => x"81c8fc51",
          7576 => x"fef3a73f",
          7577 => x"8251fef2",
          7578 => x"8f3ffbec",
          7579 => x"3981c994",
          7580 => x"51fef396",
          7581 => x"3fa251fe",
          7582 => x"f1e23ffb",
          7583 => x"db398480",
          7584 => x"810b87c0",
          7585 => x"94840c84",
          7586 => x"80810b87",
          7587 => x"c094940c",
          7588 => x"81c9ac51",
          7589 => x"fef2f33f",
          7590 => x"fbbe3981",
          7591 => x"c9c051fe",
          7592 => x"f2e83f8c",
          7593 => x"80830b87",
          7594 => x"c094840c",
          7595 => x"8c80830b",
          7596 => x"87c09494",
          7597 => x"0cfba139",
          7598 => x"b43dfef4",
          7599 => x"1153fef8",
          7600 => x"0551fefa",
          7601 => x"ca3f81d3",
          7602 => x"ac08802e",
          7603 => x"fb8a3860",
          7604 => x"5281c9d4",
          7605 => x"51fef8ac",
          7606 => x"3f605978",
          7607 => x"04b43dfe",
          7608 => x"f41153fe",
          7609 => x"f80551fe",
          7610 => x"faa53f81",
          7611 => x"d3ac0880",
          7612 => x"2efae538",
          7613 => x"605281c9",
          7614 => x"f051fef8",
          7615 => x"873f6059",
          7616 => x"782d81d3",
          7617 => x"ac085e81",
          7618 => x"d3ac0880",
          7619 => x"2efac938",
          7620 => x"81d3ac08",
          7621 => x"5281ca8c",
          7622 => x"51fef7e8",
          7623 => x"3ffab939",
          7624 => x"81caa851",
          7625 => x"fef1e33f",
          7626 => x"fed1d53f",
          7627 => x"faaa3981",
          7628 => x"cac451fe",
          7629 => x"f1d43f80",
          7630 => x"59ffa039",
          7631 => x"feed843f",
          7632 => x"fa963961",
          7633 => x"70335159",
          7634 => x"78802efa",
          7635 => x"8b387c7c",
          7636 => x"06597880",
          7637 => x"2e80cb38",
          7638 => x"b43dfef8",
          7639 => x"0551fee1",
          7640 => x"873f81ca",
          7641 => x"d85681d3",
          7642 => x"ac085581",
          7643 => x"cadc5480",
          7644 => x"5381cae0",
          7645 => x"52a03d70",
          7646 => x"5259fef7",
          7647 => x"9d3f81cb",
          7648 => x"a85881d3",
          7649 => x"e0578056",
          7650 => x"61810542",
          7651 => x"61558054",
          7652 => x"83808053",
          7653 => x"83808052",
          7654 => x"7851f4a6",
          7655 => x"3f81d3ac",
          7656 => x"085e7c81",
          7657 => x"327c8132",
          7658 => x"0759788a",
          7659 => x"387dff2e",
          7660 => x"098106f9",
          7661 => x"a33881ca",
          7662 => x"f051fef6",
          7663 => x"c73ff998",
          7664 => x"39803d0d",
          7665 => x"800b81d3",
          7666 => x"e0349b90",
          7667 => x"86e40b87",
          7668 => x"c0948c0c",
          7669 => x"9b9086e4",
          7670 => x"0b87c094",
          7671 => x"9c0c8c80",
          7672 => x"830b87c0",
          7673 => x"94840c8c",
          7674 => x"80830b87",
          7675 => x"c094940c",
          7676 => x"93f40b81",
          7677 => x"d3bc0c96",
          7678 => x"e70b81d3",
          7679 => x"c00cfee8",
          7680 => x"893ffeee",
          7681 => x"cf3f81cb",
          7682 => x"8051fee5",
          7683 => x"cb3f81cb",
          7684 => x"8c51feef",
          7685 => x"f53f81a4",
          7686 => x"c951feee",
          7687 => x"b23f8151",
          7688 => x"f3e73ff7",
          7689 => x"da3f8004",
          7690 => x"00000f44",
          7691 => x"00000f17",
          7692 => x"00000f20",
          7693 => x"00000f29",
          7694 => x"00000f32",
          7695 => x"00000f3b",
          7696 => x"000011b6",
          7697 => x"000011a7",
          7698 => x"000011be",
          7699 => x"000011c6",
          7700 => x"000011c6",
          7701 => x"000011c6",
          7702 => x"000011c6",
          7703 => x"000011c6",
          7704 => x"000011c6",
          7705 => x"000011c6",
          7706 => x"000011c6",
          7707 => x"000011c6",
          7708 => x"000011c6",
          7709 => x"000011ba",
          7710 => x"000011c6",
          7711 => x"000011c6",
          7712 => x"000011c6",
          7713 => x"0000113a",
          7714 => x"000011c6",
          7715 => x"000011be",
          7716 => x"000011c6",
          7717 => x"000011c6",
          7718 => x"000011c2",
          7719 => x"000050a6",
          7720 => x"00004fda",
          7721 => x"00004fe5",
          7722 => x"00004ff0",
          7723 => x"00004ffb",
          7724 => x"00005006",
          7725 => x"00005011",
          7726 => x"0000501c",
          7727 => x"00005027",
          7728 => x"00005032",
          7729 => x"0000503d",
          7730 => x"00005048",
          7731 => x"00005053",
          7732 => x"0000505e",
          7733 => x"00005069",
          7734 => x"00005074",
          7735 => x"0000507e",
          7736 => x"00005088",
          7737 => x"00005092",
          7738 => x"0000509c",
          7739 => x"00005458",
          7740 => x"00005743",
          7741 => x"000054a0",
          7742 => x"00005743",
          7743 => x"0000550e",
          7744 => x"00005743",
          7745 => x"00005743",
          7746 => x"00005743",
          7747 => x"00005743",
          7748 => x"00005743",
          7749 => x"00005743",
          7750 => x"00005743",
          7751 => x"00005743",
          7752 => x"00005743",
          7753 => x"00005743",
          7754 => x"00005743",
          7755 => x"00005743",
          7756 => x"00005743",
          7757 => x"00005743",
          7758 => x"00005743",
          7759 => x"00005543",
          7760 => x"00005743",
          7761 => x"00005743",
          7762 => x"00005743",
          7763 => x"00005743",
          7764 => x"00005743",
          7765 => x"00005743",
          7766 => x"00005743",
          7767 => x"00005743",
          7768 => x"00005743",
          7769 => x"00005743",
          7770 => x"00005743",
          7771 => x"00005743",
          7772 => x"00005743",
          7773 => x"00005743",
          7774 => x"00005743",
          7775 => x"00005743",
          7776 => x"00005743",
          7777 => x"00005743",
          7778 => x"00005743",
          7779 => x"00005743",
          7780 => x"00005743",
          7781 => x"00005743",
          7782 => x"000055bb",
          7783 => x"00005743",
          7784 => x"00005743",
          7785 => x"00005743",
          7786 => x"00005743",
          7787 => x"000055f4",
          7788 => x"00005743",
          7789 => x"00005743",
          7790 => x"00005743",
          7791 => x"00005743",
          7792 => x"00005743",
          7793 => x"00005743",
          7794 => x"00005743",
          7795 => x"00005743",
          7796 => x"00005743",
          7797 => x"00005743",
          7798 => x"00005743",
          7799 => x"00005743",
          7800 => x"00005743",
          7801 => x"00005743",
          7802 => x"00005743",
          7803 => x"00005743",
          7804 => x"00005743",
          7805 => x"00005743",
          7806 => x"00005743",
          7807 => x"00005743",
          7808 => x"00005743",
          7809 => x"00005743",
          7810 => x"00005743",
          7811 => x"00005743",
          7812 => x"00005743",
          7813 => x"00005743",
          7814 => x"00005743",
          7815 => x"00005743",
          7816 => x"00005743",
          7817 => x"00005743",
          7818 => x"00005743",
          7819 => x"0000565c",
          7820 => x"0000566d",
          7821 => x"00005743",
          7822 => x"00005743",
          7823 => x"0000567e",
          7824 => x"0000569b",
          7825 => x"00005743",
          7826 => x"00005743",
          7827 => x"00005743",
          7828 => x"00005743",
          7829 => x"00005743",
          7830 => x"00005743",
          7831 => x"00005743",
          7832 => x"00005743",
          7833 => x"00005743",
          7834 => x"00005743",
          7835 => x"00005743",
          7836 => x"00005743",
          7837 => x"00005743",
          7838 => x"00005743",
          7839 => x"00005743",
          7840 => x"00005743",
          7841 => x"00005743",
          7842 => x"00005743",
          7843 => x"00005743",
          7844 => x"00005743",
          7845 => x"00005743",
          7846 => x"00005743",
          7847 => x"00005743",
          7848 => x"00005743",
          7849 => x"00005743",
          7850 => x"00005743",
          7851 => x"00005743",
          7852 => x"00005743",
          7853 => x"00005743",
          7854 => x"00005743",
          7855 => x"00005743",
          7856 => x"00005743",
          7857 => x"00005743",
          7858 => x"00005743",
          7859 => x"000056b8",
          7860 => x"000056dd",
          7861 => x"00005743",
          7862 => x"00005743",
          7863 => x"00005743",
          7864 => x"00005743",
          7865 => x"00005743",
          7866 => x"00005743",
          7867 => x"00005743",
          7868 => x"00005743",
          7869 => x"00005720",
          7870 => x"0000572f",
          7871 => x"00005743",
          7872 => x"0000573c",
          7873 => x"00005743",
          7874 => x"00005458",
          7875 => x"25642f25",
          7876 => x"642f2564",
          7877 => x"2025643a",
          7878 => x"25643a25",
          7879 => x"642e2564",
          7880 => x"25640a00",
          7881 => x"536f4320",
          7882 => x"436f6e66",
          7883 => x"69677572",
          7884 => x"6174696f",
          7885 => x"6e000000",
          7886 => x"20286672",
          7887 => x"6f6d2053",
          7888 => x"6f432063",
          7889 => x"6f6e6669",
          7890 => x"67290000",
          7891 => x"3a0a4465",
          7892 => x"76696365",
          7893 => x"7320696d",
          7894 => x"706c656d",
          7895 => x"656e7465",
          7896 => x"643a0a00",
          7897 => x"20202020",
          7898 => x"494e534e",
          7899 => x"20425241",
          7900 => x"4d202853",
          7901 => x"74617274",
          7902 => x"3d253038",
          7903 => x"582c2053",
          7904 => x"697a653d",
          7905 => x"25303858",
          7906 => x"292e0a00",
          7907 => x"20202020",
          7908 => x"4252414d",
          7909 => x"20285374",
          7910 => x"6172743d",
          7911 => x"25303858",
          7912 => x"2c205369",
          7913 => x"7a653d25",
          7914 => x"30385829",
          7915 => x"2e0a0000",
          7916 => x"20202020",
          7917 => x"52414d20",
          7918 => x"28537461",
          7919 => x"72743d25",
          7920 => x"3038582c",
          7921 => x"2053697a",
          7922 => x"653d2530",
          7923 => x"3858292e",
          7924 => x"0a000000",
          7925 => x"20202020",
          7926 => x"494f4354",
          7927 => x"4c0a0000",
          7928 => x"20202020",
          7929 => x"5053320a",
          7930 => x"00000000",
          7931 => x"20202020",
          7932 => x"5350490a",
          7933 => x"00000000",
          7934 => x"20202020",
          7935 => x"53442043",
          7936 => x"61726420",
          7937 => x"28446576",
          7938 => x"69636573",
          7939 => x"3d253032",
          7940 => x"58292e0a",
          7941 => x"00000000",
          7942 => x"20202020",
          7943 => x"494e5445",
          7944 => x"52525550",
          7945 => x"5420434f",
          7946 => x"4e54524f",
          7947 => x"4c4c4552",
          7948 => x"0a000000",
          7949 => x"20202020",
          7950 => x"54494d45",
          7951 => x"52312028",
          7952 => x"54696d65",
          7953 => x"72733d25",
          7954 => x"30315829",
          7955 => x"2e0a0000",
          7956 => x"41646472",
          7957 => x"65737365",
          7958 => x"733a0a00",
          7959 => x"20202020",
          7960 => x"43505520",
          7961 => x"52657365",
          7962 => x"74205665",
          7963 => x"63746f72",
          7964 => x"20416464",
          7965 => x"72657373",
          7966 => x"203d2025",
          7967 => x"3038580a",
          7968 => x"00000000",
          7969 => x"20202020",
          7970 => x"43505520",
          7971 => x"4d656d6f",
          7972 => x"72792053",
          7973 => x"74617274",
          7974 => x"20416464",
          7975 => x"72657373",
          7976 => x"203d2025",
          7977 => x"3038580a",
          7978 => x"00000000",
          7979 => x"20202020",
          7980 => x"53746163",
          7981 => x"6b205374",
          7982 => x"61727420",
          7983 => x"41646472",
          7984 => x"65737320",
          7985 => x"20202020",
          7986 => x"203d2025",
          7987 => x"3038580a",
          7988 => x"00000000",
          7989 => x"20202020",
          7990 => x"5a505520",
          7991 => x"49642020",
          7992 => x"20202020",
          7993 => x"20202020",
          7994 => x"20202020",
          7995 => x"20202020",
          7996 => x"203d2025",
          7997 => x"3038580a",
          7998 => x"00000000",
          7999 => x"20202020",
          8000 => x"53797374",
          8001 => x"656d2043",
          8002 => x"6c6f636b",
          8003 => x"20467265",
          8004 => x"71202020",
          8005 => x"20202020",
          8006 => x"203d2025",
          8007 => x"3038580a",
          8008 => x"00000000",
          8009 => x"536d616c",
          8010 => x"6c000000",
          8011 => x"4d656469",
          8012 => x"756d0000",
          8013 => x"466c6578",
          8014 => x"00000000",
          8015 => x"45564f00",
          8016 => x"45564f6d",
          8017 => x"696e0000",
          8018 => x"556e6b6e",
          8019 => x"6f776e00",
          8020 => x"53440000",
          8021 => x"222a2b2c",
          8022 => x"3a3b3c3d",
          8023 => x"3e3f5b5d",
          8024 => x"7c7f0000",
          8025 => x"46415400",
          8026 => x"46415433",
          8027 => x"32000000",
          8028 => x"300a0000",
          8029 => x"310a0000",
          8030 => x"320a0000",
          8031 => x"330a0000",
          8032 => x"350a0000",
          8033 => x"360a0000",
          8034 => x"370a0000",
          8035 => x"380a0000",
          8036 => x"390a0000",
          8037 => x"31300a00",
          8038 => x"ebfe904d",
          8039 => x"53444f53",
          8040 => x"352e3000",
          8041 => x"4e4f204e",
          8042 => x"414d4520",
          8043 => x"20202046",
          8044 => x"41543332",
          8045 => x"20202000",
          8046 => x"4e4f204e",
          8047 => x"414d4520",
          8048 => x"20202046",
          8049 => x"41542020",
          8050 => x"20202000",
          8051 => x"00005d50",
          8052 => x"00000000",
          8053 => x"00000000",
          8054 => x"00000000",
          8055 => x"809a4541",
          8056 => x"8e418f80",
          8057 => x"45454549",
          8058 => x"49498e8f",
          8059 => x"9092924f",
          8060 => x"994f5555",
          8061 => x"59999a9b",
          8062 => x"9c9d9e9f",
          8063 => x"41494f55",
          8064 => x"a5a5a6a7",
          8065 => x"a8a9aaab",
          8066 => x"acadaeaf",
          8067 => x"b0b1b2b3",
          8068 => x"b4b5b6b7",
          8069 => x"b8b9babb",
          8070 => x"bcbdbebf",
          8071 => x"c0c1c2c3",
          8072 => x"c4c5c6c7",
          8073 => x"c8c9cacb",
          8074 => x"cccdcecf",
          8075 => x"d0d1d2d3",
          8076 => x"d4d5d6d7",
          8077 => x"d8d9dadb",
          8078 => x"dcdddedf",
          8079 => x"e0e1e2e3",
          8080 => x"e4e5e6e7",
          8081 => x"e8e9eaeb",
          8082 => x"ecedeeef",
          8083 => x"f0f1f2f3",
          8084 => x"f4f5f6f7",
          8085 => x"f8f9fafb",
          8086 => x"fcfdfeff",
          8087 => x"2b2e2c3b",
          8088 => x"3d5b5d2f",
          8089 => x"5c222a3a",
          8090 => x"3c3e3f7c",
          8091 => x"7f000000",
          8092 => x"00010004",
          8093 => x"00100040",
          8094 => x"01000200",
          8095 => x"00000000",
          8096 => x"00010002",
          8097 => x"00040008",
          8098 => x"00100020",
          8099 => x"00000000",
          8100 => x"46415431",
          8101 => x"32000000",
          8102 => x"46415431",
          8103 => x"36000000",
          8104 => x"65784641",
          8105 => x"54000000",
          8106 => x"4449534b",
          8107 => x"20494f20",
          8108 => x"434f4e54",
          8109 => x"524f4c53",
          8110 => x"00000000",
          8111 => x"4449534b",
          8112 => x"20425546",
          8113 => x"46455220",
          8114 => x"434f4e54",
          8115 => x"524f4c53",
          8116 => x"00000000",
          8117 => x"46494c45",
          8118 => x"53595354",
          8119 => x"454d2043",
          8120 => x"4f4e5452",
          8121 => x"4f4c5300",
          8122 => x"4d454d4f",
          8123 => x"52590000",
          8124 => x"48415244",
          8125 => x"57415245",
          8126 => x"00000000",
          8127 => x"54455354",
          8128 => x"494e4700",
          8129 => x"45584543",
          8130 => x"5554494f",
          8131 => x"4e000000",
          8132 => x"4d495343",
          8133 => x"20434f4d",
          8134 => x"4d414e44",
          8135 => x"53000000",
          8136 => x"6464756d",
          8137 => x"70000000",
          8138 => x"64696e69",
          8139 => x"74000000",
          8140 => x"64737461",
          8141 => x"74000000",
          8142 => x"64696f63",
          8143 => x"746c0000",
          8144 => x"6264756d",
          8145 => x"70000000",
          8146 => x"62656469",
          8147 => x"74000000",
          8148 => x"62726561",
          8149 => x"64000000",
          8150 => x"62777269",
          8151 => x"74650000",
          8152 => x"6266696c",
          8153 => x"6c000000",
          8154 => x"626c656e",
          8155 => x"00000000",
          8156 => x"66696e69",
          8157 => x"74000000",
          8158 => x"666f7065",
          8159 => x"6e000000",
          8160 => x"66636c6f",
          8161 => x"73650000",
          8162 => x"66736565",
          8163 => x"6b000000",
          8164 => x"66726561",
          8165 => x"64000000",
          8166 => x"66696e73",
          8167 => x"70656374",
          8168 => x"00000000",
          8169 => x"66777269",
          8170 => x"74650000",
          8171 => x"66747275",
          8172 => x"6e630000",
          8173 => x"66616c6c",
          8174 => x"6f630000",
          8175 => x"66617474",
          8176 => x"72000000",
          8177 => x"6674696d",
          8178 => x"65000000",
          8179 => x"6672656e",
          8180 => x"616d6500",
          8181 => x"6664656c",
          8182 => x"00000000",
          8183 => x"666d6b64",
          8184 => x"69720000",
          8185 => x"66737461",
          8186 => x"74000000",
          8187 => x"66646972",
          8188 => x"00000000",
          8189 => x"66636174",
          8190 => x"00000000",
          8191 => x"66637000",
          8192 => x"66636f6e",
          8193 => x"63617400",
          8194 => x"66787472",
          8195 => x"61637400",
          8196 => x"666c6f61",
          8197 => x"64000000",
          8198 => x"66657865",
          8199 => x"63000000",
          8200 => x"66736176",
          8201 => x"65000000",
          8202 => x"6664756d",
          8203 => x"70000000",
          8204 => x"66636400",
          8205 => x"66647269",
          8206 => x"76650000",
          8207 => x"6673686f",
          8208 => x"77646972",
          8209 => x"00000000",
          8210 => x"666c6162",
          8211 => x"656c0000",
          8212 => x"666d6b66",
          8213 => x"73000000",
          8214 => x"6d636c72",
          8215 => x"00000000",
          8216 => x"6d64756d",
          8217 => x"70000000",
          8218 => x"6d656200",
          8219 => x"6d656800",
          8220 => x"6d657700",
          8221 => x"68696400",
          8222 => x"68696500",
          8223 => x"68720000",
          8224 => x"68740000",
          8225 => x"68666400",
          8226 => x"68666500",
          8227 => x"64687279",
          8228 => x"00000000",
          8229 => x"636f7265",
          8230 => x"6d61726b",
          8231 => x"00000000",
          8232 => x"63616c6c",
          8233 => x"00000000",
          8234 => x"6a6d7000",
          8235 => x"72657374",
          8236 => x"61727400",
          8237 => x"72657365",
          8238 => x"74000000",
          8239 => x"68656c70",
          8240 => x"00000000",
          8241 => x"696e666f",
          8242 => x"00000000",
          8243 => x"74696d65",
          8244 => x"00000000",
          8245 => x"74657374",
          8246 => x"00000000",
          8247 => x"4469736b",
          8248 => x"20457272",
          8249 => x"6f720a00",
          8250 => x"496e7465",
          8251 => x"726e616c",
          8252 => x"20657272",
          8253 => x"6f722e0a",
          8254 => x"00000000",
          8255 => x"4469736b",
          8256 => x"206e6f74",
          8257 => x"20726561",
          8258 => x"64792e0a",
          8259 => x"00000000",
          8260 => x"4e6f2066",
          8261 => x"696c6520",
          8262 => x"666f756e",
          8263 => x"642e0a00",
          8264 => x"4e6f2070",
          8265 => x"61746820",
          8266 => x"666f756e",
          8267 => x"642e0a00",
          8268 => x"496e7661",
          8269 => x"6c696420",
          8270 => x"66696c65",
          8271 => x"6e616d65",
          8272 => x"2e0a0000",
          8273 => x"41636365",
          8274 => x"73732064",
          8275 => x"656e6965",
          8276 => x"642e0a00",
          8277 => x"46696c65",
          8278 => x"20616c72",
          8279 => x"65616479",
          8280 => x"20657869",
          8281 => x"7374732e",
          8282 => x"0a000000",
          8283 => x"46696c65",
          8284 => x"2068616e",
          8285 => x"646c6520",
          8286 => x"696e7661",
          8287 => x"6c69642e",
          8288 => x"0a000000",
          8289 => x"53442069",
          8290 => x"73207772",
          8291 => x"69746520",
          8292 => x"70726f74",
          8293 => x"65637465",
          8294 => x"642e0a00",
          8295 => x"44726976",
          8296 => x"65206e75",
          8297 => x"6d626572",
          8298 => x"20697320",
          8299 => x"696e7661",
          8300 => x"6c69642e",
          8301 => x"0a000000",
          8302 => x"4469736b",
          8303 => x"206e6f74",
          8304 => x"20656e61",
          8305 => x"626c6564",
          8306 => x"2e0a0000",
          8307 => x"4e6f2063",
          8308 => x"6f6d7061",
          8309 => x"7469626c",
          8310 => x"65206669",
          8311 => x"6c657379",
          8312 => x"7374656d",
          8313 => x"20666f75",
          8314 => x"6e64206f",
          8315 => x"6e206469",
          8316 => x"736b2e0a",
          8317 => x"00000000",
          8318 => x"466f726d",
          8319 => x"61742061",
          8320 => x"626f7274",
          8321 => x"65642e0a",
          8322 => x"00000000",
          8323 => x"54696d65",
          8324 => x"6f75742c",
          8325 => x"206f7065",
          8326 => x"72617469",
          8327 => x"6f6e2063",
          8328 => x"616e6365",
          8329 => x"6c6c6564",
          8330 => x"2e0a0000",
          8331 => x"46696c65",
          8332 => x"20697320",
          8333 => x"6c6f636b",
          8334 => x"65642e0a",
          8335 => x"00000000",
          8336 => x"496e7375",
          8337 => x"66666963",
          8338 => x"69656e74",
          8339 => x"206d656d",
          8340 => x"6f72792e",
          8341 => x"0a000000",
          8342 => x"546f6f20",
          8343 => x"6d616e79",
          8344 => x"206f7065",
          8345 => x"6e206669",
          8346 => x"6c65732e",
          8347 => x"0a000000",
          8348 => x"50617261",
          8349 => x"6d657465",
          8350 => x"72732069",
          8351 => x"6e636f72",
          8352 => x"72656374",
          8353 => x"2e0a0000",
          8354 => x"53756363",
          8355 => x"6573732e",
          8356 => x"0a000000",
          8357 => x"556e6b6e",
          8358 => x"6f776e20",
          8359 => x"6572726f",
          8360 => x"722e0a00",
          8361 => x"0a256c75",
          8362 => x"20627974",
          8363 => x"65732025",
          8364 => x"73206174",
          8365 => x"20256c75",
          8366 => x"20627974",
          8367 => x"65732f73",
          8368 => x"65632e0a",
          8369 => x"00000000",
          8370 => x"72656164",
          8371 => x"00000000",
          8372 => x"5a505554",
          8373 => x"41000000",
          8374 => x"0a2a2a20",
          8375 => x"25732028",
          8376 => x"00000000",
          8377 => x"31382f30",
          8378 => x"372f3230",
          8379 => x"31390000",
          8380 => x"76312e33",
          8381 => x"00000000",
          8382 => x"205a5055",
          8383 => x"2c207265",
          8384 => x"76202530",
          8385 => x"32782920",
          8386 => x"25732025",
          8387 => x"73202a2a",
          8388 => x"0a0a0000",
          8389 => x"5a505554",
          8390 => x"4120496e",
          8391 => x"74657272",
          8392 => x"75707420",
          8393 => x"48616e64",
          8394 => x"6c65720a",
          8395 => x"00000000",
          8396 => x"54696d65",
          8397 => x"7220696e",
          8398 => x"74657272",
          8399 => x"7570740a",
          8400 => x"00000000",
          8401 => x"50533220",
          8402 => x"696e7465",
          8403 => x"72727570",
          8404 => x"740a0000",
          8405 => x"494f4354",
          8406 => x"4c205244",
          8407 => x"20696e74",
          8408 => x"65727275",
          8409 => x"70740a00",
          8410 => x"494f4354",
          8411 => x"4c205752",
          8412 => x"20696e74",
          8413 => x"65727275",
          8414 => x"70740a00",
          8415 => x"55415254",
          8416 => x"30205258",
          8417 => x"20696e74",
          8418 => x"65727275",
          8419 => x"70740a00",
          8420 => x"55415254",
          8421 => x"30205458",
          8422 => x"20696e74",
          8423 => x"65727275",
          8424 => x"70740a00",
          8425 => x"55415254",
          8426 => x"31205258",
          8427 => x"20696e74",
          8428 => x"65727275",
          8429 => x"70740a00",
          8430 => x"55415254",
          8431 => x"31205458",
          8432 => x"20696e74",
          8433 => x"65727275",
          8434 => x"70740a00",
          8435 => x"53657474",
          8436 => x"696e6720",
          8437 => x"75702074",
          8438 => x"696d6572",
          8439 => x"2e2e2e0a",
          8440 => x"00000000",
          8441 => x"456e6162",
          8442 => x"6c696e67",
          8443 => x"2074696d",
          8444 => x"65722e2e",
          8445 => x"2e0a0000",
          8446 => x"303a0000",
          8447 => x"4661696c",
          8448 => x"65642074",
          8449 => x"6f20696e",
          8450 => x"69746961",
          8451 => x"6c697365",
          8452 => x"20736420",
          8453 => x"63617264",
          8454 => x"20302c20",
          8455 => x"706c6561",
          8456 => x"73652069",
          8457 => x"6e697420",
          8458 => x"6d616e75",
          8459 => x"616c6c79",
          8460 => x"2e0a0000",
          8461 => x"2a200000",
          8462 => x"42616420",
          8463 => x"6469736b",
          8464 => x"20696421",
          8465 => x"0a000000",
          8466 => x"496e6974",
          8467 => x"69616c69",
          8468 => x"7365642e",
          8469 => x"0a000000",
          8470 => x"4661696c",
          8471 => x"65642074",
          8472 => x"6f20696e",
          8473 => x"69746961",
          8474 => x"6c697365",
          8475 => x"2e0a0000",
          8476 => x"72633d25",
          8477 => x"640a0000",
          8478 => x"25753a00",
          8479 => x"44697361",
          8480 => x"626c696e",
          8481 => x"6720696e",
          8482 => x"74657272",
          8483 => x"75707473",
          8484 => x"0a000000",
          8485 => x"456e6162",
          8486 => x"6c696e67",
          8487 => x"20696e74",
          8488 => x"65727275",
          8489 => x"7074730a",
          8490 => x"00000000",
          8491 => x"44697361",
          8492 => x"626c6564",
          8493 => x"20756172",
          8494 => x"74206669",
          8495 => x"666f0a00",
          8496 => x"456e6162",
          8497 => x"6c696e67",
          8498 => x"20756172",
          8499 => x"74206669",
          8500 => x"666f0a00",
          8501 => x"45786563",
          8502 => x"7574696e",
          8503 => x"6720636f",
          8504 => x"64652040",
          8505 => x"20253038",
          8506 => x"78202e2e",
          8507 => x"2e0a0000",
          8508 => x"43616c6c",
          8509 => x"696e6720",
          8510 => x"636f6465",
          8511 => x"20402025",
          8512 => x"30387820",
          8513 => x"2e2e2e0a",
          8514 => x"00000000",
          8515 => x"43616c6c",
          8516 => x"20726574",
          8517 => x"75726e65",
          8518 => x"6420636f",
          8519 => x"64652028",
          8520 => x"2564292e",
          8521 => x"0a000000",
          8522 => x"52657374",
          8523 => x"61727469",
          8524 => x"6e672061",
          8525 => x"70706c69",
          8526 => x"63617469",
          8527 => x"6f6e2e2e",
          8528 => x"2e0a0000",
          8529 => x"436f6c64",
          8530 => x"20726562",
          8531 => x"6f6f7469",
          8532 => x"6e672e2e",
          8533 => x"2e0a0000",
          8534 => x"5a505500",
          8535 => x"62696e00",
          8536 => x"25643a5c",
          8537 => x"25735c25",
          8538 => x"732e2573",
          8539 => x"00000000",
          8540 => x"42616420",
          8541 => x"636f6d6d",
          8542 => x"616e642e",
          8543 => x"0a000000",
          8544 => x"52756e6e",
          8545 => x"696e672e",
          8546 => x"2e2e0a00",
          8547 => x"456e6162",
          8548 => x"6c696e67",
          8549 => x"20696e74",
          8550 => x"65727275",
          8551 => x"7074732e",
          8552 => x"2e2e0a00",
          8553 => x"00000000",
          8554 => x"00000000",
          8555 => x"00007fff",
          8556 => x"00000000",
          8557 => x"00007fff",
          8558 => x"00010000",
          8559 => x"00007fff",
          8560 => x"00000000",
          8561 => x"00000000",
          8562 => x"00007800",
          8563 => x"00000000",
          8564 => x"05f5e100",
          8565 => x"00010101",
          8566 => x"01010101",
          8567 => x"80010101",
          8568 => x"01000000",
          8569 => x"00000000",
          8570 => x"01000000",
          8571 => x"00005f20",
          8572 => x"00010100",
          8573 => x"00000000",
          8574 => x"00000000",
          8575 => x"00005f28",
          8576 => x"01020100",
          8577 => x"00000000",
          8578 => x"00000000",
          8579 => x"00005f30",
          8580 => x"00030100",
          8581 => x"00000000",
          8582 => x"00000000",
          8583 => x"00005f38",
          8584 => x"01040100",
          8585 => x"00000000",
          8586 => x"00000000",
          8587 => x"00005f40",
          8588 => x"000a0200",
          8589 => x"00000000",
          8590 => x"00000000",
          8591 => x"00005f48",
          8592 => x"000b0200",
          8593 => x"00000000",
          8594 => x"00000000",
          8595 => x"00005f50",
          8596 => x"000c0200",
          8597 => x"00000000",
          8598 => x"00000000",
          8599 => x"00005f58",
          8600 => x"000d0200",
          8601 => x"00000000",
          8602 => x"00000000",
          8603 => x"00005f60",
          8604 => x"000e0200",
          8605 => x"00000000",
          8606 => x"00000000",
          8607 => x"00005f68",
          8608 => x"000f0200",
          8609 => x"00000000",
          8610 => x"00000000",
          8611 => x"00005f70",
          8612 => x"01140300",
          8613 => x"00000000",
          8614 => x"00000000",
          8615 => x"00005f78",
          8616 => x"00170300",
          8617 => x"00000000",
          8618 => x"00000000",
          8619 => x"00005f80",
          8620 => x"00180300",
          8621 => x"00000000",
          8622 => x"00000000",
          8623 => x"00005f88",
          8624 => x"00190300",
          8625 => x"00000000",
          8626 => x"00000000",
          8627 => x"00005f90",
          8628 => x"001a0300",
          8629 => x"00000000",
          8630 => x"00000000",
          8631 => x"00005f98",
          8632 => x"001c0300",
          8633 => x"00000000",
          8634 => x"00000000",
          8635 => x"00005fa4",
          8636 => x"001d0300",
          8637 => x"00000000",
          8638 => x"00000000",
          8639 => x"00005fac",
          8640 => x"001e0300",
          8641 => x"00000000",
          8642 => x"00000000",
          8643 => x"00005fb4",
          8644 => x"00220300",
          8645 => x"00000000",
          8646 => x"00000000",
          8647 => x"00005fbc",
          8648 => x"00230300",
          8649 => x"00000000",
          8650 => x"00000000",
          8651 => x"00005fc4",
          8652 => x"00240300",
          8653 => x"00000000",
          8654 => x"00000000",
          8655 => x"00005fcc",
          8656 => x"001f0300",
          8657 => x"00000000",
          8658 => x"00000000",
          8659 => x"00005fd4",
          8660 => x"00200300",
          8661 => x"00000000",
          8662 => x"00000000",
          8663 => x"00005fdc",
          8664 => x"00210300",
          8665 => x"00000000",
          8666 => x"00000000",
          8667 => x"00005fe4",
          8668 => x"00150300",
          8669 => x"00000000",
          8670 => x"00000000",
          8671 => x"00005fec",
          8672 => x"00160300",
          8673 => x"00000000",
          8674 => x"00000000",
          8675 => x"00005ff4",
          8676 => x"001b0300",
          8677 => x"00000000",
          8678 => x"00000000",
          8679 => x"00005ffc",
          8680 => x"00250300",
          8681 => x"00000000",
          8682 => x"00000000",
          8683 => x"00006000",
          8684 => x"002d0300",
          8685 => x"00000000",
          8686 => x"00000000",
          8687 => x"00006008",
          8688 => x"002e0300",
          8689 => x"00000000",
          8690 => x"00000000",
          8691 => x"00006010",
          8692 => x"012b0300",
          8693 => x"00000000",
          8694 => x"00000000",
          8695 => x"00006018",
          8696 => x"01300300",
          8697 => x"00000000",
          8698 => x"00000000",
          8699 => x"00006020",
          8700 => x"002f0300",
          8701 => x"00000000",
          8702 => x"00000000",
          8703 => x"00006028",
          8704 => x"002c0300",
          8705 => x"00000000",
          8706 => x"00000000",
          8707 => x"00006030",
          8708 => x"00260300",
          8709 => x"00000000",
          8710 => x"00000000",
          8711 => x"00006034",
          8712 => x"00270300",
          8713 => x"00000000",
          8714 => x"00000000",
          8715 => x"0000603c",
          8716 => x"00280300",
          8717 => x"00000000",
          8718 => x"00000000",
          8719 => x"00006048",
          8720 => x"00290300",
          8721 => x"00000000",
          8722 => x"00000000",
          8723 => x"00006050",
          8724 => x"002a0300",
          8725 => x"00000000",
          8726 => x"00000000",
          8727 => x"00006058",
          8728 => x"003c0400",
          8729 => x"00000000",
          8730 => x"00000000",
          8731 => x"00006060",
          8732 => x"003d0400",
          8733 => x"00000000",
          8734 => x"00000000",
          8735 => x"00006068",
          8736 => x"003e0400",
          8737 => x"00000000",
          8738 => x"00000000",
          8739 => x"0000606c",
          8740 => x"003f0400",
          8741 => x"00000000",
          8742 => x"00000000",
          8743 => x"00006070",
          8744 => x"00400400",
          8745 => x"00000000",
          8746 => x"00000000",
          8747 => x"00006074",
          8748 => x"01500500",
          8749 => x"00000000",
          8750 => x"00000000",
          8751 => x"00006078",
          8752 => x"01510500",
          8753 => x"00000000",
          8754 => x"00000000",
          8755 => x"0000607c",
          8756 => x"00520500",
          8757 => x"00000000",
          8758 => x"00000000",
          8759 => x"00006080",
          8760 => x"00530500",
          8761 => x"00000000",
          8762 => x"00000000",
          8763 => x"00006084",
          8764 => x"01540500",
          8765 => x"00000000",
          8766 => x"00000000",
          8767 => x"00006088",
          8768 => x"01550500",
          8769 => x"00000000",
          8770 => x"00000000",
          8771 => x"0000608c",
          8772 => x"00640600",
          8773 => x"00000000",
          8774 => x"00000000",
          8775 => x"00006094",
          8776 => x"00650600",
          8777 => x"00000000",
          8778 => x"00000000",
          8779 => x"000060a0",
          8780 => x"01790700",
          8781 => x"00000000",
          8782 => x"00000000",
          8783 => x"000060a8",
          8784 => x"01780700",
          8785 => x"00000000",
          8786 => x"00000000",
          8787 => x"000060ac",
          8788 => x"01820800",
          8789 => x"00000000",
          8790 => x"00000000",
          8791 => x"000060b4",
          8792 => x"01830800",
          8793 => x"00000000",
          8794 => x"00000000",
          8795 => x"000060bc",
          8796 => x"00840800",
          8797 => x"00000000",
          8798 => x"00000000",
          8799 => x"000060c4",
          8800 => x"01850800",
          8801 => x"00000000",
          8802 => x"00000000",
          8803 => x"000060cc",
          8804 => x"00860800",
          8805 => x"00000000",
          8806 => x"00000000",
          8807 => x"000060d4",
          8808 => x"01870800",
          8809 => x"00000000",
          8810 => x"00000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_BIT_BRAM_32BIT_RANGE))));
        end if;
    end if;
end process;


end arch;

