-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b87ff",
             1 => x"f80d0b0b",
             2 => x"0b93b904",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90088880",
            10 => x"082d900c",
            11 => x"8c0c880c",
            12 => x"04000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b93",
            73 => x"9d040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b9380",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b82ae",
           162 => x"e4738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"93850400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b80c3",
           171 => x"f42d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b80c5",
           179 => x"e02d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d04ff",
           251 => x"ffffffff",
           252 => x"ffffffff",
           253 => x"ffffffff",
           254 => x"ffffffff",
           255 => x"ffffffff",
           256 => x"00000600",
           257 => x"ffffffff",
           258 => x"ffffffff",
           259 => x"ffffffff",
           260 => x"ffffffff",
           261 => x"ffffffff",
           262 => x"ffffffff",
           263 => x"ffffffff",
           264 => x"0b0b0b8c",
           265 => x"81040b0b",
           266 => x"0b8c8504",
           267 => x"0b0b0b8c",
           268 => x"95040b0b",
           269 => x"0b8ca404",
           270 => x"0b0b0b8c",
           271 => x"b3040b0b",
           272 => x"0b8cc204",
           273 => x"0b0b0b8c",
           274 => x"d1040b0b",
           275 => x"0b8ce004",
           276 => x"0b0b0b8c",
           277 => x"f0040b0b",
           278 => x"0b8d8004",
           279 => x"0b0b0b8d",
           280 => x"8f040b0b",
           281 => x"0b8d9e04",
           282 => x"0b0b0b8d",
           283 => x"ad040b0b",
           284 => x"0b8dbd04",
           285 => x"0b0b0b8d",
           286 => x"cd040b0b",
           287 => x"0b8ddd04",
           288 => x"0b0b0b8d",
           289 => x"ed040b0b",
           290 => x"0b8dfd04",
           291 => x"0b0b0b8e",
           292 => x"8d040b0b",
           293 => x"0b8e9d04",
           294 => x"0b0b0b8e",
           295 => x"ad040b0b",
           296 => x"0b8ebd04",
           297 => x"0b0b0b8e",
           298 => x"cd040b0b",
           299 => x"0b8edd04",
           300 => x"0b0b0b8e",
           301 => x"ed040b0b",
           302 => x"0b8efd04",
           303 => x"0b0b0b8f",
           304 => x"8d040b0b",
           305 => x"0b8f9d04",
           306 => x"0b0b0b8f",
           307 => x"ad040b0b",
           308 => x"0b8fbd04",
           309 => x"0b0b0b8f",
           310 => x"cd040b0b",
           311 => x"0b8fdd04",
           312 => x"0b0b0b8f",
           313 => x"ed040b0b",
           314 => x"0b8ffd04",
           315 => x"0b0b0b90",
           316 => x"8d040b0b",
           317 => x"0b909d04",
           318 => x"0b0b0b90",
           319 => x"ad040b0b",
           320 => x"0b90bd04",
           321 => x"0b0b0b90",
           322 => x"cd040b0b",
           323 => x"0b90dd04",
           324 => x"0b0b0b90",
           325 => x"ed040b0b",
           326 => x"0b90fd04",
           327 => x"0b0b0b91",
           328 => x"8d040b0b",
           329 => x"0b919d04",
           330 => x"0b0b0b91",
           331 => x"ad040b0b",
           332 => x"0b91bd04",
           333 => x"0b0b0b91",
           334 => x"cd040b0b",
           335 => x"0b91dd04",
           336 => x"0b0b0b91",
           337 => x"ed040b0b",
           338 => x"0b91fd04",
           339 => x"0b0b0b92",
           340 => x"8d040b0b",
           341 => x"0b929d04",
           342 => x"0b0b0b92",
           343 => x"ad040b0b",
           344 => x"0b92bd04",
           345 => x"0b0b0b92",
           346 => x"cd04ffff",
           347 => x"ffffffff",
           348 => x"ffffffff",
           349 => x"ffffffff",
           350 => x"ffffffff",
           351 => x"ffffffff",
           352 => x"ffffffff",
           353 => x"ffffffff",
           354 => x"ffffffff",
           355 => x"ffffffff",
           356 => x"ffffffff",
           357 => x"ffffffff",
           358 => x"ffffffff",
           359 => x"ffffffff",
           360 => x"ffffffff",
           361 => x"ffffffff",
           362 => x"ffffffff",
           363 => x"ffffffff",
           364 => x"ffffffff",
           365 => x"ffffffff",
           366 => x"ffffffff",
           367 => x"ffffffff",
           368 => x"ffffffff",
           369 => x"ffffffff",
           370 => x"ffffffff",
           371 => x"ffffffff",
           372 => x"ffffffff",
           373 => x"ffffffff",
           374 => x"ffffffff",
           375 => x"ffffffff",
           376 => x"ffffffff",
           377 => x"ffffffff",
           378 => x"ffffffff",
           379 => x"ffffffff",
           380 => x"ffffffff",
           381 => x"ffffffff",
           382 => x"ffffffff",
           383 => x"ffffffff",
           384 => x"04008c81",
           385 => x"0482d8d4",
           386 => x"0c80f9b3",
           387 => x"2d82d8d4",
           388 => x"08848090",
           389 => x"0482d8d4",
           390 => x"0cb3b22d",
           391 => x"82d8d408",
           392 => x"84809004",
           393 => x"82d8d40c",
           394 => x"afe32d82",
           395 => x"d8d40884",
           396 => x"80900482",
           397 => x"d8d40caf",
           398 => x"ad2d82d8",
           399 => x"d4088480",
           400 => x"900482d8",
           401 => x"d40c94ad",
           402 => x"2d82d8d4",
           403 => x"08848090",
           404 => x"0482d8d4",
           405 => x"0cb1c22d",
           406 => x"82d8d408",
           407 => x"84809004",
           408 => x"82d8d40c",
           409 => x"80cfcc2d",
           410 => x"82d8d408",
           411 => x"84809004",
           412 => x"82d8d40c",
           413 => x"80c9fb2d",
           414 => x"82d8d408",
           415 => x"84809004",
           416 => x"82d8d40c",
           417 => x"93d82d82",
           418 => x"d8d40884",
           419 => x"80900482",
           420 => x"d8d40c96",
           421 => x"c02d82d8",
           422 => x"d4088480",
           423 => x"900482d8",
           424 => x"d40c97cd",
           425 => x"2d82d8d4",
           426 => x"08848090",
           427 => x"0482d8d4",
           428 => x"0c80fcdd",
           429 => x"2d82d8d4",
           430 => x"08848090",
           431 => x"0482d8d4",
           432 => x"0c80fdbb",
           433 => x"2d82d8d4",
           434 => x"08848090",
           435 => x"0482d8d4",
           436 => x"0c80f4f8",
           437 => x"2d82d8d4",
           438 => x"08848090",
           439 => x"0482d8d4",
           440 => x"0c80f6ef",
           441 => x"2d82d8d4",
           442 => x"08848090",
           443 => x"0482d8d4",
           444 => x"0c80f8a2",
           445 => x"2d82d8d4",
           446 => x"08848090",
           447 => x"0482d8d4",
           448 => x"0c81eec7",
           449 => x"2d82d8d4",
           450 => x"08848090",
           451 => x"0482d8d4",
           452 => x"0c81fbc6",
           453 => x"2d82d8d4",
           454 => x"08848090",
           455 => x"0482d8d4",
           456 => x"0c81f3ac",
           457 => x"2d82d8d4",
           458 => x"08848090",
           459 => x"0482d8d4",
           460 => x"0c81f6ac",
           461 => x"2d82d8d4",
           462 => x"08848090",
           463 => x"0482d8d4",
           464 => x"0c828184",
           465 => x"2d82d8d4",
           466 => x"08848090",
           467 => x"0482d8d4",
           468 => x"0c8289ed",
           469 => x"2d82d8d4",
           470 => x"08848090",
           471 => x"0482d8d4",
           472 => x"0c81faa3",
           473 => x"2d82d8d4",
           474 => x"08848090",
           475 => x"0482d8d4",
           476 => x"0c8284a7",
           477 => x"2d82d8d4",
           478 => x"08848090",
           479 => x"0482d8d4",
           480 => x"0c8285c7",
           481 => x"2d82d8d4",
           482 => x"08848090",
           483 => x"0482d8d4",
           484 => x"0c8285e6",
           485 => x"2d82d8d4",
           486 => x"08848090",
           487 => x"0482d8d4",
           488 => x"0c828dda",
           489 => x"2d82d8d4",
           490 => x"08848090",
           491 => x"0482d8d4",
           492 => x"0c828bbc",
           493 => x"2d82d8d4",
           494 => x"08848090",
           495 => x"0482d8d4",
           496 => x"0c8290b6",
           497 => x"2d82d8d4",
           498 => x"08848090",
           499 => x"0482d8d4",
           500 => x"0c8286ec",
           501 => x"2d82d8d4",
           502 => x"08848090",
           503 => x"0482d8d4",
           504 => x"0c8293bb",
           505 => x"2d82d8d4",
           506 => x"08848090",
           507 => x"0482d8d4",
           508 => x"0c8294bc",
           509 => x"2d82d8d4",
           510 => x"08848090",
           511 => x"0482d8d4",
           512 => x"0c81fca6",
           513 => x"2d82d8d4",
           514 => x"08848090",
           515 => x"0482d8d4",
           516 => x"0c81fbff",
           517 => x"2d82d8d4",
           518 => x"08848090",
           519 => x"0482d8d4",
           520 => x"0c81fdaa",
           521 => x"2d82d8d4",
           522 => x"08848090",
           523 => x"0482d8d4",
           524 => x"0c8287c3",
           525 => x"2d82d8d4",
           526 => x"08848090",
           527 => x"0482d8d4",
           528 => x"0c8295ad",
           529 => x"2d82d8d4",
           530 => x"08848090",
           531 => x"0482d8d4",
           532 => x"0c8297b8",
           533 => x"2d82d8d4",
           534 => x"08848090",
           535 => x"0482d8d4",
           536 => x"0c829abf",
           537 => x"2d82d8d4",
           538 => x"08848090",
           539 => x"0482d8d4",
           540 => x"0c81ede6",
           541 => x"2d82d8d4",
           542 => x"08848090",
           543 => x"0482d8d4",
           544 => x"0c829dab",
           545 => x"2d82d8d4",
           546 => x"08848090",
           547 => x"0482d8d4",
           548 => x"0c82abe0",
           549 => x"2d82d8d4",
           550 => x"08848090",
           551 => x"0482d8d4",
           552 => x"0c82a9cc",
           553 => x"2d82d8d4",
           554 => x"08848090",
           555 => x"0482d8d4",
           556 => x"0c81adee",
           557 => x"2d82d8d4",
           558 => x"08848090",
           559 => x"0482d8d4",
           560 => x"0c81afd8",
           561 => x"2d82d8d4",
           562 => x"08848090",
           563 => x"0482d8d4",
           564 => x"0c81b1bc",
           565 => x"2d82d8d4",
           566 => x"08848090",
           567 => x"0482d8d4",
           568 => x"0c80f5a1",
           569 => x"2d82d8d4",
           570 => x"08848090",
           571 => x"0482d8d4",
           572 => x"0c80f6c5",
           573 => x"2d82d8d4",
           574 => x"08848090",
           575 => x"0482d8d4",
           576 => x"0c80faa8",
           577 => x"2d82d8d4",
           578 => x"08848090",
           579 => x"0482d8d4",
           580 => x"0c80d698",
           581 => x"2d82d8d4",
           582 => x"08848090",
           583 => x"0482d8d4",
           584 => x"0c81a882",
           585 => x"2d82d8d4",
           586 => x"08848090",
           587 => x"0482d8d4",
           588 => x"0c81a8aa",
           589 => x"2d82d8d4",
           590 => x"08848090",
           591 => x"0482d8d4",
           592 => x"0c81aca2",
           593 => x"2d82d8d4",
           594 => x"08848090",
           595 => x"0482d8d4",
           596 => x"0c81a4ec",
           597 => x"2d82d8d4",
           598 => x"08848090",
           599 => x"043c0400",
           600 => x"00101010",
           601 => x"10101010",
           602 => x"10101010",
           603 => x"10101010",
           604 => x"10101010",
           605 => x"10101010",
           606 => x"10101010",
           607 => x"10101010",
           608 => x"53510400",
           609 => x"007381ff",
           610 => x"06738306",
           611 => x"09810583",
           612 => x"05101010",
           613 => x"2b0772fc",
           614 => x"060c5151",
           615 => x"04727280",
           616 => x"728106ff",
           617 => x"05097206",
           618 => x"05711052",
           619 => x"720a100a",
           620 => x"5372ed38",
           621 => x"51515351",
           622 => x"0482d8c8",
           623 => x"7082f4b4",
           624 => x"278e3880",
           625 => x"71708405",
           626 => x"530c0b0b",
           627 => x"0b93bc04",
           628 => x"8c815180",
           629 => x"f3bb0400",
           630 => x"82d8d408",
           631 => x"0282d8d4",
           632 => x"0cfb3d0d",
           633 => x"82d8d408",
           634 => x"8c057082",
           635 => x"d8d408fc",
           636 => x"050c82d8",
           637 => x"d408fc05",
           638 => x"085482d8",
           639 => x"d4088805",
           640 => x"085382f4",
           641 => x"ac085254",
           642 => x"849a3f82",
           643 => x"d8c80870",
           644 => x"82d8d408",
           645 => x"f8050c82",
           646 => x"d8d408f8",
           647 => x"05087082",
           648 => x"d8c80c51",
           649 => x"54873d0d",
           650 => x"82d8d40c",
           651 => x"0482d8d4",
           652 => x"080282d8",
           653 => x"d40cfb3d",
           654 => x"0d82d8d4",
           655 => x"08900508",
           656 => x"85113370",
           657 => x"81327081",
           658 => x"06515151",
           659 => x"52718f38",
           660 => x"800b82d8",
           661 => x"d4088c05",
           662 => x"08258338",
           663 => x"8d39800b",
           664 => x"82d8d408",
           665 => x"f4050c81",
           666 => x"c43982d8",
           667 => x"d4088c05",
           668 => x"08ff0582",
           669 => x"d8d4088c",
           670 => x"050c800b",
           671 => x"82d8d408",
           672 => x"f8050c82",
           673 => x"d8d40888",
           674 => x"050882d8",
           675 => x"d408fc05",
           676 => x"0c82d8d4",
           677 => x"08f80508",
           678 => x"8a2e80f6",
           679 => x"38800b82",
           680 => x"d8d4088c",
           681 => x"05082580",
           682 => x"e93882d8",
           683 => x"d4089005",
           684 => x"0851a090",
           685 => x"3f82d8c8",
           686 => x"087082d8",
           687 => x"d408f805",
           688 => x"0c5282d8",
           689 => x"d408f805",
           690 => x"08ff2e09",
           691 => x"81068d38",
           692 => x"800b82d8",
           693 => x"d408f405",
           694 => x"0c80d239",
           695 => x"82d8d408",
           696 => x"fc050882",
           697 => x"d8d408f8",
           698 => x"05085353",
           699 => x"71733482",
           700 => x"d8d4088c",
           701 => x"0508ff05",
           702 => x"82d8d408",
           703 => x"8c050c82",
           704 => x"d8d408fc",
           705 => x"05088105",
           706 => x"82d8d408",
           707 => x"fc050cff",
           708 => x"803982d8",
           709 => x"d408fc05",
           710 => x"08528072",
           711 => x"3482d8d4",
           712 => x"08880508",
           713 => x"7082d8d4",
           714 => x"08f4050c",
           715 => x"5282d8d4",
           716 => x"08f40508",
           717 => x"82d8c80c",
           718 => x"873d0d82",
           719 => x"d8d40c04",
           720 => x"82d8d408",
           721 => x"0282d8d4",
           722 => x"0cf43d0d",
           723 => x"860b82d8",
           724 => x"d408e505",
           725 => x"3482d8d4",
           726 => x"08880508",
           727 => x"82d8d408",
           728 => x"e0050cfe",
           729 => x"0a0b82d8",
           730 => x"d408e805",
           731 => x"0c82d8d4",
           732 => x"08900570",
           733 => x"82d8d408",
           734 => x"fc050c82",
           735 => x"d8d408fc",
           736 => x"05085482",
           737 => x"d8d4088c",
           738 => x"05085382",
           739 => x"d8d408e0",
           740 => x"05705351",
           741 => x"54818d3f",
           742 => x"82d8c808",
           743 => x"7082d8d4",
           744 => x"08dc050c",
           745 => x"82d8d408",
           746 => x"ec050882",
           747 => x"d8d40888",
           748 => x"05080551",
           749 => x"54807434",
           750 => x"82d8d408",
           751 => x"dc050870",
           752 => x"82d8c80c",
           753 => x"548e3d0d",
           754 => x"82d8d40c",
           755 => x"0482d8d4",
           756 => x"080282d8",
           757 => x"d40cfb3d",
           758 => x"0d82d8d4",
           759 => x"08900570",
           760 => x"82d8d408",
           761 => x"fc050c82",
           762 => x"d8d408fc",
           763 => x"05085482",
           764 => x"d8d4088c",
           765 => x"05085382",
           766 => x"d8d40888",
           767 => x"05085254",
           768 => x"a33f82d8",
           769 => x"c8087082",
           770 => x"d8d408f8",
           771 => x"050c82d8",
           772 => x"d408f805",
           773 => x"087082d8",
           774 => x"c80c5154",
           775 => x"873d0d82",
           776 => x"d8d40c04",
           777 => x"82d8d408",
           778 => x"0282d8d4",
           779 => x"0ced3d0d",
           780 => x"800b82d8",
           781 => x"d408e405",
           782 => x"2382d8d4",
           783 => x"08880508",
           784 => x"53800b8c",
           785 => x"140c82d8",
           786 => x"d4088805",
           787 => x"08851133",
           788 => x"70812a70",
           789 => x"81327081",
           790 => x"06515151",
           791 => x"51537280",
           792 => x"2e8d38ff",
           793 => x"0b82d8d4",
           794 => x"08e0050c",
           795 => x"96ac3982",
           796 => x"d8d4088c",
           797 => x"05085372",
           798 => x"33537282",
           799 => x"d8d408f8",
           800 => x"05347281",
           801 => x"ff065372",
           802 => x"802e95fa",
           803 => x"3882d8d4",
           804 => x"088c0508",
           805 => x"810582d8",
           806 => x"d4088c05",
           807 => x"0c82d8d4",
           808 => x"08e40522",
           809 => x"70810651",
           810 => x"5372802e",
           811 => x"958b3882",
           812 => x"d8d408f8",
           813 => x"053353af",
           814 => x"732781fc",
           815 => x"3882d8d4",
           816 => x"08f80533",
           817 => x"5372b926",
           818 => x"81ee3882",
           819 => x"d8d408f8",
           820 => x"05335372",
           821 => x"b02e0981",
           822 => x"0680c538",
           823 => x"82d8d408",
           824 => x"e8053370",
           825 => x"982b7098",
           826 => x"2c515153",
           827 => x"72b23882",
           828 => x"d8d408e4",
           829 => x"05227083",
           830 => x"2a708132",
           831 => x"70810651",
           832 => x"51515372",
           833 => x"802e9938",
           834 => x"82d8d408",
           835 => x"e4052270",
           836 => x"82800751",
           837 => x"537282d8",
           838 => x"d408e405",
           839 => x"23fed039",
           840 => x"82d8d408",
           841 => x"e8053370",
           842 => x"982b7098",
           843 => x"2c707083",
           844 => x"2b721173",
           845 => x"11515151",
           846 => x"53515553",
           847 => x"7282d8d4",
           848 => x"08e80534",
           849 => x"82d8d408",
           850 => x"e8053354",
           851 => x"82d8d408",
           852 => x"f8053370",
           853 => x"15d01151",
           854 => x"51537282",
           855 => x"d8d408e8",
           856 => x"053482d8",
           857 => x"d408e805",
           858 => x"3370982b",
           859 => x"70982c51",
           860 => x"51537280",
           861 => x"258b3880",
           862 => x"ff0b82d8",
           863 => x"d408e805",
           864 => x"3482d8d4",
           865 => x"08e40522",
           866 => x"70832a70",
           867 => x"81065151",
           868 => x"5372fddb",
           869 => x"3882d8d4",
           870 => x"08e80533",
           871 => x"70882b70",
           872 => x"902b7090",
           873 => x"2c70882c",
           874 => x"51515151",
           875 => x"537282d8",
           876 => x"d408ec05",
           877 => x"23fdb839",
           878 => x"82d8d408",
           879 => x"e4052270",
           880 => x"832a7081",
           881 => x"06515153",
           882 => x"72802e9d",
           883 => x"3882d8d4",
           884 => x"08e80533",
           885 => x"70982b70",
           886 => x"982c5151",
           887 => x"53728a38",
           888 => x"810b82d8",
           889 => x"d408e805",
           890 => x"3482d8d4",
           891 => x"08f80533",
           892 => x"e01182d8",
           893 => x"d408c405",
           894 => x"0c5382d8",
           895 => x"d408c405",
           896 => x"0880d826",
           897 => x"92943882",
           898 => x"d8d408c4",
           899 => x"05087082",
           900 => x"2b82b0d4",
           901 => x"11700851",
           902 => x"51515372",
           903 => x"0482d8d4",
           904 => x"08e40522",
           905 => x"70900751",
           906 => x"537282d8",
           907 => x"d408e405",
           908 => x"2382d8d4",
           909 => x"08e40522",
           910 => x"70a00751",
           911 => x"537282d8",
           912 => x"d408e405",
           913 => x"23fca839",
           914 => x"82d8d408",
           915 => x"e4052270",
           916 => x"81800751",
           917 => x"537282d8",
           918 => x"d408e405",
           919 => x"23fc9039",
           920 => x"82d8d408",
           921 => x"e4052270",
           922 => x"80c00751",
           923 => x"537282d8",
           924 => x"d408e405",
           925 => x"23fbf839",
           926 => x"82d8d408",
           927 => x"e4052270",
           928 => x"88075153",
           929 => x"7282d8d4",
           930 => x"08e40523",
           931 => x"800b82d8",
           932 => x"d408e805",
           933 => x"34fbd839",
           934 => x"82d8d408",
           935 => x"e4052270",
           936 => x"84075153",
           937 => x"7282d8d4",
           938 => x"08e40523",
           939 => x"fbc139bf",
           940 => x"0b82d8d4",
           941 => x"08fc0534",
           942 => x"82d8d408",
           943 => x"ec0522ff",
           944 => x"11515372",
           945 => x"82d8d408",
           946 => x"ec052380",
           947 => x"e30b82d8",
           948 => x"d408f805",
           949 => x"348da839",
           950 => x"82d8d408",
           951 => x"90050882",
           952 => x"d8d40890",
           953 => x"05088405",
           954 => x"82d8d408",
           955 => x"90050c70",
           956 => x"08515372",
           957 => x"82d8d408",
           958 => x"fc053482",
           959 => x"d8d408ec",
           960 => x"0522ff11",
           961 => x"51537282",
           962 => x"d8d408ec",
           963 => x"05238cef",
           964 => x"3982d8d4",
           965 => x"08900508",
           966 => x"82d8d408",
           967 => x"90050884",
           968 => x"0582d8d4",
           969 => x"0890050c",
           970 => x"700882d8",
           971 => x"d408fc05",
           972 => x"0c82d8d4",
           973 => x"08e40522",
           974 => x"70832a70",
           975 => x"81065151",
           976 => x"51537280",
           977 => x"2eab3882",
           978 => x"d8d408e8",
           979 => x"05337098",
           980 => x"2b537298",
           981 => x"2c5382d8",
           982 => x"d408fc05",
           983 => x"085253a2",
           984 => x"d83f82d8",
           985 => x"c8085372",
           986 => x"82d8d408",
           987 => x"f4052399",
           988 => x"3982d8d4",
           989 => x"08fc0508",
           990 => x"519d8a3f",
           991 => x"82d8c808",
           992 => x"537282d8",
           993 => x"d408f405",
           994 => x"2382d8d4",
           995 => x"08ec0522",
           996 => x"5382d8d4",
           997 => x"08f40522",
           998 => x"73713154",
           999 => x"547282d8",
          1000 => x"d408ec05",
          1001 => x"238bd839",
          1002 => x"82d8d408",
          1003 => x"90050882",
          1004 => x"d8d40890",
          1005 => x"05088405",
          1006 => x"82d8d408",
          1007 => x"90050c70",
          1008 => x"0882d8d4",
          1009 => x"08fc050c",
          1010 => x"82d8d408",
          1011 => x"e4052270",
          1012 => x"832a7081",
          1013 => x"06515151",
          1014 => x"5372802e",
          1015 => x"ab3882d8",
          1016 => x"d408e805",
          1017 => x"3370982b",
          1018 => x"5372982c",
          1019 => x"5382d8d4",
          1020 => x"08fc0508",
          1021 => x"5253a1c1",
          1022 => x"3f82d8c8",
          1023 => x"08537282",
          1024 => x"d8d408f4",
          1025 => x"05239939",
          1026 => x"82d8d408",
          1027 => x"fc050851",
          1028 => x"9bf33f82",
          1029 => x"d8c80853",
          1030 => x"7282d8d4",
          1031 => x"08f40523",
          1032 => x"82d8d408",
          1033 => x"ec052253",
          1034 => x"82d8d408",
          1035 => x"f4052273",
          1036 => x"71315454",
          1037 => x"7282d8d4",
          1038 => x"08ec0523",
          1039 => x"8ac13982",
          1040 => x"d8d408e4",
          1041 => x"05227082",
          1042 => x"2a708106",
          1043 => x"51515372",
          1044 => x"802ea438",
          1045 => x"82d8d408",
          1046 => x"90050882",
          1047 => x"d8d40890",
          1048 => x"05088405",
          1049 => x"82d8d408",
          1050 => x"90050c70",
          1051 => x"0882d8d4",
          1052 => x"08dc050c",
          1053 => x"53a23982",
          1054 => x"d8d40890",
          1055 => x"050882d8",
          1056 => x"d4089005",
          1057 => x"08840582",
          1058 => x"d8d40890",
          1059 => x"050c7008",
          1060 => x"82d8d408",
          1061 => x"dc050c53",
          1062 => x"82d8d408",
          1063 => x"dc050882",
          1064 => x"d8d408fc",
          1065 => x"050c82d8",
          1066 => x"d408fc05",
          1067 => x"088025a4",
          1068 => x"3882d8d4",
          1069 => x"08e40522",
          1070 => x"70820751",
          1071 => x"537282d8",
          1072 => x"d408e405",
          1073 => x"2382d8d4",
          1074 => x"08fc0508",
          1075 => x"3082d8d4",
          1076 => x"08fc050c",
          1077 => x"82d8d408",
          1078 => x"e4052270",
          1079 => x"ffbf0651",
          1080 => x"537282d8",
          1081 => x"d408e405",
          1082 => x"2381af39",
          1083 => x"880b82d8",
          1084 => x"d408f405",
          1085 => x"23a93982",
          1086 => x"d8d408e4",
          1087 => x"05227080",
          1088 => x"c0075153",
          1089 => x"7282d8d4",
          1090 => x"08e40523",
          1091 => x"80f80b82",
          1092 => x"d8d408f8",
          1093 => x"0534900b",
          1094 => x"82d8d408",
          1095 => x"f4052382",
          1096 => x"d8d408e4",
          1097 => x"05227082",
          1098 => x"2a708106",
          1099 => x"51515372",
          1100 => x"802ea438",
          1101 => x"82d8d408",
          1102 => x"90050882",
          1103 => x"d8d40890",
          1104 => x"05088405",
          1105 => x"82d8d408",
          1106 => x"90050c70",
          1107 => x"0882d8d4",
          1108 => x"08d8050c",
          1109 => x"53a23982",
          1110 => x"d8d40890",
          1111 => x"050882d8",
          1112 => x"d4089005",
          1113 => x"08840582",
          1114 => x"d8d40890",
          1115 => x"050c7008",
          1116 => x"82d8d408",
          1117 => x"d8050c53",
          1118 => x"82d8d408",
          1119 => x"d8050882",
          1120 => x"d8d408fc",
          1121 => x"050c82d8",
          1122 => x"d408e405",
          1123 => x"2270cf06",
          1124 => x"51537282",
          1125 => x"d8d408e4",
          1126 => x"052382d8",
          1127 => x"d80b82d8",
          1128 => x"d408f005",
          1129 => x"0c82d8d4",
          1130 => x"08f00508",
          1131 => x"82d8d408",
          1132 => x"f4052282",
          1133 => x"d8d408fc",
          1134 => x"05087155",
          1135 => x"70545654",
          1136 => x"55a3f33f",
          1137 => x"82d8c808",
          1138 => x"53727534",
          1139 => x"82d8d408",
          1140 => x"f0050882",
          1141 => x"d8d408d4",
          1142 => x"050c82d8",
          1143 => x"d408f005",
          1144 => x"08703351",
          1145 => x"53897327",
          1146 => x"a43882d8",
          1147 => x"d408f005",
          1148 => x"08537233",
          1149 => x"5482d8d4",
          1150 => x"08f80533",
          1151 => x"7015df11",
          1152 => x"51515372",
          1153 => x"82d8d408",
          1154 => x"d0053497",
          1155 => x"3982d8d4",
          1156 => x"08f00508",
          1157 => x"537233b0",
          1158 => x"11515372",
          1159 => x"82d8d408",
          1160 => x"d0053482",
          1161 => x"d8d408d4",
          1162 => x"05085382",
          1163 => x"d8d408d0",
          1164 => x"05337334",
          1165 => x"82d8d408",
          1166 => x"f0050881",
          1167 => x"0582d8d4",
          1168 => x"08f0050c",
          1169 => x"82d8d408",
          1170 => x"f4052270",
          1171 => x"5382d8d4",
          1172 => x"08fc0508",
          1173 => x"5253a2ab",
          1174 => x"3f82d8c8",
          1175 => x"087082d8",
          1176 => x"d408fc05",
          1177 => x"0c5382d8",
          1178 => x"d408fc05",
          1179 => x"08802e84",
          1180 => x"38feb239",
          1181 => x"82d8d408",
          1182 => x"f0050882",
          1183 => x"d8d85455",
          1184 => x"72547470",
          1185 => x"75315153",
          1186 => x"7282d8d4",
          1187 => x"08fc0534",
          1188 => x"82d8d408",
          1189 => x"e4052270",
          1190 => x"b2065153",
          1191 => x"72802e94",
          1192 => x"3882d8d4",
          1193 => x"08ec0522",
          1194 => x"ff115153",
          1195 => x"7282d8d4",
          1196 => x"08ec0523",
          1197 => x"82d8d408",
          1198 => x"e4052270",
          1199 => x"862a7081",
          1200 => x"06515153",
          1201 => x"72802e80",
          1202 => x"e73882d8",
          1203 => x"d408ec05",
          1204 => x"2270902b",
          1205 => x"82d8d408",
          1206 => x"cc050c82",
          1207 => x"d8d408cc",
          1208 => x"0508902c",
          1209 => x"82d8d408",
          1210 => x"cc050c82",
          1211 => x"d8d408f4",
          1212 => x"05225153",
          1213 => x"72902e09",
          1214 => x"81069538",
          1215 => x"82d8d408",
          1216 => x"cc0508fe",
          1217 => x"05537282",
          1218 => x"d8d408c8",
          1219 => x"05239339",
          1220 => x"82d8d408",
          1221 => x"cc0508ff",
          1222 => x"05537282",
          1223 => x"d8d408c8",
          1224 => x"052382d8",
          1225 => x"d408c805",
          1226 => x"2282d8d4",
          1227 => x"08ec0523",
          1228 => x"82d8d408",
          1229 => x"e4052270",
          1230 => x"832a7081",
          1231 => x"06515153",
          1232 => x"72802e80",
          1233 => x"d03882d8",
          1234 => x"d408e805",
          1235 => x"3370982b",
          1236 => x"70982c82",
          1237 => x"d8d408fc",
          1238 => x"05335751",
          1239 => x"51537274",
          1240 => x"24973882",
          1241 => x"d8d408e4",
          1242 => x"052270f7",
          1243 => x"06515372",
          1244 => x"82d8d408",
          1245 => x"e405239d",
          1246 => x"3982d8d4",
          1247 => x"08e80533",
          1248 => x"5382d8d4",
          1249 => x"08fc0533",
          1250 => x"73713154",
          1251 => x"547282d8",
          1252 => x"d408e805",
          1253 => x"3482d8d4",
          1254 => x"08e40522",
          1255 => x"70832a70",
          1256 => x"81065151",
          1257 => x"5372802e",
          1258 => x"b13882d8",
          1259 => x"d408e805",
          1260 => x"3370882b",
          1261 => x"70902b70",
          1262 => x"902c7088",
          1263 => x"2c515151",
          1264 => x"51537254",
          1265 => x"82d8d408",
          1266 => x"ec052270",
          1267 => x"75315153",
          1268 => x"7282d8d4",
          1269 => x"08ec0523",
          1270 => x"af3982d8",
          1271 => x"d408fc05",
          1272 => x"3370882b",
          1273 => x"70902b70",
          1274 => x"902c7088",
          1275 => x"2c515151",
          1276 => x"51537254",
          1277 => x"82d8d408",
          1278 => x"ec052270",
          1279 => x"75315153",
          1280 => x"7282d8d4",
          1281 => x"08ec0523",
          1282 => x"82d8d408",
          1283 => x"e4052270",
          1284 => x"83800651",
          1285 => x"5372b038",
          1286 => x"82d8d408",
          1287 => x"ec0522ff",
          1288 => x"11545472",
          1289 => x"82d8d408",
          1290 => x"ec052373",
          1291 => x"902b7090",
          1292 => x"2c515380",
          1293 => x"73259038",
          1294 => x"82d8d408",
          1295 => x"88050852",
          1296 => x"a0518aee",
          1297 => x"3fd23982",
          1298 => x"d8d408e4",
          1299 => x"05227081",
          1300 => x"2a708106",
          1301 => x"51515372",
          1302 => x"802e9138",
          1303 => x"82d8d408",
          1304 => x"88050852",
          1305 => x"ad518aca",
          1306 => x"3f80c739",
          1307 => x"82d8d408",
          1308 => x"e4052270",
          1309 => x"842a7081",
          1310 => x"06515153",
          1311 => x"72802e90",
          1312 => x"3882d8d4",
          1313 => x"08880508",
          1314 => x"52ab518a",
          1315 => x"a53fa339",
          1316 => x"82d8d408",
          1317 => x"e4052270",
          1318 => x"852a7081",
          1319 => x"06515153",
          1320 => x"72802e8e",
          1321 => x"3882d8d4",
          1322 => x"08880508",
          1323 => x"52a0518a",
          1324 => x"813f82d8",
          1325 => x"d408e405",
          1326 => x"2270862a",
          1327 => x"70810651",
          1328 => x"51537280",
          1329 => x"2eb13882",
          1330 => x"d8d40888",
          1331 => x"050852b0",
          1332 => x"5189df3f",
          1333 => x"82d8d408",
          1334 => x"f4052253",
          1335 => x"72902e09",
          1336 => x"81069438",
          1337 => x"82d8d408",
          1338 => x"88050852",
          1339 => x"82d8d408",
          1340 => x"f8053351",
          1341 => x"89bc3f82",
          1342 => x"d8d408e4",
          1343 => x"05227088",
          1344 => x"2a708106",
          1345 => x"51515372",
          1346 => x"802eb038",
          1347 => x"82d8d408",
          1348 => x"ec0522ff",
          1349 => x"11545472",
          1350 => x"82d8d408",
          1351 => x"ec052373",
          1352 => x"902b7090",
          1353 => x"2c515380",
          1354 => x"73259038",
          1355 => x"82d8d408",
          1356 => x"88050852",
          1357 => x"b05188fa",
          1358 => x"3fd23982",
          1359 => x"d8d408e4",
          1360 => x"05227083",
          1361 => x"2a708106",
          1362 => x"51515372",
          1363 => x"802eb038",
          1364 => x"82d8d408",
          1365 => x"e80533ff",
          1366 => x"11545472",
          1367 => x"82d8d408",
          1368 => x"e8053473",
          1369 => x"982b7098",
          1370 => x"2c515380",
          1371 => x"73259038",
          1372 => x"82d8d408",
          1373 => x"88050852",
          1374 => x"b05188b6",
          1375 => x"3fd23982",
          1376 => x"d8d408e4",
          1377 => x"05227087",
          1378 => x"2a708106",
          1379 => x"51515372",
          1380 => x"b03882d8",
          1381 => x"d408ec05",
          1382 => x"22ff1154",
          1383 => x"547282d8",
          1384 => x"d408ec05",
          1385 => x"2373902b",
          1386 => x"70902c51",
          1387 => x"53807325",
          1388 => x"903882d8",
          1389 => x"d4088805",
          1390 => x"0852a051",
          1391 => x"87f43fd2",
          1392 => x"3982d8d4",
          1393 => x"08f80533",
          1394 => x"537280e3",
          1395 => x"2e098106",
          1396 => x"973882d8",
          1397 => x"d4088805",
          1398 => x"085282d8",
          1399 => x"d408fc05",
          1400 => x"335187ce",
          1401 => x"3f81ee39",
          1402 => x"82d8d408",
          1403 => x"f8053353",
          1404 => x"7280f32e",
          1405 => x"09810680",
          1406 => x"cb3882d8",
          1407 => x"d408f405",
          1408 => x"22ff1151",
          1409 => x"537282d8",
          1410 => x"d408f405",
          1411 => x"237283ff",
          1412 => x"ff065372",
          1413 => x"83ffff2e",
          1414 => x"81bb3882",
          1415 => x"d8d40888",
          1416 => x"05085282",
          1417 => x"d8d408fc",
          1418 => x"05087033",
          1419 => x"5282d8d4",
          1420 => x"08fc0508",
          1421 => x"810582d8",
          1422 => x"d408fc05",
          1423 => x"0c5386f2",
          1424 => x"3fffb739",
          1425 => x"82d8d408",
          1426 => x"f8053353",
          1427 => x"7280d32e",
          1428 => x"09810680",
          1429 => x"cb3882d8",
          1430 => x"d408f405",
          1431 => x"22ff1151",
          1432 => x"537282d8",
          1433 => x"d408f405",
          1434 => x"237283ff",
          1435 => x"ff065372",
          1436 => x"83ffff2e",
          1437 => x"80df3882",
          1438 => x"d8d40888",
          1439 => x"05085282",
          1440 => x"d8d408fc",
          1441 => x"05087033",
          1442 => x"525386a6",
          1443 => x"3f82d8d4",
          1444 => x"08fc0508",
          1445 => x"810582d8",
          1446 => x"d408fc05",
          1447 => x"0cffb739",
          1448 => x"82d8d408",
          1449 => x"f0050882",
          1450 => x"d8d82ea9",
          1451 => x"3882d8d4",
          1452 => x"08880508",
          1453 => x"5282d8d4",
          1454 => x"08f00508",
          1455 => x"ff0582d8",
          1456 => x"d408f005",
          1457 => x"0c82d8d4",
          1458 => x"08f00508",
          1459 => x"70335253",
          1460 => x"85e03fcc",
          1461 => x"3982d8d4",
          1462 => x"08e40522",
          1463 => x"70872a70",
          1464 => x"81065151",
          1465 => x"5372802e",
          1466 => x"80c33882",
          1467 => x"d8d408ec",
          1468 => x"0522ff11",
          1469 => x"54547282",
          1470 => x"d8d408ec",
          1471 => x"05237390",
          1472 => x"2b70902c",
          1473 => x"51538073",
          1474 => x"25a33882",
          1475 => x"d8d40888",
          1476 => x"050852a0",
          1477 => x"51859b3f",
          1478 => x"d23982d8",
          1479 => x"d4088805",
          1480 => x"085282d8",
          1481 => x"d408f805",
          1482 => x"33518586",
          1483 => x"3f800b82",
          1484 => x"d8d408e4",
          1485 => x"0523eab7",
          1486 => x"3982d8d4",
          1487 => x"08f80533",
          1488 => x"5372a52e",
          1489 => x"098106a8",
          1490 => x"38810b82",
          1491 => x"d8d408e4",
          1492 => x"0523800b",
          1493 => x"82d8d408",
          1494 => x"ec052380",
          1495 => x"0b82d8d4",
          1496 => x"08e80534",
          1497 => x"8a0b82d8",
          1498 => x"d408f405",
          1499 => x"23ea8039",
          1500 => x"82d8d408",
          1501 => x"88050852",
          1502 => x"82d8d408",
          1503 => x"f8053351",
          1504 => x"84b03fe9",
          1505 => x"ea3982d8",
          1506 => x"d4088805",
          1507 => x"088c1108",
          1508 => x"7082d8d4",
          1509 => x"08e0050c",
          1510 => x"515382d8",
          1511 => x"d408e005",
          1512 => x"0882d8c8",
          1513 => x"0c953d0d",
          1514 => x"82d8d40c",
          1515 => x"0482d8d4",
          1516 => x"080282d8",
          1517 => x"d40cfd3d",
          1518 => x"0d82f4a8",
          1519 => x"085382d8",
          1520 => x"d4088c05",
          1521 => x"085282d8",
          1522 => x"d4088805",
          1523 => x"0851e4dd",
          1524 => x"3f82d8c8",
          1525 => x"087082d8",
          1526 => x"c80c5485",
          1527 => x"3d0d82d8",
          1528 => x"d40c0482",
          1529 => x"d8d40802",
          1530 => x"82d8d40c",
          1531 => x"fb3d0d80",
          1532 => x"0b82d8d4",
          1533 => x"08f8050c",
          1534 => x"82f4ac08",
          1535 => x"85113370",
          1536 => x"812a7081",
          1537 => x"32708106",
          1538 => x"51515151",
          1539 => x"5372802e",
          1540 => x"8d38ff0b",
          1541 => x"82d8d408",
          1542 => x"f4050c81",
          1543 => x"923982d8",
          1544 => x"d4088805",
          1545 => x"08537233",
          1546 => x"82d8d408",
          1547 => x"88050881",
          1548 => x"0582d8d4",
          1549 => x"0888050c",
          1550 => x"537282d8",
          1551 => x"d408fc05",
          1552 => x"347281ff",
          1553 => x"06537280",
          1554 => x"2eb03882",
          1555 => x"f4ac0882",
          1556 => x"f4ac0853",
          1557 => x"82d8d408",
          1558 => x"fc053352",
          1559 => x"90110851",
          1560 => x"53722d82",
          1561 => x"d8c80853",
          1562 => x"72802eff",
          1563 => x"b138ff0b",
          1564 => x"82d8d408",
          1565 => x"f8050cff",
          1566 => x"a53982f4",
          1567 => x"ac0882f4",
          1568 => x"ac085353",
          1569 => x"8a519013",
          1570 => x"0853722d",
          1571 => x"82d8c808",
          1572 => x"5372802e",
          1573 => x"8a38ff0b",
          1574 => x"82d8d408",
          1575 => x"f8050c82",
          1576 => x"d8d408f8",
          1577 => x"05087082",
          1578 => x"d8d408f4",
          1579 => x"050c5382",
          1580 => x"d8d408f4",
          1581 => x"050882d8",
          1582 => x"c80c873d",
          1583 => x"0d82d8d4",
          1584 => x"0c0482d8",
          1585 => x"d4080282",
          1586 => x"d8d40cfb",
          1587 => x"3d0d800b",
          1588 => x"82d8d408",
          1589 => x"f8050c82",
          1590 => x"d8d4088c",
          1591 => x"05088511",
          1592 => x"3370812a",
          1593 => x"70813270",
          1594 => x"81065151",
          1595 => x"51515372",
          1596 => x"802e8d38",
          1597 => x"ff0b82d8",
          1598 => x"d408f405",
          1599 => x"0c80f339",
          1600 => x"82d8d408",
          1601 => x"88050853",
          1602 => x"723382d8",
          1603 => x"d4088805",
          1604 => x"08810582",
          1605 => x"d8d40888",
          1606 => x"050c5372",
          1607 => x"82d8d408",
          1608 => x"fc053472",
          1609 => x"81ff0653",
          1610 => x"72802eb6",
          1611 => x"3882d8d4",
          1612 => x"088c0508",
          1613 => x"82d8d408",
          1614 => x"8c050853",
          1615 => x"82d8d408",
          1616 => x"fc053352",
          1617 => x"90110851",
          1618 => x"53722d82",
          1619 => x"d8c80853",
          1620 => x"72802eff",
          1621 => x"ab38ff0b",
          1622 => x"82d8d408",
          1623 => x"f8050cff",
          1624 => x"9f3982d8",
          1625 => x"d408f805",
          1626 => x"087082d8",
          1627 => x"d408f405",
          1628 => x"0c5382d8",
          1629 => x"d408f405",
          1630 => x"0882d8c8",
          1631 => x"0c873d0d",
          1632 => x"82d8d40c",
          1633 => x"0482d8d4",
          1634 => x"080282d8",
          1635 => x"d40cfe3d",
          1636 => x"0d82f4ac",
          1637 => x"085282d8",
          1638 => x"d4088805",
          1639 => x"0851933f",
          1640 => x"82d8c808",
          1641 => x"7082d8c8",
          1642 => x"0c53843d",
          1643 => x"0d82d8d4",
          1644 => x"0c0482d8",
          1645 => x"d4080282",
          1646 => x"d8d40cfb",
          1647 => x"3d0d82d8",
          1648 => x"d4088c05",
          1649 => x"08851133",
          1650 => x"70812a70",
          1651 => x"81327081",
          1652 => x"06515151",
          1653 => x"51537280",
          1654 => x"2e8d38ff",
          1655 => x"0b82d8d4",
          1656 => x"08fc050c",
          1657 => x"81cb3982",
          1658 => x"d8d4088c",
          1659 => x"05088511",
          1660 => x"3370822a",
          1661 => x"70810651",
          1662 => x"51515372",
          1663 => x"802e80db",
          1664 => x"3882d8d4",
          1665 => x"088c0508",
          1666 => x"82d8d408",
          1667 => x"8c050854",
          1668 => x"548c1408",
          1669 => x"88140825",
          1670 => x"9f3882d8",
          1671 => x"d4088c05",
          1672 => x"08700870",
          1673 => x"82d8d408",
          1674 => x"88050852",
          1675 => x"57545472",
          1676 => x"75347308",
          1677 => x"8105740c",
          1678 => x"82d8d408",
          1679 => x"8c05088c",
          1680 => x"11088105",
          1681 => x"8c120c82",
          1682 => x"d8d40888",
          1683 => x"05087082",
          1684 => x"d8d408fc",
          1685 => x"050c5153",
          1686 => x"80d73982",
          1687 => x"d8d4088c",
          1688 => x"050882d8",
          1689 => x"d4088c05",
          1690 => x"085382d8",
          1691 => x"d4088805",
          1692 => x"087081ff",
          1693 => x"06539012",
          1694 => x"08515454",
          1695 => x"722d82d8",
          1696 => x"c8085372",
          1697 => x"a33882d8",
          1698 => x"d4088c05",
          1699 => x"088c1108",
          1700 => x"81058c12",
          1701 => x"0c82d8d4",
          1702 => x"08880508",
          1703 => x"7082d8d4",
          1704 => x"08fc050c",
          1705 => x"51538a39",
          1706 => x"ff0b82d8",
          1707 => x"d408fc05",
          1708 => x"0c82d8d4",
          1709 => x"08fc0508",
          1710 => x"82d8c80c",
          1711 => x"873d0d82",
          1712 => x"d8d40c04",
          1713 => x"82d8d408",
          1714 => x"0282d8d4",
          1715 => x"0cf93d0d",
          1716 => x"82d8d408",
          1717 => x"88050885",
          1718 => x"11337081",
          1719 => x"32708106",
          1720 => x"51515152",
          1721 => x"71802e8d",
          1722 => x"38ff0b82",
          1723 => x"d8d408f8",
          1724 => x"050c8394",
          1725 => x"3982d8d4",
          1726 => x"08880508",
          1727 => x"85113370",
          1728 => x"862a7081",
          1729 => x"06515151",
          1730 => x"5271802e",
          1731 => x"80c53882",
          1732 => x"d8d40888",
          1733 => x"050882d8",
          1734 => x"d4088805",
          1735 => x"08535385",
          1736 => x"123370ff",
          1737 => x"bf065152",
          1738 => x"71851434",
          1739 => x"82d8d408",
          1740 => x"8805088c",
          1741 => x"11088105",
          1742 => x"8c120c82",
          1743 => x"d8d40888",
          1744 => x"05088411",
          1745 => x"337082d8",
          1746 => x"d408f805",
          1747 => x"0c515152",
          1748 => x"82b63982",
          1749 => x"d8d40888",
          1750 => x"05088511",
          1751 => x"3370822a",
          1752 => x"70810651",
          1753 => x"51515271",
          1754 => x"802e80d7",
          1755 => x"3882d8d4",
          1756 => x"08880508",
          1757 => x"70087033",
          1758 => x"82d8d408",
          1759 => x"fc050c51",
          1760 => x"5282d8d4",
          1761 => x"08fc0508",
          1762 => x"a93882d8",
          1763 => x"d4088805",
          1764 => x"0882d8d4",
          1765 => x"08880508",
          1766 => x"53538512",
          1767 => x"3370a007",
          1768 => x"51527185",
          1769 => x"1434ff0b",
          1770 => x"82d8d408",
          1771 => x"f8050c81",
          1772 => x"d73982d8",
          1773 => x"d4088805",
          1774 => x"08700881",
          1775 => x"05710c52",
          1776 => x"81a13982",
          1777 => x"d8d40888",
          1778 => x"050882d8",
          1779 => x"d4088805",
          1780 => x"08529411",
          1781 => x"08515271",
          1782 => x"2d82d8c8",
          1783 => x"087082d8",
          1784 => x"d408fc05",
          1785 => x"0c5282d8",
          1786 => x"d408fc05",
          1787 => x"08802580",
          1788 => x"f23882d8",
          1789 => x"d4088805",
          1790 => x"0882d8d4",
          1791 => x"08f4050c",
          1792 => x"82d8d408",
          1793 => x"88050885",
          1794 => x"113382d8",
          1795 => x"d408f005",
          1796 => x"0c5282d8",
          1797 => x"d408fc05",
          1798 => x"08ff2e09",
          1799 => x"81069538",
          1800 => x"82d8d408",
          1801 => x"f0050890",
          1802 => x"07527182",
          1803 => x"d8d408ec",
          1804 => x"05349339",
          1805 => x"82d8d408",
          1806 => x"f00508a0",
          1807 => x"07527182",
          1808 => x"d8d408ec",
          1809 => x"053482d8",
          1810 => x"d408f405",
          1811 => x"085282d8",
          1812 => x"d408ec05",
          1813 => x"33851334",
          1814 => x"ff0b82d8",
          1815 => x"d408f805",
          1816 => x"0ca63982",
          1817 => x"d8d40888",
          1818 => x"05088c11",
          1819 => x"0881058c",
          1820 => x"120c82d8",
          1821 => x"d408fc05",
          1822 => x"087081ff",
          1823 => x"067082d8",
          1824 => x"d408f805",
          1825 => x"0c515152",
          1826 => x"82d8d408",
          1827 => x"f8050882",
          1828 => x"d8c80c89",
          1829 => x"3d0d82d8",
          1830 => x"d40c0482",
          1831 => x"d8d40802",
          1832 => x"82d8d40c",
          1833 => x"fd3d0d82",
          1834 => x"d8d40888",
          1835 => x"050882d8",
          1836 => x"d408fc05",
          1837 => x"0c82d8d4",
          1838 => x"088c0508",
          1839 => x"82d8d408",
          1840 => x"f8050c82",
          1841 => x"d8d40890",
          1842 => x"0508802e",
          1843 => x"82a23882",
          1844 => x"d8d408f8",
          1845 => x"050882d8",
          1846 => x"d408fc05",
          1847 => x"082681ac",
          1848 => x"3882d8d4",
          1849 => x"08f80508",
          1850 => x"82d8d408",
          1851 => x"90050805",
          1852 => x"5182d8d4",
          1853 => x"08fc0508",
          1854 => x"71278190",
          1855 => x"3882d8d4",
          1856 => x"08fc0508",
          1857 => x"82d8d408",
          1858 => x"90050805",
          1859 => x"82d8d408",
          1860 => x"fc050c82",
          1861 => x"d8d408f8",
          1862 => x"050882d8",
          1863 => x"d4089005",
          1864 => x"080582d8",
          1865 => x"d408f805",
          1866 => x"0c82d8d4",
          1867 => x"08900508",
          1868 => x"810582d8",
          1869 => x"d4089005",
          1870 => x"0c82d8d4",
          1871 => x"08900508",
          1872 => x"ff0582d8",
          1873 => x"d4089005",
          1874 => x"0c82d8d4",
          1875 => x"08900508",
          1876 => x"802e819c",
          1877 => x"3882d8d4",
          1878 => x"08fc0508",
          1879 => x"ff0582d8",
          1880 => x"d408fc05",
          1881 => x"0c82d8d4",
          1882 => x"08f80508",
          1883 => x"ff0582d8",
          1884 => x"d408f805",
          1885 => x"0c82d8d4",
          1886 => x"08fc0508",
          1887 => x"82d8d408",
          1888 => x"f8050853",
          1889 => x"51713371",
          1890 => x"34ffae39",
          1891 => x"82d8d408",
          1892 => x"90050881",
          1893 => x"0582d8d4",
          1894 => x"0890050c",
          1895 => x"82d8d408",
          1896 => x"900508ff",
          1897 => x"0582d8d4",
          1898 => x"0890050c",
          1899 => x"82d8d408",
          1900 => x"90050880",
          1901 => x"2eba3882",
          1902 => x"d8d408f8",
          1903 => x"05085170",
          1904 => x"3382d8d4",
          1905 => x"08f80508",
          1906 => x"810582d8",
          1907 => x"d408f805",
          1908 => x"0c82d8d4",
          1909 => x"08fc0508",
          1910 => x"52527171",
          1911 => x"3482d8d4",
          1912 => x"08fc0508",
          1913 => x"810582d8",
          1914 => x"d408fc05",
          1915 => x"0cffad39",
          1916 => x"82d8d408",
          1917 => x"88050870",
          1918 => x"82d8c80c",
          1919 => x"51853d0d",
          1920 => x"82d8d40c",
          1921 => x"0482d8d4",
          1922 => x"080282d8",
          1923 => x"d40cfe3d",
          1924 => x"0d82d8d4",
          1925 => x"08880508",
          1926 => x"82d8d408",
          1927 => x"fc050c82",
          1928 => x"d8d408fc",
          1929 => x"05085271",
          1930 => x"3382d8d4",
          1931 => x"08fc0508",
          1932 => x"810582d8",
          1933 => x"d408fc05",
          1934 => x"0c7081ff",
          1935 => x"06515170",
          1936 => x"802e8338",
          1937 => x"da3982d8",
          1938 => x"d408fc05",
          1939 => x"08ff0582",
          1940 => x"d8d408fc",
          1941 => x"050c82d8",
          1942 => x"d408fc05",
          1943 => x"0882d8d4",
          1944 => x"08880508",
          1945 => x"317082d8",
          1946 => x"c80c5184",
          1947 => x"3d0d82d8",
          1948 => x"d40c0482",
          1949 => x"d8d40802",
          1950 => x"82d8d40c",
          1951 => x"fe3d0d82",
          1952 => x"d8d40888",
          1953 => x"050882d8",
          1954 => x"d408fc05",
          1955 => x"0c82d8d4",
          1956 => x"088c0508",
          1957 => x"52713382",
          1958 => x"d8d4088c",
          1959 => x"05088105",
          1960 => x"82d8d408",
          1961 => x"8c050c82",
          1962 => x"d8d408fc",
          1963 => x"05085351",
          1964 => x"70723482",
          1965 => x"d8d408fc",
          1966 => x"05088105",
          1967 => x"82d8d408",
          1968 => x"fc050c70",
          1969 => x"81ff0651",
          1970 => x"70802e84",
          1971 => x"38ffbe39",
          1972 => x"82d8d408",
          1973 => x"88050870",
          1974 => x"82d8c80c",
          1975 => x"51843d0d",
          1976 => x"82d8d40c",
          1977 => x"0482d8d4",
          1978 => x"080282d8",
          1979 => x"d40cfd3d",
          1980 => x"0d82d8d4",
          1981 => x"08880508",
          1982 => x"82d8d408",
          1983 => x"fc050c82",
          1984 => x"d8d4088c",
          1985 => x"050882d8",
          1986 => x"d408f805",
          1987 => x"0c82d8d4",
          1988 => x"08900508",
          1989 => x"802e80e5",
          1990 => x"3882d8d4",
          1991 => x"08900508",
          1992 => x"810582d8",
          1993 => x"d4089005",
          1994 => x"0c82d8d4",
          1995 => x"08900508",
          1996 => x"ff0582d8",
          1997 => x"d4089005",
          1998 => x"0c82d8d4",
          1999 => x"08900508",
          2000 => x"802eba38",
          2001 => x"82d8d408",
          2002 => x"f8050851",
          2003 => x"703382d8",
          2004 => x"d408f805",
          2005 => x"08810582",
          2006 => x"d8d408f8",
          2007 => x"050c82d8",
          2008 => x"d408fc05",
          2009 => x"08525271",
          2010 => x"713482d8",
          2011 => x"d408fc05",
          2012 => x"08810582",
          2013 => x"d8d408fc",
          2014 => x"050cffad",
          2015 => x"3982d8d4",
          2016 => x"08880508",
          2017 => x"7082d8c8",
          2018 => x"0c51853d",
          2019 => x"0d82d8d4",
          2020 => x"0c0482d8",
          2021 => x"d4080282",
          2022 => x"d8d40cfd",
          2023 => x"3d0d82d8",
          2024 => x"d4089005",
          2025 => x"08802e81",
          2026 => x"f43882d8",
          2027 => x"d4088c05",
          2028 => x"08527133",
          2029 => x"82d8d408",
          2030 => x"8c050881",
          2031 => x"0582d8d4",
          2032 => x"088c050c",
          2033 => x"82d8d408",
          2034 => x"88050870",
          2035 => x"337281ff",
          2036 => x"06535454",
          2037 => x"5171712e",
          2038 => x"843880ce",
          2039 => x"3982d8d4",
          2040 => x"08880508",
          2041 => x"52713382",
          2042 => x"d8d40888",
          2043 => x"05088105",
          2044 => x"82d8d408",
          2045 => x"88050c70",
          2046 => x"81ff0651",
          2047 => x"51708d38",
          2048 => x"800b82d8",
          2049 => x"d408fc05",
          2050 => x"0c819b39",
          2051 => x"82d8d408",
          2052 => x"900508ff",
          2053 => x"0582d8d4",
          2054 => x"0890050c",
          2055 => x"82d8d408",
          2056 => x"90050880",
          2057 => x"2e8438ff",
          2058 => x"813982d8",
          2059 => x"d4089005",
          2060 => x"08802e80",
          2061 => x"e83882d8",
          2062 => x"d4088805",
          2063 => x"08703352",
          2064 => x"53708d38",
          2065 => x"ff0b82d8",
          2066 => x"d408fc05",
          2067 => x"0c80d739",
          2068 => x"82d8d408",
          2069 => x"8c0508ff",
          2070 => x"0582d8d4",
          2071 => x"088c050c",
          2072 => x"82d8d408",
          2073 => x"8c050870",
          2074 => x"33525270",
          2075 => x"8c38810b",
          2076 => x"82d8d408",
          2077 => x"fc050cae",
          2078 => x"3982d8d4",
          2079 => x"08880508",
          2080 => x"703382d8",
          2081 => x"d4088c05",
          2082 => x"08703372",
          2083 => x"71317082",
          2084 => x"d8d408fc",
          2085 => x"050c5355",
          2086 => x"5252538a",
          2087 => x"39800b82",
          2088 => x"d8d408fc",
          2089 => x"050c82d8",
          2090 => x"d408fc05",
          2091 => x"0882d8c8",
          2092 => x"0c853d0d",
          2093 => x"82d8d40c",
          2094 => x"0482d8d4",
          2095 => x"080282d8",
          2096 => x"d40cfd3d",
          2097 => x"0d82d8d4",
          2098 => x"08880508",
          2099 => x"82d8d408",
          2100 => x"f8050c82",
          2101 => x"d8d4088c",
          2102 => x"05088d38",
          2103 => x"800b82d8",
          2104 => x"d408fc05",
          2105 => x"0c80ec39",
          2106 => x"82d8d408",
          2107 => x"f8050852",
          2108 => x"713382d8",
          2109 => x"d408f805",
          2110 => x"08810582",
          2111 => x"d8d408f8",
          2112 => x"050c7081",
          2113 => x"ff065151",
          2114 => x"70802e9f",
          2115 => x"3882d8d4",
          2116 => x"088c0508",
          2117 => x"ff0582d8",
          2118 => x"d4088c05",
          2119 => x"0c82d8d4",
          2120 => x"088c0508",
          2121 => x"ff2e8438",
          2122 => x"ffbe3982",
          2123 => x"d8d408f8",
          2124 => x"0508ff05",
          2125 => x"82d8d408",
          2126 => x"f8050c82",
          2127 => x"d8d408f8",
          2128 => x"050882d8",
          2129 => x"d4088805",
          2130 => x"08317082",
          2131 => x"d8d408fc",
          2132 => x"050c5182",
          2133 => x"d8d408fc",
          2134 => x"050882d8",
          2135 => x"c80c853d",
          2136 => x"0d82d8d4",
          2137 => x"0c0482d8",
          2138 => x"d4080282",
          2139 => x"d8d40cfe",
          2140 => x"3d0d82d8",
          2141 => x"d4088805",
          2142 => x"0882d8d4",
          2143 => x"08fc050c",
          2144 => x"82d8d408",
          2145 => x"90050880",
          2146 => x"2e80d438",
          2147 => x"82d8d408",
          2148 => x"90050881",
          2149 => x"0582d8d4",
          2150 => x"0890050c",
          2151 => x"82d8d408",
          2152 => x"900508ff",
          2153 => x"0582d8d4",
          2154 => x"0890050c",
          2155 => x"82d8d408",
          2156 => x"90050880",
          2157 => x"2ea93882",
          2158 => x"d8d4088c",
          2159 => x"05085170",
          2160 => x"82d8d408",
          2161 => x"fc050852",
          2162 => x"52717134",
          2163 => x"82d8d408",
          2164 => x"fc050881",
          2165 => x"0582d8d4",
          2166 => x"08fc050c",
          2167 => x"ffbe3982",
          2168 => x"d8d40888",
          2169 => x"05087082",
          2170 => x"d8c80c51",
          2171 => x"843d0d82",
          2172 => x"d8d40c04",
          2173 => x"82d8d408",
          2174 => x"0282d8d4",
          2175 => x"0cf93d0d",
          2176 => x"800b82d8",
          2177 => x"d408fc05",
          2178 => x"0c82d8d4",
          2179 => x"08880508",
          2180 => x"8025b938",
          2181 => x"82d8d408",
          2182 => x"88050830",
          2183 => x"82d8d408",
          2184 => x"88050c80",
          2185 => x"0b82d8d4",
          2186 => x"08f4050c",
          2187 => x"82d8d408",
          2188 => x"fc05088a",
          2189 => x"38810b82",
          2190 => x"d8d408f4",
          2191 => x"050c82d8",
          2192 => x"d408f405",
          2193 => x"0882d8d4",
          2194 => x"08fc050c",
          2195 => x"82d8d408",
          2196 => x"8c050880",
          2197 => x"25b93882",
          2198 => x"d8d4088c",
          2199 => x"05083082",
          2200 => x"d8d4088c",
          2201 => x"050c800b",
          2202 => x"82d8d408",
          2203 => x"f0050c82",
          2204 => x"d8d408fc",
          2205 => x"05088a38",
          2206 => x"810b82d8",
          2207 => x"d408f005",
          2208 => x"0c82d8d4",
          2209 => x"08f00508",
          2210 => x"82d8d408",
          2211 => x"fc050c80",
          2212 => x"5382d8d4",
          2213 => x"088c0508",
          2214 => x"5282d8d4",
          2215 => x"08880508",
          2216 => x"5182c53f",
          2217 => x"82d8c808",
          2218 => x"7082d8d4",
          2219 => x"08f8050c",
          2220 => x"5482d8d4",
          2221 => x"08fc0508",
          2222 => x"802e9038",
          2223 => x"82d8d408",
          2224 => x"f8050830",
          2225 => x"82d8d408",
          2226 => x"f8050c82",
          2227 => x"d8d408f8",
          2228 => x"05087082",
          2229 => x"d8c80c54",
          2230 => x"893d0d82",
          2231 => x"d8d40c04",
          2232 => x"82d8d408",
          2233 => x"0282d8d4",
          2234 => x"0cfb3d0d",
          2235 => x"800b82d8",
          2236 => x"d408fc05",
          2237 => x"0c82d8d4",
          2238 => x"08880508",
          2239 => x"80259938",
          2240 => x"82d8d408",
          2241 => x"88050830",
          2242 => x"82d8d408",
          2243 => x"88050c81",
          2244 => x"0b82d8d4",
          2245 => x"08fc050c",
          2246 => x"82d8d408",
          2247 => x"8c050880",
          2248 => x"25903882",
          2249 => x"d8d4088c",
          2250 => x"05083082",
          2251 => x"d8d4088c",
          2252 => x"050c8153",
          2253 => x"82d8d408",
          2254 => x"8c050852",
          2255 => x"82d8d408",
          2256 => x"88050851",
          2257 => x"81a23f82",
          2258 => x"d8c80870",
          2259 => x"82d8d408",
          2260 => x"f8050c54",
          2261 => x"82d8d408",
          2262 => x"fc050880",
          2263 => x"2e903882",
          2264 => x"d8d408f8",
          2265 => x"05083082",
          2266 => x"d8d408f8",
          2267 => x"050c82d8",
          2268 => x"d408f805",
          2269 => x"087082d8",
          2270 => x"c80c5487",
          2271 => x"3d0d82d8",
          2272 => x"d40c0482",
          2273 => x"d8d40802",
          2274 => x"82d8d40c",
          2275 => x"fd3d0d80",
          2276 => x"5382d8d4",
          2277 => x"088c0508",
          2278 => x"5282d8d4",
          2279 => x"08880508",
          2280 => x"5180c53f",
          2281 => x"82d8c808",
          2282 => x"7082d8c8",
          2283 => x"0c54853d",
          2284 => x"0d82d8d4",
          2285 => x"0c0482d8",
          2286 => x"d4080282",
          2287 => x"d8d40cfd",
          2288 => x"3d0d8153",
          2289 => x"82d8d408",
          2290 => x"8c050852",
          2291 => x"82d8d408",
          2292 => x"88050851",
          2293 => x"933f82d8",
          2294 => x"c8087082",
          2295 => x"d8c80c54",
          2296 => x"853d0d82",
          2297 => x"d8d40c04",
          2298 => x"82d8d408",
          2299 => x"0282d8d4",
          2300 => x"0cfd3d0d",
          2301 => x"810b82d8",
          2302 => x"d408fc05",
          2303 => x"0c800b82",
          2304 => x"d8d408f8",
          2305 => x"050c82d8",
          2306 => x"d4088c05",
          2307 => x"0882d8d4",
          2308 => x"08880508",
          2309 => x"27b93882",
          2310 => x"d8d408fc",
          2311 => x"0508802e",
          2312 => x"ae38800b",
          2313 => x"82d8d408",
          2314 => x"8c050824",
          2315 => x"a23882d8",
          2316 => x"d4088c05",
          2317 => x"081082d8",
          2318 => x"d4088c05",
          2319 => x"0c82d8d4",
          2320 => x"08fc0508",
          2321 => x"1082d8d4",
          2322 => x"08fc050c",
          2323 => x"ffb83982",
          2324 => x"d8d408fc",
          2325 => x"0508802e",
          2326 => x"80e13882",
          2327 => x"d8d4088c",
          2328 => x"050882d8",
          2329 => x"d4088805",
          2330 => x"0826ad38",
          2331 => x"82d8d408",
          2332 => x"88050882",
          2333 => x"d8d4088c",
          2334 => x"05083182",
          2335 => x"d8d40888",
          2336 => x"050c82d8",
          2337 => x"d408f805",
          2338 => x"0882d8d4",
          2339 => x"08fc0508",
          2340 => x"0782d8d4",
          2341 => x"08f8050c",
          2342 => x"82d8d408",
          2343 => x"fc050881",
          2344 => x"2a82d8d4",
          2345 => x"08fc050c",
          2346 => x"82d8d408",
          2347 => x"8c050881",
          2348 => x"2a82d8d4",
          2349 => x"088c050c",
          2350 => x"ff953982",
          2351 => x"d8d40890",
          2352 => x"0508802e",
          2353 => x"933882d8",
          2354 => x"d4088805",
          2355 => x"087082d8",
          2356 => x"d408f405",
          2357 => x"0c519139",
          2358 => x"82d8d408",
          2359 => x"f8050870",
          2360 => x"82d8d408",
          2361 => x"f4050c51",
          2362 => x"82d8d408",
          2363 => x"f4050882",
          2364 => x"d8c80c85",
          2365 => x"3d0d82d8",
          2366 => x"d40c0482",
          2367 => x"d8d40802",
          2368 => x"82d8d40c",
          2369 => x"f73d0d80",
          2370 => x"0b82d8d4",
          2371 => x"08f00534",
          2372 => x"82d8d408",
          2373 => x"8c050853",
          2374 => x"80730c82",
          2375 => x"d8d40888",
          2376 => x"05087008",
          2377 => x"51537233",
          2378 => x"537282d8",
          2379 => x"d408f805",
          2380 => x"347281ff",
          2381 => x"065372a0",
          2382 => x"2e098106",
          2383 => x"913882d8",
          2384 => x"d4088805",
          2385 => x"08700881",
          2386 => x"05710c53",
          2387 => x"ce3982d8",
          2388 => x"d408f805",
          2389 => x"335372ad",
          2390 => x"2e098106",
          2391 => x"a438810b",
          2392 => x"82d8d408",
          2393 => x"f0053482",
          2394 => x"d8d40888",
          2395 => x"05087008",
          2396 => x"8105710c",
          2397 => x"70085153",
          2398 => x"723382d8",
          2399 => x"d408f805",
          2400 => x"3482d8d4",
          2401 => x"08f80533",
          2402 => x"5372b02e",
          2403 => x"09810681",
          2404 => x"dc3882d8",
          2405 => x"d4088805",
          2406 => x"08700881",
          2407 => x"05710c70",
          2408 => x"08515372",
          2409 => x"3382d8d4",
          2410 => x"08f80534",
          2411 => x"82d8d408",
          2412 => x"f8053382",
          2413 => x"d8d408e8",
          2414 => x"050c82d8",
          2415 => x"d408e805",
          2416 => x"0880e22e",
          2417 => x"b63882d8",
          2418 => x"d408e805",
          2419 => x"0880f82e",
          2420 => x"843880cd",
          2421 => x"39900b82",
          2422 => x"d8d408f4",
          2423 => x"053482d8",
          2424 => x"d4088805",
          2425 => x"08700881",
          2426 => x"05710c70",
          2427 => x"08515372",
          2428 => x"3382d8d4",
          2429 => x"08f80534",
          2430 => x"81a43982",
          2431 => x"0b82d8d4",
          2432 => x"08f40534",
          2433 => x"82d8d408",
          2434 => x"88050870",
          2435 => x"08810571",
          2436 => x"0c700851",
          2437 => x"53723382",
          2438 => x"d8d408f8",
          2439 => x"053480fe",
          2440 => x"3982d8d4",
          2441 => x"08f80533",
          2442 => x"5372a026",
          2443 => x"8d38810b",
          2444 => x"82d8d408",
          2445 => x"ec050c83",
          2446 => x"803982d8",
          2447 => x"d408f805",
          2448 => x"3353af73",
          2449 => x"27903882",
          2450 => x"d8d408f8",
          2451 => x"05335372",
          2452 => x"b9268338",
          2453 => x"8d39800b",
          2454 => x"82d8d408",
          2455 => x"ec050c82",
          2456 => x"d839880b",
          2457 => x"82d8d408",
          2458 => x"f40534b2",
          2459 => x"3982d8d4",
          2460 => x"08f80533",
          2461 => x"53af7327",
          2462 => x"903882d8",
          2463 => x"d408f805",
          2464 => x"335372b9",
          2465 => x"2683388d",
          2466 => x"39800b82",
          2467 => x"d8d408ec",
          2468 => x"050c82a5",
          2469 => x"398a0b82",
          2470 => x"d8d408f4",
          2471 => x"0534800b",
          2472 => x"82d8d408",
          2473 => x"fc050c82",
          2474 => x"d8d408f8",
          2475 => x"053353a0",
          2476 => x"732781cf",
          2477 => x"3882d8d4",
          2478 => x"08f80533",
          2479 => x"5380e073",
          2480 => x"27943882",
          2481 => x"d8d408f8",
          2482 => x"0533e011",
          2483 => x"51537282",
          2484 => x"d8d408f8",
          2485 => x"053482d8",
          2486 => x"d408f805",
          2487 => x"33d01151",
          2488 => x"537282d8",
          2489 => x"d408f805",
          2490 => x"3482d8d4",
          2491 => x"08f80533",
          2492 => x"53907327",
          2493 => x"ad3882d8",
          2494 => x"d408f805",
          2495 => x"33f91151",
          2496 => x"537282d8",
          2497 => x"d408f805",
          2498 => x"3482d8d4",
          2499 => x"08f80533",
          2500 => x"53728926",
          2501 => x"8d38800b",
          2502 => x"82d8d408",
          2503 => x"ec050c81",
          2504 => x"983982d8",
          2505 => x"d408f805",
          2506 => x"3382d8d4",
          2507 => x"08f40533",
          2508 => x"54547274",
          2509 => x"268d3880",
          2510 => x"0b82d8d4",
          2511 => x"08ec050c",
          2512 => x"80f73982",
          2513 => x"d8d408f4",
          2514 => x"05337082",
          2515 => x"d8d408fc",
          2516 => x"05082982",
          2517 => x"d8d408f8",
          2518 => x"05337012",
          2519 => x"82d8d408",
          2520 => x"fc050c82",
          2521 => x"d8d40888",
          2522 => x"05087008",
          2523 => x"8105710c",
          2524 => x"70085151",
          2525 => x"52555372",
          2526 => x"3382d8d4",
          2527 => x"08f80534",
          2528 => x"fea53982",
          2529 => x"d8d408f0",
          2530 => x"05335372",
          2531 => x"802e9038",
          2532 => x"82d8d408",
          2533 => x"fc050830",
          2534 => x"82d8d408",
          2535 => x"fc050c82",
          2536 => x"d8d4088c",
          2537 => x"050882d8",
          2538 => x"d408fc05",
          2539 => x"08710c53",
          2540 => x"810b82d8",
          2541 => x"d408ec05",
          2542 => x"0c82d8d4",
          2543 => x"08ec0508",
          2544 => x"82d8c80c",
          2545 => x"8b3d0d82",
          2546 => x"d8d40c04",
          2547 => x"82d8d408",
          2548 => x"0282d8d4",
          2549 => x"0cf73d0d",
          2550 => x"800b82d8",
          2551 => x"d408f005",
          2552 => x"3482d8d4",
          2553 => x"088c0508",
          2554 => x"5380730c",
          2555 => x"82d8d408",
          2556 => x"88050870",
          2557 => x"08515372",
          2558 => x"33537282",
          2559 => x"d8d408f8",
          2560 => x"05347281",
          2561 => x"ff065372",
          2562 => x"a02e0981",
          2563 => x"06913882",
          2564 => x"d8d40888",
          2565 => x"05087008",
          2566 => x"8105710c",
          2567 => x"53ce3982",
          2568 => x"d8d408f8",
          2569 => x"05335372",
          2570 => x"ad2e0981",
          2571 => x"06a43881",
          2572 => x"0b82d8d4",
          2573 => x"08f00534",
          2574 => x"82d8d408",
          2575 => x"88050870",
          2576 => x"08810571",
          2577 => x"0c700851",
          2578 => x"53723382",
          2579 => x"d8d408f8",
          2580 => x"053482d8",
          2581 => x"d408f805",
          2582 => x"335372b0",
          2583 => x"2e098106",
          2584 => x"81dc3882",
          2585 => x"d8d40888",
          2586 => x"05087008",
          2587 => x"8105710c",
          2588 => x"70085153",
          2589 => x"723382d8",
          2590 => x"d408f805",
          2591 => x"3482d8d4",
          2592 => x"08f80533",
          2593 => x"82d8d408",
          2594 => x"e8050c82",
          2595 => x"d8d408e8",
          2596 => x"050880e2",
          2597 => x"2eb63882",
          2598 => x"d8d408e8",
          2599 => x"050880f8",
          2600 => x"2e843880",
          2601 => x"cd39900b",
          2602 => x"82d8d408",
          2603 => x"f4053482",
          2604 => x"d8d40888",
          2605 => x"05087008",
          2606 => x"8105710c",
          2607 => x"70085153",
          2608 => x"723382d8",
          2609 => x"d408f805",
          2610 => x"3481a439",
          2611 => x"820b82d8",
          2612 => x"d408f405",
          2613 => x"3482d8d4",
          2614 => x"08880508",
          2615 => x"70088105",
          2616 => x"710c7008",
          2617 => x"51537233",
          2618 => x"82d8d408",
          2619 => x"f8053480",
          2620 => x"fe3982d8",
          2621 => x"d408f805",
          2622 => x"335372a0",
          2623 => x"268d3881",
          2624 => x"0b82d8d4",
          2625 => x"08ec050c",
          2626 => x"83803982",
          2627 => x"d8d408f8",
          2628 => x"053353af",
          2629 => x"73279038",
          2630 => x"82d8d408",
          2631 => x"f8053353",
          2632 => x"72b92683",
          2633 => x"388d3980",
          2634 => x"0b82d8d4",
          2635 => x"08ec050c",
          2636 => x"82d83988",
          2637 => x"0b82d8d4",
          2638 => x"08f40534",
          2639 => x"b23982d8",
          2640 => x"d408f805",
          2641 => x"3353af73",
          2642 => x"27903882",
          2643 => x"d8d408f8",
          2644 => x"05335372",
          2645 => x"b9268338",
          2646 => x"8d39800b",
          2647 => x"82d8d408",
          2648 => x"ec050c82",
          2649 => x"a5398a0b",
          2650 => x"82d8d408",
          2651 => x"f4053480",
          2652 => x"0b82d8d4",
          2653 => x"08fc050c",
          2654 => x"82d8d408",
          2655 => x"f8053353",
          2656 => x"a0732781",
          2657 => x"cf3882d8",
          2658 => x"d408f805",
          2659 => x"335380e0",
          2660 => x"73279438",
          2661 => x"82d8d408",
          2662 => x"f80533e0",
          2663 => x"11515372",
          2664 => x"82d8d408",
          2665 => x"f8053482",
          2666 => x"d8d408f8",
          2667 => x"0533d011",
          2668 => x"51537282",
          2669 => x"d8d408f8",
          2670 => x"053482d8",
          2671 => x"d408f805",
          2672 => x"33539073",
          2673 => x"27ad3882",
          2674 => x"d8d408f8",
          2675 => x"0533f911",
          2676 => x"51537282",
          2677 => x"d8d408f8",
          2678 => x"053482d8",
          2679 => x"d408f805",
          2680 => x"33537289",
          2681 => x"268d3880",
          2682 => x"0b82d8d4",
          2683 => x"08ec050c",
          2684 => x"81983982",
          2685 => x"d8d408f8",
          2686 => x"053382d8",
          2687 => x"d408f405",
          2688 => x"33545472",
          2689 => x"74268d38",
          2690 => x"800b82d8",
          2691 => x"d408ec05",
          2692 => x"0c80f739",
          2693 => x"82d8d408",
          2694 => x"f4053370",
          2695 => x"82d8d408",
          2696 => x"fc050829",
          2697 => x"82d8d408",
          2698 => x"f8053370",
          2699 => x"1282d8d4",
          2700 => x"08fc050c",
          2701 => x"82d8d408",
          2702 => x"88050870",
          2703 => x"08810571",
          2704 => x"0c700851",
          2705 => x"51525553",
          2706 => x"723382d8",
          2707 => x"d408f805",
          2708 => x"34fea539",
          2709 => x"82d8d408",
          2710 => x"f0053353",
          2711 => x"72802e90",
          2712 => x"3882d8d4",
          2713 => x"08fc0508",
          2714 => x"3082d8d4",
          2715 => x"08fc050c",
          2716 => x"82d8d408",
          2717 => x"8c050882",
          2718 => x"d8d408fc",
          2719 => x"0508710c",
          2720 => x"53810b82",
          2721 => x"d8d408ec",
          2722 => x"050c82d8",
          2723 => x"d408ec05",
          2724 => x"0882d8c8",
          2725 => x"0c8b3d0d",
          2726 => x"82d8d40c",
          2727 => x"04f93d0d",
          2728 => x"79700870",
          2729 => x"56565874",
          2730 => x"802e80e3",
          2731 => x"38953975",
          2732 => x"0851e6d1",
          2733 => x"3f82d8c8",
          2734 => x"0815780c",
          2735 => x"85163354",
          2736 => x"80cd3974",
          2737 => x"335473a0",
          2738 => x"2e098106",
          2739 => x"86388115",
          2740 => x"55f13980",
          2741 => x"57769029",
          2742 => x"82d3c805",
          2743 => x"70085256",
          2744 => x"e6a33f82",
          2745 => x"d8c80853",
          2746 => x"74527508",
          2747 => x"51e9a33f",
          2748 => x"82d8c808",
          2749 => x"8b388416",
          2750 => x"33547381",
          2751 => x"2effb038",
          2752 => x"81177081",
          2753 => x"ff065854",
          2754 => x"997727c9",
          2755 => x"38ff5473",
          2756 => x"82d8c80c",
          2757 => x"893d0d04",
          2758 => x"ff3d0d73",
          2759 => x"52719326",
          2760 => x"818e3871",
          2761 => x"842982ae",
          2762 => x"f4055271",
          2763 => x"080482b4",
          2764 => x"e4518180",
          2765 => x"3982b4f0",
          2766 => x"5180f939",
          2767 => x"82b58051",
          2768 => x"80f23982",
          2769 => x"b5905180",
          2770 => x"eb3982b5",
          2771 => x"a05180e4",
          2772 => x"3982b5b0",
          2773 => x"5180dd39",
          2774 => x"82b5c451",
          2775 => x"80d63982",
          2776 => x"b5d45180",
          2777 => x"cf3982b5",
          2778 => x"ec5180c8",
          2779 => x"3982b684",
          2780 => x"5180c139",
          2781 => x"82b69c51",
          2782 => x"bb3982b6",
          2783 => x"b851b539",
          2784 => x"82b6cc51",
          2785 => x"af3982b6",
          2786 => x"f451a939",
          2787 => x"82b78451",
          2788 => x"a33982b7",
          2789 => x"a4519d39",
          2790 => x"82b7b451",
          2791 => x"973982b7",
          2792 => x"cc519139",
          2793 => x"82b7e451",
          2794 => x"8b3982b7",
          2795 => x"fc518539",
          2796 => x"82b88851",
          2797 => x"d8ad3f83",
          2798 => x"3d0d04fb",
          2799 => x"3d0d7779",
          2800 => x"56567487",
          2801 => x"e7268a38",
          2802 => x"74527587",
          2803 => x"e8295190",
          2804 => x"3987e852",
          2805 => x"7451efab",
          2806 => x"3f82d8c8",
          2807 => x"08527551",
          2808 => x"efa13f82",
          2809 => x"d8c80854",
          2810 => x"79537552",
          2811 => x"82b89851",
          2812 => x"ffbbe53f",
          2813 => x"873d0d04",
          2814 => x"ec3d0d66",
          2815 => x"02840580",
          2816 => x"e305335b",
          2817 => x"57806878",
          2818 => x"30707a07",
          2819 => x"73255157",
          2820 => x"59597856",
          2821 => x"7787ff26",
          2822 => x"83388156",
          2823 => x"74760770",
          2824 => x"81ff0651",
          2825 => x"55935674",
          2826 => x"81823881",
          2827 => x"5376528c",
          2828 => x"3d705256",
          2829 => x"8196903f",
          2830 => x"82d8c808",
          2831 => x"5782d8c8",
          2832 => x"08b93882",
          2833 => x"d8c80887",
          2834 => x"c098880c",
          2835 => x"82d8c808",
          2836 => x"59963dd4",
          2837 => x"05548480",
          2838 => x"53775275",
          2839 => x"51819acc",
          2840 => x"3f82d8c8",
          2841 => x"085782d8",
          2842 => x"c8089038",
          2843 => x"7a557480",
          2844 => x"2e893874",
          2845 => x"19751959",
          2846 => x"59d73996",
          2847 => x"3dd80551",
          2848 => x"81a2c33f",
          2849 => x"76307078",
          2850 => x"0780257b",
          2851 => x"30709f2a",
          2852 => x"72065157",
          2853 => x"51567480",
          2854 => x"2e903882",
          2855 => x"b8bc5387",
          2856 => x"c0988808",
          2857 => x"527851fe",
          2858 => x"923f7656",
          2859 => x"7582d8c8",
          2860 => x"0c963d0d",
          2861 => x"04f73d0d",
          2862 => x"7d028405",
          2863 => x"bb053359",
          2864 => x"5aff5980",
          2865 => x"537c527b",
          2866 => x"51fead3f",
          2867 => x"82d8c808",
          2868 => x"80cb3877",
          2869 => x"802e8838",
          2870 => x"77812ebf",
          2871 => x"38bf3982",
          2872 => x"f4a85782",
          2873 => x"f4a85682",
          2874 => x"f4a85582",
          2875 => x"f4b00854",
          2876 => x"82f4ac08",
          2877 => x"5382f4a8",
          2878 => x"085282b8",
          2879 => x"c451ffb9",
          2880 => x"d73f82f4",
          2881 => x"a8566255",
          2882 => x"615482d8",
          2883 => x"c8536052",
          2884 => x"7f51792d",
          2885 => x"82d8c808",
          2886 => x"59833979",
          2887 => x"047882d8",
          2888 => x"c80c8b3d",
          2889 => x"0d04f33d",
          2890 => x"0d7f6163",
          2891 => x"028c0580",
          2892 => x"cf053373",
          2893 => x"73156841",
          2894 => x"5f5c5c5e",
          2895 => x"5e5e7a52",
          2896 => x"82b8f851",
          2897 => x"ffb9913f",
          2898 => x"82b98051",
          2899 => x"ffb9893f",
          2900 => x"80557479",
          2901 => x"27818038",
          2902 => x"7b902e89",
          2903 => x"387ba02e",
          2904 => x"a73880c6",
          2905 => x"39741853",
          2906 => x"727a278e",
          2907 => x"38722252",
          2908 => x"82b98451",
          2909 => x"ffb8e13f",
          2910 => x"893982b9",
          2911 => x"9051ffb8",
          2912 => x"d73f8215",
          2913 => x"5580c339",
          2914 => x"74185372",
          2915 => x"7a278e38",
          2916 => x"72085282",
          2917 => x"b8f851ff",
          2918 => x"b8be3f89",
          2919 => x"3982b98c",
          2920 => x"51ffb8b4",
          2921 => x"3f841555",
          2922 => x"a1397418",
          2923 => x"53727a27",
          2924 => x"8e387233",
          2925 => x"5282b998",
          2926 => x"51ffb89c",
          2927 => x"3f893982",
          2928 => x"b9a051ff",
          2929 => x"b8923f81",
          2930 => x"155582f4",
          2931 => x"ac0852a0",
          2932 => x"51d7df3f",
          2933 => x"fefc3982",
          2934 => x"b9a451ff",
          2935 => x"b7fa3f80",
          2936 => x"55747927",
          2937 => x"80c63874",
          2938 => x"18703355",
          2939 => x"53805672",
          2940 => x"7a278338",
          2941 => x"81568053",
          2942 => x"9f742783",
          2943 => x"38815375",
          2944 => x"73067081",
          2945 => x"ff065153",
          2946 => x"72802e90",
          2947 => x"387380fe",
          2948 => x"268a3882",
          2949 => x"f4ac0852",
          2950 => x"73518839",
          2951 => x"82f4ac08",
          2952 => x"52a051d7",
          2953 => x"8d3f8115",
          2954 => x"55ffb639",
          2955 => x"82b9a851",
          2956 => x"d3b13f78",
          2957 => x"18791c5c",
          2958 => x"58a1803f",
          2959 => x"82d8c808",
          2960 => x"982b7098",
          2961 => x"2c515776",
          2962 => x"a02e0981",
          2963 => x"06aa38a0",
          2964 => x"ea3f82d8",
          2965 => x"c808982b",
          2966 => x"70982c70",
          2967 => x"a0327030",
          2968 => x"729b3270",
          2969 => x"30707207",
          2970 => x"73750706",
          2971 => x"51585859",
          2972 => x"57515780",
          2973 => x"7324d838",
          2974 => x"769b2e09",
          2975 => x"81068538",
          2976 => x"80538c39",
          2977 => x"7c1e5372",
          2978 => x"7826fdb2",
          2979 => x"38ff5372",
          2980 => x"82d8c80c",
          2981 => x"8f3d0d04",
          2982 => x"fc3d0d02",
          2983 => x"9b053382",
          2984 => x"b9ac5382",
          2985 => x"b9b45255",
          2986 => x"ffb6ad3f",
          2987 => x"82d7a022",
          2988 => x"51a9d93f",
          2989 => x"82b9c054",
          2990 => x"82b9cc53",
          2991 => x"82d7a133",
          2992 => x"5282b9d4",
          2993 => x"51ffb690",
          2994 => x"3f74802e",
          2995 => x"8438a58d",
          2996 => x"3f863d0d",
          2997 => x"04fe3d0d",
          2998 => x"87c09680",
          2999 => x"0853aab6",
          3000 => x"3f81519c",
          3001 => x"c33f82b9",
          3002 => x"f0519dd8",
          3003 => x"3f80519c",
          3004 => x"b73f7281",
          3005 => x"2a708106",
          3006 => x"51527180",
          3007 => x"2e923881",
          3008 => x"519ca53f",
          3009 => x"82ba8851",
          3010 => x"9dba3f80",
          3011 => x"519c993f",
          3012 => x"72822a70",
          3013 => x"81065152",
          3014 => x"71802e92",
          3015 => x"3881519c",
          3016 => x"873f82ba",
          3017 => x"98519d9c",
          3018 => x"3f80519b",
          3019 => x"fb3f7283",
          3020 => x"2a708106",
          3021 => x"51527180",
          3022 => x"2e923881",
          3023 => x"519be93f",
          3024 => x"82baa851",
          3025 => x"9cfe3f80",
          3026 => x"519bdd3f",
          3027 => x"72842a70",
          3028 => x"81065152",
          3029 => x"71802e92",
          3030 => x"3881519b",
          3031 => x"cb3f82ba",
          3032 => x"bc519ce0",
          3033 => x"3f80519b",
          3034 => x"bf3f7285",
          3035 => x"2a708106",
          3036 => x"51527180",
          3037 => x"2e923881",
          3038 => x"519bad3f",
          3039 => x"82bad051",
          3040 => x"9cc23f80",
          3041 => x"519ba13f",
          3042 => x"72862a70",
          3043 => x"81065152",
          3044 => x"71802e92",
          3045 => x"3881519b",
          3046 => x"8f3f82ba",
          3047 => x"e4519ca4",
          3048 => x"3f80519b",
          3049 => x"833f7287",
          3050 => x"2a708106",
          3051 => x"51527180",
          3052 => x"2e923881",
          3053 => x"519af13f",
          3054 => x"82baf851",
          3055 => x"9c863f80",
          3056 => x"519ae53f",
          3057 => x"72882a70",
          3058 => x"81065152",
          3059 => x"71802e92",
          3060 => x"3881519a",
          3061 => x"d33f82bb",
          3062 => x"8c519be8",
          3063 => x"3f80519a",
          3064 => x"c73fa8ba",
          3065 => x"3f843d0d",
          3066 => x"04fb3d0d",
          3067 => x"77028405",
          3068 => x"a3053370",
          3069 => x"55565680",
          3070 => x"527551e2",
          3071 => x"e93f0b0b",
          3072 => x"82d3c433",
          3073 => x"5473a938",
          3074 => x"815382bb",
          3075 => x"c85282ef",
          3076 => x"d851818e",
          3077 => x"b23f82d8",
          3078 => x"c8083070",
          3079 => x"82d8c808",
          3080 => x"07802582",
          3081 => x"71315151",
          3082 => x"54730b0b",
          3083 => x"82d3c434",
          3084 => x"0b0b82d3",
          3085 => x"c4335473",
          3086 => x"812e0981",
          3087 => x"06af3882",
          3088 => x"efd85374",
          3089 => x"52755181",
          3090 => x"c9823f82",
          3091 => x"d8c80880",
          3092 => x"2e8b3882",
          3093 => x"d8c80851",
          3094 => x"cf893f91",
          3095 => x"3982efd8",
          3096 => x"51819ae2",
          3097 => x"3f820b0b",
          3098 => x"0b82d3c4",
          3099 => x"340b0b82",
          3100 => x"d3c43354",
          3101 => x"73822e09",
          3102 => x"81068c38",
          3103 => x"82bbd853",
          3104 => x"74527551",
          3105 => x"aeb23f80",
          3106 => x"0b82d8c8",
          3107 => x"0c873d0d",
          3108 => x"04ce3d0d",
          3109 => x"80707182",
          3110 => x"efd40c5f",
          3111 => x"5d81527c",
          3112 => x"5180cbcb",
          3113 => x"3f82d8c8",
          3114 => x"0881ff06",
          3115 => x"59787d2e",
          3116 => x"098106a3",
          3117 => x"38963d59",
          3118 => x"835382bb",
          3119 => x"e4527851",
          3120 => x"dca33f7c",
          3121 => x"53785282",
          3122 => x"d9f45181",
          3123 => x"8c983f82",
          3124 => x"d8c8087d",
          3125 => x"2e883882",
          3126 => x"bbe85191",
          3127 => x"d7398170",
          3128 => x"5f5d82bc",
          3129 => x"a051ffb1",
          3130 => x"ef3f963d",
          3131 => x"70465a80",
          3132 => x"f8527951",
          3133 => x"fdf33fb4",
          3134 => x"3dff8405",
          3135 => x"51f39e3f",
          3136 => x"82d8c808",
          3137 => x"902b7090",
          3138 => x"2c515978",
          3139 => x"80c12e89",
          3140 => x"d4387880",
          3141 => x"c12480d9",
          3142 => x"3878ab2e",
          3143 => x"83b93878",
          3144 => x"ab24a438",
          3145 => x"78822e81",
          3146 => x"b3387882",
          3147 => x"248a3878",
          3148 => x"802effae",
          3149 => x"388f8239",
          3150 => x"78842e82",
          3151 => x"83387894",
          3152 => x"2e82ad38",
          3153 => x"8ef33978",
          3154 => x"bd2e84fc",
          3155 => x"3878bd24",
          3156 => x"903878b0",
          3157 => x"2e83a638",
          3158 => x"78bc2e84",
          3159 => x"84388ed9",
          3160 => x"3978bf2e",
          3161 => x"85c43878",
          3162 => x"80c02e86",
          3163 => x"bd388ec9",
          3164 => x"397880d5",
          3165 => x"2e8da238",
          3166 => x"7880d524",
          3167 => x"b0387880",
          3168 => x"d02e8cd9",
          3169 => x"387880d0",
          3170 => x"24923878",
          3171 => x"80c22e89",
          3172 => x"fc387880",
          3173 => x"c32e8ba5",
          3174 => x"388e9e39",
          3175 => x"7880d12e",
          3176 => x"8cca3878",
          3177 => x"80d42e8c",
          3178 => x"d3388e8d",
          3179 => x"39788182",
          3180 => x"2e8de438",
          3181 => x"78818224",
          3182 => x"92387880",
          3183 => x"f82e8cf6",
          3184 => x"387880f9",
          3185 => x"2e8d9338",
          3186 => x"8def3978",
          3187 => x"81832e8d",
          3188 => x"d5387881",
          3189 => x"852e8ddb",
          3190 => x"388dde39",
          3191 => x"b43dff80",
          3192 => x"1153ff84",
          3193 => x"0551ebe4",
          3194 => x"3f82d8c8",
          3195 => x"08883882",
          3196 => x"bca4518f",
          3197 => x"bf39b43d",
          3198 => x"fefc1153",
          3199 => x"ff840551",
          3200 => x"ebca3f82",
          3201 => x"d8c80880",
          3202 => x"2e883881",
          3203 => x"63258338",
          3204 => x"80430280",
          3205 => x"cb053352",
          3206 => x"0280cf05",
          3207 => x"335180c8",
          3208 => x"ce3f82d8",
          3209 => x"c80881ff",
          3210 => x"0659788d",
          3211 => x"3882bcb4",
          3212 => x"51cbb03f",
          3213 => x"815efdaa",
          3214 => x"3982bcc4",
          3215 => x"518ef539",
          3216 => x"b43dff80",
          3217 => x"1153ff84",
          3218 => x"0551eb80",
          3219 => x"3f82d8c8",
          3220 => x"08802efd",
          3221 => x"8d388053",
          3222 => x"80520280",
          3223 => x"cf053351",
          3224 => x"80ccd93f",
          3225 => x"82d8c808",
          3226 => x"5282bcdc",
          3227 => x"518ca139",
          3228 => x"b43dff80",
          3229 => x"1153ff84",
          3230 => x"0551ead0",
          3231 => x"3f82d8c8",
          3232 => x"08802e87",
          3233 => x"38638926",
          3234 => x"fcd838b4",
          3235 => x"3dfefc11",
          3236 => x"53ff8405",
          3237 => x"51eab53f",
          3238 => x"82d8c808",
          3239 => x"863882d8",
          3240 => x"c8084363",
          3241 => x"5382bce4",
          3242 => x"527951ff",
          3243 => x"b1923f02",
          3244 => x"80cb0533",
          3245 => x"53795263",
          3246 => x"84b82982",
          3247 => x"d9f40551",
          3248 => x"8188a33f",
          3249 => x"82d8c808",
          3250 => x"818c3882",
          3251 => x"bcb451ca",
          3252 => x"923f815d",
          3253 => x"fc8c39b4",
          3254 => x"3dff8405",
          3255 => x"518fc23f",
          3256 => x"82d8c808",
          3257 => x"b53dff84",
          3258 => x"05525b90",
          3259 => x"d83f8153",
          3260 => x"82d8c808",
          3261 => x"527a51f1",
          3262 => x"ff3f80d1",
          3263 => x"39b43dff",
          3264 => x"8405518f",
          3265 => x"9c3f82d8",
          3266 => x"c808b53d",
          3267 => x"ff840552",
          3268 => x"5b90b23f",
          3269 => x"82d8c808",
          3270 => x"b53dff84",
          3271 => x"05525a90",
          3272 => x"a43f82d8",
          3273 => x"c808b53d",
          3274 => x"ff840552",
          3275 => x"5990963f",
          3276 => x"82d6ec58",
          3277 => x"82d8f857",
          3278 => x"80568055",
          3279 => x"82d8c808",
          3280 => x"81ff0654",
          3281 => x"78537952",
          3282 => x"7a51f2e9",
          3283 => x"3f82d8c8",
          3284 => x"08802efb",
          3285 => x"8d3882d8",
          3286 => x"c80851ef",
          3287 => x"bb3ffb82",
          3288 => x"39b43dff",
          3289 => x"801153ff",
          3290 => x"840551e8",
          3291 => x"df3f82d8",
          3292 => x"c808802e",
          3293 => x"faec38b4",
          3294 => x"3dfefc11",
          3295 => x"53ff8405",
          3296 => x"51e8c93f",
          3297 => x"82d8c808",
          3298 => x"802efad6",
          3299 => x"38b43dfe",
          3300 => x"f81153ff",
          3301 => x"840551e8",
          3302 => x"b33f82d8",
          3303 => x"c8088638",
          3304 => x"82d8c808",
          3305 => x"4282bce8",
          3306 => x"51ffacac",
          3307 => x"3f63635c",
          3308 => x"5a797b27",
          3309 => x"81ec3861",
          3310 => x"59787a70",
          3311 => x"84055c0c",
          3312 => x"7a7a26f5",
          3313 => x"3881db39",
          3314 => x"b43dff80",
          3315 => x"1153ff84",
          3316 => x"0551e7f8",
          3317 => x"3f82d8c8",
          3318 => x"08802efa",
          3319 => x"8538b43d",
          3320 => x"fefc1153",
          3321 => x"ff840551",
          3322 => x"e7e23f82",
          3323 => x"d8c80880",
          3324 => x"2ef9ef38",
          3325 => x"b43dfef8",
          3326 => x"1153ff84",
          3327 => x"0551e7cc",
          3328 => x"3f82d8c8",
          3329 => x"08802ef9",
          3330 => x"d93882bc",
          3331 => x"f851ffab",
          3332 => x"c73f635a",
          3333 => x"79632781",
          3334 => x"89386159",
          3335 => x"79708105",
          3336 => x"5b337934",
          3337 => x"61810542",
          3338 => x"eb39b43d",
          3339 => x"ff801153",
          3340 => x"ff840551",
          3341 => x"e7963f82",
          3342 => x"d8c80880",
          3343 => x"2ef9a338",
          3344 => x"b43dfefc",
          3345 => x"1153ff84",
          3346 => x"0551e780",
          3347 => x"3f82d8c8",
          3348 => x"08802ef9",
          3349 => x"8d38b43d",
          3350 => x"fef81153",
          3351 => x"ff840551",
          3352 => x"e6ea3f82",
          3353 => x"d8c80880",
          3354 => x"2ef8f738",
          3355 => x"82bd8451",
          3356 => x"ffaae53f",
          3357 => x"635a7963",
          3358 => x"27a83861",
          3359 => x"70337b33",
          3360 => x"5e5a5b78",
          3361 => x"7c2e9238",
          3362 => x"78557a54",
          3363 => x"79335379",
          3364 => x"5282bd94",
          3365 => x"51ffaac0",
          3366 => x"3f811a62",
          3367 => x"8105435a",
          3368 => x"d5398a51",
          3369 => x"c9df3ff8",
          3370 => x"b939b43d",
          3371 => x"ff801153",
          3372 => x"ff840551",
          3373 => x"e6963f82",
          3374 => x"d8c80880",
          3375 => x"df3882d7",
          3376 => x"b4335978",
          3377 => x"802e8938",
          3378 => x"82d6ec08",
          3379 => x"4480cd39",
          3380 => x"82d7b533",
          3381 => x"5978802e",
          3382 => x"883882d6",
          3383 => x"f40844bc",
          3384 => x"3982d7b6",
          3385 => x"33597880",
          3386 => x"2e883882",
          3387 => x"d6fc0844",
          3388 => x"ab3982d7",
          3389 => x"b7335978",
          3390 => x"802e8838",
          3391 => x"82d78408",
          3392 => x"449a3982",
          3393 => x"d7b23359",
          3394 => x"78802e88",
          3395 => x"3882d78c",
          3396 => x"08448939",
          3397 => x"82d79c08",
          3398 => x"fc800544",
          3399 => x"b43dfefc",
          3400 => x"1153ff84",
          3401 => x"0551e5a4",
          3402 => x"3f82d8c8",
          3403 => x"0880de38",
          3404 => x"82d7b433",
          3405 => x"5978802e",
          3406 => x"893882d6",
          3407 => x"f0084380",
          3408 => x"cc3982d7",
          3409 => x"b5335978",
          3410 => x"802e8838",
          3411 => x"82d6f808",
          3412 => x"43bb3982",
          3413 => x"d7b63359",
          3414 => x"78802e88",
          3415 => x"3882d780",
          3416 => x"0843aa39",
          3417 => x"82d7b733",
          3418 => x"5978802e",
          3419 => x"883882d7",
          3420 => x"88084399",
          3421 => x"3982d7b2",
          3422 => x"33597880",
          3423 => x"2e883882",
          3424 => x"d7900843",
          3425 => x"883982d7",
          3426 => x"9c088805",
          3427 => x"43b43dfe",
          3428 => x"f81153ff",
          3429 => x"840551e4",
          3430 => x"b33f82d8",
          3431 => x"c808802e",
          3432 => x"a7388062",
          3433 => x"5c5c7a88",
          3434 => x"2e833881",
          3435 => x"5c7a9032",
          3436 => x"70307072",
          3437 => x"079f2a70",
          3438 => x"7f065151",
          3439 => x"5a5a7880",
          3440 => x"2e88387a",
          3441 => x"a02e8338",
          3442 => x"884282bd",
          3443 => x"b051c493",
          3444 => x"3fa05563",
          3445 => x"54615362",
          3446 => x"526351ee",
          3447 => x"c93f82bd",
          3448 => x"bc5187d0",
          3449 => x"39b43dff",
          3450 => x"801153ff",
          3451 => x"840551e3",
          3452 => x"db3f82d8",
          3453 => x"c808802e",
          3454 => x"f5e838b4",
          3455 => x"3dfefc11",
          3456 => x"53ff8405",
          3457 => x"51e3c53f",
          3458 => x"82d8c808",
          3459 => x"802ea438",
          3460 => x"63590280",
          3461 => x"cb053379",
          3462 => x"34638105",
          3463 => x"44b43dfe",
          3464 => x"fc1153ff",
          3465 => x"840551e3",
          3466 => x"a33f82d8",
          3467 => x"c808e138",
          3468 => x"f5b03963",
          3469 => x"70335452",
          3470 => x"82bdc851",
          3471 => x"ffa7993f",
          3472 => x"82f4a808",
          3473 => x"5380f852",
          3474 => x"7951ffa7",
          3475 => x"e03f7945",
          3476 => x"79335978",
          3477 => x"ae2ef58a",
          3478 => x"389f7927",
          3479 => x"9f38b43d",
          3480 => x"fefc1153",
          3481 => x"ff840551",
          3482 => x"e2e23f82",
          3483 => x"d8c80880",
          3484 => x"2e913863",
          3485 => x"590280cb",
          3486 => x"05337934",
          3487 => x"63810544",
          3488 => x"ffb13982",
          3489 => x"bdd451c2",
          3490 => x"da3fffa7",
          3491 => x"39b43dfe",
          3492 => x"f41153ff",
          3493 => x"840551dc",
          3494 => x"e23f82d8",
          3495 => x"c808802e",
          3496 => x"f4c038b4",
          3497 => x"3dfef011",
          3498 => x"53ff8405",
          3499 => x"51dccc3f",
          3500 => x"82d8c808",
          3501 => x"802ea538",
          3502 => x"605902be",
          3503 => x"05227970",
          3504 => x"82055b23",
          3505 => x"7841b43d",
          3506 => x"fef01153",
          3507 => x"ff840551",
          3508 => x"dca93f82",
          3509 => x"d8c808e0",
          3510 => x"38f48739",
          3511 => x"60702254",
          3512 => x"5282bdd8",
          3513 => x"51ffa5f0",
          3514 => x"3f82f4a8",
          3515 => x"085380f8",
          3516 => x"527951ff",
          3517 => x"a6b73f79",
          3518 => x"45793359",
          3519 => x"78ae2ef3",
          3520 => x"e138789f",
          3521 => x"26873860",
          3522 => x"820541d0",
          3523 => x"39b43dfe",
          3524 => x"f01153ff",
          3525 => x"840551db",
          3526 => x"e23f82d8",
          3527 => x"c808802e",
          3528 => x"92386059",
          3529 => x"02be0522",
          3530 => x"79708205",
          3531 => x"5b237841",
          3532 => x"ffaa3982",
          3533 => x"bdd451c1",
          3534 => x"aa3fffa0",
          3535 => x"39b43dfe",
          3536 => x"f41153ff",
          3537 => x"840551db",
          3538 => x"b23f82d8",
          3539 => x"c808802e",
          3540 => x"f39038b4",
          3541 => x"3dfef011",
          3542 => x"53ff8405",
          3543 => x"51db9c3f",
          3544 => x"82d8c808",
          3545 => x"802ea038",
          3546 => x"6060710c",
          3547 => x"59608405",
          3548 => x"41b43dfe",
          3549 => x"f01153ff",
          3550 => x"840551da",
          3551 => x"fe3f82d8",
          3552 => x"c808e538",
          3553 => x"f2dc3960",
          3554 => x"70085452",
          3555 => x"82bde451",
          3556 => x"ffa4c53f",
          3557 => x"82f4a808",
          3558 => x"5380f852",
          3559 => x"7951ffa5",
          3560 => x"8c3f7945",
          3561 => x"79335978",
          3562 => x"ae2ef2b6",
          3563 => x"389f7927",
          3564 => x"9b38b43d",
          3565 => x"fef01153",
          3566 => x"ff840551",
          3567 => x"dabd3f82",
          3568 => x"d8c80880",
          3569 => x"2e8d3860",
          3570 => x"60710c59",
          3571 => x"60840541",
          3572 => x"ffb53982",
          3573 => x"bdd451c0",
          3574 => x"8a3fffab",
          3575 => x"3982bdf4",
          3576 => x"51c0803f",
          3577 => x"82519889",
          3578 => x"3ff1f739",
          3579 => x"82be8c51",
          3580 => x"ffbff03f",
          3581 => x"a25197dd",
          3582 => x"3ff1e739",
          3583 => x"82bea051",
          3584 => x"ffbfe03f",
          3585 => x"8480810b",
          3586 => x"87c09484",
          3587 => x"0c848081",
          3588 => x"0b87c094",
          3589 => x"940cf1ca",
          3590 => x"3982beb4",
          3591 => x"51ffbfc3",
          3592 => x"3f8c8083",
          3593 => x"0b87c094",
          3594 => x"840c8c80",
          3595 => x"830b87c0",
          3596 => x"94940cf1",
          3597 => x"ad39b43d",
          3598 => x"ff801153",
          3599 => x"ff840551",
          3600 => x"df8a3f82",
          3601 => x"d8c80880",
          3602 => x"2ef19738",
          3603 => x"635282be",
          3604 => x"c851ffa3",
          3605 => x"833f6359",
          3606 => x"7804b43d",
          3607 => x"ff801153",
          3608 => x"ff840551",
          3609 => x"dee63f82",
          3610 => x"d8c80880",
          3611 => x"2ef0f338",
          3612 => x"635282be",
          3613 => x"e451ffa2",
          3614 => x"df3f6359",
          3615 => x"782d82d8",
          3616 => x"c808802e",
          3617 => x"f0dc3882",
          3618 => x"d8c80852",
          3619 => x"82bf8051",
          3620 => x"ffa2c53f",
          3621 => x"f0cc3982",
          3622 => x"bf9c51ff",
          3623 => x"bec53fff",
          3624 => x"a2973ff0",
          3625 => x"bd3982bf",
          3626 => x"b851ffbe",
          3627 => x"b63f8059",
          3628 => x"ffa63991",
          3629 => x"a83ff0aa",
          3630 => x"39794579",
          3631 => x"33597880",
          3632 => x"2ef09f38",
          3633 => x"7d7d0659",
          3634 => x"78802e81",
          3635 => x"cf38b43d",
          3636 => x"ff840551",
          3637 => x"83cb3f82",
          3638 => x"d8c8085b",
          3639 => x"815c7b82",
          3640 => x"2eb2387b",
          3641 => x"82248938",
          3642 => x"7b812e8c",
          3643 => x"3880ca39",
          3644 => x"7b832ead",
          3645 => x"3880c239",
          3646 => x"82bfcc56",
          3647 => x"7a5582bf",
          3648 => x"d0548053",
          3649 => x"82bfd452",
          3650 => x"b43dffb0",
          3651 => x"0551ffa4",
          3652 => x"af3fb839",
          3653 => x"7a52b43d",
          3654 => x"ffb00551",
          3655 => x"cad53fab",
          3656 => x"397a5582",
          3657 => x"bfd05480",
          3658 => x"5382bfe4",
          3659 => x"52b43dff",
          3660 => x"b00551ff",
          3661 => x"a48a3f93",
          3662 => x"397a5480",
          3663 => x"5382bff0",
          3664 => x"52b43dff",
          3665 => x"b00551ff",
          3666 => x"a3f63f82",
          3667 => x"d6ec5882",
          3668 => x"d8f85780",
          3669 => x"56645580",
          3670 => x"54848080",
          3671 => x"53848080",
          3672 => x"52b43dff",
          3673 => x"b00551e6",
          3674 => x"cc3f82d8",
          3675 => x"c80882d8",
          3676 => x"c8080970",
          3677 => x"30707207",
          3678 => x"8025515b",
          3679 => x"5b5f805a",
          3680 => x"7b832683",
          3681 => x"38815a78",
          3682 => x"7a065978",
          3683 => x"802e8d38",
          3684 => x"811c7081",
          3685 => x"ff065d59",
          3686 => x"7bfec338",
          3687 => x"7d81327d",
          3688 => x"81320759",
          3689 => x"788a387e",
          3690 => x"ff2e0981",
          3691 => x"06eeb338",
          3692 => x"82bff851",
          3693 => x"ffbcac3f",
          3694 => x"eea839f5",
          3695 => x"3d0d800b",
          3696 => x"82d8f834",
          3697 => x"87c0948c",
          3698 => x"70085455",
          3699 => x"87848052",
          3700 => x"7251d3af",
          3701 => x"3f82d8c8",
          3702 => x"08902b75",
          3703 => x"08555387",
          3704 => x"84805273",
          3705 => x"51d39c3f",
          3706 => x"7282d8c8",
          3707 => x"0807750c",
          3708 => x"87c0949c",
          3709 => x"70085455",
          3710 => x"87848052",
          3711 => x"7251d383",
          3712 => x"3f82d8c8",
          3713 => x"08902b75",
          3714 => x"08555387",
          3715 => x"84805273",
          3716 => x"51d2f03f",
          3717 => x"7282d8c8",
          3718 => x"0807750c",
          3719 => x"8c80830b",
          3720 => x"87c09484",
          3721 => x"0c8c8083",
          3722 => x"0b87c094",
          3723 => x"940c80fa",
          3724 => x"c05a80fd",
          3725 => x"ac5b8302",
          3726 => x"84059905",
          3727 => x"34805c82",
          3728 => x"f4a80b87",
          3729 => x"3d708813",
          3730 => x"0c70720c",
          3731 => x"82f4ac0c",
          3732 => x"5489be3f",
          3733 => x"93c03f82",
          3734 => x"c08851ff",
          3735 => x"bb853f82",
          3736 => x"c09451ff",
          3737 => x"bafd3f80",
          3738 => x"ddd55192",
          3739 => x"e33f8151",
          3740 => x"e8a63fec",
          3741 => x"9c3f8004",
          3742 => x"fe3d0d80",
          3743 => x"52835371",
          3744 => x"882b5287",
          3745 => x"d83f82d8",
          3746 => x"c80881ff",
          3747 => x"067207ff",
          3748 => x"14545272",
          3749 => x"8025e838",
          3750 => x"7182d8c8",
          3751 => x"0c843d0d",
          3752 => x"04fc3d0d",
          3753 => x"76700854",
          3754 => x"55807352",
          3755 => x"5472742e",
          3756 => x"818a3872",
          3757 => x"335170a0",
          3758 => x"2e098106",
          3759 => x"86388113",
          3760 => x"53f13972",
          3761 => x"335170a2",
          3762 => x"2e098106",
          3763 => x"86388113",
          3764 => x"53815472",
          3765 => x"5273812e",
          3766 => x"0981069f",
          3767 => x"38843981",
          3768 => x"12528072",
          3769 => x"33525470",
          3770 => x"a22e8338",
          3771 => x"81547080",
          3772 => x"2e9d3873",
          3773 => x"ea389839",
          3774 => x"81125280",
          3775 => x"72335254",
          3776 => x"70a02e83",
          3777 => x"38815470",
          3778 => x"802e8438",
          3779 => x"73ea3880",
          3780 => x"72335254",
          3781 => x"70a02e09",
          3782 => x"81068338",
          3783 => x"815470a2",
          3784 => x"32703070",
          3785 => x"80257607",
          3786 => x"51515170",
          3787 => x"802e8838",
          3788 => x"80727081",
          3789 => x"05543471",
          3790 => x"750c7251",
          3791 => x"7082d8c8",
          3792 => x"0c863d0d",
          3793 => x"04fc3d0d",
          3794 => x"76537208",
          3795 => x"802e9138",
          3796 => x"863dfc05",
          3797 => x"527251d3",
          3798 => x"a23f82d8",
          3799 => x"c8088538",
          3800 => x"80538339",
          3801 => x"74537282",
          3802 => x"d8c80c86",
          3803 => x"3d0d04fc",
          3804 => x"3d0d7682",
          3805 => x"1133ff05",
          3806 => x"52538152",
          3807 => x"708b2681",
          3808 => x"98388313",
          3809 => x"33ff0551",
          3810 => x"8252709e",
          3811 => x"26818a38",
          3812 => x"84133351",
          3813 => x"83527097",
          3814 => x"2680fe38",
          3815 => x"85133351",
          3816 => x"845270bb",
          3817 => x"2680f238",
          3818 => x"86133351",
          3819 => x"855270bb",
          3820 => x"2680e638",
          3821 => x"88132255",
          3822 => x"86527487",
          3823 => x"e72680d9",
          3824 => x"388a1322",
          3825 => x"54875273",
          3826 => x"87e72680",
          3827 => x"cc38810b",
          3828 => x"87c0989c",
          3829 => x"0c722287",
          3830 => x"c098bc0c",
          3831 => x"82133387",
          3832 => x"c098b80c",
          3833 => x"83133387",
          3834 => x"c098b40c",
          3835 => x"84133387",
          3836 => x"c098b00c",
          3837 => x"85133387",
          3838 => x"c098ac0c",
          3839 => x"86133387",
          3840 => x"c098a80c",
          3841 => x"7487c098",
          3842 => x"a40c7387",
          3843 => x"c098a00c",
          3844 => x"800b87c0",
          3845 => x"989c0c80",
          3846 => x"527182d8",
          3847 => x"c80c863d",
          3848 => x"0d04f33d",
          3849 => x"0d7f5b87",
          3850 => x"c0989c5d",
          3851 => x"817d0c87",
          3852 => x"c098bc08",
          3853 => x"5e7d7b23",
          3854 => x"87c098b8",
          3855 => x"085a7982",
          3856 => x"1c3487c0",
          3857 => x"98b4085a",
          3858 => x"79831c34",
          3859 => x"87c098b0",
          3860 => x"085a7984",
          3861 => x"1c3487c0",
          3862 => x"98ac085a",
          3863 => x"79851c34",
          3864 => x"87c098a8",
          3865 => x"085a7986",
          3866 => x"1c3487c0",
          3867 => x"98a4085c",
          3868 => x"7b881c23",
          3869 => x"87c098a0",
          3870 => x"085a798a",
          3871 => x"1c23807d",
          3872 => x"0c7983ff",
          3873 => x"ff06597b",
          3874 => x"83ffff06",
          3875 => x"58861b33",
          3876 => x"57851b33",
          3877 => x"56841b33",
          3878 => x"55831b33",
          3879 => x"54821b33",
          3880 => x"537d83ff",
          3881 => x"ff065282",
          3882 => x"c0ac51ff",
          3883 => x"9aaa3f8f",
          3884 => x"3d0d04fb",
          3885 => x"3d0d029f",
          3886 => x"053382d6",
          3887 => x"e8337081",
          3888 => x"ff065855",
          3889 => x"5587c094",
          3890 => x"84517580",
          3891 => x"2e863887",
          3892 => x"c0949451",
          3893 => x"70087096",
          3894 => x"2a708106",
          3895 => x"53545270",
          3896 => x"802e8c38",
          3897 => x"71912a70",
          3898 => x"81065151",
          3899 => x"70d73872",
          3900 => x"81327081",
          3901 => x"06515170",
          3902 => x"802e8d38",
          3903 => x"71932a70",
          3904 => x"81065151",
          3905 => x"70ffbe38",
          3906 => x"7381ff06",
          3907 => x"5187c094",
          3908 => x"80527080",
          3909 => x"2e863887",
          3910 => x"c0949052",
          3911 => x"74720c74",
          3912 => x"82d8c80c",
          3913 => x"873d0d04",
          3914 => x"ff3d0d02",
          3915 => x"8f053370",
          3916 => x"30709f2a",
          3917 => x"51525270",
          3918 => x"82d6e834",
          3919 => x"833d0d04",
          3920 => x"f93d0d02",
          3921 => x"a7053358",
          3922 => x"778a2e09",
          3923 => x"81068738",
          3924 => x"7a528d51",
          3925 => x"eb3f82d6",
          3926 => x"e8337081",
          3927 => x"ff065856",
          3928 => x"87c09484",
          3929 => x"5376802e",
          3930 => x"863887c0",
          3931 => x"94945372",
          3932 => x"0870962a",
          3933 => x"70810655",
          3934 => x"56547280",
          3935 => x"2e8c3873",
          3936 => x"912a7081",
          3937 => x"06515372",
          3938 => x"d7387481",
          3939 => x"32708106",
          3940 => x"51537280",
          3941 => x"2e8d3873",
          3942 => x"932a7081",
          3943 => x"06515372",
          3944 => x"ffbe3875",
          3945 => x"81ff0653",
          3946 => x"87c09480",
          3947 => x"5472802e",
          3948 => x"863887c0",
          3949 => x"94905477",
          3950 => x"740c800b",
          3951 => x"82d8c80c",
          3952 => x"893d0d04",
          3953 => x"f93d0d79",
          3954 => x"54807433",
          3955 => x"7081ff06",
          3956 => x"53535770",
          3957 => x"772e80fc",
          3958 => x"387181ff",
          3959 => x"06811582",
          3960 => x"d6e83370",
          3961 => x"81ff0659",
          3962 => x"57555887",
          3963 => x"c0948451",
          3964 => x"75802e86",
          3965 => x"3887c094",
          3966 => x"94517008",
          3967 => x"70962a70",
          3968 => x"81065354",
          3969 => x"5270802e",
          3970 => x"8c387191",
          3971 => x"2a708106",
          3972 => x"515170d7",
          3973 => x"38728132",
          3974 => x"70810651",
          3975 => x"5170802e",
          3976 => x"8d387193",
          3977 => x"2a708106",
          3978 => x"515170ff",
          3979 => x"be387481",
          3980 => x"ff065187",
          3981 => x"c0948052",
          3982 => x"70802e86",
          3983 => x"3887c094",
          3984 => x"90527772",
          3985 => x"0c811774",
          3986 => x"337081ff",
          3987 => x"06535357",
          3988 => x"70ff8638",
          3989 => x"7682d8c8",
          3990 => x"0c893d0d",
          3991 => x"04fe3d0d",
          3992 => x"82d6e833",
          3993 => x"7081ff06",
          3994 => x"545287c0",
          3995 => x"94845172",
          3996 => x"802e8638",
          3997 => x"87c09494",
          3998 => x"51700870",
          3999 => x"822a7081",
          4000 => x"06515151",
          4001 => x"70802ee2",
          4002 => x"387181ff",
          4003 => x"065187c0",
          4004 => x"94805270",
          4005 => x"802e8638",
          4006 => x"87c09490",
          4007 => x"52710870",
          4008 => x"81ff0682",
          4009 => x"d8c80c51",
          4010 => x"843d0d04",
          4011 => x"ffaf3f82",
          4012 => x"d8c80881",
          4013 => x"ff0682d8",
          4014 => x"c80c04fe",
          4015 => x"3d0d82d6",
          4016 => x"e8337081",
          4017 => x"ff065253",
          4018 => x"87c09484",
          4019 => x"5270802e",
          4020 => x"863887c0",
          4021 => x"94945271",
          4022 => x"0870822a",
          4023 => x"70810651",
          4024 => x"5151ff52",
          4025 => x"70802ea0",
          4026 => x"387281ff",
          4027 => x"065187c0",
          4028 => x"94805270",
          4029 => x"802e8638",
          4030 => x"87c09490",
          4031 => x"52710870",
          4032 => x"982b7098",
          4033 => x"2c515351",
          4034 => x"7182d8c8",
          4035 => x"0c843d0d",
          4036 => x"04ff3d0d",
          4037 => x"87c09e80",
          4038 => x"08709c2a",
          4039 => x"8a065151",
          4040 => x"70802e84",
          4041 => x"b43887c0",
          4042 => x"9ea40882",
          4043 => x"d6ec0c87",
          4044 => x"c09ea808",
          4045 => x"82d6f00c",
          4046 => x"87c09e94",
          4047 => x"0882d6f4",
          4048 => x"0c87c09e",
          4049 => x"980882d6",
          4050 => x"f80c87c0",
          4051 => x"9e9c0882",
          4052 => x"d6fc0c87",
          4053 => x"c09ea008",
          4054 => x"82d7800c",
          4055 => x"87c09eac",
          4056 => x"0882d784",
          4057 => x"0c87c09e",
          4058 => x"b00882d7",
          4059 => x"880c87c0",
          4060 => x"9eb40882",
          4061 => x"d78c0c87",
          4062 => x"c09eb808",
          4063 => x"82d7900c",
          4064 => x"87c09ebc",
          4065 => x"0882d794",
          4066 => x"0c87c09e",
          4067 => x"c00882d7",
          4068 => x"980c87c0",
          4069 => x"9ec40882",
          4070 => x"d79c0c87",
          4071 => x"c09e8008",
          4072 => x"517082d7",
          4073 => x"a02387c0",
          4074 => x"9e840882",
          4075 => x"d7a40c87",
          4076 => x"c09e8808",
          4077 => x"82d7a80c",
          4078 => x"87c09e8c",
          4079 => x"0882d7ac",
          4080 => x"0c810b82",
          4081 => x"d7b03480",
          4082 => x"0b87c09e",
          4083 => x"90087084",
          4084 => x"800a0651",
          4085 => x"52527080",
          4086 => x"2e833881",
          4087 => x"527182d7",
          4088 => x"b134800b",
          4089 => x"87c09e90",
          4090 => x"08708880",
          4091 => x"0a065152",
          4092 => x"5270802e",
          4093 => x"83388152",
          4094 => x"7182d7b2",
          4095 => x"34800b87",
          4096 => x"c09e9008",
          4097 => x"7090800a",
          4098 => x"06515252",
          4099 => x"70802e83",
          4100 => x"38815271",
          4101 => x"82d7b334",
          4102 => x"800b87c0",
          4103 => x"9e900870",
          4104 => x"88808006",
          4105 => x"51525270",
          4106 => x"802e8338",
          4107 => x"81527182",
          4108 => x"d7b43480",
          4109 => x"0b87c09e",
          4110 => x"900870a0",
          4111 => x"80800651",
          4112 => x"52527080",
          4113 => x"2e833881",
          4114 => x"527182d7",
          4115 => x"b534800b",
          4116 => x"87c09e90",
          4117 => x"08709080",
          4118 => x"80065152",
          4119 => x"5270802e",
          4120 => x"83388152",
          4121 => x"7182d7b6",
          4122 => x"34800b87",
          4123 => x"c09e9008",
          4124 => x"70848080",
          4125 => x"06515252",
          4126 => x"70802e83",
          4127 => x"38815271",
          4128 => x"82d7b734",
          4129 => x"800b87c0",
          4130 => x"9e900870",
          4131 => x"82808006",
          4132 => x"51525270",
          4133 => x"802e8338",
          4134 => x"81527182",
          4135 => x"d7b83480",
          4136 => x"0b87c09e",
          4137 => x"90087081",
          4138 => x"80800651",
          4139 => x"52527080",
          4140 => x"2e833881",
          4141 => x"527182d7",
          4142 => x"b934800b",
          4143 => x"87c09e90",
          4144 => x"087080c0",
          4145 => x"80065152",
          4146 => x"5270802e",
          4147 => x"83388152",
          4148 => x"7182d7ba",
          4149 => x"34800b87",
          4150 => x"c09e9008",
          4151 => x"70a08006",
          4152 => x"51525270",
          4153 => x"802e8338",
          4154 => x"81527182",
          4155 => x"d7bb3487",
          4156 => x"c09e9008",
          4157 => x"70988006",
          4158 => x"708a2a51",
          4159 => x"51517082",
          4160 => x"d7bc3480",
          4161 => x"0b87c09e",
          4162 => x"90087084",
          4163 => x"80065152",
          4164 => x"5270802e",
          4165 => x"83388152",
          4166 => x"7182d7bd",
          4167 => x"3487c09e",
          4168 => x"90087083",
          4169 => x"f0067084",
          4170 => x"2a515151",
          4171 => x"7082d7be",
          4172 => x"34800b87",
          4173 => x"c09e9008",
          4174 => x"70880651",
          4175 => x"52527080",
          4176 => x"2e833881",
          4177 => x"527182d7",
          4178 => x"bf3487c0",
          4179 => x"9e900870",
          4180 => x"87065151",
          4181 => x"7082d7c0",
          4182 => x"34833d0d",
          4183 => x"04fb3d0d",
          4184 => x"82c0c451",
          4185 => x"ff90f13f",
          4186 => x"82d7b033",
          4187 => x"5473802e",
          4188 => x"893882c0",
          4189 => x"d851ff90",
          4190 => x"df3f82c0",
          4191 => x"ec51ffac",
          4192 => x"e23f82d7",
          4193 => x"b2335473",
          4194 => x"802e9438",
          4195 => x"82d78c08",
          4196 => x"82d79008",
          4197 => x"11545282",
          4198 => x"c18451ff",
          4199 => x"90ba3f82",
          4200 => x"d7b73354",
          4201 => x"73802e94",
          4202 => x"3882d784",
          4203 => x"0882d788",
          4204 => x"08115452",
          4205 => x"82c1a051",
          4206 => x"ff909d3f",
          4207 => x"82d7b433",
          4208 => x"5473802e",
          4209 => x"943882d6",
          4210 => x"ec0882d6",
          4211 => x"f0081154",
          4212 => x"5282c1bc",
          4213 => x"51ff9080",
          4214 => x"3f82d7b5",
          4215 => x"33547380",
          4216 => x"2e943882",
          4217 => x"d6f40882",
          4218 => x"d6f80811",
          4219 => x"545282c1",
          4220 => x"d851ff8f",
          4221 => x"e33f82d7",
          4222 => x"b6335473",
          4223 => x"802e9438",
          4224 => x"82d6fc08",
          4225 => x"82d78008",
          4226 => x"11545282",
          4227 => x"c1f451ff",
          4228 => x"8fc63f82",
          4229 => x"d7bb3354",
          4230 => x"73802e8e",
          4231 => x"3882d7bc",
          4232 => x"335282c2",
          4233 => x"9051ff8f",
          4234 => x"af3f82d7",
          4235 => x"bf335473",
          4236 => x"802e8e38",
          4237 => x"82d7c033",
          4238 => x"5282c2b0",
          4239 => x"51ff8f98",
          4240 => x"3f82d7bd",
          4241 => x"33547380",
          4242 => x"2e8e3882",
          4243 => x"d7be3352",
          4244 => x"82c2d051",
          4245 => x"ff8f813f",
          4246 => x"82d7b133",
          4247 => x"5473802e",
          4248 => x"893882c2",
          4249 => x"f051ffaa",
          4250 => x"fa3f82d7",
          4251 => x"b3335473",
          4252 => x"802e8938",
          4253 => x"82c38451",
          4254 => x"ffaae83f",
          4255 => x"82d7b833",
          4256 => x"5473802e",
          4257 => x"893882c3",
          4258 => x"9051ffaa",
          4259 => x"d63f82d7",
          4260 => x"b9335473",
          4261 => x"802e8938",
          4262 => x"82c39c51",
          4263 => x"ffaac43f",
          4264 => x"82d7ba33",
          4265 => x"5473802e",
          4266 => x"893882c3",
          4267 => x"a451ffaa",
          4268 => x"b23f82c3",
          4269 => x"ac51ffaa",
          4270 => x"aa3f82d7",
          4271 => x"94085282",
          4272 => x"c3b851ff",
          4273 => x"8e923f82",
          4274 => x"d7980852",
          4275 => x"82c3e051",
          4276 => x"ff8e853f",
          4277 => x"82d79c08",
          4278 => x"5282c488",
          4279 => x"51ff8df8",
          4280 => x"3f82c4b0",
          4281 => x"51ffa9fb",
          4282 => x"3f82d7a0",
          4283 => x"225282c4",
          4284 => x"b851ff8d",
          4285 => x"e33f82d7",
          4286 => x"a40856bd",
          4287 => x"84c05275",
          4288 => x"51c1803f",
          4289 => x"82d8c808",
          4290 => x"bd84c029",
          4291 => x"76713154",
          4292 => x"5482d8c8",
          4293 => x"085282c4",
          4294 => x"e051ff8d",
          4295 => x"bb3f82d7",
          4296 => x"b7335473",
          4297 => x"802ea938",
          4298 => x"82d7a808",
          4299 => x"56bd84c0",
          4300 => x"527551c0",
          4301 => x"ce3f82d8",
          4302 => x"c808bd84",
          4303 => x"c0297671",
          4304 => x"31545482",
          4305 => x"d8c80852",
          4306 => x"82c58c51",
          4307 => x"ff8d893f",
          4308 => x"82d7b233",
          4309 => x"5473802e",
          4310 => x"a93882d7",
          4311 => x"ac0856bd",
          4312 => x"84c05275",
          4313 => x"51c09c3f",
          4314 => x"82d8c808",
          4315 => x"bd84c029",
          4316 => x"76713154",
          4317 => x"5482d8c8",
          4318 => x"085282c5",
          4319 => x"b851ff8c",
          4320 => x"d73f8a51",
          4321 => x"ffabfe3f",
          4322 => x"873d0d04",
          4323 => x"fe3d0d02",
          4324 => x"920533ff",
          4325 => x"05527184",
          4326 => x"26aa3871",
          4327 => x"842982af",
          4328 => x"c4055271",
          4329 => x"080482c5",
          4330 => x"e4519d39",
          4331 => x"82c5ec51",
          4332 => x"973982c5",
          4333 => x"f4519139",
          4334 => x"82c5fc51",
          4335 => x"8b3982c6",
          4336 => x"80518539",
          4337 => x"82c68851",
          4338 => x"ff8c8d3f",
          4339 => x"843d0d04",
          4340 => x"7188800c",
          4341 => x"04ff3d0d",
          4342 => x"87c09684",
          4343 => x"70085252",
          4344 => x"80720c70",
          4345 => x"74077082",
          4346 => x"d7c40c72",
          4347 => x"0c833d0d",
          4348 => x"04ff3d0d",
          4349 => x"87c09684",
          4350 => x"700882d7",
          4351 => x"c40c5280",
          4352 => x"720c7309",
          4353 => x"7082d7c4",
          4354 => x"08067082",
          4355 => x"d7c40c73",
          4356 => x"0c51833d",
          4357 => x"0d04800b",
          4358 => x"87c09684",
          4359 => x"0c0482d7",
          4360 => x"c40887c0",
          4361 => x"96840c04",
          4362 => x"fd3d0d76",
          4363 => x"982b7098",
          4364 => x"2c79982b",
          4365 => x"70982c72",
          4366 => x"10137082",
          4367 => x"2b515351",
          4368 => x"54515180",
          4369 => x"0b82c694",
          4370 => x"12335553",
          4371 => x"7174259c",
          4372 => x"3882c690",
          4373 => x"11081202",
          4374 => x"84059705",
          4375 => x"33713352",
          4376 => x"52527072",
          4377 => x"2e098106",
          4378 => x"83388153",
          4379 => x"7282d8c8",
          4380 => x"0c853d0d",
          4381 => x"04fb3d0d",
          4382 => x"79028405",
          4383 => x"a3053371",
          4384 => x"33555654",
          4385 => x"72802eb1",
          4386 => x"3882f4ac",
          4387 => x"08528851",
          4388 => x"ffaa9f3f",
          4389 => x"82f4ac08",
          4390 => x"52a051ff",
          4391 => x"aa943f82",
          4392 => x"f4ac0852",
          4393 => x"8851ffaa",
          4394 => x"893f7333",
          4395 => x"ff055372",
          4396 => x"74347281",
          4397 => x"ff0653cc",
          4398 => x"397751ff",
          4399 => x"8a9a3f74",
          4400 => x"7434873d",
          4401 => x"0d04f63d",
          4402 => x"0d7c0284",
          4403 => x"05b70533",
          4404 => x"028805bb",
          4405 => x"053382d8",
          4406 => x"a0337084",
          4407 => x"2982d7c8",
          4408 => x"05700851",
          4409 => x"59595a58",
          4410 => x"5974802e",
          4411 => x"86387451",
          4412 => x"9afa3f82",
          4413 => x"d8a03370",
          4414 => x"842982d7",
          4415 => x"c8058119",
          4416 => x"70545856",
          4417 => x"5a9dfb3f",
          4418 => x"82d8c808",
          4419 => x"750c82d8",
          4420 => x"a0337084",
          4421 => x"2982d7c8",
          4422 => x"05700851",
          4423 => x"565a7480",
          4424 => x"2ea73875",
          4425 => x"53785274",
          4426 => x"51ffb3b9",
          4427 => x"3f82d8a0",
          4428 => x"33810555",
          4429 => x"7482d8a0",
          4430 => x"347481ff",
          4431 => x"06559375",
          4432 => x"27873880",
          4433 => x"0b82d8a0",
          4434 => x"3477802e",
          4435 => x"b63882d8",
          4436 => x"9c085675",
          4437 => x"802eac38",
          4438 => x"82d89833",
          4439 => x"5574a438",
          4440 => x"8c3dfc05",
          4441 => x"54765378",
          4442 => x"52755180",
          4443 => x"ebbe3f82",
          4444 => x"d89c0852",
          4445 => x"8a5181a0",
          4446 => x"e73f82d8",
          4447 => x"9c085180",
          4448 => x"efa13f8c",
          4449 => x"3d0d04fd",
          4450 => x"3d0d82d7",
          4451 => x"c8539354",
          4452 => x"72085271",
          4453 => x"802e8938",
          4454 => x"715199d0",
          4455 => x"3f80730c",
          4456 => x"ff148414",
          4457 => x"54547380",
          4458 => x"25e63880",
          4459 => x"0b82d8a0",
          4460 => x"3482d89c",
          4461 => x"08527180",
          4462 => x"2e953871",
          4463 => x"5180f086",
          4464 => x"3f82d89c",
          4465 => x"085199a4",
          4466 => x"3f800b82",
          4467 => x"d89c0c85",
          4468 => x"3d0d04dc",
          4469 => x"3d0d8157",
          4470 => x"805282d8",
          4471 => x"9c085180",
          4472 => x"f5a23f82",
          4473 => x"d8c80880",
          4474 => x"d33882d8",
          4475 => x"9c085380",
          4476 => x"f852883d",
          4477 => x"70525681",
          4478 => x"9dd23f82",
          4479 => x"d8c80880",
          4480 => x"2eba3875",
          4481 => x"51ffaffd",
          4482 => x"3f82d8c8",
          4483 => x"0855800b",
          4484 => x"82d8c808",
          4485 => x"259d3882",
          4486 => x"d8c808ff",
          4487 => x"05701755",
          4488 => x"55807434",
          4489 => x"75537652",
          4490 => x"811782c9",
          4491 => x"845257ff",
          4492 => x"87a63f74",
          4493 => x"ff2e0981",
          4494 => x"06ffaf38",
          4495 => x"a63d0d04",
          4496 => x"d93d0daa",
          4497 => x"3d08ad3d",
          4498 => x"085a5a81",
          4499 => x"70585880",
          4500 => x"5282d89c",
          4501 => x"085180f4",
          4502 => x"ab3f82d8",
          4503 => x"c8088195",
          4504 => x"38ff0b82",
          4505 => x"d89c0854",
          4506 => x"5580f852",
          4507 => x"8b3d7052",
          4508 => x"56819cd8",
          4509 => x"3f82d8c8",
          4510 => x"08802ea5",
          4511 => x"387551ff",
          4512 => x"af833f82",
          4513 => x"d8c80881",
          4514 => x"18585580",
          4515 => x"0b82d8c8",
          4516 => x"08258e38",
          4517 => x"82d8c808",
          4518 => x"ff057017",
          4519 => x"55558074",
          4520 => x"34740970",
          4521 => x"30707207",
          4522 => x"9f2a5155",
          4523 => x"5578772e",
          4524 => x"853873ff",
          4525 => x"ac3882d8",
          4526 => x"9c088c11",
          4527 => x"08535180",
          4528 => x"f3c23f82",
          4529 => x"d8c80880",
          4530 => x"2e893882",
          4531 => x"c99051ff",
          4532 => x"86863f78",
          4533 => x"772e0981",
          4534 => x"069b3875",
          4535 => x"527951ff",
          4536 => x"af913f79",
          4537 => x"51ffae9d",
          4538 => x"3fab3d08",
          4539 => x"5482d8c8",
          4540 => x"08743480",
          4541 => x"587782d8",
          4542 => x"c80ca93d",
          4543 => x"0d04f63d",
          4544 => x"0d7c7e71",
          4545 => x"5c717233",
          4546 => x"57595a58",
          4547 => x"73a02e09",
          4548 => x"8106a238",
          4549 => x"78337805",
          4550 => x"56777627",
          4551 => x"98388117",
          4552 => x"705b7071",
          4553 => x"33565855",
          4554 => x"73a02e09",
          4555 => x"81068638",
          4556 => x"757526ea",
          4557 => x"38805473",
          4558 => x"882982d8",
          4559 => x"a4057008",
          4560 => x"5255ffad",
          4561 => x"c03f82d8",
          4562 => x"c8085379",
          4563 => x"52740851",
          4564 => x"ffb0bf3f",
          4565 => x"82d8c808",
          4566 => x"80c53884",
          4567 => x"15335574",
          4568 => x"812e8838",
          4569 => x"74822e88",
          4570 => x"38b539fc",
          4571 => x"e63fac39",
          4572 => x"811a5a8c",
          4573 => x"3dfc1153",
          4574 => x"f80551c0",
          4575 => x"cf3f82d8",
          4576 => x"c808802e",
          4577 => x"9a38ff1b",
          4578 => x"53785277",
          4579 => x"51fdb13f",
          4580 => x"82d8c808",
          4581 => x"81ff0655",
          4582 => x"74853874",
          4583 => x"54913981",
          4584 => x"147081ff",
          4585 => x"06515482",
          4586 => x"7427ff8b",
          4587 => x"38805473",
          4588 => x"82d8c80c",
          4589 => x"8c3d0d04",
          4590 => x"d33d0db0",
          4591 => x"3d08b23d",
          4592 => x"08b43d08",
          4593 => x"595f5a80",
          4594 => x"0baf3d34",
          4595 => x"82d8a033",
          4596 => x"82d89c08",
          4597 => x"555b7381",
          4598 => x"cb387382",
          4599 => x"d8983355",
          4600 => x"55738338",
          4601 => x"81557680",
          4602 => x"2e81bc38",
          4603 => x"81707606",
          4604 => x"55567380",
          4605 => x"2e81ad38",
          4606 => x"a8519886",
          4607 => x"3f82d8c8",
          4608 => x"0882d89c",
          4609 => x"0c82d8c8",
          4610 => x"08802e81",
          4611 => x"92389353",
          4612 => x"765282d8",
          4613 => x"c8085180",
          4614 => x"dead3f82",
          4615 => x"d8c80880",
          4616 => x"2e8c3882",
          4617 => x"c9bc51ff",
          4618 => x"9fb93f80",
          4619 => x"f73982d8",
          4620 => x"c8085b82",
          4621 => x"d89c0853",
          4622 => x"80f85290",
          4623 => x"3d705254",
          4624 => x"8199893f",
          4625 => x"82d8c808",
          4626 => x"5682d8c8",
          4627 => x"08742e09",
          4628 => x"810680d0",
          4629 => x"3882d8c8",
          4630 => x"0851ffab",
          4631 => x"a83f82d8",
          4632 => x"c8085580",
          4633 => x"0b82d8c8",
          4634 => x"0825a938",
          4635 => x"82d8c808",
          4636 => x"ff057017",
          4637 => x"55558074",
          4638 => x"34805374",
          4639 => x"81ff0652",
          4640 => x"7551f8c2",
          4641 => x"3f811b70",
          4642 => x"81ff065c",
          4643 => x"54937b27",
          4644 => x"8338805b",
          4645 => x"74ff2e09",
          4646 => x"8106ff97",
          4647 => x"38863975",
          4648 => x"82d89834",
          4649 => x"768c3882",
          4650 => x"d89c0880",
          4651 => x"2e8438f9",
          4652 => x"d63f8f3d",
          4653 => x"5dec843f",
          4654 => x"82d8c808",
          4655 => x"982b7098",
          4656 => x"2c515978",
          4657 => x"ff2eee38",
          4658 => x"7881ff06",
          4659 => x"82f08433",
          4660 => x"70982b70",
          4661 => x"982c82f0",
          4662 => x"80337098",
          4663 => x"2b70972c",
          4664 => x"71982c05",
          4665 => x"70842982",
          4666 => x"c6900570",
          4667 => x"08157033",
          4668 => x"51515151",
          4669 => x"59595159",
          4670 => x"5d588156",
          4671 => x"73782e80",
          4672 => x"e9387774",
          4673 => x"27b43874",
          4674 => x"81800a29",
          4675 => x"81ff0a05",
          4676 => x"70982c51",
          4677 => x"55807524",
          4678 => x"80ce3876",
          4679 => x"53745277",
          4680 => x"51f6853f",
          4681 => x"82d8c808",
          4682 => x"81ff0654",
          4683 => x"73802ed7",
          4684 => x"387482f0",
          4685 => x"80348156",
          4686 => x"b1397481",
          4687 => x"800a2981",
          4688 => x"800a0570",
          4689 => x"982c7081",
          4690 => x"ff065651",
          4691 => x"55739526",
          4692 => x"97387653",
          4693 => x"74527751",
          4694 => x"f5ce3f82",
          4695 => x"d8c80881",
          4696 => x"ff065473",
          4697 => x"cc38d339",
          4698 => x"80567580",
          4699 => x"2e80ca38",
          4700 => x"811c5574",
          4701 => x"82f08434",
          4702 => x"74982b70",
          4703 => x"982c82f0",
          4704 => x"80337098",
          4705 => x"2b70982c",
          4706 => x"70101170",
          4707 => x"822b82c6",
          4708 => x"9411335e",
          4709 => x"51515157",
          4710 => x"58515574",
          4711 => x"772e0981",
          4712 => x"06fe9238",
          4713 => x"82c69814",
          4714 => x"087d0c80",
          4715 => x"0b82f084",
          4716 => x"34800b82",
          4717 => x"f0803492",
          4718 => x"397582f0",
          4719 => x"84347582",
          4720 => x"f0803478",
          4721 => x"af3d3475",
          4722 => x"7d0c7e54",
          4723 => x"739526fd",
          4724 => x"e1387384",
          4725 => x"2982afd8",
          4726 => x"05547308",
          4727 => x"0482f08c",
          4728 => x"3354737e",
          4729 => x"2efdcb38",
          4730 => x"82f08833",
          4731 => x"55737527",
          4732 => x"ab387498",
          4733 => x"2b70982c",
          4734 => x"51557375",
          4735 => x"249e3874",
          4736 => x"1a547333",
          4737 => x"81153474",
          4738 => x"81800a29",
          4739 => x"81ff0a05",
          4740 => x"70982c82",
          4741 => x"f08c3356",
          4742 => x"5155df39",
          4743 => x"82f08c33",
          4744 => x"81115654",
          4745 => x"7482f08c",
          4746 => x"34731a54",
          4747 => x"ae3d3374",
          4748 => x"3482f088",
          4749 => x"3354737e",
          4750 => x"25893881",
          4751 => x"14547382",
          4752 => x"f0883482",
          4753 => x"f08c3370",
          4754 => x"81800a29",
          4755 => x"81ff0a05",
          4756 => x"70982c82",
          4757 => x"f088335a",
          4758 => x"51565674",
          4759 => x"7725a838",
          4760 => x"82f4ac08",
          4761 => x"52741a70",
          4762 => x"335254ff",
          4763 => x"9ec43f74",
          4764 => x"81800a29",
          4765 => x"81800a05",
          4766 => x"70982c82",
          4767 => x"f0883356",
          4768 => x"51557375",
          4769 => x"24da3882",
          4770 => x"f08c3370",
          4771 => x"982b7098",
          4772 => x"2c82f088",
          4773 => x"335a5156",
          4774 => x"56747725",
          4775 => x"fc943882",
          4776 => x"f4ac0852",
          4777 => x"8851ff9e",
          4778 => x"893f7481",
          4779 => x"800a2981",
          4780 => x"800a0570",
          4781 => x"982c82f0",
          4782 => x"88335651",
          4783 => x"55737524",
          4784 => x"de38fbee",
          4785 => x"39837a34",
          4786 => x"800b811b",
          4787 => x"3482f08c",
          4788 => x"53805282",
          4789 => x"b8b851f3",
          4790 => x"9c3f81fd",
          4791 => x"3982f08c",
          4792 => x"337081ff",
          4793 => x"06555573",
          4794 => x"802efbc6",
          4795 => x"3882f088",
          4796 => x"33ff0554",
          4797 => x"7382f088",
          4798 => x"34ff1554",
          4799 => x"7382f08c",
          4800 => x"3482f4ac",
          4801 => x"08528851",
          4802 => x"ff9da73f",
          4803 => x"82f08c33",
          4804 => x"70982b70",
          4805 => x"982c82f0",
          4806 => x"88335751",
          4807 => x"56577474",
          4808 => x"25ad3874",
          4809 => x"1a548114",
          4810 => x"33743482",
          4811 => x"f4ac0852",
          4812 => x"733351ff",
          4813 => x"9cfc3f74",
          4814 => x"81800a29",
          4815 => x"81800a05",
          4816 => x"70982c82",
          4817 => x"f0883358",
          4818 => x"51557575",
          4819 => x"24d53882",
          4820 => x"f4ac0852",
          4821 => x"a051ff9c",
          4822 => x"d93f82f0",
          4823 => x"8c337098",
          4824 => x"2b70982c",
          4825 => x"82f08833",
          4826 => x"57515657",
          4827 => x"747424fa",
          4828 => x"c13882f4",
          4829 => x"ac085288",
          4830 => x"51ff9cb6",
          4831 => x"3f748180",
          4832 => x"0a298180",
          4833 => x"0a057098",
          4834 => x"2c82f088",
          4835 => x"33585155",
          4836 => x"757525de",
          4837 => x"38fa9b39",
          4838 => x"82f08833",
          4839 => x"7a055480",
          4840 => x"743482f4",
          4841 => x"ac08528a",
          4842 => x"51ff9c86",
          4843 => x"3f82f088",
          4844 => x"527951f6",
          4845 => x"c93f82d8",
          4846 => x"c80881ff",
          4847 => x"06547396",
          4848 => x"3882f088",
          4849 => x"33547380",
          4850 => x"2e8f3881",
          4851 => x"53735279",
          4852 => x"51f1f33f",
          4853 => x"8439807a",
          4854 => x"34800b82",
          4855 => x"f08c3480",
          4856 => x"0b82f088",
          4857 => x"347982d8",
          4858 => x"c80caf3d",
          4859 => x"0d0482f0",
          4860 => x"8c335473",
          4861 => x"802ef9ba",
          4862 => x"3882f4ac",
          4863 => x"08528851",
          4864 => x"ff9baf3f",
          4865 => x"82f08c33",
          4866 => x"ff055473",
          4867 => x"82f08c34",
          4868 => x"7381ff06",
          4869 => x"54dd3982",
          4870 => x"f08c3382",
          4871 => x"f0883355",
          4872 => x"5573752e",
          4873 => x"f98c38ff",
          4874 => x"14547382",
          4875 => x"f0883474",
          4876 => x"982b7098",
          4877 => x"2c7581ff",
          4878 => x"06565155",
          4879 => x"747425ad",
          4880 => x"38741a54",
          4881 => x"81143374",
          4882 => x"3482f4ac",
          4883 => x"08527333",
          4884 => x"51ff9ade",
          4885 => x"3f748180",
          4886 => x"0a298180",
          4887 => x"0a057098",
          4888 => x"2c82f088",
          4889 => x"33585155",
          4890 => x"757524d5",
          4891 => x"3882f4ac",
          4892 => x"0852a051",
          4893 => x"ff9abb3f",
          4894 => x"82f08c33",
          4895 => x"70982b70",
          4896 => x"982c82f0",
          4897 => x"88335751",
          4898 => x"56577474",
          4899 => x"24f8a338",
          4900 => x"82f4ac08",
          4901 => x"528851ff",
          4902 => x"9a983f74",
          4903 => x"81800a29",
          4904 => x"81800a05",
          4905 => x"70982c82",
          4906 => x"f0883358",
          4907 => x"51557575",
          4908 => x"25de38f7",
          4909 => x"fd3982f0",
          4910 => x"8c337081",
          4911 => x"ff0682f0",
          4912 => x"88335956",
          4913 => x"54747727",
          4914 => x"f7e83882",
          4915 => x"f4ac0852",
          4916 => x"81145473",
          4917 => x"82f08c34",
          4918 => x"741a7033",
          4919 => x"5254ff99",
          4920 => x"d13f82f0",
          4921 => x"8c337081",
          4922 => x"ff0682f0",
          4923 => x"88335856",
          4924 => x"54757526",
          4925 => x"d638f7ba",
          4926 => x"3982f08c",
          4927 => x"53805282",
          4928 => x"b8b851ee",
          4929 => x"f03f800b",
          4930 => x"82f08c34",
          4931 => x"800b82f0",
          4932 => x"8834f79e",
          4933 => x"397ab038",
          4934 => x"82d89408",
          4935 => x"5574802e",
          4936 => x"a6387451",
          4937 => x"ffa1de3f",
          4938 => x"82d8c808",
          4939 => x"82f08834",
          4940 => x"82d8c808",
          4941 => x"81ff0681",
          4942 => x"05537452",
          4943 => x"7951ffa3",
          4944 => x"a43f935b",
          4945 => x"81c0397a",
          4946 => x"842982d7",
          4947 => x"c805fc11",
          4948 => x"08565474",
          4949 => x"802ea738",
          4950 => x"7451ffa1",
          4951 => x"a83f82d8",
          4952 => x"c80882f0",
          4953 => x"883482d8",
          4954 => x"c80881ff",
          4955 => x"06810553",
          4956 => x"74527951",
          4957 => x"ffa2ee3f",
          4958 => x"ff1b5480",
          4959 => x"fa397308",
          4960 => x"5574802e",
          4961 => x"f6ac3874",
          4962 => x"51ffa0f9",
          4963 => x"3f99397a",
          4964 => x"932e0981",
          4965 => x"06ae3882",
          4966 => x"d7c80855",
          4967 => x"74802ea4",
          4968 => x"387451ff",
          4969 => x"a0df3f82",
          4970 => x"d8c80882",
          4971 => x"f0883482",
          4972 => x"d8c80881",
          4973 => x"ff068105",
          4974 => x"53745279",
          4975 => x"51ffa2a5",
          4976 => x"3f80c339",
          4977 => x"7a842982",
          4978 => x"d7cc0570",
          4979 => x"08565474",
          4980 => x"802eab38",
          4981 => x"7451ffa0",
          4982 => x"ac3f82d8",
          4983 => x"c80882f0",
          4984 => x"883482d8",
          4985 => x"c80881ff",
          4986 => x"06810553",
          4987 => x"74527951",
          4988 => x"ffa1f23f",
          4989 => x"811b5473",
          4990 => x"81ff065b",
          4991 => x"89397482",
          4992 => x"f0883474",
          4993 => x"7a3482f0",
          4994 => x"8c5382f0",
          4995 => x"88335279",
          4996 => x"51ece23f",
          4997 => x"f59c3982",
          4998 => x"f08c3370",
          4999 => x"81ff0682",
          5000 => x"f0883359",
          5001 => x"56547477",
          5002 => x"27f58738",
          5003 => x"82f4ac08",
          5004 => x"52811454",
          5005 => x"7382f08c",
          5006 => x"34741a70",
          5007 => x"335254ff",
          5008 => x"96f03ff4",
          5009 => x"ed3982f0",
          5010 => x"8c335473",
          5011 => x"802ef4e2",
          5012 => x"3882f4ac",
          5013 => x"08528851",
          5014 => x"ff96d73f",
          5015 => x"82f08c33",
          5016 => x"ff055473",
          5017 => x"82f08c34",
          5018 => x"f4c839f9",
          5019 => x"3d0d83c0",
          5020 => x"800b82d8",
          5021 => x"c00c8480",
          5022 => x"0b82d8bc",
          5023 => x"23a08053",
          5024 => x"805283c0",
          5025 => x"8051ffa5",
          5026 => x"dd3f82d8",
          5027 => x"c0085480",
          5028 => x"58777434",
          5029 => x"81577681",
          5030 => x"153482d8",
          5031 => x"c0085477",
          5032 => x"84153476",
          5033 => x"85153482",
          5034 => x"d8c00854",
          5035 => x"77861534",
          5036 => x"76871534",
          5037 => x"82d8c008",
          5038 => x"82d8bc22",
          5039 => x"ff05fe80",
          5040 => x"80077083",
          5041 => x"ffff0670",
          5042 => x"882a5851",
          5043 => x"55567488",
          5044 => x"17347389",
          5045 => x"173482d8",
          5046 => x"bc227088",
          5047 => x"2982d8c0",
          5048 => x"0805f811",
          5049 => x"51555577",
          5050 => x"82153476",
          5051 => x"83153489",
          5052 => x"3d0d04ff",
          5053 => x"3d0d7352",
          5054 => x"81518472",
          5055 => x"278f38fb",
          5056 => x"12832a82",
          5057 => x"117083ff",
          5058 => x"ff065151",
          5059 => x"517082d8",
          5060 => x"c80c833d",
          5061 => x"0d04f93d",
          5062 => x"0d02a605",
          5063 => x"22028405",
          5064 => x"aa052271",
          5065 => x"0582d8c0",
          5066 => x"0871832b",
          5067 => x"71117483",
          5068 => x"2b731170",
          5069 => x"33811233",
          5070 => x"71882b07",
          5071 => x"02a405ae",
          5072 => x"05227181",
          5073 => x"ffff0607",
          5074 => x"70882a53",
          5075 => x"51525954",
          5076 => x"5b5b5753",
          5077 => x"54557177",
          5078 => x"34708118",
          5079 => x"3482d8c0",
          5080 => x"08147588",
          5081 => x"2a525470",
          5082 => x"82153474",
          5083 => x"83153482",
          5084 => x"d8c00870",
          5085 => x"17703381",
          5086 => x"12337188",
          5087 => x"2b077083",
          5088 => x"2b8ffff8",
          5089 => x"06515256",
          5090 => x"52710573",
          5091 => x"83ffff06",
          5092 => x"70882a54",
          5093 => x"54517182",
          5094 => x"12347281",
          5095 => x"ff065372",
          5096 => x"83123482",
          5097 => x"d8c00816",
          5098 => x"56717634",
          5099 => x"72811734",
          5100 => x"893d0d04",
          5101 => x"fb3d0d82",
          5102 => x"d8c00802",
          5103 => x"84059e05",
          5104 => x"2270832b",
          5105 => x"72118611",
          5106 => x"33871233",
          5107 => x"718b2b71",
          5108 => x"832b0758",
          5109 => x"5b595255",
          5110 => x"52720584",
          5111 => x"12338513",
          5112 => x"3371882b",
          5113 => x"0770882a",
          5114 => x"54565652",
          5115 => x"70841334",
          5116 => x"73851334",
          5117 => x"82d8c008",
          5118 => x"70148411",
          5119 => x"33851233",
          5120 => x"718b2b71",
          5121 => x"832b0756",
          5122 => x"59575272",
          5123 => x"05861233",
          5124 => x"87133371",
          5125 => x"882b0770",
          5126 => x"882a5456",
          5127 => x"56527086",
          5128 => x"13347387",
          5129 => x"133482d8",
          5130 => x"c0081370",
          5131 => x"33811233",
          5132 => x"71882b07",
          5133 => x"7081ffff",
          5134 => x"0670882a",
          5135 => x"53515353",
          5136 => x"53717334",
          5137 => x"70811434",
          5138 => x"873d0d04",
          5139 => x"fa3d0d02",
          5140 => x"a2052282",
          5141 => x"d8c00871",
          5142 => x"832b7111",
          5143 => x"70338112",
          5144 => x"3371882b",
          5145 => x"07708829",
          5146 => x"15703381",
          5147 => x"12337198",
          5148 => x"2b71902b",
          5149 => x"07535f53",
          5150 => x"55525a56",
          5151 => x"57535471",
          5152 => x"802580f6",
          5153 => x"387251fe",
          5154 => x"ab3f82d8",
          5155 => x"c0087016",
          5156 => x"70338112",
          5157 => x"33718b2b",
          5158 => x"71832b07",
          5159 => x"74117033",
          5160 => x"81123371",
          5161 => x"882b0770",
          5162 => x"832b8fff",
          5163 => x"f8065152",
          5164 => x"5451535a",
          5165 => x"58537205",
          5166 => x"74882a54",
          5167 => x"52728213",
          5168 => x"34738313",
          5169 => x"3482d8c0",
          5170 => x"08701670",
          5171 => x"33811233",
          5172 => x"718b2b71",
          5173 => x"832b0756",
          5174 => x"59575572",
          5175 => x"05703381",
          5176 => x"12337188",
          5177 => x"2b077081",
          5178 => x"ffff0670",
          5179 => x"882a5751",
          5180 => x"52585272",
          5181 => x"74347181",
          5182 => x"1534883d",
          5183 => x"0d04fb3d",
          5184 => x"0d82d8c0",
          5185 => x"08028405",
          5186 => x"9e052270",
          5187 => x"832b7211",
          5188 => x"82113383",
          5189 => x"1233718b",
          5190 => x"2b71832b",
          5191 => x"07595b59",
          5192 => x"52565273",
          5193 => x"05713381",
          5194 => x"13337188",
          5195 => x"2b07028c",
          5196 => x"05a20522",
          5197 => x"71077088",
          5198 => x"2a535153",
          5199 => x"53537173",
          5200 => x"34708114",
          5201 => x"3482d8c0",
          5202 => x"08701570",
          5203 => x"33811233",
          5204 => x"718b2b71",
          5205 => x"832b0756",
          5206 => x"59575272",
          5207 => x"05821233",
          5208 => x"83133371",
          5209 => x"882b0770",
          5210 => x"882a5455",
          5211 => x"56527082",
          5212 => x"13347283",
          5213 => x"133482d8",
          5214 => x"c0081482",
          5215 => x"11338312",
          5216 => x"3371882b",
          5217 => x"0782d8c8",
          5218 => x"0c525487",
          5219 => x"3d0d04f7",
          5220 => x"3d0d7b82",
          5221 => x"d8c00831",
          5222 => x"832a7083",
          5223 => x"ffff0670",
          5224 => x"535753fd",
          5225 => x"a73f82d8",
          5226 => x"c0087683",
          5227 => x"2b711182",
          5228 => x"11338312",
          5229 => x"33718b2b",
          5230 => x"71832b07",
          5231 => x"75117033",
          5232 => x"81123371",
          5233 => x"982b7190",
          5234 => x"2b075342",
          5235 => x"4051535b",
          5236 => x"58555954",
          5237 => x"7280258d",
          5238 => x"38828080",
          5239 => x"527551fe",
          5240 => x"9d3f8184",
          5241 => x"39841433",
          5242 => x"85153371",
          5243 => x"8b2b7183",
          5244 => x"2b077611",
          5245 => x"79882a53",
          5246 => x"51555855",
          5247 => x"76861434",
          5248 => x"7581ff06",
          5249 => x"56758714",
          5250 => x"3482d8c0",
          5251 => x"08701984",
          5252 => x"12338513",
          5253 => x"3371882b",
          5254 => x"0770882a",
          5255 => x"54575b56",
          5256 => x"53728416",
          5257 => x"34738516",
          5258 => x"3482d8c0",
          5259 => x"08185380",
          5260 => x"0b861434",
          5261 => x"800b8714",
          5262 => x"3482d8c0",
          5263 => x"08537684",
          5264 => x"14347585",
          5265 => x"143482d8",
          5266 => x"c0081870",
          5267 => x"33811233",
          5268 => x"71882b07",
          5269 => x"70828080",
          5270 => x"0770882a",
          5271 => x"53515556",
          5272 => x"54747434",
          5273 => x"72811534",
          5274 => x"8b3d0d04",
          5275 => x"ff3d0d73",
          5276 => x"5282d8c0",
          5277 => x"088438f7",
          5278 => x"f23f7180",
          5279 => x"2e863871",
          5280 => x"51fe8c3f",
          5281 => x"833d0d04",
          5282 => x"f53d0d80",
          5283 => x"7e5258f8",
          5284 => x"e23f82d8",
          5285 => x"c80883ff",
          5286 => x"ff0682d8",
          5287 => x"c0088411",
          5288 => x"33851233",
          5289 => x"71882b07",
          5290 => x"705f5956",
          5291 => x"585a81ff",
          5292 => x"ff597578",
          5293 => x"2e80cb38",
          5294 => x"75882917",
          5295 => x"70338112",
          5296 => x"3371882b",
          5297 => x"077081ff",
          5298 => x"ff067931",
          5299 => x"7083ffff",
          5300 => x"06707f27",
          5301 => x"52535156",
          5302 => x"59557779",
          5303 => x"278a3873",
          5304 => x"802e8538",
          5305 => x"75785a5b",
          5306 => x"84153385",
          5307 => x"16337188",
          5308 => x"2b075754",
          5309 => x"75c23878",
          5310 => x"81ffff2e",
          5311 => x"85387a79",
          5312 => x"59568076",
          5313 => x"832b82d8",
          5314 => x"c0081170",
          5315 => x"33811233",
          5316 => x"71882b07",
          5317 => x"7081ffff",
          5318 => x"0651525a",
          5319 => x"565c5573",
          5320 => x"752e8338",
          5321 => x"81558054",
          5322 => x"79782681",
          5323 => x"cc387454",
          5324 => x"74802e81",
          5325 => x"c438777a",
          5326 => x"2e098106",
          5327 => x"89387551",
          5328 => x"f8f23f81",
          5329 => x"ac398280",
          5330 => x"80537952",
          5331 => x"7551f7c6",
          5332 => x"3f82d8c0",
          5333 => x"08701c86",
          5334 => x"11338712",
          5335 => x"33718b2b",
          5336 => x"71832b07",
          5337 => x"535a5e55",
          5338 => x"74057a17",
          5339 => x"7083ffff",
          5340 => x"0670882a",
          5341 => x"5c595654",
          5342 => x"78841534",
          5343 => x"7681ff06",
          5344 => x"57768515",
          5345 => x"3482d8c0",
          5346 => x"0875832b",
          5347 => x"7111721e",
          5348 => x"86113387",
          5349 => x"12337188",
          5350 => x"2b077088",
          5351 => x"2a535b5e",
          5352 => x"535a5654",
          5353 => x"73861934",
          5354 => x"75871934",
          5355 => x"82d8c008",
          5356 => x"701c8411",
          5357 => x"33851233",
          5358 => x"718b2b71",
          5359 => x"832b0753",
          5360 => x"5d5a5574",
          5361 => x"05547886",
          5362 => x"15347687",
          5363 => x"153482d8",
          5364 => x"c0087016",
          5365 => x"711d8411",
          5366 => x"33851233",
          5367 => x"71882b07",
          5368 => x"70882a53",
          5369 => x"5a5f5256",
          5370 => x"54738416",
          5371 => x"34758516",
          5372 => x"3482d8c0",
          5373 => x"081b8405",
          5374 => x"547382d8",
          5375 => x"c80c8d3d",
          5376 => x"0d04fe3d",
          5377 => x"0d745282",
          5378 => x"d8c00884",
          5379 => x"38f4dc3f",
          5380 => x"71537180",
          5381 => x"2e8b3871",
          5382 => x"51fced3f",
          5383 => x"82d8c808",
          5384 => x"537282d8",
          5385 => x"c80c843d",
          5386 => x"0d04ee3d",
          5387 => x"0d646640",
          5388 => x"5c807042",
          5389 => x"4082d8c0",
          5390 => x"08602e09",
          5391 => x"81068438",
          5392 => x"f4a93f7b",
          5393 => x"8e387e51",
          5394 => x"ffb83f82",
          5395 => x"d8c80854",
          5396 => x"83c7397e",
          5397 => x"8b387b51",
          5398 => x"fc923f7e",
          5399 => x"5483ba39",
          5400 => x"7e51f58f",
          5401 => x"3f82d8c8",
          5402 => x"0883ffff",
          5403 => x"0682d8c0",
          5404 => x"087d7131",
          5405 => x"832a7083",
          5406 => x"ffff0670",
          5407 => x"832b7311",
          5408 => x"70338112",
          5409 => x"3371882b",
          5410 => x"07707531",
          5411 => x"7083ffff",
          5412 => x"06708829",
          5413 => x"fc057388",
          5414 => x"291a7033",
          5415 => x"81123371",
          5416 => x"882b0770",
          5417 => x"902b5344",
          5418 => x"4e534841",
          5419 => x"525c545b",
          5420 => x"415c565b",
          5421 => x"5b738025",
          5422 => x"8f387681",
          5423 => x"ffff0675",
          5424 => x"317083ff",
          5425 => x"ff064254",
          5426 => x"82163383",
          5427 => x"17337188",
          5428 => x"2b077088",
          5429 => x"291c7033",
          5430 => x"81123371",
          5431 => x"982b7190",
          5432 => x"2b075347",
          5433 => x"45525654",
          5434 => x"7380258b",
          5435 => x"38787531",
          5436 => x"7083ffff",
          5437 => x"06415477",
          5438 => x"7b2781fe",
          5439 => x"38601854",
          5440 => x"737b2e09",
          5441 => x"81068f38",
          5442 => x"7851f6c0",
          5443 => x"3f7a83ff",
          5444 => x"ff065881",
          5445 => x"e5397f8e",
          5446 => x"387a7424",
          5447 => x"89387851",
          5448 => x"f6aa3f81",
          5449 => x"a5397f18",
          5450 => x"557a7524",
          5451 => x"80c83879",
          5452 => x"1d821133",
          5453 => x"83123371",
          5454 => x"882b0753",
          5455 => x"5754f4f4",
          5456 => x"3f805278",
          5457 => x"51f7b73f",
          5458 => x"82d8c808",
          5459 => x"83ffff06",
          5460 => x"7e547c53",
          5461 => x"70832b82",
          5462 => x"d8c00811",
          5463 => x"84055355",
          5464 => x"59ff8eb7",
          5465 => x"3f82d8c0",
          5466 => x"08148405",
          5467 => x"7583ffff",
          5468 => x"06595c81",
          5469 => x"85396015",
          5470 => x"547a7424",
          5471 => x"80d43878",
          5472 => x"51f5c93f",
          5473 => x"82d8c008",
          5474 => x"1d821133",
          5475 => x"83123371",
          5476 => x"882b0753",
          5477 => x"4354f49c",
          5478 => x"3f805278",
          5479 => x"51f6df3f",
          5480 => x"82d8c808",
          5481 => x"83ffff06",
          5482 => x"7e547c53",
          5483 => x"70832b82",
          5484 => x"d8c00811",
          5485 => x"84055355",
          5486 => x"59ff8ddf",
          5487 => x"3f82d8c0",
          5488 => x"08148405",
          5489 => x"60620519",
          5490 => x"555c7383",
          5491 => x"ffff0658",
          5492 => x"a9397b7f",
          5493 => x"5254f9b0",
          5494 => x"3f82d8c8",
          5495 => x"085c82d8",
          5496 => x"c808802e",
          5497 => x"93387d53",
          5498 => x"735282d8",
          5499 => x"c80851ff",
          5500 => x"91f33f73",
          5501 => x"51f7983f",
          5502 => x"7a587a78",
          5503 => x"27993880",
          5504 => x"537a5278",
          5505 => x"51f28f3f",
          5506 => x"7a19832b",
          5507 => x"82d8c008",
          5508 => x"05840551",
          5509 => x"f6f93f7b",
          5510 => x"547382d8",
          5511 => x"c80c943d",
          5512 => x"0d04fc3d",
          5513 => x"0d777729",
          5514 => x"705254fb",
          5515 => x"d53f82d8",
          5516 => x"c8085582",
          5517 => x"d8c80880",
          5518 => x"2e8e3873",
          5519 => x"53805282",
          5520 => x"d8c80851",
          5521 => x"ff969f3f",
          5522 => x"7482d8c8",
          5523 => x"0c863d0d",
          5524 => x"04ff3d0d",
          5525 => x"028f0533",
          5526 => x"51815270",
          5527 => x"72268738",
          5528 => x"82d8c411",
          5529 => x"33527182",
          5530 => x"d8c80c83",
          5531 => x"3d0d04fc",
          5532 => x"3d0d029b",
          5533 => x"05330284",
          5534 => x"059f0533",
          5535 => x"56538351",
          5536 => x"72812680",
          5537 => x"e0387284",
          5538 => x"2b87c092",
          5539 => x"8c115351",
          5540 => x"88547480",
          5541 => x"2e843881",
          5542 => x"88547372",
          5543 => x"0c87c092",
          5544 => x"8c115181",
          5545 => x"710c850b",
          5546 => x"87c0988c",
          5547 => x"0c705271",
          5548 => x"08708206",
          5549 => x"51517080",
          5550 => x"2e8a3887",
          5551 => x"c0988c08",
          5552 => x"5170ec38",
          5553 => x"7108fc80",
          5554 => x"80065271",
          5555 => x"923887c0",
          5556 => x"988c0851",
          5557 => x"70802e87",
          5558 => x"387182d8",
          5559 => x"c4143482",
          5560 => x"d8c41333",
          5561 => x"517082d8",
          5562 => x"c80c863d",
          5563 => x"0d04f33d",
          5564 => x"0d606264",
          5565 => x"028c05bf",
          5566 => x"05335740",
          5567 => x"585b8374",
          5568 => x"525afecd",
          5569 => x"3f82d8c8",
          5570 => x"0881067a",
          5571 => x"54527181",
          5572 => x"be387172",
          5573 => x"75842b87",
          5574 => x"c0928011",
          5575 => x"87c0928c",
          5576 => x"1287c092",
          5577 => x"8413415a",
          5578 => x"40575a58",
          5579 => x"850b87c0",
          5580 => x"988c0c76",
          5581 => x"7d0c8476",
          5582 => x"0c750870",
          5583 => x"852a7081",
          5584 => x"06515354",
          5585 => x"71802e8e",
          5586 => x"387b0852",
          5587 => x"717b7081",
          5588 => x"055d3481",
          5589 => x"19598074",
          5590 => x"a2065353",
          5591 => x"71732e83",
          5592 => x"38815378",
          5593 => x"83ff268f",
          5594 => x"3872802e",
          5595 => x"8a3887c0",
          5596 => x"988c0852",
          5597 => x"71c33887",
          5598 => x"c0988c08",
          5599 => x"5271802e",
          5600 => x"87387884",
          5601 => x"802e9938",
          5602 => x"81760c87",
          5603 => x"c0928c15",
          5604 => x"53720870",
          5605 => x"82065152",
          5606 => x"71f738ff",
          5607 => x"1a5a8d39",
          5608 => x"84801781",
          5609 => x"197081ff",
          5610 => x"065a5357",
          5611 => x"79802e90",
          5612 => x"3873fc80",
          5613 => x"80065271",
          5614 => x"87387d78",
          5615 => x"26feed38",
          5616 => x"73fc8080",
          5617 => x"06527180",
          5618 => x"2e833881",
          5619 => x"52715372",
          5620 => x"82d8c80c",
          5621 => x"8f3d0d04",
          5622 => x"f33d0d60",
          5623 => x"6264028c",
          5624 => x"05bf0533",
          5625 => x"5740585b",
          5626 => x"83598074",
          5627 => x"5258fce1",
          5628 => x"3f82d8c8",
          5629 => x"08810679",
          5630 => x"54527178",
          5631 => x"2e098106",
          5632 => x"81b13877",
          5633 => x"74842b87",
          5634 => x"c0928011",
          5635 => x"87c0928c",
          5636 => x"1287c092",
          5637 => x"84134059",
          5638 => x"5f565a85",
          5639 => x"0b87c098",
          5640 => x"8c0c767d",
          5641 => x"0c82760c",
          5642 => x"80587508",
          5643 => x"70842a70",
          5644 => x"81065153",
          5645 => x"5471802e",
          5646 => x"8c387a70",
          5647 => x"81055c33",
          5648 => x"7c0c8118",
          5649 => x"5873812a",
          5650 => x"70810651",
          5651 => x"5271802e",
          5652 => x"8a3887c0",
          5653 => x"988c0852",
          5654 => x"71d03887",
          5655 => x"c0988c08",
          5656 => x"5271802e",
          5657 => x"87387784",
          5658 => x"802e9938",
          5659 => x"81760c87",
          5660 => x"c0928c15",
          5661 => x"53720870",
          5662 => x"82065152",
          5663 => x"71f738ff",
          5664 => x"19598d39",
          5665 => x"811a7081",
          5666 => x"ff068480",
          5667 => x"19595b52",
          5668 => x"78802e90",
          5669 => x"3873fc80",
          5670 => x"80065271",
          5671 => x"87387d7a",
          5672 => x"26fef838",
          5673 => x"73fc8080",
          5674 => x"06527180",
          5675 => x"2e833881",
          5676 => x"52715372",
          5677 => x"82d8c80c",
          5678 => x"8f3d0d04",
          5679 => x"fa3d0d7a",
          5680 => x"028405a3",
          5681 => x"05330288",
          5682 => x"05a70533",
          5683 => x"71545456",
          5684 => x"57fafe3f",
          5685 => x"82d8c808",
          5686 => x"81065383",
          5687 => x"547280fe",
          5688 => x"38850b87",
          5689 => x"c0988c0c",
          5690 => x"81567176",
          5691 => x"2e80dc38",
          5692 => x"71762493",
          5693 => x"3874842b",
          5694 => x"87c0928c",
          5695 => x"11545471",
          5696 => x"802e8d38",
          5697 => x"80d43971",
          5698 => x"832e80c6",
          5699 => x"3880cb39",
          5700 => x"72087081",
          5701 => x"2a708106",
          5702 => x"51515271",
          5703 => x"802e8a38",
          5704 => x"87c0988c",
          5705 => x"085271e8",
          5706 => x"3887c098",
          5707 => x"8c085271",
          5708 => x"96388173",
          5709 => x"0c87c092",
          5710 => x"8c145372",
          5711 => x"08708206",
          5712 => x"515271f7",
          5713 => x"38963980",
          5714 => x"56923988",
          5715 => x"800a770c",
          5716 => x"85398180",
          5717 => x"770c7256",
          5718 => x"83398456",
          5719 => x"75547382",
          5720 => x"d8c80c88",
          5721 => x"3d0d04fe",
          5722 => x"3d0d7481",
          5723 => x"11337133",
          5724 => x"71882b07",
          5725 => x"82d8c80c",
          5726 => x"5351843d",
          5727 => x"0d04fd3d",
          5728 => x"0d758311",
          5729 => x"33821233",
          5730 => x"71902b71",
          5731 => x"882b0781",
          5732 => x"14337072",
          5733 => x"07882b75",
          5734 => x"33710782",
          5735 => x"d8c80c52",
          5736 => x"53545654",
          5737 => x"52853d0d",
          5738 => x"04ff3d0d",
          5739 => x"73028405",
          5740 => x"92052252",
          5741 => x"52707270",
          5742 => x"81055434",
          5743 => x"70882a51",
          5744 => x"70723483",
          5745 => x"3d0d04ff",
          5746 => x"3d0d7375",
          5747 => x"52527072",
          5748 => x"70810554",
          5749 => x"3470882a",
          5750 => x"51707270",
          5751 => x"81055434",
          5752 => x"70882a51",
          5753 => x"70727081",
          5754 => x"05543470",
          5755 => x"882a5170",
          5756 => x"7234833d",
          5757 => x"0d04fe3d",
          5758 => x"0d767577",
          5759 => x"54545170",
          5760 => x"802e9238",
          5761 => x"71708105",
          5762 => x"53337370",
          5763 => x"81055534",
          5764 => x"ff1151eb",
          5765 => x"39843d0d",
          5766 => x"04fe3d0d",
          5767 => x"75777654",
          5768 => x"52537272",
          5769 => x"70810554",
          5770 => x"34ff1151",
          5771 => x"70f43884",
          5772 => x"3d0d04fc",
          5773 => x"3d0d7877",
          5774 => x"79565653",
          5775 => x"74708105",
          5776 => x"56337470",
          5777 => x"81055633",
          5778 => x"717131ff",
          5779 => x"16565252",
          5780 => x"5272802e",
          5781 => x"86387180",
          5782 => x"2ee23871",
          5783 => x"82d8c80c",
          5784 => x"863d0d04",
          5785 => x"fe3d0d74",
          5786 => x"76545189",
          5787 => x"3971732e",
          5788 => x"8a388111",
          5789 => x"51703352",
          5790 => x"71f33870",
          5791 => x"3382d8c8",
          5792 => x"0c843d0d",
          5793 => x"04800b82",
          5794 => x"d8c80c04",
          5795 => x"fb3d0d77",
          5796 => x"70087070",
          5797 => x"81055233",
          5798 => x"70545555",
          5799 => x"56e73fff",
          5800 => x"5582d8c8",
          5801 => x"08a23872",
          5802 => x"802e9838",
          5803 => x"83b55272",
          5804 => x"5180f7b6",
          5805 => x"3f82d8c8",
          5806 => x"0883ffff",
          5807 => x"06537280",
          5808 => x"2e863873",
          5809 => x"760c7255",
          5810 => x"7482d8c8",
          5811 => x"0c873d0d",
          5812 => x"04f73d0d",
          5813 => x"7b56800b",
          5814 => x"83173356",
          5815 => x"5a747a2e",
          5816 => x"80d63881",
          5817 => x"54b41608",
          5818 => x"53b81670",
          5819 => x"53811733",
          5820 => x"5259f9e4",
          5821 => x"3f82d8c8",
          5822 => x"087a2e09",
          5823 => x"8106b738",
          5824 => x"82d8c808",
          5825 => x"831734b4",
          5826 => x"160870a8",
          5827 => x"180831a0",
          5828 => x"18085956",
          5829 => x"58747727",
          5830 => x"9f388216",
          5831 => x"33557482",
          5832 => x"2e098106",
          5833 => x"93388154",
          5834 => x"76185378",
          5835 => x"52811633",
          5836 => x"51f9a53f",
          5837 => x"8339815a",
          5838 => x"7982d8c8",
          5839 => x"0c8b3d0d",
          5840 => x"04fa3d0d",
          5841 => x"787a5656",
          5842 => x"805774b4",
          5843 => x"17082eaf",
          5844 => x"387551fe",
          5845 => x"fc3f82d8",
          5846 => x"c8085782",
          5847 => x"d8c8089f",
          5848 => x"38815474",
          5849 => x"53b81652",
          5850 => x"81163351",
          5851 => x"f7803f82",
          5852 => x"d8c80880",
          5853 => x"2e8538ff",
          5854 => x"55815774",
          5855 => x"b4170c76",
          5856 => x"82d8c80c",
          5857 => x"883d0d04",
          5858 => x"f83d0d7a",
          5859 => x"705257fe",
          5860 => x"c03f82d8",
          5861 => x"c8085882",
          5862 => x"d8c80881",
          5863 => x"91387633",
          5864 => x"5574832e",
          5865 => x"09810680",
          5866 => x"f0388417",
          5867 => x"33597881",
          5868 => x"2e098106",
          5869 => x"80e33884",
          5870 => x"805382d8",
          5871 => x"c80852b8",
          5872 => x"17705256",
          5873 => x"fcd33f82",
          5874 => x"d4d55284",
          5875 => x"b61751fb",
          5876 => x"d83f848b",
          5877 => x"85a4d252",
          5878 => x"7551fbeb",
          5879 => x"3f868a85",
          5880 => x"e4f25284",
          5881 => x"9c1751fb",
          5882 => x"de3f9417",
          5883 => x"085284a0",
          5884 => x"1751fbd3",
          5885 => x"3f901708",
          5886 => x"5284a417",
          5887 => x"51fbc83f",
          5888 => x"a4170881",
          5889 => x"0570b419",
          5890 => x"0c795553",
          5891 => x"75528117",
          5892 => x"3351f7c4",
          5893 => x"3f778418",
          5894 => x"34805380",
          5895 => x"52811733",
          5896 => x"51f9993f",
          5897 => x"82d8c808",
          5898 => x"802e8338",
          5899 => x"81587782",
          5900 => x"d8c80c8a",
          5901 => x"3d0d04fb",
          5902 => x"3d0d77fe",
          5903 => x"1a9c1208",
          5904 => x"fe055556",
          5905 => x"54805674",
          5906 => x"73278d38",
          5907 => x"8a142275",
          5908 => x"7129b016",
          5909 => x"08055753",
          5910 => x"7582d8c8",
          5911 => x"0c873d0d",
          5912 => x"04f93d0d",
          5913 => x"7a7a7008",
          5914 => x"56545781",
          5915 => x"772781df",
          5916 => x"38769c15",
          5917 => x"082781d7",
          5918 => x"38ff7433",
          5919 => x"54587282",
          5920 => x"2e80f538",
          5921 => x"72822489",
          5922 => x"3872812e",
          5923 => x"8d3881bf",
          5924 => x"3972832e",
          5925 => x"818e3881",
          5926 => x"b6397681",
          5927 => x"2a177089",
          5928 => x"2aa81608",
          5929 => x"05537452",
          5930 => x"55fd963f",
          5931 => x"82d8c808",
          5932 => x"819f3874",
          5933 => x"83ff0614",
          5934 => x"b8113381",
          5935 => x"1770892a",
          5936 => x"a8180805",
          5937 => x"55765457",
          5938 => x"5753fcf5",
          5939 => x"3f82d8c8",
          5940 => x"0880fe38",
          5941 => x"7483ff06",
          5942 => x"14b81133",
          5943 => x"70882b78",
          5944 => x"07798106",
          5945 => x"71842a5c",
          5946 => x"52585153",
          5947 => x"7280e238",
          5948 => x"759fff06",
          5949 => x"5880da39",
          5950 => x"76882aa8",
          5951 => x"15080552",
          5952 => x"7351fcbd",
          5953 => x"3f82d8c8",
          5954 => x"0880c638",
          5955 => x"761083fe",
          5956 => x"067405b8",
          5957 => x"0551f8cf",
          5958 => x"3f82d8c8",
          5959 => x"0883ffff",
          5960 => x"0658ae39",
          5961 => x"76872aa8",
          5962 => x"15080552",
          5963 => x"7351fc91",
          5964 => x"3f82d8c8",
          5965 => x"089b3876",
          5966 => x"822b83fc",
          5967 => x"067405b8",
          5968 => x"0551f8ba",
          5969 => x"3f82d8c8",
          5970 => x"08f00a06",
          5971 => x"58833981",
          5972 => x"587782d8",
          5973 => x"c80c893d",
          5974 => x"0d04f83d",
          5975 => x"0d7a7c7e",
          5976 => x"5a585682",
          5977 => x"59817727",
          5978 => x"829e3876",
          5979 => x"9c170827",
          5980 => x"82963875",
          5981 => x"33537279",
          5982 => x"2e819d38",
          5983 => x"72792489",
          5984 => x"3872812e",
          5985 => x"8d388280",
          5986 => x"3972832e",
          5987 => x"81b83881",
          5988 => x"f7397681",
          5989 => x"2a177089",
          5990 => x"2aa81808",
          5991 => x"05537652",
          5992 => x"55fb9e3f",
          5993 => x"82d8c808",
          5994 => x"5982d8c8",
          5995 => x"0881d938",
          5996 => x"7483ff06",
          5997 => x"16b80581",
          5998 => x"16788106",
          5999 => x"59565477",
          6000 => x"5376802e",
          6001 => x"8f387784",
          6002 => x"2b9ff006",
          6003 => x"74338f06",
          6004 => x"71075153",
          6005 => x"72743481",
          6006 => x"0b831734",
          6007 => x"74892aa8",
          6008 => x"17080552",
          6009 => x"7551fad9",
          6010 => x"3f82d8c8",
          6011 => x"085982d8",
          6012 => x"c8088194",
          6013 => x"387483ff",
          6014 => x"0616b805",
          6015 => x"78842a54",
          6016 => x"54768f38",
          6017 => x"77882a74",
          6018 => x"3381f006",
          6019 => x"718f0607",
          6020 => x"51537274",
          6021 => x"3480ec39",
          6022 => x"76882aa8",
          6023 => x"17080552",
          6024 => x"7551fa9d",
          6025 => x"3f82d8c8",
          6026 => x"085982d8",
          6027 => x"c80880d8",
          6028 => x"387783ff",
          6029 => x"ff065276",
          6030 => x"1083fe06",
          6031 => x"7605b805",
          6032 => x"51f6e63f",
          6033 => x"be397687",
          6034 => x"2aa81708",
          6035 => x"05527551",
          6036 => x"f9ef3f82",
          6037 => x"d8c80859",
          6038 => x"82d8c808",
          6039 => x"ab3877f0",
          6040 => x"0a067782",
          6041 => x"2b83fc06",
          6042 => x"7018b805",
          6043 => x"70545154",
          6044 => x"54f68b3f",
          6045 => x"82d8c808",
          6046 => x"8f0a0674",
          6047 => x"07527251",
          6048 => x"f6c53f81",
          6049 => x"0b831734",
          6050 => x"7882d8c8",
          6051 => x"0c8a3d0d",
          6052 => x"04f83d0d",
          6053 => x"7a7c7e72",
          6054 => x"08595656",
          6055 => x"59817527",
          6056 => x"a438749c",
          6057 => x"1708279d",
          6058 => x"3873802e",
          6059 => x"aa38ff53",
          6060 => x"73527551",
          6061 => x"fda43f82",
          6062 => x"d8c80854",
          6063 => x"82d8c808",
          6064 => x"80f23893",
          6065 => x"39825480",
          6066 => x"eb398154",
          6067 => x"80e63982",
          6068 => x"d8c80854",
          6069 => x"80de3974",
          6070 => x"527851fb",
          6071 => x"843f82d8",
          6072 => x"c8085882",
          6073 => x"d8c80880",
          6074 => x"2e80c738",
          6075 => x"82d8c808",
          6076 => x"812ed238",
          6077 => x"82d8c808",
          6078 => x"ff2ecf38",
          6079 => x"80537452",
          6080 => x"7551fcd6",
          6081 => x"3f82d8c8",
          6082 => x"08c5389c",
          6083 => x"1608fe11",
          6084 => x"94180857",
          6085 => x"55577474",
          6086 => x"27903881",
          6087 => x"1594170c",
          6088 => x"84163381",
          6089 => x"07547384",
          6090 => x"17347755",
          6091 => x"767826ff",
          6092 => x"a6388054",
          6093 => x"7382d8c8",
          6094 => x"0c8a3d0d",
          6095 => x"04f63d0d",
          6096 => x"7c7e7108",
          6097 => x"595b5b79",
          6098 => x"95389017",
          6099 => x"08587780",
          6100 => x"2e88389c",
          6101 => x"17087826",
          6102 => x"b2388158",
          6103 => x"ae397952",
          6104 => x"7a51f9fd",
          6105 => x"3f815574",
          6106 => x"82d8c808",
          6107 => x"2782e038",
          6108 => x"82d8c808",
          6109 => x"5582d8c8",
          6110 => x"08ff2e82",
          6111 => x"d2389c17",
          6112 => x"0882d8c8",
          6113 => x"082682c7",
          6114 => x"38795894",
          6115 => x"17087056",
          6116 => x"5473802e",
          6117 => x"82b93877",
          6118 => x"7a2e0981",
          6119 => x"0680e238",
          6120 => x"811a569c",
          6121 => x"17087626",
          6122 => x"83388256",
          6123 => x"75527a51",
          6124 => x"f9af3f80",
          6125 => x"5982d8c8",
          6126 => x"08812e09",
          6127 => x"81068638",
          6128 => x"82d8c808",
          6129 => x"5982d8c8",
          6130 => x"08097030",
          6131 => x"70720780",
          6132 => x"25707c07",
          6133 => x"82d8c808",
          6134 => x"54515155",
          6135 => x"557381ef",
          6136 => x"3882d8c8",
          6137 => x"08802e95",
          6138 => x"38901708",
          6139 => x"54817427",
          6140 => x"9038739c",
          6141 => x"18082789",
          6142 => x"38735885",
          6143 => x"397580db",
          6144 => x"38775681",
          6145 => x"16569c17",
          6146 => x"08762689",
          6147 => x"38825675",
          6148 => x"782681ac",
          6149 => x"3875527a",
          6150 => x"51f8c63f",
          6151 => x"82d8c808",
          6152 => x"802eb838",
          6153 => x"805982d8",
          6154 => x"c808812e",
          6155 => x"09810686",
          6156 => x"3882d8c8",
          6157 => x"085982d8",
          6158 => x"c8080970",
          6159 => x"30707207",
          6160 => x"8025707c",
          6161 => x"07515155",
          6162 => x"557380f8",
          6163 => x"3875782e",
          6164 => x"098106ff",
          6165 => x"ae387355",
          6166 => x"80f539ff",
          6167 => x"53755276",
          6168 => x"51f9f73f",
          6169 => x"82d8c808",
          6170 => x"82d8c808",
          6171 => x"307082d8",
          6172 => x"c8080780",
          6173 => x"25515555",
          6174 => x"79802e94",
          6175 => x"3873802e",
          6176 => x"8f387553",
          6177 => x"79527651",
          6178 => x"f9d03f82",
          6179 => x"d8c80855",
          6180 => x"74a53875",
          6181 => x"90180c9c",
          6182 => x"1708fe05",
          6183 => x"94180856",
          6184 => x"54747426",
          6185 => x"8638ff15",
          6186 => x"94180c84",
          6187 => x"17338107",
          6188 => x"54738418",
          6189 => x"349739ff",
          6190 => x"5674812e",
          6191 => x"90388c39",
          6192 => x"80558c39",
          6193 => x"82d8c808",
          6194 => x"55853981",
          6195 => x"56755574",
          6196 => x"82d8c80c",
          6197 => x"8c3d0d04",
          6198 => x"f83d0d7a",
          6199 => x"705255f3",
          6200 => x"f03f82d8",
          6201 => x"c8085881",
          6202 => x"5682d8c8",
          6203 => x"0880d838",
          6204 => x"7b527451",
          6205 => x"f6c13f82",
          6206 => x"d8c80882",
          6207 => x"d8c808b4",
          6208 => x"170c5984",
          6209 => x"80537752",
          6210 => x"b8157052",
          6211 => x"57f28a3f",
          6212 => x"77568439",
          6213 => x"8116568a",
          6214 => x"15225875",
          6215 => x"78279738",
          6216 => x"81547519",
          6217 => x"53765281",
          6218 => x"153351ed",
          6219 => x"ab3f82d8",
          6220 => x"c808802e",
          6221 => x"df388a15",
          6222 => x"22763270",
          6223 => x"30707207",
          6224 => x"709f2a53",
          6225 => x"51565675",
          6226 => x"82d8c80c",
          6227 => x"8a3d0d04",
          6228 => x"f83d0d7a",
          6229 => x"7c710858",
          6230 => x"565774f0",
          6231 => x"800a2680",
          6232 => x"f138749f",
          6233 => x"06537280",
          6234 => x"e9387490",
          6235 => x"180c8817",
          6236 => x"085473aa",
          6237 => x"38753353",
          6238 => x"82732788",
          6239 => x"38ac1608",
          6240 => x"54739b38",
          6241 => x"74852a53",
          6242 => x"820b8817",
          6243 => x"225a5872",
          6244 => x"792780fe",
          6245 => x"38ac1608",
          6246 => x"98180c80",
          6247 => x"cd398a16",
          6248 => x"2270892b",
          6249 => x"54587275",
          6250 => x"26b23873",
          6251 => x"527651f5",
          6252 => x"b03f82d8",
          6253 => x"c8085482",
          6254 => x"d8c808ff",
          6255 => x"2ebd3881",
          6256 => x"0b82d8c8",
          6257 => x"08278b38",
          6258 => x"9c160882",
          6259 => x"d8c80826",
          6260 => x"85388258",
          6261 => x"bd397473",
          6262 => x"3155cb39",
          6263 => x"73527551",
          6264 => x"f4d53f82",
          6265 => x"d8c80898",
          6266 => x"180c7394",
          6267 => x"180c9817",
          6268 => x"08538258",
          6269 => x"72802e9a",
          6270 => x"38853981",
          6271 => x"58943974",
          6272 => x"892a1398",
          6273 => x"180c7483",
          6274 => x"ff0616b8",
          6275 => x"059c180c",
          6276 => x"80587782",
          6277 => x"d8c80c8a",
          6278 => x"3d0d04f8",
          6279 => x"3d0d7a70",
          6280 => x"08901208",
          6281 => x"a0055957",
          6282 => x"54f0800a",
          6283 => x"77278638",
          6284 => x"800b9815",
          6285 => x"0c981408",
          6286 => x"53845572",
          6287 => x"802e81cb",
          6288 => x"387683ff",
          6289 => x"06587781",
          6290 => x"b5388113",
          6291 => x"98150c94",
          6292 => x"14085574",
          6293 => x"92387685",
          6294 => x"2a881722",
          6295 => x"56537473",
          6296 => x"26819b38",
          6297 => x"80c0398a",
          6298 => x"1622ff05",
          6299 => x"77892a06",
          6300 => x"5372818a",
          6301 => x"38745273",
          6302 => x"51f3e63f",
          6303 => x"82d8c808",
          6304 => x"53825581",
          6305 => x"0b82d8c8",
          6306 => x"082780ff",
          6307 => x"38815582",
          6308 => x"d8c808ff",
          6309 => x"2e80f438",
          6310 => x"9c160882",
          6311 => x"d8c80826",
          6312 => x"80ca387b",
          6313 => x"8a387798",
          6314 => x"150c8455",
          6315 => x"80dd3994",
          6316 => x"14085273",
          6317 => x"51f9863f",
          6318 => x"82d8c808",
          6319 => x"53875582",
          6320 => x"d8c80880",
          6321 => x"2e80c438",
          6322 => x"825582d8",
          6323 => x"c808812e",
          6324 => x"ba388155",
          6325 => x"82d8c808",
          6326 => x"ff2eb038",
          6327 => x"82d8c808",
          6328 => x"527551fb",
          6329 => x"f33f82d8",
          6330 => x"c808a038",
          6331 => x"7294150c",
          6332 => x"72527551",
          6333 => x"f2c13f82",
          6334 => x"d8c80898",
          6335 => x"150c7690",
          6336 => x"150c7716",
          6337 => x"b8059c15",
          6338 => x"0c805574",
          6339 => x"82d8c80c",
          6340 => x"8a3d0d04",
          6341 => x"f73d0d7b",
          6342 => x"7d71085b",
          6343 => x"5b578052",
          6344 => x"7651fcac",
          6345 => x"3f82d8c8",
          6346 => x"085482d8",
          6347 => x"c80880ec",
          6348 => x"3882d8c8",
          6349 => x"08569817",
          6350 => x"08527851",
          6351 => x"f0833f82",
          6352 => x"d8c80854",
          6353 => x"82d8c808",
          6354 => x"80d23882",
          6355 => x"d8c8089c",
          6356 => x"18087033",
          6357 => x"51545872",
          6358 => x"81e52e09",
          6359 => x"81068338",
          6360 => x"815882d8",
          6361 => x"c8085572",
          6362 => x"83388155",
          6363 => x"77750753",
          6364 => x"72802e8e",
          6365 => x"38811656",
          6366 => x"757a2e09",
          6367 => x"81068838",
          6368 => x"a53982d8",
          6369 => x"c8085681",
          6370 => x"527651fd",
          6371 => x"8e3f82d8",
          6372 => x"c8085482",
          6373 => x"d8c80880",
          6374 => x"2eff9b38",
          6375 => x"73842e09",
          6376 => x"81068338",
          6377 => x"87547382",
          6378 => x"d8c80c8b",
          6379 => x"3d0d04fd",
          6380 => x"3d0d769a",
          6381 => x"115254eb",
          6382 => x"ae3f82d8",
          6383 => x"c80883ff",
          6384 => x"ff067670",
          6385 => x"33515353",
          6386 => x"71832e09",
          6387 => x"81069038",
          6388 => x"941451eb",
          6389 => x"923f82d8",
          6390 => x"c808902b",
          6391 => x"73075372",
          6392 => x"82d8c80c",
          6393 => x"853d0d04",
          6394 => x"fc3d0d77",
          6395 => x"797083ff",
          6396 => x"ff06549a",
          6397 => x"12535555",
          6398 => x"ebaf3f76",
          6399 => x"70335153",
          6400 => x"72832e09",
          6401 => x"81068b38",
          6402 => x"73902a52",
          6403 => x"941551eb",
          6404 => x"983f863d",
          6405 => x"0d04fd3d",
          6406 => x"0d755480",
          6407 => x"518b5370",
          6408 => x"812a7181",
          6409 => x"80290574",
          6410 => x"70810556",
          6411 => x"33710570",
          6412 => x"81ff06ff",
          6413 => x"16565151",
          6414 => x"5172e438",
          6415 => x"7082d8c8",
          6416 => x"0c853d0d",
          6417 => x"04f23d0d",
          6418 => x"60624059",
          6419 => x"8479085f",
          6420 => x"5b81ff70",
          6421 => x"5d5d9819",
          6422 => x"08802e83",
          6423 => x"80389819",
          6424 => x"08527d51",
          6425 => x"eddb3f82",
          6426 => x"d8c8085b",
          6427 => x"82d8c808",
          6428 => x"82eb389c",
          6429 => x"19087033",
          6430 => x"55557386",
          6431 => x"38845b82",
          6432 => x"dc398b15",
          6433 => x"33bf0670",
          6434 => x"81ff0658",
          6435 => x"5372861a",
          6436 => x"3482d8c8",
          6437 => x"08567381",
          6438 => x"e52e0981",
          6439 => x"06833881",
          6440 => x"5682d8c8",
          6441 => x"085373ae",
          6442 => x"2e098106",
          6443 => x"83388153",
          6444 => x"75730753",
          6445 => x"72993882",
          6446 => x"d8c80877",
          6447 => x"df065456",
          6448 => x"72882e09",
          6449 => x"81068338",
          6450 => x"8156757f",
          6451 => x"2e873881",
          6452 => x"ff5c81ef",
          6453 => x"39768f2e",
          6454 => x"09810681",
          6455 => x"ca387386",
          6456 => x"2a708106",
          6457 => x"51537280",
          6458 => x"2e92388d",
          6459 => x"15337481",
          6460 => x"bf067090",
          6461 => x"1c08ac1d",
          6462 => x"0c565d5d",
          6463 => x"737c2e09",
          6464 => x"8106819c",
          6465 => x"388d1533",
          6466 => x"537c732e",
          6467 => x"09810681",
          6468 => x"8f388c1e",
          6469 => x"089a1652",
          6470 => x"5ae8cc3f",
          6471 => x"82d8c808",
          6472 => x"83ffff06",
          6473 => x"537280f8",
          6474 => x"38743370",
          6475 => x"81bf068d",
          6476 => x"29f30551",
          6477 => x"54817b58",
          6478 => x"5882cad0",
          6479 => x"17337505",
          6480 => x"51e8a43f",
          6481 => x"82d8c808",
          6482 => x"83ffff06",
          6483 => x"5677802e",
          6484 => x"96387381",
          6485 => x"fe2680c8",
          6486 => x"3873101a",
          6487 => x"76595375",
          6488 => x"73238114",
          6489 => x"548b3975",
          6490 => x"83ffff2e",
          6491 => x"098106b0",
          6492 => x"38811757",
          6493 => x"8c7727c1",
          6494 => x"38743370",
          6495 => x"862a7081",
          6496 => x"06515455",
          6497 => x"72802e8e",
          6498 => x"387381fe",
          6499 => x"26923873",
          6500 => x"101a5380",
          6501 => x"7323ff1c",
          6502 => x"7081ff06",
          6503 => x"51538439",
          6504 => x"81ff5372",
          6505 => x"5c9d397b",
          6506 => x"93387451",
          6507 => x"fce83f82",
          6508 => x"d8c80881",
          6509 => x"ff065372",
          6510 => x"7d2ea738",
          6511 => x"ff0bac1a",
          6512 => x"0ca03980",
          6513 => x"527851f8",
          6514 => x"d23f82d8",
          6515 => x"c8085b82",
          6516 => x"d8c80889",
          6517 => x"38981908",
          6518 => x"fd843886",
          6519 => x"39800b98",
          6520 => x"1a0c7a82",
          6521 => x"d8c80c90",
          6522 => x"3d0d04f2",
          6523 => x"3d0d6070",
          6524 => x"08405980",
          6525 => x"527851f6",
          6526 => x"d73f82d8",
          6527 => x"c8085882",
          6528 => x"d8c80883",
          6529 => x"a43881ff",
          6530 => x"705f5cff",
          6531 => x"0bac1a0c",
          6532 => x"98190852",
          6533 => x"7e51eaa9",
          6534 => x"3f82d8c8",
          6535 => x"085882d8",
          6536 => x"c8088385",
          6537 => x"389c1908",
          6538 => x"70335757",
          6539 => x"75863884",
          6540 => x"5882f639",
          6541 => x"8b1733bf",
          6542 => x"067081ff",
          6543 => x"06565473",
          6544 => x"861a3475",
          6545 => x"81e52e82",
          6546 => x"c3387483",
          6547 => x"2a708106",
          6548 => x"5154748f",
          6549 => x"2e8e3873",
          6550 => x"82b23874",
          6551 => x"8f2e0981",
          6552 => x"0681f738",
          6553 => x"ab193370",
          6554 => x"862a7081",
          6555 => x"06515555",
          6556 => x"7382a138",
          6557 => x"75862a70",
          6558 => x"81065154",
          6559 => x"73802e92",
          6560 => x"388d1733",
          6561 => x"7681bf06",
          6562 => x"70901c08",
          6563 => x"ac1d0c58",
          6564 => x"5d5e757c",
          6565 => x"2e098106",
          6566 => x"81b9388d",
          6567 => x"1733567d",
          6568 => x"762e0981",
          6569 => x"0681ac38",
          6570 => x"8c1f089a",
          6571 => x"18525de5",
          6572 => x"b63f82d8",
          6573 => x"c80883ff",
          6574 => x"ff065574",
          6575 => x"81953876",
          6576 => x"3370bf06",
          6577 => x"8d29f305",
          6578 => x"59568175",
          6579 => x"5c5a82ca",
          6580 => x"d01b3377",
          6581 => x"0551e58f",
          6582 => x"3f82d8c8",
          6583 => x"0883ffff",
          6584 => x"06567980",
          6585 => x"2eb13877",
          6586 => x"81fe2680",
          6587 => x"e6387551",
          6588 => x"80dfb43f",
          6589 => x"82d8c808",
          6590 => x"78101e70",
          6591 => x"22535581",
          6592 => x"19595580",
          6593 => x"dfa13f74",
          6594 => x"82d8c808",
          6595 => x"2e098106",
          6596 => x"80c13875",
          6597 => x"5a8b3975",
          6598 => x"83ffff2e",
          6599 => x"098106b3",
          6600 => x"38811b5b",
          6601 => x"8c7b27ff",
          6602 => x"a5387633",
          6603 => x"70862a70",
          6604 => x"81065155",
          6605 => x"5779802e",
          6606 => x"90387380",
          6607 => x"2e8b3877",
          6608 => x"101d7022",
          6609 => x"5154738b",
          6610 => x"38ff1c70",
          6611 => x"81ff0651",
          6612 => x"54843981",
          6613 => x"ff54735c",
          6614 => x"bb397b93",
          6615 => x"387651f9",
          6616 => x"b53f82d8",
          6617 => x"c80881ff",
          6618 => x"0654737e",
          6619 => x"2ebb38ab",
          6620 => x"19338106",
          6621 => x"54739538",
          6622 => x"8b53a019",
          6623 => x"529c1908",
          6624 => x"51e5b03f",
          6625 => x"82d8c808",
          6626 => x"802e9e38",
          6627 => x"81ff5cff",
          6628 => x"0bac1a0c",
          6629 => x"80527851",
          6630 => x"f5813f82",
          6631 => x"d8c80858",
          6632 => x"82d8c808",
          6633 => x"802efce8",
          6634 => x"387782d8",
          6635 => x"c80c903d",
          6636 => x"0d04ee3d",
          6637 => x"0d647008",
          6638 => x"ab123381",
          6639 => x"a006565d",
          6640 => x"5a865573",
          6641 => x"85b53873",
          6642 => x"8c1d0870",
          6643 => x"2256565d",
          6644 => x"73802e8d",
          6645 => x"38811d70",
          6646 => x"10167022",
          6647 => x"51555df0",
          6648 => x"398c53a0",
          6649 => x"1a705392",
          6650 => x"3d70535f",
          6651 => x"59e4873f",
          6652 => x"0280cb05",
          6653 => x"33810654",
          6654 => x"73802e82",
          6655 => x"a83880c0",
          6656 => x"0bab1b34",
          6657 => x"815b8c1c",
          6658 => x"087b5658",
          6659 => x"8b537d52",
          6660 => x"7851e3e2",
          6661 => x"3f857b27",
          6662 => x"80c6387a",
          6663 => x"56772270",
          6664 => x"83ffff06",
          6665 => x"55557380",
          6666 => x"2eb43874",
          6667 => x"83ffff06",
          6668 => x"82195955",
          6669 => x"8f577481",
          6670 => x"06761007",
          6671 => x"75812a71",
          6672 => x"902a7081",
          6673 => x"06515656",
          6674 => x"5673802e",
          6675 => x"87387584",
          6676 => x"a0a13256",
          6677 => x"ff175776",
          6678 => x"8025db38",
          6679 => x"c0397555",
          6680 => x"87028405",
          6681 => x"bf055757",
          6682 => x"74b007bf",
          6683 => x"0654b974",
          6684 => x"27843887",
          6685 => x"14547376",
          6686 => x"34ff16ff",
          6687 => x"1876842a",
          6688 => x"57585674",
          6689 => x"e338943d",
          6690 => x"ec051754",
          6691 => x"80fe7434",
          6692 => x"807727b5",
          6693 => x"38783354",
          6694 => x"73a02ead",
          6695 => x"38741970",
          6696 => x"335254e3",
          6697 => x"e03f82d8",
          6698 => x"c808802e",
          6699 => x"8c38ff17",
          6700 => x"5474742e",
          6701 => x"94388115",
          6702 => x"55811555",
          6703 => x"74772789",
          6704 => x"38741970",
          6705 => x"335154d0",
          6706 => x"39943d77",
          6707 => x"05eb0554",
          6708 => x"78158116",
          6709 => x"5658a056",
          6710 => x"7687268a",
          6711 => x"38811781",
          6712 => x"15703358",
          6713 => x"55577578",
          6714 => x"34877527",
          6715 => x"e3387951",
          6716 => x"f9f93f82",
          6717 => x"d8c8088b",
          6718 => x"38811b5b",
          6719 => x"80e37b27",
          6720 => x"fe843887",
          6721 => x"557a80e4",
          6722 => x"2e82f038",
          6723 => x"82d8c808",
          6724 => x"5582d8c8",
          6725 => x"08842e09",
          6726 => x"810682df",
          6727 => x"380280cb",
          6728 => x"0533ab1b",
          6729 => x"340280cb",
          6730 => x"05337081",
          6731 => x"2a708106",
          6732 => x"51555e81",
          6733 => x"5973802e",
          6734 => x"90388d52",
          6735 => x"8c1d51fe",
          6736 => x"f4c13f82",
          6737 => x"d8c80819",
          6738 => x"59785279",
          6739 => x"51f3c53f",
          6740 => x"82d8c808",
          6741 => x"5782d8c8",
          6742 => x"08829e38",
          6743 => x"ff195978",
          6744 => x"802e81d4",
          6745 => x"3878852b",
          6746 => x"901b0871",
          6747 => x"31535479",
          6748 => x"51efdd3f",
          6749 => x"82d8c808",
          6750 => x"5782d8c8",
          6751 => x"0881fa38",
          6752 => x"a01a51f5",
          6753 => x"913f82d8",
          6754 => x"c80881ff",
          6755 => x"065d981a",
          6756 => x"08527b51",
          6757 => x"e3ab3f82",
          6758 => x"d8c80857",
          6759 => x"82d8c808",
          6760 => x"81d7388c",
          6761 => x"1c089c1b",
          6762 => x"087a81ff",
          6763 => x"065a575b",
          6764 => x"7c8d1734",
          6765 => x"8f0b8b17",
          6766 => x"3482d8c8",
          6767 => x"088c1734",
          6768 => x"82d8c808",
          6769 => x"529a1651",
          6770 => x"dfdf3f77",
          6771 => x"8d29f305",
          6772 => x"77555573",
          6773 => x"83ffff2e",
          6774 => x"8b387410",
          6775 => x"1b702281",
          6776 => x"17575154",
          6777 => x"735282ca",
          6778 => x"d0173376",
          6779 => x"0551dfb9",
          6780 => x"3f738538",
          6781 => x"83ffff54",
          6782 => x"8117578c",
          6783 => x"7727d438",
          6784 => x"7383ffff",
          6785 => x"2e8b3874",
          6786 => x"101b7022",
          6787 => x"51547386",
          6788 => x"387780c0",
          6789 => x"07587776",
          6790 => x"34810b83",
          6791 => x"1d348052",
          6792 => x"7951eff7",
          6793 => x"3f82d8c8",
          6794 => x"085782d8",
          6795 => x"c80880c9",
          6796 => x"38ff1959",
          6797 => x"78fed738",
          6798 => x"981a0852",
          6799 => x"7b51e281",
          6800 => x"3f82d8c8",
          6801 => x"085782d8",
          6802 => x"c808ae38",
          6803 => x"a05382d8",
          6804 => x"c808529c",
          6805 => x"1a0851df",
          6806 => x"c03f8b53",
          6807 => x"a01a529c",
          6808 => x"1a0851df",
          6809 => x"913f9c1a",
          6810 => x"08ab1b33",
          6811 => x"98065555",
          6812 => x"738c1634",
          6813 => x"810b831d",
          6814 => x"34765574",
          6815 => x"82d8c80c",
          6816 => x"943d0d04",
          6817 => x"fa3d0d78",
          6818 => x"70089012",
          6819 => x"08ac1308",
          6820 => x"56595755",
          6821 => x"72ff2e94",
          6822 => x"38725274",
          6823 => x"51edb13f",
          6824 => x"82d8c808",
          6825 => x"5482d8c8",
          6826 => x"0880c938",
          6827 => x"98150852",
          6828 => x"7551e18d",
          6829 => x"3f82d8c8",
          6830 => x"085482d8",
          6831 => x"c808ab38",
          6832 => x"9c150853",
          6833 => x"e5733481",
          6834 => x"0b831734",
          6835 => x"90150877",
          6836 => x"27a23882",
          6837 => x"d8c80852",
          6838 => x"7451eebf",
          6839 => x"3f82d8c8",
          6840 => x"085482d8",
          6841 => x"c808802e",
          6842 => x"c3387384",
          6843 => x"2e098106",
          6844 => x"83388254",
          6845 => x"7382d8c8",
          6846 => x"0c883d0d",
          6847 => x"04f43d0d",
          6848 => x"7e607108",
          6849 => x"5f595c80",
          6850 => x"0b961934",
          6851 => x"981c0880",
          6852 => x"2e83e238",
          6853 => x"ac1c08ff",
          6854 => x"2e81bb38",
          6855 => x"8070717f",
          6856 => x"8c050870",
          6857 => x"2257575b",
          6858 => x"5c577277",
          6859 => x"2e819d38",
          6860 => x"78101470",
          6861 => x"22811b5b",
          6862 => x"56537a97",
          6863 => x"3880d080",
          6864 => x"157083ff",
          6865 => x"ff065153",
          6866 => x"728fff26",
          6867 => x"8638745b",
          6868 => x"80df3976",
          6869 => x"18961181",
          6870 => x"ff793158",
          6871 => x"5b5483b5",
          6872 => x"527a902b",
          6873 => x"75075180",
          6874 => x"d5983f82",
          6875 => x"d8c80883",
          6876 => x"ffff0655",
          6877 => x"81ff7527",
          6878 => x"95388176",
          6879 => x"27a53874",
          6880 => x"882a5372",
          6881 => x"7a347497",
          6882 => x"15348255",
          6883 => x"9f397430",
          6884 => x"76307078",
          6885 => x"07802572",
          6886 => x"80250752",
          6887 => x"54547380",
          6888 => x"2e853880",
          6889 => x"579a3974",
          6890 => x"7a348155",
          6891 => x"74175780",
          6892 => x"5b8c1d08",
          6893 => x"79101170",
          6894 => x"22515454",
          6895 => x"72fef138",
          6896 => x"7a307080",
          6897 => x"25703079",
          6898 => x"06595153",
          6899 => x"77179405",
          6900 => x"53800b82",
          6901 => x"14348070",
          6902 => x"891a585a",
          6903 => x"579c1c08",
          6904 => x"19703381",
          6905 => x"1b5b5653",
          6906 => x"74a02eb7",
          6907 => x"3874852e",
          6908 => x"09810684",
          6909 => x"3881e555",
          6910 => x"78893270",
          6911 => x"30707207",
          6912 => x"80255154",
          6913 => x"54768b26",
          6914 => x"90387280",
          6915 => x"2e8b38ae",
          6916 => x"76708105",
          6917 => x"58348117",
          6918 => x"57747670",
          6919 => x"81055834",
          6920 => x"8117578a",
          6921 => x"7927ffb5",
          6922 => x"38771788",
          6923 => x"0553800b",
          6924 => x"81143496",
          6925 => x"18335372",
          6926 => x"81873876",
          6927 => x"8b38bf0b",
          6928 => x"96193481",
          6929 => x"5780e139",
          6930 => x"7273891a",
          6931 => x"33555a57",
          6932 => x"72802e80",
          6933 => x"d3389618",
          6934 => x"89195556",
          6935 => x"7333ffbf",
          6936 => x"11545572",
          6937 => x"9926aa38",
          6938 => x"9c1c088c",
          6939 => x"11335153",
          6940 => x"88792787",
          6941 => x"3872842a",
          6942 => x"53853972",
          6943 => x"832a5372",
          6944 => x"81065372",
          6945 => x"802e8a38",
          6946 => x"a0157083",
          6947 => x"ffff0656",
          6948 => x"53747670",
          6949 => x"81055834",
          6950 => x"81198115",
          6951 => x"81197133",
          6952 => x"56595559",
          6953 => x"72ffb538",
          6954 => x"77179405",
          6955 => x"53800b82",
          6956 => x"14349c1c",
          6957 => x"088c1133",
          6958 => x"51537285",
          6959 => x"38728919",
          6960 => x"349c1c08",
          6961 => x"538b1333",
          6962 => x"8819349c",
          6963 => x"1c089c11",
          6964 => x"5253d9aa",
          6965 => x"3f82d8c8",
          6966 => x"08780c96",
          6967 => x"1351d987",
          6968 => x"3f82d8c8",
          6969 => x"08861923",
          6970 => x"981351d8",
          6971 => x"fa3f82d8",
          6972 => x"c8088419",
          6973 => x"238e3d0d",
          6974 => x"04f03d0d",
          6975 => x"62700841",
          6976 => x"5e806470",
          6977 => x"33515555",
          6978 => x"73af2e83",
          6979 => x"38815573",
          6980 => x"80dc2e92",
          6981 => x"3874802e",
          6982 => x"8d387f98",
          6983 => x"0508881f",
          6984 => x"0caa3981",
          6985 => x"15448064",
          6986 => x"70335656",
          6987 => x"5673af2e",
          6988 => x"09810683",
          6989 => x"38815673",
          6990 => x"80dc3270",
          6991 => x"30708025",
          6992 => x"78075151",
          6993 => x"5473dc38",
          6994 => x"73881f0c",
          6995 => x"63703351",
          6996 => x"54739f26",
          6997 => x"9638ff80",
          6998 => x"0bab1f34",
          6999 => x"80527d51",
          7000 => x"e7ee3f82",
          7001 => x"d8c80856",
          7002 => x"87e13963",
          7003 => x"417d088c",
          7004 => x"11085b54",
          7005 => x"8059923d",
          7006 => x"fc0551da",
          7007 => x"8f3f82d8",
          7008 => x"c808ff2e",
          7009 => x"82b13883",
          7010 => x"ffff0b82",
          7011 => x"d8c80827",
          7012 => x"92387810",
          7013 => x"1a82d8c8",
          7014 => x"08902a55",
          7015 => x"55737523",
          7016 => x"81195982",
          7017 => x"d8c80883",
          7018 => x"ffff0670",
          7019 => x"af327030",
          7020 => x"9f732771",
          7021 => x"80250751",
          7022 => x"51555673",
          7023 => x"b4387580",
          7024 => x"dc2eae38",
          7025 => x"7580ff26",
          7026 => x"91387552",
          7027 => x"82c9ec51",
          7028 => x"d9923f82",
          7029 => x"d8c80881",
          7030 => x"de387881",
          7031 => x"fe2681d7",
          7032 => x"3878101a",
          7033 => x"54757423",
          7034 => x"811959ff",
          7035 => x"89398115",
          7036 => x"41806170",
          7037 => x"33565657",
          7038 => x"73af2e09",
          7039 => x"81068338",
          7040 => x"81577380",
          7041 => x"dc327030",
          7042 => x"70802579",
          7043 => x"07515154",
          7044 => x"73dc3874",
          7045 => x"449f7627",
          7046 => x"822b5778",
          7047 => x"812e0981",
          7048 => x"068c3879",
          7049 => x"225473ae",
          7050 => x"2ea53880",
          7051 => x"d2397882",
          7052 => x"2e098106",
          7053 => x"80c93882",
          7054 => x"1a225473",
          7055 => x"ae2e0981",
          7056 => x"0680c138",
          7057 => x"79225473",
          7058 => x"ae2e0981",
          7059 => x"06b63878",
          7060 => x"101a5480",
          7061 => x"7423800b",
          7062 => x"a01f5658",
          7063 => x"ae547878",
          7064 => x"268338a0",
          7065 => x"54737570",
          7066 => x"81055734",
          7067 => x"8118588a",
          7068 => x"7827e938",
          7069 => x"76a00754",
          7070 => x"73ab1f34",
          7071 => x"84c43978",
          7072 => x"802ea838",
          7073 => x"78101afe",
          7074 => x"05557422",
          7075 => x"fe167172",
          7076 => x"a0327030",
          7077 => x"709f2a51",
          7078 => x"51535856",
          7079 => x"5475ae2e",
          7080 => x"84387387",
          7081 => x"38ff1959",
          7082 => x"78e03878",
          7083 => x"197a1155",
          7084 => x"56807423",
          7085 => x"788d3886",
          7086 => x"56859039",
          7087 => x"76830757",
          7088 => x"83993980",
          7089 => x"7a227083",
          7090 => x"ffff0656",
          7091 => x"565d73a0",
          7092 => x"2e098106",
          7093 => x"9338811d",
          7094 => x"70101b70",
          7095 => x"2251555d",
          7096 => x"73a02ef2",
          7097 => x"387c8f38",
          7098 => x"7483ffff",
          7099 => x"065473ae",
          7100 => x"2e098106",
          7101 => x"85387683",
          7102 => x"07577880",
          7103 => x"2eaa3879",
          7104 => x"16fe0570",
          7105 => x"22515473",
          7106 => x"ae2e9d38",
          7107 => x"78101afe",
          7108 => x"0555ff19",
          7109 => x"5978802e",
          7110 => x"8f38fe15",
          7111 => x"70225555",
          7112 => x"73ae2e09",
          7113 => x"8106eb38",
          7114 => x"8b53a052",
          7115 => x"a01e51d5",
          7116 => x"e83f8070",
          7117 => x"595c885f",
          7118 => x"7c101a70",
          7119 => x"22811f5f",
          7120 => x"57547580",
          7121 => x"2e829438",
          7122 => x"75a02e96",
          7123 => x"3875ae32",
          7124 => x"70307080",
          7125 => x"25515154",
          7126 => x"7c792e8c",
          7127 => x"3873802e",
          7128 => x"89387683",
          7129 => x"0757d139",
          7130 => x"8054735b",
          7131 => x"7e782683",
          7132 => x"38815b7c",
          7133 => x"79327030",
          7134 => x"70720780",
          7135 => x"25707e07",
          7136 => x"51515555",
          7137 => x"73802ea6",
          7138 => x"387e8b2e",
          7139 => x"feae387c",
          7140 => x"792e8b38",
          7141 => x"76830757",
          7142 => x"7c792681",
          7143 => x"be38785d",
          7144 => x"88588b7c",
          7145 => x"822b81fc",
          7146 => x"065d5fff",
          7147 => x"8b3980ff",
          7148 => x"7627af38",
          7149 => x"76820757",
          7150 => x"83b55275",
          7151 => x"5180ccc2",
          7152 => x"3f82d8c8",
          7153 => x"0883ffff",
          7154 => x"0670872a",
          7155 => x"70810651",
          7156 => x"55567380",
          7157 => x"2e8c3875",
          7158 => x"80ff0682",
          7159 => x"cae01133",
          7160 => x"575481ff",
          7161 => x"7627a438",
          7162 => x"ff1f5473",
          7163 => x"78268a38",
          7164 => x"7683077f",
          7165 => x"5957fec0",
          7166 => x"397d18a0",
          7167 => x"0576882a",
          7168 => x"55557375",
          7169 => x"34811858",
          7170 => x"80c33975",
          7171 => x"802e9238",
          7172 => x"755282c9",
          7173 => x"f851d4cc",
          7174 => x"3f82d8c8",
          7175 => x"08802e8a",
          7176 => x"3880df77",
          7177 => x"83075856",
          7178 => x"a439ffbf",
          7179 => x"16547399",
          7180 => x"2685387b",
          7181 => x"82075cff",
          7182 => x"9f165473",
          7183 => x"99268e38",
          7184 => x"7b8107e0",
          7185 => x"177083ff",
          7186 => x"ff065855",
          7187 => x"5c7d18a0",
          7188 => x"05547574",
          7189 => x"34811858",
          7190 => x"fdde39a0",
          7191 => x"1e335473",
          7192 => x"81e52e09",
          7193 => x"81068638",
          7194 => x"850ba01f",
          7195 => x"347e882e",
          7196 => x"09810688",
          7197 => x"387b822b",
          7198 => x"81fc065c",
          7199 => x"7b8c0654",
          7200 => x"738c2e8d",
          7201 => x"387b8306",
          7202 => x"5473832e",
          7203 => x"09810685",
          7204 => x"38768207",
          7205 => x"5776812a",
          7206 => x"70810651",
          7207 => x"54739f38",
          7208 => x"7b810654",
          7209 => x"73802e85",
          7210 => x"38769007",
          7211 => x"577b822a",
          7212 => x"70810651",
          7213 => x"5473802e",
          7214 => x"85387688",
          7215 => x"075776ab",
          7216 => x"1f347d51",
          7217 => x"eaa53f82",
          7218 => x"d8c808ab",
          7219 => x"1f335656",
          7220 => x"82d8c808",
          7221 => x"802ebe38",
          7222 => x"82d8c808",
          7223 => x"842e0981",
          7224 => x"0680e838",
          7225 => x"74852a70",
          7226 => x"81067682",
          7227 => x"2a575154",
          7228 => x"73802e96",
          7229 => x"38748106",
          7230 => x"5473802e",
          7231 => x"f8ed38ff",
          7232 => x"800bab1f",
          7233 => x"34805680",
          7234 => x"c2397481",
          7235 => x"065473bb",
          7236 => x"388556b7",
          7237 => x"3974822a",
          7238 => x"70810651",
          7239 => x"5473ac38",
          7240 => x"861e3370",
          7241 => x"842a7081",
          7242 => x"06515555",
          7243 => x"73802ee1",
          7244 => x"38901e08",
          7245 => x"83ff0660",
          7246 => x"05b80552",
          7247 => x"7f51e4ef",
          7248 => x"3f82d8c8",
          7249 => x"08881f0c",
          7250 => x"f8a13975",
          7251 => x"82d8c80c",
          7252 => x"923d0d04",
          7253 => x"f63d0d7c",
          7254 => x"5bff7b08",
          7255 => x"70717355",
          7256 => x"595c5559",
          7257 => x"73802e81",
          7258 => x"c6387570",
          7259 => x"81055733",
          7260 => x"709f2652",
          7261 => x"5271ba2e",
          7262 => x"8d3870ee",
          7263 => x"3871ba2e",
          7264 => x"09810681",
          7265 => x"a5387333",
          7266 => x"d0117081",
          7267 => x"ff065152",
          7268 => x"53708926",
          7269 => x"91388214",
          7270 => x"7381ff06",
          7271 => x"d0055652",
          7272 => x"71762e80",
          7273 => x"f738800b",
          7274 => x"82cac059",
          7275 => x"5577087a",
          7276 => x"55577670",
          7277 => x"81055833",
          7278 => x"74708105",
          7279 => x"5633ff9f",
          7280 => x"12535353",
          7281 => x"70992689",
          7282 => x"38e01370",
          7283 => x"81ff0654",
          7284 => x"51ff9f12",
          7285 => x"51709926",
          7286 => x"8938e012",
          7287 => x"7081ff06",
          7288 => x"53517230",
          7289 => x"709f2a51",
          7290 => x"5172722e",
          7291 => x"09810685",
          7292 => x"3870ffbe",
          7293 => x"38723074",
          7294 => x"77327030",
          7295 => x"7072079f",
          7296 => x"2a739f2a",
          7297 => x"07535454",
          7298 => x"5170802e",
          7299 => x"8f388115",
          7300 => x"84195955",
          7301 => x"837525ff",
          7302 => x"94388b39",
          7303 => x"74832486",
          7304 => x"3874767c",
          7305 => x"0c597851",
          7306 => x"863982f0",
          7307 => x"a4335170",
          7308 => x"82d8c80c",
          7309 => x"8c3d0d04",
          7310 => x"fa3d0d78",
          7311 => x"56800b83",
          7312 => x"1734ff0b",
          7313 => x"b4170c79",
          7314 => x"527551d1",
          7315 => x"f43f8455",
          7316 => x"82d8c808",
          7317 => x"81803884",
          7318 => x"b61651ce",
          7319 => x"8a3f82d8",
          7320 => x"c80883ff",
          7321 => x"ff065483",
          7322 => x"557382d4",
          7323 => x"d52e0981",
          7324 => x"0680e338",
          7325 => x"800bb817",
          7326 => x"33565774",
          7327 => x"81e92e09",
          7328 => x"81068338",
          7329 => x"81577481",
          7330 => x"eb327030",
          7331 => x"70802579",
          7332 => x"07515154",
          7333 => x"738a3874",
          7334 => x"81e82e09",
          7335 => x"8106b538",
          7336 => x"835382ca",
          7337 => x"805280ee",
          7338 => x"1651cf87",
          7339 => x"3f82d8c8",
          7340 => x"085582d8",
          7341 => x"c808802e",
          7342 => x"9d388553",
          7343 => x"82ca8452",
          7344 => x"818a1651",
          7345 => x"ceed3f82",
          7346 => x"d8c80855",
          7347 => x"82d8c808",
          7348 => x"802e8338",
          7349 => x"82557482",
          7350 => x"d8c80c88",
          7351 => x"3d0d04f2",
          7352 => x"3d0d6102",
          7353 => x"840580cb",
          7354 => x"05335855",
          7355 => x"80750c60",
          7356 => x"51fce13f",
          7357 => x"82d8c808",
          7358 => x"588b5680",
          7359 => x"0b82d8c8",
          7360 => x"08248784",
          7361 => x"3882d8c8",
          7362 => x"08842982",
          7363 => x"f0900570",
          7364 => x"0855538c",
          7365 => x"5673802e",
          7366 => x"86ee3873",
          7367 => x"750c7681",
          7368 => x"fe067433",
          7369 => x"54577280",
          7370 => x"2eae3881",
          7371 => x"143351c6",
          7372 => x"a03f82d8",
          7373 => x"c80881ff",
          7374 => x"06708106",
          7375 => x"54557298",
          7376 => x"3876802e",
          7377 => x"86c03874",
          7378 => x"822a7081",
          7379 => x"0651538a",
          7380 => x"567286b4",
          7381 => x"3886af39",
          7382 => x"80743477",
          7383 => x"81153481",
          7384 => x"52811433",
          7385 => x"51c6883f",
          7386 => x"82d8c808",
          7387 => x"81ff0670",
          7388 => x"81065455",
          7389 => x"83567286",
          7390 => x"8f387680",
          7391 => x"2e8f3874",
          7392 => x"822a7081",
          7393 => x"0651538a",
          7394 => x"567285fc",
          7395 => x"38807053",
          7396 => x"74525bfd",
          7397 => x"a33f82d8",
          7398 => x"c80881ff",
          7399 => x"06577682",
          7400 => x"2e098106",
          7401 => x"80e2388c",
          7402 => x"3d745658",
          7403 => x"835683fa",
          7404 => x"15337058",
          7405 => x"5372802e",
          7406 => x"8d3883fe",
          7407 => x"1551cbbe",
          7408 => x"3f82d8c8",
          7409 => x"08577678",
          7410 => x"7084055a",
          7411 => x"0cff1690",
          7412 => x"16565675",
          7413 => x"8025d738",
          7414 => x"800b8d3d",
          7415 => x"54567270",
          7416 => x"84055408",
          7417 => x"5b83577a",
          7418 => x"802e9538",
          7419 => x"7a527351",
          7420 => x"fcc63f82",
          7421 => x"d8c80881",
          7422 => x"ff065781",
          7423 => x"77278938",
          7424 => x"81165683",
          7425 => x"7627d738",
          7426 => x"81567684",
          7427 => x"2e84f938",
          7428 => x"8d567681",
          7429 => x"2684f138",
          7430 => x"80c31451",
          7431 => x"cac93f82",
          7432 => x"d8c80883",
          7433 => x"ffff0653",
          7434 => x"7284802e",
          7435 => x"09810684",
          7436 => x"d73880ce",
          7437 => x"1451caaf",
          7438 => x"3f82d8c8",
          7439 => x"0883ffff",
          7440 => x"0658778d",
          7441 => x"3880dc14",
          7442 => x"51cab33f",
          7443 => x"82d8c808",
          7444 => x"5877a015",
          7445 => x"0c80c814",
          7446 => x"33821534",
          7447 => x"80c81433",
          7448 => x"ff117081",
          7449 => x"ff065154",
          7450 => x"558d5672",
          7451 => x"81268498",
          7452 => x"387481ff",
          7453 => x"06787129",
          7454 => x"80c51633",
          7455 => x"52595372",
          7456 => x"8a152372",
          7457 => x"802e8b38",
          7458 => x"ff137306",
          7459 => x"5372802e",
          7460 => x"86388d56",
          7461 => x"83f23980",
          7462 => x"c91451c9",
          7463 => x"ca3f82d8",
          7464 => x"c8085382",
          7465 => x"d8c80888",
          7466 => x"1523728f",
          7467 => x"06578d56",
          7468 => x"7683d538",
          7469 => x"80cb1451",
          7470 => x"c9ad3f82",
          7471 => x"d8c80883",
          7472 => x"ffff0655",
          7473 => x"748d3880",
          7474 => x"d81451c9",
          7475 => x"b13f82d8",
          7476 => x"c8085580",
          7477 => x"c61451c9",
          7478 => x"8e3f82d8",
          7479 => x"c80883ff",
          7480 => x"ff06538d",
          7481 => x"5672802e",
          7482 => x"839e3888",
          7483 => x"14227814",
          7484 => x"71842a05",
          7485 => x"5a5a7875",
          7486 => x"26838d38",
          7487 => x"8a142252",
          7488 => x"74793151",
          7489 => x"fedcfc3f",
          7490 => x"82d8c808",
          7491 => x"5582d8c8",
          7492 => x"08802e82",
          7493 => x"f33882d8",
          7494 => x"c80880ff",
          7495 => x"fffff526",
          7496 => x"83388357",
          7497 => x"7483fff5",
          7498 => x"26833882",
          7499 => x"57749ff5",
          7500 => x"26853881",
          7501 => x"5789398d",
          7502 => x"5676802e",
          7503 => x"82ca3882",
          7504 => x"15709c16",
          7505 => x"0c7ba416",
          7506 => x"0c731c70",
          7507 => x"a8170c7a",
          7508 => x"1db0170c",
          7509 => x"54557683",
          7510 => x"2e098106",
          7511 => x"af3880e2",
          7512 => x"1451c883",
          7513 => x"3f82d8c8",
          7514 => x"0883ffff",
          7515 => x"06538d56",
          7516 => x"72829538",
          7517 => x"79829138",
          7518 => x"80e41451",
          7519 => x"c8803f82",
          7520 => x"d8c808ac",
          7521 => x"150c7482",
          7522 => x"2b53a239",
          7523 => x"8d567980",
          7524 => x"2e81f538",
          7525 => x"7713ac15",
          7526 => x"0c741553",
          7527 => x"76822e8d",
          7528 => x"38741015",
          7529 => x"70812a76",
          7530 => x"81060551",
          7531 => x"5383ff13",
          7532 => x"892a538d",
          7533 => x"5672a015",
          7534 => x"082681cc",
          7535 => x"38ff0b94",
          7536 => x"150cff0b",
          7537 => x"90150cff",
          7538 => x"800b8415",
          7539 => x"3476832e",
          7540 => x"09810681",
          7541 => x"923880e8",
          7542 => x"1451c78b",
          7543 => x"3f82d8c8",
          7544 => x"0883ffff",
          7545 => x"06537281",
          7546 => x"2e098106",
          7547 => x"80f93881",
          7548 => x"1b527351",
          7549 => x"cacb3f82",
          7550 => x"d8c80880",
          7551 => x"ea3882d8",
          7552 => x"c8088415",
          7553 => x"3484b614",
          7554 => x"51c6dc3f",
          7555 => x"82d8c808",
          7556 => x"83ffff06",
          7557 => x"537282d4",
          7558 => x"d52e0981",
          7559 => x"0680c838",
          7560 => x"b81451c6",
          7561 => x"d93f82d8",
          7562 => x"c808848b",
          7563 => x"85a4d22e",
          7564 => x"098106b3",
          7565 => x"38849c14",
          7566 => x"51c6c33f",
          7567 => x"82d8c808",
          7568 => x"868a85e4",
          7569 => x"f22e0981",
          7570 => x"069d3884",
          7571 => x"a01451c6",
          7572 => x"ad3f82d8",
          7573 => x"c8089415",
          7574 => x"0c84a414",
          7575 => x"51c69f3f",
          7576 => x"82d8c808",
          7577 => x"90150c76",
          7578 => x"743482f0",
          7579 => x"a0228105",
          7580 => x"537282f0",
          7581 => x"a0237286",
          7582 => x"152382f0",
          7583 => x"a80b8c15",
          7584 => x"0c800b98",
          7585 => x"150c8056",
          7586 => x"7582d8c8",
          7587 => x"0c903d0d",
          7588 => x"04fb3d0d",
          7589 => x"77548955",
          7590 => x"73802eba",
          7591 => x"38730853",
          7592 => x"72802eb2",
          7593 => x"38723352",
          7594 => x"71802eaa",
          7595 => x"38861322",
          7596 => x"84152257",
          7597 => x"5271762e",
          7598 => x"0981069a",
          7599 => x"38811333",
          7600 => x"51ffbf8d",
          7601 => x"3f82d8c8",
          7602 => x"08810652",
          7603 => x"71883871",
          7604 => x"74085455",
          7605 => x"83398053",
          7606 => x"7873710c",
          7607 => x"527482d8",
          7608 => x"c80c873d",
          7609 => x"0d04fa3d",
          7610 => x"0d02ab05",
          7611 => x"337a5889",
          7612 => x"3dfc0552",
          7613 => x"56f4dd3f",
          7614 => x"8b54800b",
          7615 => x"82d8c808",
          7616 => x"24bc3882",
          7617 => x"d8c80884",
          7618 => x"2982f090",
          7619 => x"05700855",
          7620 => x"5573802e",
          7621 => x"84388074",
          7622 => x"34785473",
          7623 => x"802e8438",
          7624 => x"80743478",
          7625 => x"750c7554",
          7626 => x"75802e92",
          7627 => x"38805389",
          7628 => x"3d705384",
          7629 => x"0551f7a7",
          7630 => x"3f82d8c8",
          7631 => x"08547382",
          7632 => x"d8c80c88",
          7633 => x"3d0d04ea",
          7634 => x"3d0d6802",
          7635 => x"840580eb",
          7636 => x"05335959",
          7637 => x"89547880",
          7638 => x"2e84c838",
          7639 => x"77bf0670",
          7640 => x"54993dcc",
          7641 => x"05539a3d",
          7642 => x"84055258",
          7643 => x"f6f13f82",
          7644 => x"d8c80855",
          7645 => x"82d8c808",
          7646 => x"84a4387a",
          7647 => x"5c69528c",
          7648 => x"3d705256",
          7649 => x"eaf33f82",
          7650 => x"d8c80855",
          7651 => x"82d8c808",
          7652 => x"92380280",
          7653 => x"d7053370",
          7654 => x"982b5557",
          7655 => x"73802583",
          7656 => x"38865577",
          7657 => x"9c065473",
          7658 => x"802e81ab",
          7659 => x"3874802e",
          7660 => x"95387484",
          7661 => x"2e098106",
          7662 => x"aa387551",
          7663 => x"dff43f82",
          7664 => x"d8c80855",
          7665 => x"9e3902b2",
          7666 => x"05339106",
          7667 => x"547381b8",
          7668 => x"3877822a",
          7669 => x"70810651",
          7670 => x"5473802e",
          7671 => x"8e388855",
          7672 => x"83bc3977",
          7673 => x"88075874",
          7674 => x"83b43877",
          7675 => x"832a7081",
          7676 => x"06515473",
          7677 => x"802e81af",
          7678 => x"3862527a",
          7679 => x"51d7b03f",
          7680 => x"82d8c808",
          7681 => x"568288b2",
          7682 => x"0a52628e",
          7683 => x"0551c3b7",
          7684 => x"3f6254a0",
          7685 => x"0b8b1534",
          7686 => x"80536252",
          7687 => x"7a51d7c8",
          7688 => x"3f805262",
          7689 => x"9c0551c3",
          7690 => x"9e3f7a54",
          7691 => x"810b8315",
          7692 => x"3475802e",
          7693 => x"80f1387a",
          7694 => x"b4110851",
          7695 => x"54805375",
          7696 => x"52983dd0",
          7697 => x"0551ccc9",
          7698 => x"3f82d8c8",
          7699 => x"085582d8",
          7700 => x"c80882ca",
          7701 => x"38b73974",
          7702 => x"82c43802",
          7703 => x"b2053370",
          7704 => x"842a7081",
          7705 => x"06515556",
          7706 => x"73802e86",
          7707 => x"38845582",
          7708 => x"ad397781",
          7709 => x"2a708106",
          7710 => x"51547380",
          7711 => x"2ea93875",
          7712 => x"81065473",
          7713 => x"802ea038",
          7714 => x"87558292",
          7715 => x"3973527a",
          7716 => x"51c5ae3f",
          7717 => x"82d8c808",
          7718 => x"7bff1890",
          7719 => x"120c5555",
          7720 => x"82d8c808",
          7721 => x"81f83877",
          7722 => x"832a7081",
          7723 => x"06515473",
          7724 => x"802e8638",
          7725 => x"7780c007",
          7726 => x"587ab411",
          7727 => x"08a01b0c",
          7728 => x"63a41b0c",
          7729 => x"63537052",
          7730 => x"57d5e43f",
          7731 => x"82d8c808",
          7732 => x"82d8c808",
          7733 => x"881b0c63",
          7734 => x"9c05525a",
          7735 => x"c1a03f82",
          7736 => x"d8c80882",
          7737 => x"d8c8088c",
          7738 => x"1b0c777a",
          7739 => x"0c568617",
          7740 => x"22841a23",
          7741 => x"77901a34",
          7742 => x"800b911a",
          7743 => x"34800b9c",
          7744 => x"1a0c800b",
          7745 => x"941a0c77",
          7746 => x"852a7081",
          7747 => x"06515473",
          7748 => x"802e818d",
          7749 => x"3882d8c8",
          7750 => x"08802e81",
          7751 => x"843882d8",
          7752 => x"c808941a",
          7753 => x"0c8a1722",
          7754 => x"70892b7b",
          7755 => x"525957a8",
          7756 => x"39765278",
          7757 => x"51c6aa3f",
          7758 => x"82d8c808",
          7759 => x"5782d8c8",
          7760 => x"08812683",
          7761 => x"38825582",
          7762 => x"d8c808ff",
          7763 => x"2e098106",
          7764 => x"83387955",
          7765 => x"75783156",
          7766 => x"74307076",
          7767 => x"07802551",
          7768 => x"54777627",
          7769 => x"8a388170",
          7770 => x"7506555a",
          7771 => x"73c33876",
          7772 => x"981a0c74",
          7773 => x"a9387583",
          7774 => x"ff065473",
          7775 => x"802ea238",
          7776 => x"76527a51",
          7777 => x"c5b13f82",
          7778 => x"d8c80885",
          7779 => x"3882558e",
          7780 => x"3975892a",
          7781 => x"82d8c808",
          7782 => x"059c1a0c",
          7783 => x"84398079",
          7784 => x"0c745473",
          7785 => x"82d8c80c",
          7786 => x"983d0d04",
          7787 => x"f23d0d60",
          7788 => x"63656440",
          7789 => x"405d5980",
          7790 => x"7e0c903d",
          7791 => x"fc055278",
          7792 => x"51f9ce3f",
          7793 => x"82d8c808",
          7794 => x"5582d8c8",
          7795 => x"088a3891",
          7796 => x"19335574",
          7797 => x"802e8638",
          7798 => x"745682c7",
          7799 => x"39901933",
          7800 => x"81065587",
          7801 => x"5674802e",
          7802 => x"82b93895",
          7803 => x"39820b91",
          7804 => x"1a348256",
          7805 => x"82ad3981",
          7806 => x"0b911a34",
          7807 => x"815682a3",
          7808 => x"398c1908",
          7809 => x"941a0831",
          7810 => x"55747c27",
          7811 => x"8338745c",
          7812 => x"7b802e82",
          7813 => x"8c389419",
          7814 => x"087083ff",
          7815 => x"06565674",
          7816 => x"81b4387e",
          7817 => x"8a1122ff",
          7818 => x"0577892a",
          7819 => x"065b5579",
          7820 => x"a8387587",
          7821 => x"38881908",
          7822 => x"558f3998",
          7823 => x"19085278",
          7824 => x"51c49e3f",
          7825 => x"82d8c808",
          7826 => x"55817527",
          7827 => x"ff9f3874",
          7828 => x"ff2effa3",
          7829 => x"3874981a",
          7830 => x"0c981908",
          7831 => x"527e51c3",
          7832 => x"d63f82d8",
          7833 => x"c808802e",
          7834 => x"ff833882",
          7835 => x"d8c8081a",
          7836 => x"7c892a59",
          7837 => x"5777802e",
          7838 => x"80d83877",
          7839 => x"1a7f8a11",
          7840 => x"22585c55",
          7841 => x"75752785",
          7842 => x"38757a31",
          7843 => x"58775476",
          7844 => x"537c5281",
          7845 => x"1b3351ff",
          7846 => x"b8d43f82",
          7847 => x"d8c808fe",
          7848 => x"d6387e83",
          7849 => x"11335656",
          7850 => x"74802ea0",
          7851 => x"38b41608",
          7852 => x"77315574",
          7853 => x"78279538",
          7854 => x"848053b8",
          7855 => x"1652b416",
          7856 => x"08773189",
          7857 => x"2b7d0551",
          7858 => x"ffbeab3f",
          7859 => x"77892b56",
          7860 => x"ba39769c",
          7861 => x"1a0c9419",
          7862 => x"0883ff06",
          7863 => x"84807131",
          7864 => x"57557b76",
          7865 => x"2783387b",
          7866 => x"569c1908",
          7867 => x"527e51c0",
          7868 => x"d03f82d8",
          7869 => x"c808fdff",
          7870 => x"38755394",
          7871 => x"190883ff",
          7872 => x"061fb805",
          7873 => x"527c51ff",
          7874 => x"bdec3f7b",
          7875 => x"76317e08",
          7876 => x"177f0c76",
          7877 => x"1e941b08",
          7878 => x"18941c0c",
          7879 => x"5e5cfdf0",
          7880 => x"39805675",
          7881 => x"82d8c80c",
          7882 => x"903d0d04",
          7883 => x"f23d0d60",
          7884 => x"63656440",
          7885 => x"405d5880",
          7886 => x"7e0c903d",
          7887 => x"fc055277",
          7888 => x"51f6ce3f",
          7889 => x"82d8c808",
          7890 => x"5582d8c8",
          7891 => x"088a3891",
          7892 => x"18335574",
          7893 => x"802e8638",
          7894 => x"745683be",
          7895 => x"39901833",
          7896 => x"70812a70",
          7897 => x"81065156",
          7898 => x"56875674",
          7899 => x"802e83aa",
          7900 => x"38953982",
          7901 => x"0b911934",
          7902 => x"8256839e",
          7903 => x"39810b91",
          7904 => x"19348156",
          7905 => x"83943994",
          7906 => x"18087c11",
          7907 => x"56567476",
          7908 => x"27843875",
          7909 => x"095c7b80",
          7910 => x"2e82f238",
          7911 => x"94180870",
          7912 => x"83ff0656",
          7913 => x"56748281",
          7914 => x"387e8a11",
          7915 => x"22ff0577",
          7916 => x"892a065c",
          7917 => x"557abf38",
          7918 => x"758c3888",
          7919 => x"18085574",
          7920 => x"9c387a52",
          7921 => x"85399818",
          7922 => x"08527751",
          7923 => x"c6ef3f82",
          7924 => x"d8c80855",
          7925 => x"82d8c808",
          7926 => x"802e82b1",
          7927 => x"3874812e",
          7928 => x"ff913874",
          7929 => x"ff2eff95",
          7930 => x"38749819",
          7931 => x"0c881808",
          7932 => x"85387488",
          7933 => x"190c7e55",
          7934 => x"b415089c",
          7935 => x"19082e09",
          7936 => x"81068e38",
          7937 => x"7451ffbd",
          7938 => x"c83f82d8",
          7939 => x"c808feed",
          7940 => x"38981808",
          7941 => x"527e51c0",
          7942 => x"9e3f82d8",
          7943 => x"c808802e",
          7944 => x"fed13882",
          7945 => x"d8c8081b",
          7946 => x"7c892a5a",
          7947 => x"5778802e",
          7948 => x"80d73878",
          7949 => x"1b7f8a11",
          7950 => x"22585b55",
          7951 => x"75752785",
          7952 => x"38757b31",
          7953 => x"59785476",
          7954 => x"537c5281",
          7955 => x"1a3351ff",
          7956 => x"b7863f82",
          7957 => x"d8c808fe",
          7958 => x"a4387eb4",
          7959 => x"11087831",
          7960 => x"56567479",
          7961 => x"279c3884",
          7962 => x"8053b416",
          7963 => x"08773189",
          7964 => x"2b7d0552",
          7965 => x"b81651ff",
          7966 => x"bafc3f7e",
          7967 => x"55800b83",
          7968 => x"16347889",
          7969 => x"2b5680de",
          7970 => x"398c1808",
          7971 => x"94190826",
          7972 => x"94387e51",
          7973 => x"ffbcba3f",
          7974 => x"82d8c808",
          7975 => x"fddf387e",
          7976 => x"77b4120c",
          7977 => x"55769c19",
          7978 => x"0c941808",
          7979 => x"83ff0684",
          7980 => x"80713157",
          7981 => x"557b7627",
          7982 => x"83387b56",
          7983 => x"9c180852",
          7984 => x"7e51ffbc",
          7985 => x"fc3f82d8",
          7986 => x"c808fdb1",
          7987 => x"3875537c",
          7988 => x"52941808",
          7989 => x"83ff061f",
          7990 => x"b80551ff",
          7991 => x"ba983f7e",
          7992 => x"55810b83",
          7993 => x"16347b76",
          7994 => x"317e0817",
          7995 => x"7f0c761e",
          7996 => x"941a0818",
          7997 => x"70941c0c",
          7998 => x"8c1b0858",
          7999 => x"585e5c74",
          8000 => x"76278338",
          8001 => x"7555748c",
          8002 => x"190cfd8a",
          8003 => x"39901833",
          8004 => x"80c00755",
          8005 => x"74901934",
          8006 => x"80567582",
          8007 => x"d8c80c90",
          8008 => x"3d0d04f8",
          8009 => x"3d0d7a8b",
          8010 => x"3dfc0553",
          8011 => x"705256f2",
          8012 => x"e03f82d8",
          8013 => x"c8085782",
          8014 => x"d8c80881",
          8015 => x"80389016",
          8016 => x"3370862a",
          8017 => x"70810651",
          8018 => x"55557380",
          8019 => x"2e80ee38",
          8020 => x"a0160852",
          8021 => x"7851ffbb",
          8022 => x"e83f82d8",
          8023 => x"c8085782",
          8024 => x"d8c80880",
          8025 => x"d838a416",
          8026 => x"088b1133",
          8027 => x"a0075555",
          8028 => x"738b1634",
          8029 => x"88160853",
          8030 => x"74527508",
          8031 => x"51cce93f",
          8032 => x"8c160852",
          8033 => x"9c1551ff",
          8034 => x"b8bd3f82",
          8035 => x"88b20a52",
          8036 => x"961551ff",
          8037 => x"b8b13f76",
          8038 => x"52921551",
          8039 => x"ffb88a3f",
          8040 => x"7854810b",
          8041 => x"83153478",
          8042 => x"51ffbbdc",
          8043 => x"3f82d8c8",
          8044 => x"08901733",
          8045 => x"81bf0655",
          8046 => x"57739017",
          8047 => x"347682d8",
          8048 => x"c80c8a3d",
          8049 => x"0d04fc3d",
          8050 => x"0d767052",
          8051 => x"54fed43f",
          8052 => x"82d8c808",
          8053 => x"5382d8c8",
          8054 => x"089c3886",
          8055 => x"3dfc0552",
          8056 => x"7351f1ad",
          8057 => x"3f82d8c8",
          8058 => x"085382d8",
          8059 => x"c8088738",
          8060 => x"82d8c808",
          8061 => x"740c7282",
          8062 => x"d8c80c86",
          8063 => x"3d0d04ff",
          8064 => x"3d0d843d",
          8065 => x"51e6cd3f",
          8066 => x"8b52800b",
          8067 => x"82d8c808",
          8068 => x"248b3882",
          8069 => x"d8c80882",
          8070 => x"f0a43480",
          8071 => x"527182d8",
          8072 => x"c80c833d",
          8073 => x"0d04ee3d",
          8074 => x"0d805394",
          8075 => x"3dcc0552",
          8076 => x"953d51e9",
          8077 => x"aa3f82d8",
          8078 => x"c8085582",
          8079 => x"d8c80880",
          8080 => x"e0387658",
          8081 => x"6452943d",
          8082 => x"d00551dd",
          8083 => x"ac3f82d8",
          8084 => x"c8085582",
          8085 => x"d8c808bc",
          8086 => x"380280c7",
          8087 => x"05337098",
          8088 => x"2b555673",
          8089 => x"80258938",
          8090 => x"767a9812",
          8091 => x"0c54b239",
          8092 => x"02a20533",
          8093 => x"70842a70",
          8094 => x"81065155",
          8095 => x"5673802e",
          8096 => x"9e38767f",
          8097 => x"53705254",
          8098 => x"caa53f82",
          8099 => x"d8c80898",
          8100 => x"150c8e39",
          8101 => x"82d8c808",
          8102 => x"842e0981",
          8103 => x"06833885",
          8104 => x"557482d8",
          8105 => x"c80c943d",
          8106 => x"0d04ffa3",
          8107 => x"3d0d80e1",
          8108 => x"3d0880e1",
          8109 => x"3d085b5b",
          8110 => x"807a3480",
          8111 => x"5380df3d",
          8112 => x"fdb40552",
          8113 => x"80e03d51",
          8114 => x"e8953f82",
          8115 => x"d8c80857",
          8116 => x"82d8c808",
          8117 => x"83a1387b",
          8118 => x"80d43d0c",
          8119 => x"7a7c9811",
          8120 => x"0880d83d",
          8121 => x"0c555880",
          8122 => x"d53d0854",
          8123 => x"73802e82",
          8124 => x"8338a052",
          8125 => x"80d33d70",
          8126 => x"5255c4d4",
          8127 => x"3f82d8c8",
          8128 => x"085782d8",
          8129 => x"c80882ef",
          8130 => x"3880d93d",
          8131 => x"08527b51",
          8132 => x"ffb8ae3f",
          8133 => x"82d8c808",
          8134 => x"5782d8c8",
          8135 => x"0882d838",
          8136 => x"80da3d08",
          8137 => x"527b51c9",
          8138 => x"863f82d8",
          8139 => x"c80880d6",
          8140 => x"3d0c7652",
          8141 => x"7451c498",
          8142 => x"3f82d8c8",
          8143 => x"085782d8",
          8144 => x"c80882b3",
          8145 => x"38805274",
          8146 => x"51c9fa3f",
          8147 => x"82d8c808",
          8148 => x"5782d8c8",
          8149 => x"08a73880",
          8150 => x"da3d0852",
          8151 => x"7b51c8cf",
          8152 => x"3f7382d8",
          8153 => x"c8082ea6",
          8154 => x"38765274",
          8155 => x"51c5ac3f",
          8156 => x"82d8c808",
          8157 => x"5782d8c8",
          8158 => x"08802ec9",
          8159 => x"3876842e",
          8160 => x"09810686",
          8161 => x"38825781",
          8162 => x"ee397681",
          8163 => x"ea3880df",
          8164 => x"3dfdb805",
          8165 => x"527451d6",
          8166 => x"e43f7693",
          8167 => x"3d781182",
          8168 => x"11335156",
          8169 => x"5a567380",
          8170 => x"2e923802",
          8171 => x"80c60555",
          8172 => x"81168116",
          8173 => x"70335656",
          8174 => x"5673f538",
          8175 => x"81165473",
          8176 => x"78268199",
          8177 => x"3875802e",
          8178 => x"9c387816",
          8179 => x"820555ff",
          8180 => x"1880e13d",
          8181 => x"0811ff18",
          8182 => x"ff185858",
          8183 => x"55587433",
          8184 => x"743475eb",
          8185 => x"38ff1880",
          8186 => x"e13d0811",
          8187 => x"5558af74",
          8188 => x"34fdf439",
          8189 => x"777b2e09",
          8190 => x"81068d38",
          8191 => x"ff1880e1",
          8192 => x"3d081155",
          8193 => x"58af7434",
          8194 => x"800b82f0",
          8195 => x"a4337084",
          8196 => x"2982cac0",
          8197 => x"05700870",
          8198 => x"33525c56",
          8199 => x"56567376",
          8200 => x"2e8d3881",
          8201 => x"16701a70",
          8202 => x"33515556",
          8203 => x"73f53882",
          8204 => x"16547378",
          8205 => x"26a73880",
          8206 => x"55747627",
          8207 => x"91387419",
          8208 => x"5473337a",
          8209 => x"7081055c",
          8210 => x"34811555",
          8211 => x"ec39ba7a",
          8212 => x"7081055c",
          8213 => x"3474ff2e",
          8214 => x"09810685",
          8215 => x"38915797",
          8216 => x"3980e03d",
          8217 => x"08188119",
          8218 => x"59547333",
          8219 => x"7a708105",
          8220 => x"5c347a78",
          8221 => x"26eb3880",
          8222 => x"7a347682",
          8223 => x"d8c80c80",
          8224 => x"df3d0d04",
          8225 => x"f73d0d7b",
          8226 => x"7d8d3dfc",
          8227 => x"05547153",
          8228 => x"5755ebfd",
          8229 => x"3f82d8c8",
          8230 => x"085382d8",
          8231 => x"c80882fe",
          8232 => x"38911533",
          8233 => x"537282f6",
          8234 => x"388c1508",
          8235 => x"54737627",
          8236 => x"92389015",
          8237 => x"3370812a",
          8238 => x"70810651",
          8239 => x"54577283",
          8240 => x"38735694",
          8241 => x"15085480",
          8242 => x"7094170c",
          8243 => x"5875782e",
          8244 => x"829b3879",
          8245 => x"8a112270",
          8246 => x"892b5951",
          8247 => x"5373782e",
          8248 => x"b7387652",
          8249 => x"ff1651fe",
          8250 => x"c5993f82",
          8251 => x"d8c808ff",
          8252 => x"15785470",
          8253 => x"535553fe",
          8254 => x"c5893f82",
          8255 => x"d8c80873",
          8256 => x"26963876",
          8257 => x"30707506",
          8258 => x"7094180c",
          8259 => x"77713198",
          8260 => x"18085758",
          8261 => x"5153b239",
          8262 => x"88150854",
          8263 => x"73a73873",
          8264 => x"527451ff",
          8265 => x"bc973f82",
          8266 => x"d8c80854",
          8267 => x"82d8c808",
          8268 => x"812e819d",
          8269 => x"3882d8c8",
          8270 => x"08ff2e81",
          8271 => x"9e3882d8",
          8272 => x"c8088816",
          8273 => x"0c739816",
          8274 => x"0c73802e",
          8275 => x"819f3876",
          8276 => x"762780de",
          8277 => x"38757731",
          8278 => x"94160818",
          8279 => x"94170c90",
          8280 => x"16337081",
          8281 => x"2a708106",
          8282 => x"51555a56",
          8283 => x"72802e9b",
          8284 => x"38735274",
          8285 => x"51ffbbc5",
          8286 => x"3f82d8c8",
          8287 => x"085482d8",
          8288 => x"c8089538",
          8289 => x"82d8c808",
          8290 => x"56a83973",
          8291 => x"527451ff",
          8292 => x"b5cf3f82",
          8293 => x"d8c80854",
          8294 => x"73ff2ebf",
          8295 => x"38817427",
          8296 => x"b0387953",
          8297 => x"739c1408",
          8298 => x"27a73873",
          8299 => x"98160cff",
          8300 => x"9e399415",
          8301 => x"08169416",
          8302 => x"0c7583ff",
          8303 => x"06537280",
          8304 => x"2eab3873",
          8305 => x"527951ff",
          8306 => x"b4ed3f82",
          8307 => x"d8c80894",
          8308 => x"38820b91",
          8309 => x"16348253",
          8310 => x"80c43981",
          8311 => x"0b911634",
          8312 => x"8153bb39",
          8313 => x"75892a82",
          8314 => x"d8c80805",
          8315 => x"58941508",
          8316 => x"548c1508",
          8317 => x"74279038",
          8318 => x"738c160c",
          8319 => x"90153380",
          8320 => x"c0075372",
          8321 => x"90163473",
          8322 => x"83ff0653",
          8323 => x"72802e8c",
          8324 => x"38779c16",
          8325 => x"082e8538",
          8326 => x"779c160c",
          8327 => x"80537282",
          8328 => x"d8c80c8b",
          8329 => x"3d0d04f9",
          8330 => x"3d0d7956",
          8331 => x"89547580",
          8332 => x"2e818b38",
          8333 => x"8053893d",
          8334 => x"fc05528a",
          8335 => x"3d840551",
          8336 => x"e19d3f82",
          8337 => x"d8c80855",
          8338 => x"82d8c808",
          8339 => x"80eb3877",
          8340 => x"760c7a52",
          8341 => x"7551d5a1",
          8342 => x"3f82d8c8",
          8343 => x"085582d8",
          8344 => x"c80880c4",
          8345 => x"38ab1633",
          8346 => x"70982b55",
          8347 => x"57807424",
          8348 => x"a2388616",
          8349 => x"3370842a",
          8350 => x"70810651",
          8351 => x"55577380",
          8352 => x"2eae389c",
          8353 => x"16085277",
          8354 => x"51c2a43f",
          8355 => x"82d8c808",
          8356 => x"88170c77",
          8357 => x"54861422",
          8358 => x"84172374",
          8359 => x"527551ff",
          8360 => x"bdae3f82",
          8361 => x"d8c80855",
          8362 => x"74842e09",
          8363 => x"81068538",
          8364 => x"85558639",
          8365 => x"74802e84",
          8366 => x"3880760c",
          8367 => x"74547382",
          8368 => x"d8c80c89",
          8369 => x"3d0d04fc",
          8370 => x"3d0d7687",
          8371 => x"3dfc0553",
          8372 => x"705253e7",
          8373 => x"bc3f82d8",
          8374 => x"c8088738",
          8375 => x"82d8c808",
          8376 => x"730c863d",
          8377 => x"0d04fb3d",
          8378 => x"0d777989",
          8379 => x"3dfc0554",
          8380 => x"71535654",
          8381 => x"e79b3f82",
          8382 => x"d8c80853",
          8383 => x"82d8c808",
          8384 => x"80e13874",
          8385 => x"943882d8",
          8386 => x"c8085273",
          8387 => x"51ffbcc0",
          8388 => x"3f82d8c8",
          8389 => x"085380cb",
          8390 => x"3982d8c8",
          8391 => x"08527351",
          8392 => x"c2a33f82",
          8393 => x"d8c80853",
          8394 => x"82d8c808",
          8395 => x"842e0981",
          8396 => x"06853880",
          8397 => x"53873982",
          8398 => x"d8c808a7",
          8399 => x"38745273",
          8400 => x"51cfba3f",
          8401 => x"72527351",
          8402 => x"ffbdd03f",
          8403 => x"82d8c808",
          8404 => x"84327030",
          8405 => x"7072079f",
          8406 => x"2c7082d8",
          8407 => x"c8080651",
          8408 => x"51545472",
          8409 => x"82d8c80c",
          8410 => x"873d0d04",
          8411 => x"ed3d0d66",
          8412 => x"57805389",
          8413 => x"3d705397",
          8414 => x"3d5256de",
          8415 => x"e23f82d8",
          8416 => x"c8085582",
          8417 => x"d8c808b2",
          8418 => x"38655275",
          8419 => x"51d2ea3f",
          8420 => x"82d8c808",
          8421 => x"5582d8c8",
          8422 => x"08a03802",
          8423 => x"80cb0533",
          8424 => x"70982b55",
          8425 => x"58738025",
          8426 => x"85388655",
          8427 => x"8d397680",
          8428 => x"2e883876",
          8429 => x"527551ce",
          8430 => x"c43f7482",
          8431 => x"d8c80c95",
          8432 => x"3d0d04f0",
          8433 => x"3d0d6365",
          8434 => x"555c8053",
          8435 => x"923dec05",
          8436 => x"52933d51",
          8437 => x"de893f82",
          8438 => x"d8c8085b",
          8439 => x"82d8c808",
          8440 => x"8282387c",
          8441 => x"740c7308",
          8442 => x"9c1108fe",
          8443 => x"11941308",
          8444 => x"59565855",
          8445 => x"75742691",
          8446 => x"38757c0c",
          8447 => x"81e63981",
          8448 => x"5b81ce39",
          8449 => x"825b81c9",
          8450 => x"3982d8c8",
          8451 => x"08753355",
          8452 => x"5973812e",
          8453 => x"09810680",
          8454 => x"c0388275",
          8455 => x"5f577652",
          8456 => x"923df005",
          8457 => x"51ffb0b9",
          8458 => x"3f82d8c8",
          8459 => x"08ff2ecf",
          8460 => x"3882d8c8",
          8461 => x"08812ecc",
          8462 => x"3882d8c8",
          8463 => x"08307082",
          8464 => x"d8c80807",
          8465 => x"80257a05",
          8466 => x"81197f53",
          8467 => x"595a549c",
          8468 => x"14087726",
          8469 => x"c93880f9",
          8470 => x"39a81508",
          8471 => x"82d8c808",
          8472 => x"57587598",
          8473 => x"38775281",
          8474 => x"187d5258",
          8475 => x"ffadd23f",
          8476 => x"82d8c808",
          8477 => x"5b82d8c8",
          8478 => x"0880d638",
          8479 => x"7c703377",
          8480 => x"12ff1a5d",
          8481 => x"52565474",
          8482 => x"822e0981",
          8483 => x"069e38b8",
          8484 => x"1451ffa9",
          8485 => x"d23f82d8",
          8486 => x"c80883ff",
          8487 => x"ff067030",
          8488 => x"7080251b",
          8489 => x"8219595b",
          8490 => x"51549b39",
          8491 => x"b81451ff",
          8492 => x"a9cc3f82",
          8493 => x"d8c808f0",
          8494 => x"0a067030",
          8495 => x"7080251b",
          8496 => x"8419595b",
          8497 => x"51547583",
          8498 => x"ff067a58",
          8499 => x"5679ff92",
          8500 => x"38787c0c",
          8501 => x"7c799412",
          8502 => x"0c841133",
          8503 => x"81075654",
          8504 => x"74841534",
          8505 => x"7a82d8c8",
          8506 => x"0c923d0d",
          8507 => x"04f93d0d",
          8508 => x"798a3dfc",
          8509 => x"05537052",
          8510 => x"57e3963f",
          8511 => x"82d8c808",
          8512 => x"5682d8c8",
          8513 => x"0881aa38",
          8514 => x"91173356",
          8515 => x"7581a238",
          8516 => x"90173370",
          8517 => x"812a7081",
          8518 => x"06515555",
          8519 => x"87557380",
          8520 => x"2e819038",
          8521 => x"94170854",
          8522 => x"738c1808",
          8523 => x"27818238",
          8524 => x"739c3882",
          8525 => x"d8c80853",
          8526 => x"88170852",
          8527 => x"7651ffb2",
          8528 => x"d03f82d8",
          8529 => x"c8087488",
          8530 => x"190c5680",
          8531 => x"ca399817",
          8532 => x"08527651",
          8533 => x"ffae8a3f",
          8534 => x"82d8c808",
          8535 => x"ff2e0981",
          8536 => x"06833881",
          8537 => x"5682d8c8",
          8538 => x"08812e09",
          8539 => x"81068538",
          8540 => x"8256a439",
          8541 => x"75a13877",
          8542 => x"5482d8c8",
          8543 => x"089c1508",
          8544 => x"27953898",
          8545 => x"17085382",
          8546 => x"d8c80852",
          8547 => x"7651ffb2",
          8548 => x"803f82d8",
          8549 => x"c8085694",
          8550 => x"17088c18",
          8551 => x"0c901733",
          8552 => x"80c00754",
          8553 => x"73901834",
          8554 => x"75802e85",
          8555 => x"38759118",
          8556 => x"34755574",
          8557 => x"82d8c80c",
          8558 => x"893d0d04",
          8559 => x"e03d0d82",
          8560 => x"53a23dff",
          8561 => x"9c0552a3",
          8562 => x"3d51da93",
          8563 => x"3f82d8c8",
          8564 => x"085582d8",
          8565 => x"c80881f9",
          8566 => x"387846a3",
          8567 => x"3d085296",
          8568 => x"3d705258",
          8569 => x"ce933f82",
          8570 => x"d8c80855",
          8571 => x"82d8c808",
          8572 => x"81df3802",
          8573 => x"80ff0533",
          8574 => x"70852a70",
          8575 => x"81065155",
          8576 => x"56865573",
          8577 => x"81cb3875",
          8578 => x"982b5480",
          8579 => x"742481c1",
          8580 => x"380280da",
          8581 => x"05337081",
          8582 => x"06585487",
          8583 => x"557681b1",
          8584 => x"386c5278",
          8585 => x"51ffbb87",
          8586 => x"3f82d8c8",
          8587 => x"0874842a",
          8588 => x"70810651",
          8589 => x"55567380",
          8590 => x"2e80d638",
          8591 => x"785482d8",
          8592 => x"c8089815",
          8593 => x"082e8189",
          8594 => x"38735a82",
          8595 => x"d8c8085c",
          8596 => x"76528a3d",
          8597 => x"705254ff",
          8598 => x"b5f63f82",
          8599 => x"d8c80855",
          8600 => x"82d8c808",
          8601 => x"80eb3882",
          8602 => x"d8c80852",
          8603 => x"7351ffbb",
          8604 => x"d43f82d8",
          8605 => x"c8085582",
          8606 => x"d8c80886",
          8607 => x"38875580",
          8608 => x"d03982d8",
          8609 => x"c808842e",
          8610 => x"883882d8",
          8611 => x"c80880c1",
          8612 => x"387751c7",
          8613 => x"ef3f82d8",
          8614 => x"c80882d8",
          8615 => x"c8083070",
          8616 => x"82d8c808",
          8617 => x"07802551",
          8618 => x"55557580",
          8619 => x"2e953873",
          8620 => x"802e9038",
          8621 => x"80537552",
          8622 => x"7751ffaf",
          8623 => x"d43f82d8",
          8624 => x"c8085574",
          8625 => x"8c387851",
          8626 => x"ffa9bd3f",
          8627 => x"82d8c808",
          8628 => x"557482d8",
          8629 => x"c80ca23d",
          8630 => x"0d04e83d",
          8631 => x"0d82539a",
          8632 => x"3dffbc05",
          8633 => x"529b3d51",
          8634 => x"d7f53f82",
          8635 => x"d8c80854",
          8636 => x"82d8c808",
          8637 => x"82b73878",
          8638 => x"5e6a528e",
          8639 => x"3d705258",
          8640 => x"cbf73f82",
          8641 => x"d8c80854",
          8642 => x"82d8c808",
          8643 => x"86388854",
          8644 => x"829b3982",
          8645 => x"d8c80884",
          8646 => x"2e098106",
          8647 => x"828f3802",
          8648 => x"80df0533",
          8649 => x"70852a81",
          8650 => x"06515586",
          8651 => x"547481fd",
          8652 => x"38785a74",
          8653 => x"528a3d70",
          8654 => x"5257ffb0",
          8655 => x"803f82d8",
          8656 => x"c8087555",
          8657 => x"5682d8c8",
          8658 => x"08833887",
          8659 => x"5482d8c8",
          8660 => x"08812e09",
          8661 => x"81068338",
          8662 => x"825482d8",
          8663 => x"c808ff2e",
          8664 => x"09810686",
          8665 => x"38815481",
          8666 => x"ba397381",
          8667 => x"b63882d8",
          8668 => x"c8085278",
          8669 => x"51ffb2e0",
          8670 => x"3f82d8c8",
          8671 => x"085482d8",
          8672 => x"c808819f",
          8673 => x"388b53a0",
          8674 => x"52b81951",
          8675 => x"ffa58a3f",
          8676 => x"7854ae0b",
          8677 => x"b8153478",
          8678 => x"54900b80",
          8679 => x"c3153482",
          8680 => x"88b20a52",
          8681 => x"80ce1951",
          8682 => x"ffa49c3f",
          8683 => x"755378b8",
          8684 => x"115351ff",
          8685 => x"b8b23fa0",
          8686 => x"5378b811",
          8687 => x"5380d805",
          8688 => x"51ffa4b2",
          8689 => x"3f7854ae",
          8690 => x"0b80d915",
          8691 => x"347f5378",
          8692 => x"80d81153",
          8693 => x"51ffb890",
          8694 => x"3f785481",
          8695 => x"0b831534",
          8696 => x"7751ffbf",
          8697 => x"cd3f82d8",
          8698 => x"c8085482",
          8699 => x"d8c808b3",
          8700 => x"388288b2",
          8701 => x"0a526496",
          8702 => x"0551ffa3",
          8703 => x"ca3f7553",
          8704 => x"64527851",
          8705 => x"ffb7e13f",
          8706 => x"6454900b",
          8707 => x"8b153478",
          8708 => x"54810b83",
          8709 => x"15347851",
          8710 => x"ffa6ed3f",
          8711 => x"82d8c808",
          8712 => x"548b3980",
          8713 => x"53755276",
          8714 => x"51fface5",
          8715 => x"3f7382d8",
          8716 => x"c80c9a3d",
          8717 => x"0d04d83d",
          8718 => x"0dab3d84",
          8719 => x"0551d294",
          8720 => x"3f8253aa",
          8721 => x"3dfefc05",
          8722 => x"52ab3d51",
          8723 => x"d5913f82",
          8724 => x"d8c80855",
          8725 => x"82d8c808",
          8726 => x"82d83878",
          8727 => x"4eab3d08",
          8728 => x"529e3d70",
          8729 => x"5258c991",
          8730 => x"3f82d8c8",
          8731 => x"085582d8",
          8732 => x"c80882be",
          8733 => x"3802819f",
          8734 => x"053381a0",
          8735 => x"06548655",
          8736 => x"7382af38",
          8737 => x"a053a53d",
          8738 => x"0852aa3d",
          8739 => x"ff800551",
          8740 => x"ffa2e33f",
          8741 => x"b0537752",
          8742 => x"923d7052",
          8743 => x"54ffa2d6",
          8744 => x"3fac3d08",
          8745 => x"527351c8",
          8746 => x"d03f82d8",
          8747 => x"c8085582",
          8748 => x"d8c80897",
          8749 => x"3863a13d",
          8750 => x"082e0981",
          8751 => x"06883865",
          8752 => x"a33d082e",
          8753 => x"92388855",
          8754 => x"81e83982",
          8755 => x"d8c80884",
          8756 => x"2e098106",
          8757 => x"81bb3873",
          8758 => x"51ffbdd6",
          8759 => x"3f82d8c8",
          8760 => x"085582d8",
          8761 => x"c80881ca",
          8762 => x"38685693",
          8763 => x"53aa3dff",
          8764 => x"8d05528d",
          8765 => x"1651ffa1",
          8766 => x"fd3f02af",
          8767 => x"05338b17",
          8768 => x"348b1633",
          8769 => x"70842a70",
          8770 => x"81065155",
          8771 => x"55738938",
          8772 => x"74a00754",
          8773 => x"738b1734",
          8774 => x"7854810b",
          8775 => x"8315348b",
          8776 => x"16337084",
          8777 => x"2a708106",
          8778 => x"51555573",
          8779 => x"802e80e7",
          8780 => x"386f642e",
          8781 => x"80e13875",
          8782 => x"527851ff",
          8783 => x"b4f13f82",
          8784 => x"d8c80852",
          8785 => x"7851ffa5",
          8786 => x"ee3f8255",
          8787 => x"82d8c808",
          8788 => x"802e80de",
          8789 => x"3882d8c8",
          8790 => x"08527851",
          8791 => x"ffa3e23f",
          8792 => x"82d8c808",
          8793 => x"7980d811",
          8794 => x"58585582",
          8795 => x"d8c80880",
          8796 => x"c1388116",
          8797 => x"335473ae",
          8798 => x"2e098106",
          8799 => x"9a386353",
          8800 => x"75527651",
          8801 => x"ffb4e13f",
          8802 => x"7854810b",
          8803 => x"83153487",
          8804 => x"3982d8c8",
          8805 => x"089c3877",
          8806 => x"51c1e93f",
          8807 => x"82d8c808",
          8808 => x"5582d8c8",
          8809 => x"088c3878",
          8810 => x"51ffa3dc",
          8811 => x"3f82d8c8",
          8812 => x"08557482",
          8813 => x"d8c80caa",
          8814 => x"3d0d04ec",
          8815 => x"3d0d0280",
          8816 => x"df053302",
          8817 => x"840580e3",
          8818 => x"05335757",
          8819 => x"8253963d",
          8820 => x"cc055297",
          8821 => x"3d51d287",
          8822 => x"3f82d8c8",
          8823 => x"085582d8",
          8824 => x"c80880cf",
          8825 => x"38785a66",
          8826 => x"52963dd0",
          8827 => x"0551c689",
          8828 => x"3f82d8c8",
          8829 => x"085582d8",
          8830 => x"c808b838",
          8831 => x"0280cf05",
          8832 => x"3381a006",
          8833 => x"54865573",
          8834 => x"aa3875a7",
          8835 => x"06617109",
          8836 => x"8b123371",
          8837 => x"067a7406",
          8838 => x"07515755",
          8839 => x"56748b15",
          8840 => x"34785481",
          8841 => x"0b831534",
          8842 => x"7851ffa2",
          8843 => x"db3f82d8",
          8844 => x"c8085574",
          8845 => x"82d8c80c",
          8846 => x"963d0d04",
          8847 => x"ee3d0d65",
          8848 => x"56825394",
          8849 => x"3dcc0552",
          8850 => x"953d51d1",
          8851 => x"923f82d8",
          8852 => x"c8085582",
          8853 => x"d8c80880",
          8854 => x"cb387658",
          8855 => x"6452943d",
          8856 => x"d00551c5",
          8857 => x"943f82d8",
          8858 => x"c8085582",
          8859 => x"d8c808b4",
          8860 => x"380280c7",
          8861 => x"053381a0",
          8862 => x"06548655",
          8863 => x"73a63884",
          8864 => x"16228617",
          8865 => x"2271902b",
          8866 => x"07535496",
          8867 => x"1f51ff9e",
          8868 => x"b63f7654",
          8869 => x"810b8315",
          8870 => x"347651ff",
          8871 => x"a1ea3f82",
          8872 => x"d8c80855",
          8873 => x"7482d8c8",
          8874 => x"0c943d0d",
          8875 => x"04e93d0d",
          8876 => x"6a6c5c5a",
          8877 => x"8053993d",
          8878 => x"cc05529a",
          8879 => x"3d51d09f",
          8880 => x"3f82d8c8",
          8881 => x"0882d8c8",
          8882 => x"08307082",
          8883 => x"d8c80807",
          8884 => x"80255155",
          8885 => x"5779802e",
          8886 => x"81863881",
          8887 => x"70750655",
          8888 => x"5573802e",
          8889 => x"80fa387b",
          8890 => x"5d805f80",
          8891 => x"528d3d70",
          8892 => x"5254ffac",
          8893 => x"db3f82d8",
          8894 => x"c8085782",
          8895 => x"d8c80880",
          8896 => x"d2387452",
          8897 => x"7351ffb2",
          8898 => x"bc3f82d8",
          8899 => x"c8085782",
          8900 => x"d8c808bf",
          8901 => x"3882d8c8",
          8902 => x"0882d8c8",
          8903 => x"08655b59",
          8904 => x"56781881",
          8905 => x"197b1856",
          8906 => x"59557433",
          8907 => x"74348116",
          8908 => x"568a7827",
          8909 => x"ec388b56",
          8910 => x"751a5480",
          8911 => x"74347580",
          8912 => x"2e9e38ff",
          8913 => x"16701b70",
          8914 => x"33515556",
          8915 => x"73a02ee8",
          8916 => x"388e3976",
          8917 => x"842e0981",
          8918 => x"06863880",
          8919 => x"7a348057",
          8920 => x"76307078",
          8921 => x"07802551",
          8922 => x"547a802e",
          8923 => x"80c13873",
          8924 => x"802ebc38",
          8925 => x"7ba41108",
          8926 => x"5351ff9f",
          8927 => x"c43f82d8",
          8928 => x"c8085782",
          8929 => x"d8c808a7",
          8930 => x"387b7033",
          8931 => x"555580c3",
          8932 => x"5673832e",
          8933 => x"8b3880e4",
          8934 => x"5673842e",
          8935 => x"8338a756",
          8936 => x"7515b805",
          8937 => x"51ff9bd6",
          8938 => x"3f82d8c8",
          8939 => x"087b0c76",
          8940 => x"82d8c80c",
          8941 => x"993d0d04",
          8942 => x"e63d0d82",
          8943 => x"539c3dff",
          8944 => x"b405529d",
          8945 => x"3d51ce97",
          8946 => x"3f82d8c8",
          8947 => x"0882d8c8",
          8948 => x"08565482",
          8949 => x"d8c80882",
          8950 => x"dd388b53",
          8951 => x"a0528a3d",
          8952 => x"705258ff",
          8953 => x"9cb33f73",
          8954 => x"6d703351",
          8955 => x"55569f74",
          8956 => x"27818638",
          8957 => x"77579d3d",
          8958 => x"51ff9d90",
          8959 => x"3f82d8c8",
          8960 => x"0883ffff",
          8961 => x"2680c438",
          8962 => x"82d8c808",
          8963 => x"5195983f",
          8964 => x"83b55282",
          8965 => x"d8c80851",
          8966 => x"93e83f82",
          8967 => x"d8c80883",
          8968 => x"ffff0655",
          8969 => x"74802ea3",
          8970 => x"38745282",
          8971 => x"cbe051ff",
          8972 => x"9cb23f82",
          8973 => x"d8c80893",
          8974 => x"3881ff75",
          8975 => x"27883875",
          8976 => x"89268838",
          8977 => x"8b398a76",
          8978 => x"27863886",
          8979 => x"5581e739",
          8980 => x"81ff7527",
          8981 => x"8f387488",
          8982 => x"2a547377",
          8983 => x"70810559",
          8984 => x"34811656",
          8985 => x"74777081",
          8986 => x"05593481",
          8987 => x"166d7033",
          8988 => x"51555673",
          8989 => x"9f26fefe",
          8990 => x"388a3d33",
          8991 => x"54865573",
          8992 => x"81e52e81",
          8993 => x"b1387580",
          8994 => x"2e993802",
          8995 => x"a3055575",
          8996 => x"15703351",
          8997 => x"5473a02e",
          8998 => x"09810687",
          8999 => x"38ff1656",
          9000 => x"75ed3878",
          9001 => x"40804280",
          9002 => x"52903d70",
          9003 => x"5255ffa9",
          9004 => x"9f3f82d8",
          9005 => x"c8085482",
          9006 => x"d8c80880",
          9007 => x"f7388152",
          9008 => x"7451ffaf",
          9009 => x"803f82d8",
          9010 => x"c8085482",
          9011 => x"d8c8088d",
          9012 => x"387580c4",
          9013 => x"386654e5",
          9014 => x"743480c6",
          9015 => x"3982d8c8",
          9016 => x"08842e09",
          9017 => x"810680cc",
          9018 => x"38805475",
          9019 => x"742e80c4",
          9020 => x"38815274",
          9021 => x"51ffac9c",
          9022 => x"3f82d8c8",
          9023 => x"085482d8",
          9024 => x"c808b138",
          9025 => x"a05382d8",
          9026 => x"c8085266",
          9027 => x"51ff9a89",
          9028 => x"3f665488",
          9029 => x"0b8b1534",
          9030 => x"8b537752",
          9031 => x"6651ff99",
          9032 => x"d53f7854",
          9033 => x"810b8315",
          9034 => x"347851ff",
          9035 => x"9cda3f82",
          9036 => x"d8c80854",
          9037 => x"73557482",
          9038 => x"d8c80c9c",
          9039 => x"3d0d04f2",
          9040 => x"3d0d6062",
          9041 => x"02880580",
          9042 => x"cb053393",
          9043 => x"3dfc0555",
          9044 => x"7254405e",
          9045 => x"5ad2ba3f",
          9046 => x"82d8c808",
          9047 => x"5882d8c8",
          9048 => x"0882bd38",
          9049 => x"911a3358",
          9050 => x"7782b538",
          9051 => x"7c802e97",
          9052 => x"388c1a08",
          9053 => x"59789038",
          9054 => x"901a3370",
          9055 => x"812a7081",
          9056 => x"06515555",
          9057 => x"73903887",
          9058 => x"54829739",
          9059 => x"82588290",
          9060 => x"39815882",
          9061 => x"8b397e8a",
          9062 => x"11227089",
          9063 => x"2b70557f",
          9064 => x"54565656",
          9065 => x"feabdc3f",
          9066 => x"ff147d06",
          9067 => x"70307072",
          9068 => x"079f2a82",
          9069 => x"d8c80805",
          9070 => x"9019087c",
          9071 => x"405a5d55",
          9072 => x"55817727",
          9073 => x"88389c16",
          9074 => x"08772683",
          9075 => x"38825776",
          9076 => x"77565980",
          9077 => x"56745279",
          9078 => x"51ff9d85",
          9079 => x"3f81157f",
          9080 => x"55559c14",
          9081 => x"08752683",
          9082 => x"38825582",
          9083 => x"d8c80881",
          9084 => x"2eff9938",
          9085 => x"82d8c808",
          9086 => x"ff2eff95",
          9087 => x"3882d8c8",
          9088 => x"088e3881",
          9089 => x"1656757b",
          9090 => x"2e098106",
          9091 => x"87389339",
          9092 => x"74598056",
          9093 => x"74772e09",
          9094 => x"8106ffb9",
          9095 => x"38875880",
          9096 => x"ff397d80",
          9097 => x"2eba3878",
          9098 => x"7b55557a",
          9099 => x"802eb438",
          9100 => x"81155673",
          9101 => x"812e0981",
          9102 => x"068338ff",
          9103 => x"56755374",
          9104 => x"527e51ff",
          9105 => x"9e943f82",
          9106 => x"d8c80858",
          9107 => x"82d8c808",
          9108 => x"80ce3874",
          9109 => x"8116ff16",
          9110 => x"56565c73",
          9111 => x"d3388439",
          9112 => x"ff195c7e",
          9113 => x"7c90120c",
          9114 => x"557d802e",
          9115 => x"b3387888",
          9116 => x"1b0c7c8c",
          9117 => x"1b0c901a",
          9118 => x"3380c007",
          9119 => x"5473901b",
          9120 => x"349c1508",
          9121 => x"fe059416",
          9122 => x"08575475",
          9123 => x"74269138",
          9124 => x"757b3194",
          9125 => x"160c8415",
          9126 => x"33810754",
          9127 => x"73841634",
          9128 => x"77547382",
          9129 => x"d8c80c90",
          9130 => x"3d0d04e9",
          9131 => x"3d0d6b6d",
          9132 => x"02880580",
          9133 => x"eb05339d",
          9134 => x"3d545a5c",
          9135 => x"59c5953f",
          9136 => x"8b56800b",
          9137 => x"82d8c808",
          9138 => x"248bf838",
          9139 => x"82d8c808",
          9140 => x"842982f0",
          9141 => x"90057008",
          9142 => x"51557480",
          9143 => x"2e843880",
          9144 => x"753482d8",
          9145 => x"c80881ff",
          9146 => x"065f8152",
          9147 => x"7e51ff8e",
          9148 => x"fe3f82d8",
          9149 => x"c80881ff",
          9150 => x"06708106",
          9151 => x"56578356",
          9152 => x"748bc038",
          9153 => x"76822a70",
          9154 => x"81065155",
          9155 => x"8a56748b",
          9156 => x"b238993d",
          9157 => x"fc055383",
          9158 => x"527e51ff",
          9159 => x"939e3f82",
          9160 => x"d8c80899",
          9161 => x"38675574",
          9162 => x"802e9238",
          9163 => x"74828080",
          9164 => x"268b38ff",
          9165 => x"15750655",
          9166 => x"74802e83",
          9167 => x"38814878",
          9168 => x"802e8738",
          9169 => x"84807926",
          9170 => x"92387881",
          9171 => x"800a268b",
          9172 => x"38ff1979",
          9173 => x"06557480",
          9174 => x"2e863893",
          9175 => x"568ae439",
          9176 => x"78892a6e",
          9177 => x"892a7089",
          9178 => x"2b775948",
          9179 => x"43597a83",
          9180 => x"38815661",
          9181 => x"30708025",
          9182 => x"77075155",
          9183 => x"9156748a",
          9184 => x"c238993d",
          9185 => x"f8055381",
          9186 => x"527e51ff",
          9187 => x"92ae3f81",
          9188 => x"5682d8c8",
          9189 => x"088aac38",
          9190 => x"77832a70",
          9191 => x"770682d8",
          9192 => x"c8084356",
          9193 => x"45748338",
          9194 => x"bf416655",
          9195 => x"8e566075",
          9196 => x"268a9038",
          9197 => x"74613170",
          9198 => x"485580ff",
          9199 => x"75278a83",
          9200 => x"38935678",
          9201 => x"81802689",
          9202 => x"fa387781",
          9203 => x"2a708106",
          9204 => x"56437480",
          9205 => x"2e953877",
          9206 => x"87065574",
          9207 => x"822e838d",
          9208 => x"38778106",
          9209 => x"5574802e",
          9210 => x"83833877",
          9211 => x"81065593",
          9212 => x"56825e74",
          9213 => x"802e89cb",
          9214 => x"38785a7d",
          9215 => x"832e0981",
          9216 => x"0680e138",
          9217 => x"78ae3866",
          9218 => x"912a5781",
          9219 => x"0b82cc84",
          9220 => x"22565a74",
          9221 => x"802e9d38",
          9222 => x"74772698",
          9223 => x"3882cc84",
          9224 => x"56791082",
          9225 => x"17702257",
          9226 => x"575a7480",
          9227 => x"2e863876",
          9228 => x"7527ee38",
          9229 => x"79526651",
          9230 => x"fea6c83f",
          9231 => x"82d8c808",
          9232 => x"84298487",
          9233 => x"0570892a",
          9234 => x"5e55a05c",
          9235 => x"800b82d8",
          9236 => x"c808fc80",
          9237 => x"8a055644",
          9238 => x"fdfff00a",
          9239 => x"752780ec",
          9240 => x"3888d339",
          9241 => x"78ae3866",
          9242 => x"8c2a5781",
          9243 => x"0b82cbf4",
          9244 => x"22565a74",
          9245 => x"802e9d38",
          9246 => x"74772698",
          9247 => x"3882cbf4",
          9248 => x"56791082",
          9249 => x"17702257",
          9250 => x"575a7480",
          9251 => x"2e863876",
          9252 => x"7527ee38",
          9253 => x"79526651",
          9254 => x"fea5e83f",
          9255 => x"82d8c808",
          9256 => x"10840557",
          9257 => x"82d8c808",
          9258 => x"9ff52696",
          9259 => x"38810b82",
          9260 => x"d8c80810",
          9261 => x"82d8c808",
          9262 => x"05711172",
          9263 => x"2a830559",
          9264 => x"565e83ff",
          9265 => x"17892a5d",
          9266 => x"815ca044",
          9267 => x"601c7d11",
          9268 => x"65056970",
          9269 => x"12ff0571",
          9270 => x"30707206",
          9271 => x"74315c52",
          9272 => x"59575940",
          9273 => x"7d832e09",
          9274 => x"81068938",
          9275 => x"761c6018",
          9276 => x"415c8439",
          9277 => x"761d5d79",
          9278 => x"90291870",
          9279 => x"62316858",
          9280 => x"51557476",
          9281 => x"2687af38",
          9282 => x"757c317d",
          9283 => x"317a5370",
          9284 => x"65315255",
          9285 => x"fea4ec3f",
          9286 => x"82d8c808",
          9287 => x"587d832e",
          9288 => x"0981069b",
          9289 => x"3882d8c8",
          9290 => x"0883fff5",
          9291 => x"2680dd38",
          9292 => x"78878338",
          9293 => x"79812a59",
          9294 => x"78fdbe38",
          9295 => x"86f8397d",
          9296 => x"822e0981",
          9297 => x"0680c538",
          9298 => x"83fff50b",
          9299 => x"82d8c808",
          9300 => x"27a03878",
          9301 => x"8f38791a",
          9302 => x"557480c0",
          9303 => x"26863874",
          9304 => x"59fd9639",
          9305 => x"62810655",
          9306 => x"74802e8f",
          9307 => x"38835efd",
          9308 => x"883982d8",
          9309 => x"c8089ff5",
          9310 => x"26923878",
          9311 => x"86b83879",
          9312 => x"1a598180",
          9313 => x"7927fcf1",
          9314 => x"3886ab39",
          9315 => x"80557d81",
          9316 => x"2e098106",
          9317 => x"83387d55",
          9318 => x"9ff57827",
          9319 => x"8b387481",
          9320 => x"06558e56",
          9321 => x"74869c38",
          9322 => x"84805380",
          9323 => x"527a51ff",
          9324 => x"90e73f8b",
          9325 => x"5382ca8c",
          9326 => x"527a51ff",
          9327 => x"90b83f84",
          9328 => x"80528b1b",
          9329 => x"51ff8fe1",
          9330 => x"3f798d1c",
          9331 => x"347b83ff",
          9332 => x"ff06528e",
          9333 => x"1b51ff8f",
          9334 => x"d03f810b",
          9335 => x"901c347d",
          9336 => x"83327030",
          9337 => x"70962a84",
          9338 => x"80065451",
          9339 => x"55911b51",
          9340 => x"ff8fb63f",
          9341 => x"66557483",
          9342 => x"ffff2690",
          9343 => x"387483ff",
          9344 => x"ff065293",
          9345 => x"1b51ff8f",
          9346 => x"a03f8a39",
          9347 => x"7452a01b",
          9348 => x"51ff8fb3",
          9349 => x"3ff80b95",
          9350 => x"1c34bf52",
          9351 => x"981b51ff",
          9352 => x"8f873f81",
          9353 => x"ff529a1b",
          9354 => x"51ff8efd",
          9355 => x"3f60529c",
          9356 => x"1b51ff8f",
          9357 => x"923f7d83",
          9358 => x"2e098106",
          9359 => x"80cb3882",
          9360 => x"88b20a52",
          9361 => x"80c31b51",
          9362 => x"ff8efc3f",
          9363 => x"7c52a41b",
          9364 => x"51ff8ef3",
          9365 => x"3f8252ac",
          9366 => x"1b51ff8e",
          9367 => x"ea3f8152",
          9368 => x"b01b51ff",
          9369 => x"8ec33f86",
          9370 => x"52b21b51",
          9371 => x"ff8eba3f",
          9372 => x"ff800b80",
          9373 => x"c01c34a9",
          9374 => x"0b80c21c",
          9375 => x"34935382",
          9376 => x"ca985280",
          9377 => x"c71b51ae",
          9378 => x"398288b2",
          9379 => x"0a52a71b",
          9380 => x"51ff8eb3",
          9381 => x"3f7c83ff",
          9382 => x"ff065296",
          9383 => x"1b51ff8e",
          9384 => x"883fff80",
          9385 => x"0ba41c34",
          9386 => x"a90ba61c",
          9387 => x"34935382",
          9388 => x"caac52ab",
          9389 => x"1b51ff8e",
          9390 => x"bd3f82d4",
          9391 => x"d55283fe",
          9392 => x"1b705259",
          9393 => x"ff8de23f",
          9394 => x"81546053",
          9395 => x"7a527e51",
          9396 => x"ff8a853f",
          9397 => x"815682d8",
          9398 => x"c80883e7",
          9399 => x"387d832e",
          9400 => x"09810680",
          9401 => x"ee387554",
          9402 => x"60860553",
          9403 => x"7a527e51",
          9404 => x"ff89e53f",
          9405 => x"84805380",
          9406 => x"527a51ff",
          9407 => x"8e9b3f84",
          9408 => x"8b85a4d2",
          9409 => x"527a51ff",
          9410 => x"8dbd3f86",
          9411 => x"8a85e4f2",
          9412 => x"5283e41b",
          9413 => x"51ff8daf",
          9414 => x"3fff1852",
          9415 => x"83e81b51",
          9416 => x"ff8da43f",
          9417 => x"825283ec",
          9418 => x"1b51ff8d",
          9419 => x"9a3f82d4",
          9420 => x"d5527851",
          9421 => x"ff8cf23f",
          9422 => x"75546087",
          9423 => x"05537a52",
          9424 => x"7e51ff89",
          9425 => x"933f7554",
          9426 => x"6016537a",
          9427 => x"527e51ff",
          9428 => x"89863f65",
          9429 => x"5380527a",
          9430 => x"51ff8dbd",
          9431 => x"3f7f5680",
          9432 => x"587d832e",
          9433 => x"0981069a",
          9434 => x"38f8527a",
          9435 => x"51ff8cd7",
          9436 => x"3fff5284",
          9437 => x"1b51ff8c",
          9438 => x"ce3ff00a",
          9439 => x"52881b51",
          9440 => x"913987ff",
          9441 => x"fff8557d",
          9442 => x"812e8338",
          9443 => x"f8557452",
          9444 => x"7a51ff8c",
          9445 => x"b23f7c55",
          9446 => x"61577462",
          9447 => x"26833874",
          9448 => x"57765475",
          9449 => x"537a527e",
          9450 => x"51ff88ac",
          9451 => x"3f82d8c8",
          9452 => x"08828738",
          9453 => x"84805382",
          9454 => x"d8c80852",
          9455 => x"7a51ff8c",
          9456 => x"d83f7616",
          9457 => x"75783156",
          9458 => x"5674cd38",
          9459 => x"81185877",
          9460 => x"802eff8d",
          9461 => x"3879557d",
          9462 => x"832e8338",
          9463 => x"63556157",
          9464 => x"74622683",
          9465 => x"38745776",
          9466 => x"5475537a",
          9467 => x"527e51ff",
          9468 => x"87e63f82",
          9469 => x"d8c80881",
          9470 => x"c1387616",
          9471 => x"75783156",
          9472 => x"5674db38",
          9473 => x"8c567d83",
          9474 => x"2e933886",
          9475 => x"566683ff",
          9476 => x"ff268a38",
          9477 => x"84567d82",
          9478 => x"2e833881",
          9479 => x"56648106",
          9480 => x"587780fe",
          9481 => x"38848053",
          9482 => x"77527a51",
          9483 => x"ff8bea3f",
          9484 => x"82d4d552",
          9485 => x"7851ff8a",
          9486 => x"f03f83be",
          9487 => x"1b557775",
          9488 => x"34810b81",
          9489 => x"1634810b",
          9490 => x"82163477",
          9491 => x"83163475",
          9492 => x"84163460",
          9493 => x"67055680",
          9494 => x"fdc15275",
          9495 => x"51fe9ea3",
          9496 => x"3ffe0b85",
          9497 => x"163482d8",
          9498 => x"c808822a",
          9499 => x"bf075675",
          9500 => x"86163482",
          9501 => x"d8c80887",
          9502 => x"16346052",
          9503 => x"83c61b51",
          9504 => x"ff8ac43f",
          9505 => x"665283ca",
          9506 => x"1b51ff8a",
          9507 => x"ba3f8154",
          9508 => x"77537a52",
          9509 => x"7e51ff86",
          9510 => x"bf3f8156",
          9511 => x"82d8c808",
          9512 => x"a2388053",
          9513 => x"80527e51",
          9514 => x"ff88913f",
          9515 => x"815682d8",
          9516 => x"c8089038",
          9517 => x"89398e56",
          9518 => x"8a398156",
          9519 => x"863982d8",
          9520 => x"c8085675",
          9521 => x"82d8c80c",
          9522 => x"993d0d04",
          9523 => x"f53d0d7d",
          9524 => x"605b5980",
          9525 => x"7960ff05",
          9526 => x"5a575776",
          9527 => x"7825b438",
          9528 => x"8d3df811",
          9529 => x"55558153",
          9530 => x"fc155279",
          9531 => x"51c9bd3f",
          9532 => x"7a812e09",
          9533 => x"81069c38",
          9534 => x"8c3d3355",
          9535 => x"748d2edb",
          9536 => x"38747670",
          9537 => x"81055834",
          9538 => x"81175774",
          9539 => x"8a2e0981",
          9540 => x"06c93880",
          9541 => x"76347855",
          9542 => x"76833876",
          9543 => x"557482d8",
          9544 => x"c80c8d3d",
          9545 => x"0d04f73d",
          9546 => x"0d7b0284",
          9547 => x"05b30533",
          9548 => x"5957778a",
          9549 => x"2e098106",
          9550 => x"87388d52",
          9551 => x"7651e73f",
          9552 => x"84170856",
          9553 => x"807624be",
          9554 => x"38881708",
          9555 => x"77178c05",
          9556 => x"56597775",
          9557 => x"34811656",
          9558 => x"bb7625a1",
          9559 => x"388b3dfc",
          9560 => x"05547553",
          9561 => x"8c175276",
          9562 => x"0851cbc0",
          9563 => x"3f797632",
          9564 => x"70307072",
          9565 => x"079f2a70",
          9566 => x"30535156",
          9567 => x"56758418",
          9568 => x"0c811988",
          9569 => x"180c8b3d",
          9570 => x"0d04f93d",
          9571 => x"0d798411",
          9572 => x"08565680",
          9573 => x"7524a738",
          9574 => x"893dfc05",
          9575 => x"5474538c",
          9576 => x"16527508",
          9577 => x"51cb853f",
          9578 => x"82d8c808",
          9579 => x"91388416",
          9580 => x"08782e09",
          9581 => x"81068738",
          9582 => x"88160855",
          9583 => x"8339ff55",
          9584 => x"7482d8c8",
          9585 => x"0c893d0d",
          9586 => x"04fd3d0d",
          9587 => x"755480cc",
          9588 => x"53805273",
          9589 => x"51ff88c1",
          9590 => x"3f76740c",
          9591 => x"853d0d04",
          9592 => x"ea3d0d02",
          9593 => x"80e30533",
          9594 => x"6a53863d",
          9595 => x"70535454",
          9596 => x"d83f7352",
          9597 => x"7251feae",
          9598 => x"3f7251ff",
          9599 => x"8d3f983d",
          9600 => x"0d04fd3d",
          9601 => x"0d750284",
          9602 => x"059a0522",
          9603 => x"55538052",
          9604 => x"7280ff26",
          9605 => x"8a387283",
          9606 => x"ffff0652",
          9607 => x"80c33983",
          9608 => x"ffff7327",
          9609 => x"517383b5",
          9610 => x"2e098106",
          9611 => x"b4387080",
          9612 => x"2eaf3882",
          9613 => x"cc942251",
          9614 => x"72712e9c",
          9615 => x"38811270",
          9616 => x"83ffff06",
          9617 => x"53517180",
          9618 => x"ff268d38",
          9619 => x"711082cc",
          9620 => x"94057022",
          9621 => x"5151e139",
          9622 => x"81801270",
          9623 => x"81ff0653",
          9624 => x"517182d8",
          9625 => x"c80c853d",
          9626 => x"0d04fe3d",
          9627 => x"0d029205",
          9628 => x"22028405",
          9629 => x"96052253",
          9630 => x"51805370",
          9631 => x"80ff2685",
          9632 => x"3870539a",
          9633 => x"397183b5",
          9634 => x"2e098106",
          9635 => x"91387081",
          9636 => x"ff268b38",
          9637 => x"701082ca",
          9638 => x"94057022",
          9639 => x"54517282",
          9640 => x"d8c80c84",
          9641 => x"3d0d04fb",
          9642 => x"3d0d7751",
          9643 => x"7083ffff",
          9644 => x"2681a738",
          9645 => x"7083ffff",
          9646 => x"0682ce94",
          9647 => x"57529fff",
          9648 => x"72278538",
          9649 => x"82d28856",
          9650 => x"75708205",
          9651 => x"57227030",
          9652 => x"70802572",
          9653 => x"75260751",
          9654 => x"52557080",
          9655 => x"fb387570",
          9656 => x"82055722",
          9657 => x"70882a71",
          9658 => x"81ff0670",
          9659 => x"18545255",
          9660 => x"53717125",
          9661 => x"80d73873",
          9662 => x"882680dc",
          9663 => x"38738429",
          9664 => x"82b0b005",
          9665 => x"51700804",
          9666 => x"71753110",
          9667 => x"76117022",
          9668 => x"54515180",
          9669 => x"c3397175",
          9670 => x"31810672",
          9671 => x"71315151",
          9672 => x"a439f012",
          9673 => x"519f39e0",
          9674 => x"12519a39",
          9675 => x"d0125195",
          9676 => x"39e61251",
          9677 => x"90398812",
          9678 => x"518b39ff",
          9679 => x"b0125185",
          9680 => x"39c7a012",
          9681 => x"517083ff",
          9682 => x"ff06528c",
          9683 => x"3973fef8",
          9684 => x"38721016",
          9685 => x"56fef139",
          9686 => x"71517082",
          9687 => x"d8c80c87",
          9688 => x"3d0d0400",
          9689 => x"00ffffff",
          9690 => x"ff00ffff",
          9691 => x"ffff00ff",
          9692 => x"ffffff00",
          9693 => x"00002baa",
          9694 => x"00002b2e",
          9695 => x"00002b35",
          9696 => x"00002b3c",
          9697 => x"00002b43",
          9698 => x"00002b4a",
          9699 => x"00002b51",
          9700 => x"00002b58",
          9701 => x"00002b5f",
          9702 => x"00002b66",
          9703 => x"00002b6d",
          9704 => x"00002b74",
          9705 => x"00002b7a",
          9706 => x"00002b80",
          9707 => x"00002b86",
          9708 => x"00002b8c",
          9709 => x"00002b92",
          9710 => x"00002b98",
          9711 => x"00002b9e",
          9712 => x"00002ba4",
          9713 => x"000043a6",
          9714 => x"000043ac",
          9715 => x"000043b2",
          9716 => x"000043b8",
          9717 => x"000043be",
          9718 => x"000049dd",
          9719 => x"00004add",
          9720 => x"00004bee",
          9721 => x"00004e46",
          9722 => x"00004ac5",
          9723 => x"000048b2",
          9724 => x"00004cb6",
          9725 => x"00004e17",
          9726 => x"00004cf9",
          9727 => x"00004d8f",
          9728 => x"00004d15",
          9729 => x"00004b98",
          9730 => x"000048b2",
          9731 => x"00004bee",
          9732 => x"00004c17",
          9733 => x"00004cb6",
          9734 => x"000048b2",
          9735 => x"000048b2",
          9736 => x"00004d15",
          9737 => x"00004d8f",
          9738 => x"00004e17",
          9739 => x"00004e46",
          9740 => x"00009708",
          9741 => x"00009716",
          9742 => x"00009722",
          9743 => x"00009727",
          9744 => x"0000972c",
          9745 => x"00009731",
          9746 => x"00009736",
          9747 => x"0000973b",
          9748 => x"00009741",
          9749 => x"00000e31",
          9750 => x"0000171a",
          9751 => x"0000171a",
          9752 => x"00000e60",
          9753 => x"0000171a",
          9754 => x"0000171a",
          9755 => x"0000171a",
          9756 => x"0000171a",
          9757 => x"0000171a",
          9758 => x"0000171a",
          9759 => x"0000171a",
          9760 => x"00000e1d",
          9761 => x"0000171a",
          9762 => x"00000e48",
          9763 => x"00000e78",
          9764 => x"0000171a",
          9765 => x"0000171a",
          9766 => x"0000171a",
          9767 => x"0000171a",
          9768 => x"0000171a",
          9769 => x"0000171a",
          9770 => x"0000171a",
          9771 => x"0000171a",
          9772 => x"0000171a",
          9773 => x"0000171a",
          9774 => x"0000171a",
          9775 => x"0000171a",
          9776 => x"0000171a",
          9777 => x"0000171a",
          9778 => x"0000171a",
          9779 => x"0000171a",
          9780 => x"0000171a",
          9781 => x"0000171a",
          9782 => x"0000171a",
          9783 => x"0000171a",
          9784 => x"0000171a",
          9785 => x"0000171a",
          9786 => x"0000171a",
          9787 => x"0000171a",
          9788 => x"0000171a",
          9789 => x"0000171a",
          9790 => x"0000171a",
          9791 => x"0000171a",
          9792 => x"0000171a",
          9793 => x"0000171a",
          9794 => x"0000171a",
          9795 => x"0000171a",
          9796 => x"0000171a",
          9797 => x"0000171a",
          9798 => x"0000171a",
          9799 => x"0000171a",
          9800 => x"00000fa8",
          9801 => x"0000171a",
          9802 => x"0000171a",
          9803 => x"0000171a",
          9804 => x"0000171a",
          9805 => x"00001116",
          9806 => x"0000171a",
          9807 => x"0000171a",
          9808 => x"0000171a",
          9809 => x"0000171a",
          9810 => x"0000171a",
          9811 => x"0000171a",
          9812 => x"0000171a",
          9813 => x"0000171a",
          9814 => x"0000171a",
          9815 => x"0000171a",
          9816 => x"00000ed8",
          9817 => x"0000103f",
          9818 => x"00000eaf",
          9819 => x"00000eaf",
          9820 => x"00000eaf",
          9821 => x"0000171a",
          9822 => x"0000103f",
          9823 => x"0000171a",
          9824 => x"0000171a",
          9825 => x"00000e98",
          9826 => x"0000171a",
          9827 => x"0000171a",
          9828 => x"000010ec",
          9829 => x"000010f7",
          9830 => x"0000171a",
          9831 => x"0000171a",
          9832 => x"00000f11",
          9833 => x"0000171a",
          9834 => x"0000111f",
          9835 => x"0000171a",
          9836 => x"0000171a",
          9837 => x"00001116",
          9838 => x"64696e69",
          9839 => x"74000000",
          9840 => x"64696f63",
          9841 => x"746c0000",
          9842 => x"66696e69",
          9843 => x"74000000",
          9844 => x"666c6f61",
          9845 => x"64000000",
          9846 => x"66657865",
          9847 => x"63000000",
          9848 => x"6d636c65",
          9849 => x"61720000",
          9850 => x"6d636f70",
          9851 => x"79000000",
          9852 => x"6d646966",
          9853 => x"66000000",
          9854 => x"6d64756d",
          9855 => x"70000000",
          9856 => x"6d656200",
          9857 => x"6d656800",
          9858 => x"6d657700",
          9859 => x"68696400",
          9860 => x"68696500",
          9861 => x"68666400",
          9862 => x"68666500",
          9863 => x"63616c6c",
          9864 => x"00000000",
          9865 => x"6a6d7000",
          9866 => x"72657374",
          9867 => x"61727400",
          9868 => x"72657365",
          9869 => x"74000000",
          9870 => x"696e666f",
          9871 => x"00000000",
          9872 => x"74657374",
          9873 => x"00000000",
          9874 => x"74626173",
          9875 => x"69630000",
          9876 => x"6d626173",
          9877 => x"69630000",
          9878 => x"6b696c6f",
          9879 => x"00000000",
          9880 => x"65640000",
          9881 => x"4469736b",
          9882 => x"20457272",
          9883 => x"6f720000",
          9884 => x"496e7465",
          9885 => x"726e616c",
          9886 => x"20657272",
          9887 => x"6f722e00",
          9888 => x"4469736b",
          9889 => x"206e6f74",
          9890 => x"20726561",
          9891 => x"64792e00",
          9892 => x"4e6f2066",
          9893 => x"696c6520",
          9894 => x"666f756e",
          9895 => x"642e0000",
          9896 => x"4e6f2070",
          9897 => x"61746820",
          9898 => x"666f756e",
          9899 => x"642e0000",
          9900 => x"496e7661",
          9901 => x"6c696420",
          9902 => x"66696c65",
          9903 => x"6e616d65",
          9904 => x"2e000000",
          9905 => x"41636365",
          9906 => x"73732064",
          9907 => x"656e6965",
          9908 => x"642e0000",
          9909 => x"46696c65",
          9910 => x"20616c72",
          9911 => x"65616479",
          9912 => x"20657869",
          9913 => x"7374732e",
          9914 => x"00000000",
          9915 => x"46696c65",
          9916 => x"2068616e",
          9917 => x"646c6520",
          9918 => x"696e7661",
          9919 => x"6c69642e",
          9920 => x"00000000",
          9921 => x"53442069",
          9922 => x"73207772",
          9923 => x"69746520",
          9924 => x"70726f74",
          9925 => x"65637465",
          9926 => x"642e0000",
          9927 => x"44726976",
          9928 => x"65206e75",
          9929 => x"6d626572",
          9930 => x"20697320",
          9931 => x"696e7661",
          9932 => x"6c69642e",
          9933 => x"00000000",
          9934 => x"4469736b",
          9935 => x"206e6f74",
          9936 => x"20656e61",
          9937 => x"626c6564",
          9938 => x"2e000000",
          9939 => x"4e6f2063",
          9940 => x"6f6d7061",
          9941 => x"7469626c",
          9942 => x"65206669",
          9943 => x"6c657379",
          9944 => x"7374656d",
          9945 => x"20666f75",
          9946 => x"6e64206f",
          9947 => x"6e206469",
          9948 => x"736b2e00",
          9949 => x"466f726d",
          9950 => x"61742061",
          9951 => x"626f7274",
          9952 => x"65642e00",
          9953 => x"54696d65",
          9954 => x"6f75742c",
          9955 => x"206f7065",
          9956 => x"72617469",
          9957 => x"6f6e2063",
          9958 => x"616e6365",
          9959 => x"6c6c6564",
          9960 => x"2e000000",
          9961 => x"46696c65",
          9962 => x"20697320",
          9963 => x"6c6f636b",
          9964 => x"65642e00",
          9965 => x"496e7375",
          9966 => x"66666963",
          9967 => x"69656e74",
          9968 => x"206d656d",
          9969 => x"6f72792e",
          9970 => x"00000000",
          9971 => x"546f6f20",
          9972 => x"6d616e79",
          9973 => x"206f7065",
          9974 => x"6e206669",
          9975 => x"6c65732e",
          9976 => x"00000000",
          9977 => x"50617261",
          9978 => x"6d657465",
          9979 => x"72732069",
          9980 => x"6e636f72",
          9981 => x"72656374",
          9982 => x"2e000000",
          9983 => x"53756363",
          9984 => x"6573732e",
          9985 => x"00000000",
          9986 => x"556e6b6e",
          9987 => x"6f776e20",
          9988 => x"6572726f",
          9989 => x"722e0000",
          9990 => x"0a256c75",
          9991 => x"20627974",
          9992 => x"65732025",
          9993 => x"73206174",
          9994 => x"20256c75",
          9995 => x"20627974",
          9996 => x"65732f73",
          9997 => x"65632e0a",
          9998 => x"00000000",
          9999 => x"72656164",
         10000 => x"00000000",
         10001 => x"303d2530",
         10002 => x"386c782c",
         10003 => x"20313d25",
         10004 => x"30386c78",
         10005 => x"2c20323d",
         10006 => x"2530386c",
         10007 => x"782c205f",
         10008 => x"494f423d",
         10009 => x"2530386c",
         10010 => x"78202530",
         10011 => x"386c7820",
         10012 => x"2530386c",
         10013 => x"780a0000",
         10014 => x"2530386c",
         10015 => x"58000000",
         10016 => x"3a202000",
         10017 => x"25303458",
         10018 => x"00000000",
         10019 => x"20202020",
         10020 => x"20202020",
         10021 => x"00000000",
         10022 => x"25303258",
         10023 => x"00000000",
         10024 => x"20200000",
         10025 => x"207c0000",
         10026 => x"7c000000",
         10027 => x"5a505554",
         10028 => x"41000000",
         10029 => x"0a2a2a20",
         10030 => x"25732028",
         10031 => x"00000000",
         10032 => x"30322f30",
         10033 => x"352f3230",
         10034 => x"32300000",
         10035 => x"76312e35",
         10036 => x"32000000",
         10037 => x"205a5055",
         10038 => x"2c207265",
         10039 => x"76202530",
         10040 => x"32782920",
         10041 => x"25732025",
         10042 => x"73202a2a",
         10043 => x"0a0a0000",
         10044 => x"5a505554",
         10045 => x"4120496e",
         10046 => x"74657272",
         10047 => x"75707420",
         10048 => x"48616e64",
         10049 => x"6c657200",
         10050 => x"54696d65",
         10051 => x"7220696e",
         10052 => x"74657272",
         10053 => x"75707400",
         10054 => x"50533220",
         10055 => x"696e7465",
         10056 => x"72727570",
         10057 => x"74000000",
         10058 => x"494f4354",
         10059 => x"4c205244",
         10060 => x"20696e74",
         10061 => x"65727275",
         10062 => x"70740000",
         10063 => x"494f4354",
         10064 => x"4c205752",
         10065 => x"20696e74",
         10066 => x"65727275",
         10067 => x"70740000",
         10068 => x"55415254",
         10069 => x"30205258",
         10070 => x"20696e74",
         10071 => x"65727275",
         10072 => x"70740000",
         10073 => x"55415254",
         10074 => x"30205458",
         10075 => x"20696e74",
         10076 => x"65727275",
         10077 => x"70740000",
         10078 => x"55415254",
         10079 => x"31205258",
         10080 => x"20696e74",
         10081 => x"65727275",
         10082 => x"70740000",
         10083 => x"55415254",
         10084 => x"31205458",
         10085 => x"20696e74",
         10086 => x"65727275",
         10087 => x"70740000",
         10088 => x"53657474",
         10089 => x"696e6720",
         10090 => x"75702074",
         10091 => x"696d6572",
         10092 => x"2e2e2e00",
         10093 => x"456e6162",
         10094 => x"6c696e67",
         10095 => x"2074696d",
         10096 => x"65722e2e",
         10097 => x"2e000000",
         10098 => x"6175746f",
         10099 => x"65786563",
         10100 => x"2e626174",
         10101 => x"00000000",
         10102 => x"7a707574",
         10103 => x"612e6873",
         10104 => x"74000000",
         10105 => x"303a0000",
         10106 => x"4661696c",
         10107 => x"65642074",
         10108 => x"6f20696e",
         10109 => x"69746961",
         10110 => x"6c697365",
         10111 => x"20736420",
         10112 => x"63617264",
         10113 => x"20302c20",
         10114 => x"706c6561",
         10115 => x"73652069",
         10116 => x"6e697420",
         10117 => x"6d616e75",
         10118 => x"616c6c79",
         10119 => x"2e000000",
         10120 => x"2a200000",
         10121 => x"42616420",
         10122 => x"6469736b",
         10123 => x"20696421",
         10124 => x"00000000",
         10125 => x"496e6974",
         10126 => x"69616c69",
         10127 => x"7365642e",
         10128 => x"00000000",
         10129 => x"4661696c",
         10130 => x"65642074",
         10131 => x"6f20696e",
         10132 => x"69746961",
         10133 => x"6c697365",
         10134 => x"2e000000",
         10135 => x"72633d25",
         10136 => x"640a0000",
         10137 => x"25753a00",
         10138 => x"436c6561",
         10139 => x"72696e67",
         10140 => x"2e2e2e2e",
         10141 => x"00000000",
         10142 => x"436f7079",
         10143 => x"696e672e",
         10144 => x"2e2e0000",
         10145 => x"436f6d70",
         10146 => x"6172696e",
         10147 => x"672e2e2e",
         10148 => x"00000000",
         10149 => x"2530386c",
         10150 => x"78282530",
         10151 => x"3878292d",
         10152 => x"3e253038",
         10153 => x"6c782825",
         10154 => x"30387829",
         10155 => x"0a000000",
         10156 => x"44756d70",
         10157 => x"204d656d",
         10158 => x"6f727900",
         10159 => x"0a436f6d",
         10160 => x"706c6574",
         10161 => x"652e0000",
         10162 => x"2530386c",
         10163 => x"58202530",
         10164 => x"32582d00",
         10165 => x"3f3f3f00",
         10166 => x"2530386c",
         10167 => x"58202530",
         10168 => x"34582d00",
         10169 => x"2530386c",
         10170 => x"58202530",
         10171 => x"386c582d",
         10172 => x"00000000",
         10173 => x"44697361",
         10174 => x"626c696e",
         10175 => x"6720696e",
         10176 => x"74657272",
         10177 => x"75707473",
         10178 => x"00000000",
         10179 => x"456e6162",
         10180 => x"6c696e67",
         10181 => x"20696e74",
         10182 => x"65727275",
         10183 => x"70747300",
         10184 => x"44697361",
         10185 => x"626c6564",
         10186 => x"20756172",
         10187 => x"74206669",
         10188 => x"666f0000",
         10189 => x"456e6162",
         10190 => x"6c696e67",
         10191 => x"20756172",
         10192 => x"74206669",
         10193 => x"666f0000",
         10194 => x"45786563",
         10195 => x"7574696e",
         10196 => x"6720636f",
         10197 => x"64652040",
         10198 => x"20253038",
         10199 => x"6c78202e",
         10200 => x"2e2e0a00",
         10201 => x"43616c6c",
         10202 => x"696e6720",
         10203 => x"636f6465",
         10204 => x"20402025",
         10205 => x"30386c78",
         10206 => x"202e2e2e",
         10207 => x"0a000000",
         10208 => x"43616c6c",
         10209 => x"20726574",
         10210 => x"75726e65",
         10211 => x"6420636f",
         10212 => x"64652028",
         10213 => x"2564292e",
         10214 => x"0a000000",
         10215 => x"52657374",
         10216 => x"61727469",
         10217 => x"6e672061",
         10218 => x"70706c69",
         10219 => x"63617469",
         10220 => x"6f6e2e2e",
         10221 => x"2e000000",
         10222 => x"436f6c64",
         10223 => x"20726562",
         10224 => x"6f6f7469",
         10225 => x"6e672e2e",
         10226 => x"2e000000",
         10227 => x"5a505500",
         10228 => x"62696e00",
         10229 => x"25643a5c",
         10230 => x"25735c25",
         10231 => x"732e2573",
         10232 => x"00000000",
         10233 => x"25643a5c",
         10234 => x"25735c25",
         10235 => x"73000000",
         10236 => x"25643a5c",
         10237 => x"25730000",
         10238 => x"42616420",
         10239 => x"636f6d6d",
         10240 => x"616e642e",
         10241 => x"00000000",
         10242 => x"52756e6e",
         10243 => x"696e672e",
         10244 => x"2e2e0000",
         10245 => x"456e6162",
         10246 => x"6c696e67",
         10247 => x"20696e74",
         10248 => x"65727275",
         10249 => x"7074732e",
         10250 => x"2e2e0000",
         10251 => x"25642f25",
         10252 => x"642f2564",
         10253 => x"2025643a",
         10254 => x"25643a25",
         10255 => x"642e2564",
         10256 => x"25640a00",
         10257 => x"536f4320",
         10258 => x"436f6e66",
         10259 => x"69677572",
         10260 => x"6174696f",
         10261 => x"6e000000",
         10262 => x"20286672",
         10263 => x"6f6d2053",
         10264 => x"6f432063",
         10265 => x"6f6e6669",
         10266 => x"67290000",
         10267 => x"3a0a4465",
         10268 => x"76696365",
         10269 => x"7320696d",
         10270 => x"706c656d",
         10271 => x"656e7465",
         10272 => x"643a0000",
         10273 => x"20202020",
         10274 => x"57422053",
         10275 => x"4452414d",
         10276 => x"20202825",
         10277 => x"3038583a",
         10278 => x"25303858",
         10279 => x"292e0a00",
         10280 => x"20202020",
         10281 => x"53445241",
         10282 => x"4d202020",
         10283 => x"20202825",
         10284 => x"3038583a",
         10285 => x"25303858",
         10286 => x"292e0a00",
         10287 => x"20202020",
         10288 => x"494e534e",
         10289 => x"20425241",
         10290 => x"4d202825",
         10291 => x"3038583a",
         10292 => x"25303858",
         10293 => x"292e0a00",
         10294 => x"20202020",
         10295 => x"4252414d",
         10296 => x"20202020",
         10297 => x"20202825",
         10298 => x"3038583a",
         10299 => x"25303858",
         10300 => x"292e0a00",
         10301 => x"20202020",
         10302 => x"52414d20",
         10303 => x"20202020",
         10304 => x"20202825",
         10305 => x"3038583a",
         10306 => x"25303858",
         10307 => x"292e0a00",
         10308 => x"20202020",
         10309 => x"53442043",
         10310 => x"41524420",
         10311 => x"20202844",
         10312 => x"65766963",
         10313 => x"6573203d",
         10314 => x"25303264",
         10315 => x"292e0a00",
         10316 => x"20202020",
         10317 => x"54494d45",
         10318 => x"52312020",
         10319 => x"20202854",
         10320 => x"696d6572",
         10321 => x"7320203d",
         10322 => x"25303264",
         10323 => x"292e0a00",
         10324 => x"20202020",
         10325 => x"494e5452",
         10326 => x"20435452",
         10327 => x"4c202843",
         10328 => x"68616e6e",
         10329 => x"656c733d",
         10330 => x"25303264",
         10331 => x"292e0a00",
         10332 => x"20202020",
         10333 => x"57495348",
         10334 => x"424f4e45",
         10335 => x"20425553",
         10336 => x"00000000",
         10337 => x"20202020",
         10338 => x"57422049",
         10339 => x"32430000",
         10340 => x"20202020",
         10341 => x"494f4354",
         10342 => x"4c000000",
         10343 => x"20202020",
         10344 => x"50533200",
         10345 => x"20202020",
         10346 => x"53504900",
         10347 => x"41646472",
         10348 => x"65737365",
         10349 => x"733a0000",
         10350 => x"20202020",
         10351 => x"43505520",
         10352 => x"52657365",
         10353 => x"74205665",
         10354 => x"63746f72",
         10355 => x"20416464",
         10356 => x"72657373",
         10357 => x"203d2025",
         10358 => x"3038580a",
         10359 => x"00000000",
         10360 => x"20202020",
         10361 => x"43505520",
         10362 => x"4d656d6f",
         10363 => x"72792053",
         10364 => x"74617274",
         10365 => x"20416464",
         10366 => x"72657373",
         10367 => x"203d2025",
         10368 => x"3038580a",
         10369 => x"00000000",
         10370 => x"20202020",
         10371 => x"53746163",
         10372 => x"6b205374",
         10373 => x"61727420",
         10374 => x"41646472",
         10375 => x"65737320",
         10376 => x"20202020",
         10377 => x"203d2025",
         10378 => x"3038580a",
         10379 => x"00000000",
         10380 => x"4d697363",
         10381 => x"3a000000",
         10382 => x"20202020",
         10383 => x"5a505520",
         10384 => x"49642020",
         10385 => x"20202020",
         10386 => x"20202020",
         10387 => x"20202020",
         10388 => x"20202020",
         10389 => x"203d2025",
         10390 => x"3034580a",
         10391 => x"00000000",
         10392 => x"20202020",
         10393 => x"53797374",
         10394 => x"656d2043",
         10395 => x"6c6f636b",
         10396 => x"20467265",
         10397 => x"71202020",
         10398 => x"20202020",
         10399 => x"203d2025",
         10400 => x"642e2530",
         10401 => x"34644d48",
         10402 => x"7a0a0000",
         10403 => x"20202020",
         10404 => x"53445241",
         10405 => x"4d20436c",
         10406 => x"6f636b20",
         10407 => x"46726571",
         10408 => x"20202020",
         10409 => x"20202020",
         10410 => x"203d2025",
         10411 => x"642e2530",
         10412 => x"34644d48",
         10413 => x"7a0a0000",
         10414 => x"20202020",
         10415 => x"57697368",
         10416 => x"626f6e65",
         10417 => x"20534452",
         10418 => x"414d2043",
         10419 => x"6c6f636b",
         10420 => x"20467265",
         10421 => x"713d2025",
         10422 => x"642e2530",
         10423 => x"34644d48",
         10424 => x"7a0a0000",
         10425 => x"536d616c",
         10426 => x"6c000000",
         10427 => x"4d656469",
         10428 => x"756d0000",
         10429 => x"466c6578",
         10430 => x"00000000",
         10431 => x"45564f00",
         10432 => x"45564f6d",
         10433 => x"00000000",
         10434 => x"556e6b6e",
         10435 => x"6f776e00",
         10436 => x"0000a46c",
         10437 => x"01000000",
         10438 => x"00000002",
         10439 => x"0000a468",
         10440 => x"01000000",
         10441 => x"00000003",
         10442 => x"0000a464",
         10443 => x"01000000",
         10444 => x"00000004",
         10445 => x"0000a460",
         10446 => x"01000000",
         10447 => x"00000005",
         10448 => x"0000a45c",
         10449 => x"01000000",
         10450 => x"00000006",
         10451 => x"0000a458",
         10452 => x"01000000",
         10453 => x"00000007",
         10454 => x"0000a454",
         10455 => x"01000000",
         10456 => x"00000001",
         10457 => x"0000a450",
         10458 => x"01000000",
         10459 => x"00000008",
         10460 => x"0000a44c",
         10461 => x"01000000",
         10462 => x"0000000b",
         10463 => x"0000a448",
         10464 => x"01000000",
         10465 => x"00000009",
         10466 => x"0000a444",
         10467 => x"01000000",
         10468 => x"0000000a",
         10469 => x"0000a440",
         10470 => x"04000000",
         10471 => x"0000000d",
         10472 => x"0000a43c",
         10473 => x"04000000",
         10474 => x"0000000c",
         10475 => x"0000a438",
         10476 => x"04000000",
         10477 => x"0000000e",
         10478 => x"0000a434",
         10479 => x"03000000",
         10480 => x"0000000f",
         10481 => x"0000a430",
         10482 => x"04000000",
         10483 => x"0000000f",
         10484 => x"0000a42c",
         10485 => x"04000000",
         10486 => x"00000010",
         10487 => x"0000a428",
         10488 => x"04000000",
         10489 => x"00000011",
         10490 => x"0000a424",
         10491 => x"03000000",
         10492 => x"00000012",
         10493 => x"0000a420",
         10494 => x"03000000",
         10495 => x"00000013",
         10496 => x"0000a41c",
         10497 => x"03000000",
         10498 => x"00000014",
         10499 => x"0000a418",
         10500 => x"03000000",
         10501 => x"00000015",
         10502 => x"1b5b4400",
         10503 => x"1b5b4300",
         10504 => x"1b5b4200",
         10505 => x"1b5b4100",
         10506 => x"1b5b367e",
         10507 => x"1b5b357e",
         10508 => x"1b5b347e",
         10509 => x"1b304600",
         10510 => x"1b5b337e",
         10511 => x"1b5b327e",
         10512 => x"1b5b317e",
         10513 => x"10000000",
         10514 => x"0e000000",
         10515 => x"0d000000",
         10516 => x"0b000000",
         10517 => x"08000000",
         10518 => x"06000000",
         10519 => x"05000000",
         10520 => x"04000000",
         10521 => x"03000000",
         10522 => x"02000000",
         10523 => x"01000000",
         10524 => x"68697374",
         10525 => x"6f727900",
         10526 => x"68697374",
         10527 => x"00000000",
         10528 => x"21000000",
         10529 => x"2530346c",
         10530 => x"75202025",
         10531 => x"730a0000",
         10532 => x"4661696c",
         10533 => x"65642074",
         10534 => x"6f207265",
         10535 => x"73657420",
         10536 => x"74686520",
         10537 => x"68697374",
         10538 => x"6f727920",
         10539 => x"66696c65",
         10540 => x"20746f20",
         10541 => x"454f462e",
         10542 => x"00000000",
         10543 => x"43616e6e",
         10544 => x"6f74206f",
         10545 => x"70656e2f",
         10546 => x"63726561",
         10547 => x"74652068",
         10548 => x"6973746f",
         10549 => x"72792066",
         10550 => x"696c652c",
         10551 => x"20646973",
         10552 => x"61626c69",
         10553 => x"6e672e00",
         10554 => x"53440000",
         10555 => x"222a3a3c",
         10556 => x"3e3f7c7f",
         10557 => x"00000000",
         10558 => x"2b2c3b3d",
         10559 => x"5b5d0000",
         10560 => x"46415400",
         10561 => x"46415433",
         10562 => x"32000000",
         10563 => x"ebfe904d",
         10564 => x"53444f53",
         10565 => x"352e3000",
         10566 => x"4e4f204e",
         10567 => x"414d4520",
         10568 => x"20202046",
         10569 => x"41543332",
         10570 => x"20202000",
         10571 => x"4e4f204e",
         10572 => x"414d4520",
         10573 => x"20202046",
         10574 => x"41542020",
         10575 => x"20202000",
         10576 => x"0000a4e8",
         10577 => x"00000000",
         10578 => x"00000000",
         10579 => x"00000000",
         10580 => x"01030507",
         10581 => x"090e1012",
         10582 => x"1416181c",
         10583 => x"1e000000",
         10584 => x"809a4541",
         10585 => x"8e418f80",
         10586 => x"45454549",
         10587 => x"49498e8f",
         10588 => x"9092924f",
         10589 => x"994f5555",
         10590 => x"59999a9b",
         10591 => x"9c9d9e9f",
         10592 => x"41494f55",
         10593 => x"a5a5a6a7",
         10594 => x"a8a9aaab",
         10595 => x"acadaeaf",
         10596 => x"b0b1b2b3",
         10597 => x"b4b5b6b7",
         10598 => x"b8b9babb",
         10599 => x"bcbdbebf",
         10600 => x"c0c1c2c3",
         10601 => x"c4c5c6c7",
         10602 => x"c8c9cacb",
         10603 => x"cccdcecf",
         10604 => x"d0d1d2d3",
         10605 => x"d4d5d6d7",
         10606 => x"d8d9dadb",
         10607 => x"dcdddedf",
         10608 => x"e0e1e2e3",
         10609 => x"e4e5e6e7",
         10610 => x"e8e9eaeb",
         10611 => x"ecedeeef",
         10612 => x"f0f1f2f3",
         10613 => x"f4f5f6f7",
         10614 => x"f8f9fafb",
         10615 => x"fcfdfeff",
         10616 => x"2b2e2c3b",
         10617 => x"3d5b5d2f",
         10618 => x"5c222a3a",
         10619 => x"3c3e3f7c",
         10620 => x"7f000000",
         10621 => x"00010004",
         10622 => x"00100040",
         10623 => x"01000200",
         10624 => x"00000000",
         10625 => x"00010002",
         10626 => x"00040008",
         10627 => x"00100020",
         10628 => x"00000000",
         10629 => x"00c700fc",
         10630 => x"00e900e2",
         10631 => x"00e400e0",
         10632 => x"00e500e7",
         10633 => x"00ea00eb",
         10634 => x"00e800ef",
         10635 => x"00ee00ec",
         10636 => x"00c400c5",
         10637 => x"00c900e6",
         10638 => x"00c600f4",
         10639 => x"00f600f2",
         10640 => x"00fb00f9",
         10641 => x"00ff00d6",
         10642 => x"00dc00a2",
         10643 => x"00a300a5",
         10644 => x"20a70192",
         10645 => x"00e100ed",
         10646 => x"00f300fa",
         10647 => x"00f100d1",
         10648 => x"00aa00ba",
         10649 => x"00bf2310",
         10650 => x"00ac00bd",
         10651 => x"00bc00a1",
         10652 => x"00ab00bb",
         10653 => x"25912592",
         10654 => x"25932502",
         10655 => x"25242561",
         10656 => x"25622556",
         10657 => x"25552563",
         10658 => x"25512557",
         10659 => x"255d255c",
         10660 => x"255b2510",
         10661 => x"25142534",
         10662 => x"252c251c",
         10663 => x"2500253c",
         10664 => x"255e255f",
         10665 => x"255a2554",
         10666 => x"25692566",
         10667 => x"25602550",
         10668 => x"256c2567",
         10669 => x"25682564",
         10670 => x"25652559",
         10671 => x"25582552",
         10672 => x"2553256b",
         10673 => x"256a2518",
         10674 => x"250c2588",
         10675 => x"2584258c",
         10676 => x"25902580",
         10677 => x"03b100df",
         10678 => x"039303c0",
         10679 => x"03a303c3",
         10680 => x"00b503c4",
         10681 => x"03a60398",
         10682 => x"03a903b4",
         10683 => x"221e03c6",
         10684 => x"03b52229",
         10685 => x"226100b1",
         10686 => x"22652264",
         10687 => x"23202321",
         10688 => x"00f72248",
         10689 => x"00b02219",
         10690 => x"00b7221a",
         10691 => x"207f00b2",
         10692 => x"25a000a0",
         10693 => x"0061031a",
         10694 => x"00e00317",
         10695 => x"00f80307",
         10696 => x"00ff0001",
         10697 => x"01780100",
         10698 => x"01300132",
         10699 => x"01060139",
         10700 => x"0110014a",
         10701 => x"012e0179",
         10702 => x"01060180",
         10703 => x"004d0243",
         10704 => x"01810182",
         10705 => x"01820184",
         10706 => x"01840186",
         10707 => x"01870187",
         10708 => x"0189018a",
         10709 => x"018b018b",
         10710 => x"018d018e",
         10711 => x"018f0190",
         10712 => x"01910191",
         10713 => x"01930194",
         10714 => x"01f60196",
         10715 => x"01970198",
         10716 => x"0198023d",
         10717 => x"019b019c",
         10718 => x"019d0220",
         10719 => x"019f01a0",
         10720 => x"01a001a2",
         10721 => x"01a201a4",
         10722 => x"01a401a6",
         10723 => x"01a701a7",
         10724 => x"01a901aa",
         10725 => x"01ab01ac",
         10726 => x"01ac01ae",
         10727 => x"01af01af",
         10728 => x"01b101b2",
         10729 => x"01b301b3",
         10730 => x"01b501b5",
         10731 => x"01b701b8",
         10732 => x"01b801ba",
         10733 => x"01bb01bc",
         10734 => x"01bc01be",
         10735 => x"01f701c0",
         10736 => x"01c101c2",
         10737 => x"01c301c4",
         10738 => x"01c501c4",
         10739 => x"01c701c8",
         10740 => x"01c701ca",
         10741 => x"01cb01ca",
         10742 => x"01cd0110",
         10743 => x"01dd0001",
         10744 => x"018e01de",
         10745 => x"011201f3",
         10746 => x"000301f1",
         10747 => x"01f401f4",
         10748 => x"01f80128",
         10749 => x"02220112",
         10750 => x"023a0009",
         10751 => x"2c65023b",
         10752 => x"023b023d",
         10753 => x"2c66023f",
         10754 => x"02400241",
         10755 => x"02410246",
         10756 => x"010a0253",
         10757 => x"00400181",
         10758 => x"01860255",
         10759 => x"0189018a",
         10760 => x"0258018f",
         10761 => x"025a0190",
         10762 => x"025c025d",
         10763 => x"025e025f",
         10764 => x"01930261",
         10765 => x"02620194",
         10766 => x"02640265",
         10767 => x"02660267",
         10768 => x"01970196",
         10769 => x"026a2c62",
         10770 => x"026c026d",
         10771 => x"026e019c",
         10772 => x"02700271",
         10773 => x"019d0273",
         10774 => x"0274019f",
         10775 => x"02760277",
         10776 => x"02780279",
         10777 => x"027a027b",
         10778 => x"027c2c64",
         10779 => x"027e027f",
         10780 => x"01a60281",
         10781 => x"028201a9",
         10782 => x"02840285",
         10783 => x"02860287",
         10784 => x"01ae0244",
         10785 => x"01b101b2",
         10786 => x"0245028d",
         10787 => x"028e028f",
         10788 => x"02900291",
         10789 => x"01b7037b",
         10790 => x"000303fd",
         10791 => x"03fe03ff",
         10792 => x"03ac0004",
         10793 => x"03860388",
         10794 => x"0389038a",
         10795 => x"03b10311",
         10796 => x"03c20002",
         10797 => x"03a303a3",
         10798 => x"03c40308",
         10799 => x"03cc0003",
         10800 => x"038c038e",
         10801 => x"038f03d8",
         10802 => x"011803f2",
         10803 => x"000a03f9",
         10804 => x"03f303f4",
         10805 => x"03f503f6",
         10806 => x"03f703f7",
         10807 => x"03f903fa",
         10808 => x"03fa0430",
         10809 => x"03200450",
         10810 => x"07100460",
         10811 => x"0122048a",
         10812 => x"013604c1",
         10813 => x"010e04cf",
         10814 => x"000104c0",
         10815 => x"04d00144",
         10816 => x"05610426",
         10817 => x"00000000",
         10818 => x"1d7d0001",
         10819 => x"2c631e00",
         10820 => x"01961ea0",
         10821 => x"015a1f00",
         10822 => x"06081f10",
         10823 => x"06061f20",
         10824 => x"06081f30",
         10825 => x"06081f40",
         10826 => x"06061f51",
         10827 => x"00071f59",
         10828 => x"1f521f5b",
         10829 => x"1f541f5d",
         10830 => x"1f561f5f",
         10831 => x"1f600608",
         10832 => x"1f70000e",
         10833 => x"1fba1fbb",
         10834 => x"1fc81fc9",
         10835 => x"1fca1fcb",
         10836 => x"1fda1fdb",
         10837 => x"1ff81ff9",
         10838 => x"1fea1feb",
         10839 => x"1ffa1ffb",
         10840 => x"1f800608",
         10841 => x"1f900608",
         10842 => x"1fa00608",
         10843 => x"1fb00004",
         10844 => x"1fb81fb9",
         10845 => x"1fb21fbc",
         10846 => x"1fcc0001",
         10847 => x"1fc31fd0",
         10848 => x"06021fe0",
         10849 => x"06021fe5",
         10850 => x"00011fec",
         10851 => x"1ff30001",
         10852 => x"1ffc214e",
         10853 => x"00012132",
         10854 => x"21700210",
         10855 => x"21840001",
         10856 => x"218324d0",
         10857 => x"051a2c30",
         10858 => x"042f2c60",
         10859 => x"01022c67",
         10860 => x"01062c75",
         10861 => x"01022c80",
         10862 => x"01642d00",
         10863 => x"0826ff41",
         10864 => x"031a0000",
         10865 => x"00000000",
         10866 => x"000099b8",
         10867 => x"01020100",
         10868 => x"00000000",
         10869 => x"00000000",
         10870 => x"000099c0",
         10871 => x"01040100",
         10872 => x"00000000",
         10873 => x"00000000",
         10874 => x"000099c8",
         10875 => x"01140300",
         10876 => x"00000000",
         10877 => x"00000000",
         10878 => x"000099d0",
         10879 => x"012b0300",
         10880 => x"00000000",
         10881 => x"00000000",
         10882 => x"000099d8",
         10883 => x"01300300",
         10884 => x"00000000",
         10885 => x"00000000",
         10886 => x"000099e0",
         10887 => x"013c0400",
         10888 => x"00000000",
         10889 => x"00000000",
         10890 => x"000099e8",
         10891 => x"013d0400",
         10892 => x"00000000",
         10893 => x"00000000",
         10894 => x"000099f0",
         10895 => x"013f0400",
         10896 => x"00000000",
         10897 => x"00000000",
         10898 => x"000099f8",
         10899 => x"01400400",
         10900 => x"00000000",
         10901 => x"00000000",
         10902 => x"00009a00",
         10903 => x"01410400",
         10904 => x"00000000",
         10905 => x"00000000",
         10906 => x"00009a04",
         10907 => x"01420400",
         10908 => x"00000000",
         10909 => x"00000000",
         10910 => x"00009a08",
         10911 => x"01430400",
         10912 => x"00000000",
         10913 => x"00000000",
         10914 => x"00009a0c",
         10915 => x"01500500",
         10916 => x"00000000",
         10917 => x"00000000",
         10918 => x"00009a10",
         10919 => x"01510500",
         10920 => x"00000000",
         10921 => x"00000000",
         10922 => x"00009a14",
         10923 => x"01540500",
         10924 => x"00000000",
         10925 => x"00000000",
         10926 => x"00009a18",
         10927 => x"01550500",
         10928 => x"00000000",
         10929 => x"00000000",
         10930 => x"00009a1c",
         10931 => x"01790700",
         10932 => x"00000000",
         10933 => x"00000000",
         10934 => x"00009a24",
         10935 => x"01780700",
         10936 => x"00000000",
         10937 => x"00000000",
         10938 => x"00009a28",
         10939 => x"01820800",
         10940 => x"00000000",
         10941 => x"00000000",
         10942 => x"00009a30",
         10943 => x"01830800",
         10944 => x"00000000",
         10945 => x"00000000",
         10946 => x"00009a38",
         10947 => x"01850800",
         10948 => x"00000000",
         10949 => x"00000000",
         10950 => x"00009a40",
         10951 => x"01870800",
         10952 => x"00000000",
         10953 => x"00000000",
         10954 => x"00009a48",
         10955 => x"018c0900",
         10956 => x"00000000",
         10957 => x"00000000",
         10958 => x"00009a50",
         10959 => x"018d0900",
         10960 => x"00000000",
         10961 => x"00000000",
         10962 => x"00009a58",
         10963 => x"018e0900",
         10964 => x"00000000",
         10965 => x"00000000",
         10966 => x"00009a60",
         10967 => x"018f0900",
         10968 => x"00000000",
         10969 => x"00000000",
         10970 => x"00000000",
         10971 => x"00000000",
         10972 => x"00007fff",
         10973 => x"00000000",
         10974 => x"00007fff",
         10975 => x"00010000",
         10976 => x"00007fff",
         10977 => x"00010000",
         10978 => x"00810000",
         10979 => x"01000000",
         10980 => x"017fffff",
         10981 => x"00000000",
         10982 => x"00000000",
         10983 => x"00007800",
         10984 => x"00000000",
         10985 => x"05f5e100",
         10986 => x"05f5e100",
         10987 => x"05f5e100",
         10988 => x"00000000",
         10989 => x"01010101",
         10990 => x"01010101",
         10991 => x"01011001",
         10992 => x"01000000",
         10993 => x"00000000",
         10994 => x"00000000",
         10995 => x"00000000",
         10996 => x"00000000",
         10997 => x"00000000",
         10998 => x"00000000",
         10999 => x"00000000",
         11000 => x"00000000",
         11001 => x"00000000",
         11002 => x"00000000",
         11003 => x"00000000",
         11004 => x"00000000",
         11005 => x"00000000",
         11006 => x"00000000",
         11007 => x"00000000",
         11008 => x"00000000",
         11009 => x"00000000",
         11010 => x"00000000",
         11011 => x"00000000",
         11012 => x"00000000",
         11013 => x"00000000",
         11014 => x"00000000",
         11015 => x"00000000",
         11016 => x"00000000",
         11017 => x"0000a470",
         11018 => x"01000000",
         11019 => x"0000a478",
         11020 => x"01000000",
         11021 => x"0000a480",
         11022 => x"02000000",
         11023 => x"00000000",
         11024 => x"00000000",
         11025 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

