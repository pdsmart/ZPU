-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBRAM;

architecture arch of SinglePortBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"84",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"84",
             9 => x"0b",
            10 => x"04",
            11 => x"84",
            12 => x"0b",
            13 => x"04",
            14 => x"84",
            15 => x"0b",
            16 => x"04",
            17 => x"84",
            18 => x"0b",
            19 => x"04",
            20 => x"84",
            21 => x"0b",
            22 => x"04",
            23 => x"85",
            24 => x"0b",
            25 => x"04",
            26 => x"85",
            27 => x"0b",
            28 => x"04",
            29 => x"85",
            30 => x"0b",
            31 => x"04",
            32 => x"86",
            33 => x"0b",
            34 => x"04",
            35 => x"86",
            36 => x"0b",
            37 => x"04",
            38 => x"86",
            39 => x"0b",
            40 => x"04",
            41 => x"86",
            42 => x"0b",
            43 => x"04",
            44 => x"87",
            45 => x"0b",
            46 => x"04",
            47 => x"87",
            48 => x"0b",
            49 => x"04",
            50 => x"87",
            51 => x"0b",
            52 => x"04",
            53 => x"87",
            54 => x"0b",
            55 => x"04",
            56 => x"88",
            57 => x"0b",
            58 => x"04",
            59 => x"88",
            60 => x"0b",
            61 => x"04",
            62 => x"88",
            63 => x"0b",
            64 => x"04",
            65 => x"88",
            66 => x"0b",
            67 => x"04",
            68 => x"89",
            69 => x"0b",
            70 => x"04",
            71 => x"89",
            72 => x"0b",
            73 => x"04",
            74 => x"89",
            75 => x"0b",
            76 => x"04",
            77 => x"8a",
            78 => x"0b",
            79 => x"04",
            80 => x"8a",
            81 => x"0b",
            82 => x"04",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"80",
           129 => x"94",
           130 => x"8f",
           131 => x"94",
           132 => x"80",
           133 => x"ca",
           134 => x"9f",
           135 => x"ca",
           136 => x"c0",
           137 => x"91",
           138 => x"90",
           139 => x"91",
           140 => x"88",
           141 => x"04",
           142 => x"0c",
           143 => x"2d",
           144 => x"08",
           145 => x"90",
           146 => x"94",
           147 => x"da",
           148 => x"94",
           149 => x"80",
           150 => x"ca",
           151 => x"a7",
           152 => x"ca",
           153 => x"c0",
           154 => x"91",
           155 => x"90",
           156 => x"91",
           157 => x"88",
           158 => x"04",
           159 => x"0c",
           160 => x"2d",
           161 => x"08",
           162 => x"90",
           163 => x"94",
           164 => x"e7",
           165 => x"94",
           166 => x"80",
           167 => x"ca",
           168 => x"a6",
           169 => x"ca",
           170 => x"c0",
           171 => x"91",
           172 => x"90",
           173 => x"91",
           174 => x"88",
           175 => x"04",
           176 => x"0c",
           177 => x"2d",
           178 => x"08",
           179 => x"90",
           180 => x"94",
           181 => x"9c",
           182 => x"94",
           183 => x"80",
           184 => x"ca",
           185 => x"97",
           186 => x"ca",
           187 => x"c0",
           188 => x"91",
           189 => x"90",
           190 => x"91",
           191 => x"88",
           192 => x"04",
           193 => x"0c",
           194 => x"2d",
           195 => x"08",
           196 => x"90",
           197 => x"94",
           198 => x"f1",
           199 => x"94",
           200 => x"80",
           201 => x"ca",
           202 => x"dc",
           203 => x"ca",
           204 => x"c0",
           205 => x"91",
           206 => x"90",
           207 => x"91",
           208 => x"88",
           209 => x"04",
           210 => x"0c",
           211 => x"2d",
           212 => x"08",
           213 => x"90",
           214 => x"94",
           215 => x"fe",
           216 => x"94",
           217 => x"80",
           218 => x"ca",
           219 => x"ee",
           220 => x"ca",
           221 => x"c0",
           222 => x"91",
           223 => x"90",
           224 => x"91",
           225 => x"88",
           226 => x"04",
           227 => x"0c",
           228 => x"2d",
           229 => x"08",
           230 => x"90",
           231 => x"94",
           232 => x"bb",
           233 => x"94",
           234 => x"80",
           235 => x"ca",
           236 => x"f2",
           237 => x"ca",
           238 => x"c0",
           239 => x"91",
           240 => x"90",
           241 => x"91",
           242 => x"88",
           243 => x"04",
           244 => x"0c",
           245 => x"2d",
           246 => x"08",
           247 => x"90",
           248 => x"94",
           249 => x"c9",
           250 => x"94",
           251 => x"80",
           252 => x"ca",
           253 => x"fd",
           254 => x"ca",
           255 => x"c0",
           256 => x"91",
           257 => x"90",
           258 => x"91",
           259 => x"88",
           260 => x"04",
           261 => x"0c",
           262 => x"2d",
           263 => x"08",
           264 => x"90",
           265 => x"94",
           266 => x"b8",
           267 => x"94",
           268 => x"80",
           269 => x"ca",
           270 => x"e9",
           271 => x"ca",
           272 => x"c0",
           273 => x"91",
           274 => x"90",
           275 => x"91",
           276 => x"88",
           277 => x"04",
           278 => x"0c",
           279 => x"2d",
           280 => x"08",
           281 => x"90",
           282 => x"94",
           283 => x"d4",
           284 => x"94",
           285 => x"80",
           286 => x"ca",
           287 => x"82",
           288 => x"ca",
           289 => x"c0",
           290 => x"91",
           291 => x"91",
           292 => x"91",
           293 => x"88",
           294 => x"04",
           295 => x"0c",
           296 => x"2d",
           297 => x"08",
           298 => x"90",
           299 => x"94",
           300 => x"bb",
           301 => x"94",
           302 => x"80",
           303 => x"ca",
           304 => x"8a",
           305 => x"ca",
           306 => x"c0",
           307 => x"91",
           308 => x"90",
           309 => x"91",
           310 => x"88",
           311 => x"04",
           312 => x"0c",
           313 => x"2d",
           314 => x"08",
           315 => x"90",
           316 => x"94",
           317 => x"c4",
           318 => x"94",
           319 => x"80",
           320 => x"ca",
           321 => x"90",
           322 => x"ca",
           323 => x"c0",
           324 => x"91",
           325 => x"90",
           326 => x"91",
           327 => x"88",
           328 => x"04",
           329 => x"0c",
           330 => x"2d",
           331 => x"08",
           332 => x"90",
           333 => x"94",
           334 => x"82",
           335 => x"94",
           336 => x"80",
           337 => x"ca",
           338 => x"e1",
           339 => x"38",
           340 => x"84",
           341 => x"0b",
           342 => x"c9",
           343 => x"80",
           344 => x"c5",
           345 => x"91",
           346 => x"02",
           347 => x"0c",
           348 => x"80",
           349 => x"94",
           350 => x"08",
           351 => x"94",
           352 => x"08",
           353 => x"3f",
           354 => x"08",
           355 => x"88",
           356 => x"3d",
           357 => x"94",
           358 => x"ca",
           359 => x"91",
           360 => x"fd",
           361 => x"53",
           362 => x"08",
           363 => x"52",
           364 => x"08",
           365 => x"51",
           366 => x"ca",
           367 => x"91",
           368 => x"54",
           369 => x"91",
           370 => x"04",
           371 => x"08",
           372 => x"94",
           373 => x"0d",
           374 => x"ca",
           375 => x"05",
           376 => x"91",
           377 => x"f8",
           378 => x"ca",
           379 => x"05",
           380 => x"94",
           381 => x"08",
           382 => x"91",
           383 => x"fc",
           384 => x"2e",
           385 => x"0b",
           386 => x"08",
           387 => x"24",
           388 => x"ca",
           389 => x"05",
           390 => x"ca",
           391 => x"05",
           392 => x"94",
           393 => x"08",
           394 => x"94",
           395 => x"0c",
           396 => x"91",
           397 => x"fc",
           398 => x"2e",
           399 => x"91",
           400 => x"8c",
           401 => x"ca",
           402 => x"05",
           403 => x"38",
           404 => x"08",
           405 => x"91",
           406 => x"8c",
           407 => x"91",
           408 => x"88",
           409 => x"ca",
           410 => x"05",
           411 => x"94",
           412 => x"08",
           413 => x"94",
           414 => x"0c",
           415 => x"08",
           416 => x"81",
           417 => x"94",
           418 => x"0c",
           419 => x"08",
           420 => x"81",
           421 => x"94",
           422 => x"0c",
           423 => x"91",
           424 => x"90",
           425 => x"2e",
           426 => x"ca",
           427 => x"05",
           428 => x"ca",
           429 => x"05",
           430 => x"39",
           431 => x"08",
           432 => x"70",
           433 => x"08",
           434 => x"51",
           435 => x"08",
           436 => x"91",
           437 => x"85",
           438 => x"ca",
           439 => x"fc",
           440 => x"79",
           441 => x"05",
           442 => x"57",
           443 => x"83",
           444 => x"38",
           445 => x"51",
           446 => x"a4",
           447 => x"52",
           448 => x"93",
           449 => x"70",
           450 => x"34",
           451 => x"71",
           452 => x"81",
           453 => x"74",
           454 => x"0c",
           455 => x"04",
           456 => x"2b",
           457 => x"71",
           458 => x"51",
           459 => x"72",
           460 => x"72",
           461 => x"05",
           462 => x"71",
           463 => x"53",
           464 => x"70",
           465 => x"0c",
           466 => x"84",
           467 => x"f0",
           468 => x"8f",
           469 => x"83",
           470 => x"38",
           471 => x"84",
           472 => x"fc",
           473 => x"83",
           474 => x"70",
           475 => x"39",
           476 => x"77",
           477 => x"07",
           478 => x"54",
           479 => x"38",
           480 => x"08",
           481 => x"71",
           482 => x"80",
           483 => x"75",
           484 => x"33",
           485 => x"06",
           486 => x"80",
           487 => x"72",
           488 => x"75",
           489 => x"06",
           490 => x"12",
           491 => x"33",
           492 => x"06",
           493 => x"52",
           494 => x"72",
           495 => x"81",
           496 => x"81",
           497 => x"71",
           498 => x"88",
           499 => x"87",
           500 => x"71",
           501 => x"fb",
           502 => x"06",
           503 => x"82",
           504 => x"51",
           505 => x"97",
           506 => x"84",
           507 => x"54",
           508 => x"75",
           509 => x"38",
           510 => x"52",
           511 => x"80",
           512 => x"88",
           513 => x"0d",
           514 => x"0d",
           515 => x"53",
           516 => x"52",
           517 => x"91",
           518 => x"81",
           519 => x"07",
           520 => x"52",
           521 => x"e8",
           522 => x"ca",
           523 => x"3d",
           524 => x"3d",
           525 => x"08",
           526 => x"56",
           527 => x"80",
           528 => x"33",
           529 => x"2e",
           530 => x"86",
           531 => x"52",
           532 => x"53",
           533 => x"13",
           534 => x"33",
           535 => x"06",
           536 => x"70",
           537 => x"38",
           538 => x"80",
           539 => x"74",
           540 => x"81",
           541 => x"70",
           542 => x"81",
           543 => x"80",
           544 => x"05",
           545 => x"76",
           546 => x"70",
           547 => x"0c",
           548 => x"04",
           549 => x"76",
           550 => x"80",
           551 => x"86",
           552 => x"52",
           553 => x"bf",
           554 => x"88",
           555 => x"80",
           556 => x"74",
           557 => x"ca",
           558 => x"3d",
           559 => x"3d",
           560 => x"11",
           561 => x"52",
           562 => x"70",
           563 => x"98",
           564 => x"33",
           565 => x"82",
           566 => x"26",
           567 => x"84",
           568 => x"83",
           569 => x"26",
           570 => x"85",
           571 => x"84",
           572 => x"26",
           573 => x"86",
           574 => x"85",
           575 => x"26",
           576 => x"88",
           577 => x"86",
           578 => x"e7",
           579 => x"38",
           580 => x"54",
           581 => x"87",
           582 => x"cc",
           583 => x"87",
           584 => x"0c",
           585 => x"c0",
           586 => x"82",
           587 => x"c0",
           588 => x"83",
           589 => x"c0",
           590 => x"84",
           591 => x"c0",
           592 => x"85",
           593 => x"c0",
           594 => x"86",
           595 => x"c0",
           596 => x"74",
           597 => x"a4",
           598 => x"c0",
           599 => x"80",
           600 => x"98",
           601 => x"52",
           602 => x"88",
           603 => x"0d",
           604 => x"0d",
           605 => x"c0",
           606 => x"81",
           607 => x"c0",
           608 => x"5e",
           609 => x"87",
           610 => x"08",
           611 => x"1c",
           612 => x"98",
           613 => x"79",
           614 => x"87",
           615 => x"08",
           616 => x"1c",
           617 => x"98",
           618 => x"79",
           619 => x"87",
           620 => x"08",
           621 => x"1c",
           622 => x"98",
           623 => x"7b",
           624 => x"87",
           625 => x"08",
           626 => x"1c",
           627 => x"0c",
           628 => x"ff",
           629 => x"83",
           630 => x"58",
           631 => x"57",
           632 => x"56",
           633 => x"55",
           634 => x"54",
           635 => x"53",
           636 => x"ff",
           637 => x"b3",
           638 => x"84",
           639 => x"0d",
           640 => x"0d",
           641 => x"33",
           642 => x"9f",
           643 => x"52",
           644 => x"91",
           645 => x"83",
           646 => x"fb",
           647 => x"0b",
           648 => x"e0",
           649 => x"ff",
           650 => x"56",
           651 => x"84",
           652 => x"2e",
           653 => x"c0",
           654 => x"70",
           655 => x"2a",
           656 => x"53",
           657 => x"80",
           658 => x"71",
           659 => x"81",
           660 => x"70",
           661 => x"81",
           662 => x"06",
           663 => x"80",
           664 => x"71",
           665 => x"81",
           666 => x"70",
           667 => x"73",
           668 => x"51",
           669 => x"80",
           670 => x"2e",
           671 => x"c0",
           672 => x"75",
           673 => x"91",
           674 => x"87",
           675 => x"fb",
           676 => x"9f",
           677 => x"0b",
           678 => x"33",
           679 => x"06",
           680 => x"87",
           681 => x"51",
           682 => x"86",
           683 => x"94",
           684 => x"08",
           685 => x"70",
           686 => x"54",
           687 => x"2e",
           688 => x"91",
           689 => x"06",
           690 => x"d7",
           691 => x"32",
           692 => x"51",
           693 => x"2e",
           694 => x"93",
           695 => x"06",
           696 => x"ff",
           697 => x"81",
           698 => x"87",
           699 => x"52",
           700 => x"86",
           701 => x"94",
           702 => x"72",
           703 => x"0d",
           704 => x"0d",
           705 => x"74",
           706 => x"ff",
           707 => x"57",
           708 => x"80",
           709 => x"81",
           710 => x"15",
           711 => x"c6",
           712 => x"81",
           713 => x"57",
           714 => x"c0",
           715 => x"75",
           716 => x"38",
           717 => x"94",
           718 => x"70",
           719 => x"81",
           720 => x"52",
           721 => x"8c",
           722 => x"2a",
           723 => x"51",
           724 => x"38",
           725 => x"70",
           726 => x"51",
           727 => x"8d",
           728 => x"2a",
           729 => x"51",
           730 => x"be",
           731 => x"ff",
           732 => x"c0",
           733 => x"70",
           734 => x"38",
           735 => x"90",
           736 => x"0c",
           737 => x"33",
           738 => x"06",
           739 => x"70",
           740 => x"76",
           741 => x"0c",
           742 => x"04",
           743 => x"0b",
           744 => x"e0",
           745 => x"ff",
           746 => x"87",
           747 => x"51",
           748 => x"86",
           749 => x"94",
           750 => x"08",
           751 => x"70",
           752 => x"51",
           753 => x"2e",
           754 => x"81",
           755 => x"87",
           756 => x"52",
           757 => x"86",
           758 => x"94",
           759 => x"08",
           760 => x"06",
           761 => x"0c",
           762 => x"0d",
           763 => x"0d",
           764 => x"c6",
           765 => x"81",
           766 => x"53",
           767 => x"84",
           768 => x"2e",
           769 => x"c0",
           770 => x"71",
           771 => x"2a",
           772 => x"51",
           773 => x"52",
           774 => x"a0",
           775 => x"ff",
           776 => x"c0",
           777 => x"70",
           778 => x"38",
           779 => x"90",
           780 => x"70",
           781 => x"98",
           782 => x"51",
           783 => x"88",
           784 => x"0d",
           785 => x"0d",
           786 => x"80",
           787 => x"2a",
           788 => x"51",
           789 => x"83",
           790 => x"c0",
           791 => x"91",
           792 => x"87",
           793 => x"08",
           794 => x"0c",
           795 => x"8c",
           796 => x"ec",
           797 => x"9e",
           798 => x"c6",
           799 => x"c0",
           800 => x"91",
           801 => x"87",
           802 => x"08",
           803 => x"0c",
           804 => x"a4",
           805 => x"fc",
           806 => x"9e",
           807 => x"c7",
           808 => x"c0",
           809 => x"91",
           810 => x"87",
           811 => x"08",
           812 => x"c7",
           813 => x"c0",
           814 => x"91",
           815 => x"81",
           816 => x"90",
           817 => x"87",
           818 => x"08",
           819 => x"06",
           820 => x"70",
           821 => x"38",
           822 => x"91",
           823 => x"80",
           824 => x"9e",
           825 => x"81",
           826 => x"51",
           827 => x"80",
           828 => x"81",
           829 => x"c7",
           830 => x"0b",
           831 => x"88",
           832 => x"c0",
           833 => x"52",
           834 => x"2e",
           835 => x"52",
           836 => x"93",
           837 => x"87",
           838 => x"08",
           839 => x"06",
           840 => x"70",
           841 => x"38",
           842 => x"91",
           843 => x"80",
           844 => x"9e",
           845 => x"88",
           846 => x"52",
           847 => x"2e",
           848 => x"52",
           849 => x"95",
           850 => x"87",
           851 => x"08",
           852 => x"06",
           853 => x"70",
           854 => x"38",
           855 => x"91",
           856 => x"80",
           857 => x"9e",
           858 => x"82",
           859 => x"52",
           860 => x"2e",
           861 => x"52",
           862 => x"97",
           863 => x"87",
           864 => x"08",
           865 => x"06",
           866 => x"70",
           867 => x"38",
           868 => x"91",
           869 => x"87",
           870 => x"08",
           871 => x"06",
           872 => x"51",
           873 => x"91",
           874 => x"80",
           875 => x"9e",
           876 => x"90",
           877 => x"52",
           878 => x"83",
           879 => x"71",
           880 => x"34",
           881 => x"c0",
           882 => x"70",
           883 => x"52",
           884 => x"2e",
           885 => x"52",
           886 => x"9b",
           887 => x"9e",
           888 => x"87",
           889 => x"70",
           890 => x"34",
           891 => x"04",
           892 => x"91",
           893 => x"84",
           894 => x"c7",
           895 => x"73",
           896 => x"38",
           897 => x"51",
           898 => x"91",
           899 => x"84",
           900 => x"c7",
           901 => x"73",
           902 => x"38",
           903 => x"08",
           904 => x"e4",
           905 => x"b4",
           906 => x"d4",
           907 => x"92",
           908 => x"80",
           909 => x"91",
           910 => x"53",
           911 => x"08",
           912 => x"ec",
           913 => x"3f",
           914 => x"33",
           915 => x"38",
           916 => x"33",
           917 => x"2e",
           918 => x"c6",
           919 => x"91",
           920 => x"52",
           921 => x"51",
           922 => x"91",
           923 => x"54",
           924 => x"88",
           925 => x"b4",
           926 => x"3f",
           927 => x"33",
           928 => x"2e",
           929 => x"b5",
           930 => x"90",
           931 => x"97",
           932 => x"80",
           933 => x"91",
           934 => x"82",
           935 => x"c7",
           936 => x"73",
           937 => x"38",
           938 => x"33",
           939 => x"d8",
           940 => x"3f",
           941 => x"33",
           942 => x"2e",
           943 => x"b5",
           944 => x"d8",
           945 => x"9b",
           946 => x"80",
           947 => x"91",
           948 => x"52",
           949 => x"51",
           950 => x"91",
           951 => x"82",
           952 => x"c6",
           953 => x"91",
           954 => x"88",
           955 => x"c7",
           956 => x"91",
           957 => x"88",
           958 => x"c7",
           959 => x"91",
           960 => x"87",
           961 => x"c7",
           962 => x"91",
           963 => x"87",
           964 => x"c7",
           965 => x"91",
           966 => x"87",
           967 => x"3d",
           968 => x"3d",
           969 => x"05",
           970 => x"52",
           971 => x"ac",
           972 => x"29",
           973 => x"b3",
           974 => x"71",
           975 => x"b8",
           976 => x"39",
           977 => x"51",
           978 => x"b8",
           979 => x"39",
           980 => x"51",
           981 => x"b8",
           982 => x"39",
           983 => x"51",
           984 => x"84",
           985 => x"71",
           986 => x"04",
           987 => x"c0",
           988 => x"04",
           989 => x"87",
           990 => x"70",
           991 => x"80",
           992 => x"74",
           993 => x"c7",
           994 => x"0c",
           995 => x"04",
           996 => x"87",
           997 => x"70",
           998 => x"a0",
           999 => x"72",
          1000 => x"70",
          1001 => x"08",
          1002 => x"c7",
          1003 => x"0c",
          1004 => x"0d",
          1005 => x"a0",
          1006 => x"96",
          1007 => x"fe",
          1008 => x"93",
          1009 => x"72",
          1010 => x"81",
          1011 => x"8d",
          1012 => x"91",
          1013 => x"52",
          1014 => x"90",
          1015 => x"34",
          1016 => x"08",
          1017 => x"ca",
          1018 => x"39",
          1019 => x"08",
          1020 => x"2e",
          1021 => x"51",
          1022 => x"3d",
          1023 => x"3d",
          1024 => x"05",
          1025 => x"98",
          1026 => x"ca",
          1027 => x"51",
          1028 => x"72",
          1029 => x"0c",
          1030 => x"04",
          1031 => x"75",
          1032 => x"70",
          1033 => x"53",
          1034 => x"2e",
          1035 => x"81",
          1036 => x"81",
          1037 => x"87",
          1038 => x"85",
          1039 => x"fc",
          1040 => x"91",
          1041 => x"78",
          1042 => x"0c",
          1043 => x"33",
          1044 => x"06",
          1045 => x"80",
          1046 => x"72",
          1047 => x"51",
          1048 => x"fe",
          1049 => x"39",
          1050 => x"98",
          1051 => x"0d",
          1052 => x"0d",
          1053 => x"59",
          1054 => x"05",
          1055 => x"75",
          1056 => x"f8",
          1057 => x"2e",
          1058 => x"82",
          1059 => x"70",
          1060 => x"05",
          1061 => x"5b",
          1062 => x"2e",
          1063 => x"85",
          1064 => x"8b",
          1065 => x"2e",
          1066 => x"8a",
          1067 => x"78",
          1068 => x"5a",
          1069 => x"aa",
          1070 => x"06",
          1071 => x"84",
          1072 => x"7b",
          1073 => x"5d",
          1074 => x"59",
          1075 => x"d0",
          1076 => x"89",
          1077 => x"7a",
          1078 => x"10",
          1079 => x"d0",
          1080 => x"81",
          1081 => x"57",
          1082 => x"75",
          1083 => x"70",
          1084 => x"07",
          1085 => x"80",
          1086 => x"30",
          1087 => x"80",
          1088 => x"53",
          1089 => x"55",
          1090 => x"2e",
          1091 => x"84",
          1092 => x"81",
          1093 => x"57",
          1094 => x"2e",
          1095 => x"75",
          1096 => x"76",
          1097 => x"e0",
          1098 => x"ff",
          1099 => x"73",
          1100 => x"81",
          1101 => x"80",
          1102 => x"38",
          1103 => x"2e",
          1104 => x"73",
          1105 => x"8b",
          1106 => x"c2",
          1107 => x"38",
          1108 => x"73",
          1109 => x"81",
          1110 => x"8f",
          1111 => x"d5",
          1112 => x"38",
          1113 => x"24",
          1114 => x"80",
          1115 => x"38",
          1116 => x"73",
          1117 => x"80",
          1118 => x"ef",
          1119 => x"19",
          1120 => x"59",
          1121 => x"33",
          1122 => x"75",
          1123 => x"81",
          1124 => x"70",
          1125 => x"55",
          1126 => x"79",
          1127 => x"90",
          1128 => x"16",
          1129 => x"7b",
          1130 => x"a0",
          1131 => x"3f",
          1132 => x"53",
          1133 => x"e9",
          1134 => x"fc",
          1135 => x"81",
          1136 => x"72",
          1137 => x"b0",
          1138 => x"fb",
          1139 => x"39",
          1140 => x"83",
          1141 => x"59",
          1142 => x"82",
          1143 => x"88",
          1144 => x"8a",
          1145 => x"90",
          1146 => x"75",
          1147 => x"3f",
          1148 => x"79",
          1149 => x"81",
          1150 => x"72",
          1151 => x"38",
          1152 => x"59",
          1153 => x"84",
          1154 => x"58",
          1155 => x"80",
          1156 => x"30",
          1157 => x"80",
          1158 => x"55",
          1159 => x"25",
          1160 => x"80",
          1161 => x"74",
          1162 => x"07",
          1163 => x"0b",
          1164 => x"57",
          1165 => x"51",
          1166 => x"91",
          1167 => x"81",
          1168 => x"53",
          1169 => x"e6",
          1170 => x"ca",
          1171 => x"89",
          1172 => x"38",
          1173 => x"75",
          1174 => x"84",
          1175 => x"53",
          1176 => x"06",
          1177 => x"53",
          1178 => x"81",
          1179 => x"81",
          1180 => x"70",
          1181 => x"2a",
          1182 => x"76",
          1183 => x"38",
          1184 => x"38",
          1185 => x"70",
          1186 => x"53",
          1187 => x"8e",
          1188 => x"77",
          1189 => x"53",
          1190 => x"81",
          1191 => x"7a",
          1192 => x"55",
          1193 => x"83",
          1194 => x"79",
          1195 => x"81",
          1196 => x"72",
          1197 => x"17",
          1198 => x"27",
          1199 => x"51",
          1200 => x"75",
          1201 => x"72",
          1202 => x"81",
          1203 => x"7a",
          1204 => x"38",
          1205 => x"05",
          1206 => x"ff",
          1207 => x"70",
          1208 => x"57",
          1209 => x"76",
          1210 => x"81",
          1211 => x"72",
          1212 => x"84",
          1213 => x"f9",
          1214 => x"39",
          1215 => x"04",
          1216 => x"86",
          1217 => x"84",
          1218 => x"55",
          1219 => x"fa",
          1220 => x"3d",
          1221 => x"3d",
          1222 => x"ca",
          1223 => x"3d",
          1224 => x"75",
          1225 => x"3f",
          1226 => x"08",
          1227 => x"34",
          1228 => x"ca",
          1229 => x"3d",
          1230 => x"3d",
          1231 => x"98",
          1232 => x"ca",
          1233 => x"3d",
          1234 => x"77",
          1235 => x"a1",
          1236 => x"ca",
          1237 => x"3d",
          1238 => x"3d",
          1239 => x"91",
          1240 => x"70",
          1241 => x"55",
          1242 => x"80",
          1243 => x"38",
          1244 => x"08",
          1245 => x"91",
          1246 => x"81",
          1247 => x"72",
          1248 => x"cb",
          1249 => x"2e",
          1250 => x"88",
          1251 => x"70",
          1252 => x"51",
          1253 => x"2e",
          1254 => x"80",
          1255 => x"ff",
          1256 => x"39",
          1257 => x"c8",
          1258 => x"52",
          1259 => x"c0",
          1260 => x"52",
          1261 => x"81",
          1262 => x"51",
          1263 => x"ff",
          1264 => x"15",
          1265 => x"34",
          1266 => x"f3",
          1267 => x"72",
          1268 => x"0c",
          1269 => x"04",
          1270 => x"91",
          1271 => x"75",
          1272 => x"0c",
          1273 => x"52",
          1274 => x"3f",
          1275 => x"9c",
          1276 => x"0d",
          1277 => x"0d",
          1278 => x"56",
          1279 => x"0c",
          1280 => x"70",
          1281 => x"73",
          1282 => x"81",
          1283 => x"81",
          1284 => x"ed",
          1285 => x"2e",
          1286 => x"8e",
          1287 => x"08",
          1288 => x"76",
          1289 => x"56",
          1290 => x"b0",
          1291 => x"06",
          1292 => x"75",
          1293 => x"76",
          1294 => x"70",
          1295 => x"73",
          1296 => x"8b",
          1297 => x"73",
          1298 => x"85",
          1299 => x"82",
          1300 => x"76",
          1301 => x"70",
          1302 => x"ac",
          1303 => x"a0",
          1304 => x"fa",
          1305 => x"53",
          1306 => x"57",
          1307 => x"98",
          1308 => x"39",
          1309 => x"80",
          1310 => x"26",
          1311 => x"86",
          1312 => x"80",
          1313 => x"57",
          1314 => x"74",
          1315 => x"38",
          1316 => x"27",
          1317 => x"14",
          1318 => x"06",
          1319 => x"14",
          1320 => x"06",
          1321 => x"74",
          1322 => x"f9",
          1323 => x"ff",
          1324 => x"89",
          1325 => x"38",
          1326 => x"c5",
          1327 => x"29",
          1328 => x"81",
          1329 => x"76",
          1330 => x"56",
          1331 => x"ba",
          1332 => x"2e",
          1333 => x"30",
          1334 => x"0c",
          1335 => x"91",
          1336 => x"8a",
          1337 => x"f8",
          1338 => x"7c",
          1339 => x"70",
          1340 => x"75",
          1341 => x"55",
          1342 => x"2e",
          1343 => x"87",
          1344 => x"76",
          1345 => x"73",
          1346 => x"81",
          1347 => x"81",
          1348 => x"77",
          1349 => x"70",
          1350 => x"58",
          1351 => x"09",
          1352 => x"c2",
          1353 => x"81",
          1354 => x"75",
          1355 => x"55",
          1356 => x"e2",
          1357 => x"90",
          1358 => x"f8",
          1359 => x"8f",
          1360 => x"81",
          1361 => x"75",
          1362 => x"55",
          1363 => x"81",
          1364 => x"27",
          1365 => x"d0",
          1366 => x"55",
          1367 => x"73",
          1368 => x"80",
          1369 => x"14",
          1370 => x"72",
          1371 => x"e0",
          1372 => x"80",
          1373 => x"39",
          1374 => x"55",
          1375 => x"80",
          1376 => x"e0",
          1377 => x"38",
          1378 => x"81",
          1379 => x"53",
          1380 => x"81",
          1381 => x"53",
          1382 => x"8e",
          1383 => x"70",
          1384 => x"55",
          1385 => x"27",
          1386 => x"77",
          1387 => x"74",
          1388 => x"76",
          1389 => x"77",
          1390 => x"70",
          1391 => x"55",
          1392 => x"77",
          1393 => x"38",
          1394 => x"74",
          1395 => x"55",
          1396 => x"88",
          1397 => x"0d",
          1398 => x"0d",
          1399 => x"33",
          1400 => x"70",
          1401 => x"38",
          1402 => x"11",
          1403 => x"91",
          1404 => x"83",
          1405 => x"fc",
          1406 => x"9b",
          1407 => x"84",
          1408 => x"33",
          1409 => x"51",
          1410 => x"80",
          1411 => x"84",
          1412 => x"92",
          1413 => x"51",
          1414 => x"80",
          1415 => x"81",
          1416 => x"72",
          1417 => x"92",
          1418 => x"81",
          1419 => x"0b",
          1420 => x"8c",
          1421 => x"71",
          1422 => x"06",
          1423 => x"80",
          1424 => x"87",
          1425 => x"08",
          1426 => x"38",
          1427 => x"80",
          1428 => x"71",
          1429 => x"c0",
          1430 => x"51",
          1431 => x"87",
          1432 => x"c7",
          1433 => x"91",
          1434 => x"33",
          1435 => x"ca",
          1436 => x"3d",
          1437 => x"3d",
          1438 => x"64",
          1439 => x"bf",
          1440 => x"40",
          1441 => x"74",
          1442 => x"cd",
          1443 => x"88",
          1444 => x"7a",
          1445 => x"81",
          1446 => x"72",
          1447 => x"87",
          1448 => x"11",
          1449 => x"8c",
          1450 => x"92",
          1451 => x"5a",
          1452 => x"58",
          1453 => x"c0",
          1454 => x"76",
          1455 => x"76",
          1456 => x"70",
          1457 => x"81",
          1458 => x"54",
          1459 => x"8e",
          1460 => x"52",
          1461 => x"81",
          1462 => x"81",
          1463 => x"74",
          1464 => x"53",
          1465 => x"83",
          1466 => x"78",
          1467 => x"8f",
          1468 => x"2e",
          1469 => x"c0",
          1470 => x"52",
          1471 => x"87",
          1472 => x"08",
          1473 => x"2e",
          1474 => x"84",
          1475 => x"38",
          1476 => x"87",
          1477 => x"15",
          1478 => x"70",
          1479 => x"52",
          1480 => x"ff",
          1481 => x"39",
          1482 => x"81",
          1483 => x"ff",
          1484 => x"57",
          1485 => x"90",
          1486 => x"80",
          1487 => x"71",
          1488 => x"78",
          1489 => x"38",
          1490 => x"80",
          1491 => x"80",
          1492 => x"81",
          1493 => x"72",
          1494 => x"0c",
          1495 => x"04",
          1496 => x"60",
          1497 => x"8c",
          1498 => x"33",
          1499 => x"5b",
          1500 => x"74",
          1501 => x"e1",
          1502 => x"88",
          1503 => x"79",
          1504 => x"78",
          1505 => x"06",
          1506 => x"77",
          1507 => x"87",
          1508 => x"11",
          1509 => x"8c",
          1510 => x"92",
          1511 => x"59",
          1512 => x"85",
          1513 => x"98",
          1514 => x"7d",
          1515 => x"0c",
          1516 => x"08",
          1517 => x"70",
          1518 => x"53",
          1519 => x"2e",
          1520 => x"70",
          1521 => x"33",
          1522 => x"18",
          1523 => x"2a",
          1524 => x"51",
          1525 => x"2e",
          1526 => x"c0",
          1527 => x"52",
          1528 => x"87",
          1529 => x"08",
          1530 => x"2e",
          1531 => x"84",
          1532 => x"38",
          1533 => x"87",
          1534 => x"15",
          1535 => x"70",
          1536 => x"52",
          1537 => x"ff",
          1538 => x"39",
          1539 => x"81",
          1540 => x"80",
          1541 => x"52",
          1542 => x"90",
          1543 => x"80",
          1544 => x"71",
          1545 => x"7a",
          1546 => x"38",
          1547 => x"80",
          1548 => x"80",
          1549 => x"81",
          1550 => x"72",
          1551 => x"0c",
          1552 => x"04",
          1553 => x"7e",
          1554 => x"b3",
          1555 => x"88",
          1556 => x"33",
          1557 => x"56",
          1558 => x"3f",
          1559 => x"08",
          1560 => x"83",
          1561 => x"fe",
          1562 => x"87",
          1563 => x"0c",
          1564 => x"76",
          1565 => x"38",
          1566 => x"93",
          1567 => x"2b",
          1568 => x"8c",
          1569 => x"71",
          1570 => x"38",
          1571 => x"71",
          1572 => x"c6",
          1573 => x"39",
          1574 => x"81",
          1575 => x"06",
          1576 => x"71",
          1577 => x"38",
          1578 => x"8c",
          1579 => x"e8",
          1580 => x"98",
          1581 => x"71",
          1582 => x"73",
          1583 => x"92",
          1584 => x"72",
          1585 => x"06",
          1586 => x"f7",
          1587 => x"80",
          1588 => x"88",
          1589 => x"0c",
          1590 => x"80",
          1591 => x"56",
          1592 => x"56",
          1593 => x"91",
          1594 => x"8c",
          1595 => x"fe",
          1596 => x"81",
          1597 => x"33",
          1598 => x"07",
          1599 => x"0c",
          1600 => x"3d",
          1601 => x"3d",
          1602 => x"11",
          1603 => x"33",
          1604 => x"71",
          1605 => x"81",
          1606 => x"72",
          1607 => x"75",
          1608 => x"91",
          1609 => x"52",
          1610 => x"54",
          1611 => x"0d",
          1612 => x"0d",
          1613 => x"05",
          1614 => x"52",
          1615 => x"70",
          1616 => x"34",
          1617 => x"51",
          1618 => x"83",
          1619 => x"ff",
          1620 => x"75",
          1621 => x"72",
          1622 => x"54",
          1623 => x"2a",
          1624 => x"70",
          1625 => x"34",
          1626 => x"51",
          1627 => x"81",
          1628 => x"70",
          1629 => x"70",
          1630 => x"3d",
          1631 => x"3d",
          1632 => x"77",
          1633 => x"70",
          1634 => x"38",
          1635 => x"05",
          1636 => x"70",
          1637 => x"34",
          1638 => x"eb",
          1639 => x"0d",
          1640 => x"0d",
          1641 => x"54",
          1642 => x"72",
          1643 => x"54",
          1644 => x"51",
          1645 => x"84",
          1646 => x"fc",
          1647 => x"77",
          1648 => x"53",
          1649 => x"05",
          1650 => x"70",
          1651 => x"33",
          1652 => x"ff",
          1653 => x"52",
          1654 => x"2e",
          1655 => x"80",
          1656 => x"71",
          1657 => x"0c",
          1658 => x"04",
          1659 => x"74",
          1660 => x"89",
          1661 => x"2e",
          1662 => x"11",
          1663 => x"52",
          1664 => x"70",
          1665 => x"88",
          1666 => x"0d",
          1667 => x"91",
          1668 => x"04",
          1669 => x"ca",
          1670 => x"f7",
          1671 => x"56",
          1672 => x"17",
          1673 => x"74",
          1674 => x"d6",
          1675 => x"b0",
          1676 => x"b4",
          1677 => x"81",
          1678 => x"59",
          1679 => x"91",
          1680 => x"7a",
          1681 => x"06",
          1682 => x"ca",
          1683 => x"17",
          1684 => x"08",
          1685 => x"08",
          1686 => x"08",
          1687 => x"74",
          1688 => x"38",
          1689 => x"55",
          1690 => x"09",
          1691 => x"38",
          1692 => x"18",
          1693 => x"81",
          1694 => x"f9",
          1695 => x"39",
          1696 => x"91",
          1697 => x"8b",
          1698 => x"fa",
          1699 => x"7a",
          1700 => x"57",
          1701 => x"08",
          1702 => x"75",
          1703 => x"3f",
          1704 => x"08",
          1705 => x"88",
          1706 => x"81",
          1707 => x"b4",
          1708 => x"16",
          1709 => x"be",
          1710 => x"88",
          1711 => x"85",
          1712 => x"81",
          1713 => x"17",
          1714 => x"ca",
          1715 => x"3d",
          1716 => x"3d",
          1717 => x"52",
          1718 => x"3f",
          1719 => x"08",
          1720 => x"88",
          1721 => x"38",
          1722 => x"74",
          1723 => x"81",
          1724 => x"38",
          1725 => x"59",
          1726 => x"09",
          1727 => x"e3",
          1728 => x"53",
          1729 => x"08",
          1730 => x"70",
          1731 => x"91",
          1732 => x"d5",
          1733 => x"17",
          1734 => x"3f",
          1735 => x"a4",
          1736 => x"51",
          1737 => x"86",
          1738 => x"f2",
          1739 => x"17",
          1740 => x"3f",
          1741 => x"52",
          1742 => x"51",
          1743 => x"8c",
          1744 => x"84",
          1745 => x"fc",
          1746 => x"17",
          1747 => x"70",
          1748 => x"79",
          1749 => x"52",
          1750 => x"51",
          1751 => x"77",
          1752 => x"80",
          1753 => x"81",
          1754 => x"f9",
          1755 => x"ca",
          1756 => x"2e",
          1757 => x"58",
          1758 => x"88",
          1759 => x"0d",
          1760 => x"0d",
          1761 => x"98",
          1762 => x"05",
          1763 => x"80",
          1764 => x"27",
          1765 => x"14",
          1766 => x"29",
          1767 => x"05",
          1768 => x"91",
          1769 => x"87",
          1770 => x"f9",
          1771 => x"7a",
          1772 => x"54",
          1773 => x"27",
          1774 => x"76",
          1775 => x"27",
          1776 => x"ff",
          1777 => x"58",
          1778 => x"80",
          1779 => x"82",
          1780 => x"72",
          1781 => x"38",
          1782 => x"72",
          1783 => x"8e",
          1784 => x"39",
          1785 => x"17",
          1786 => x"a4",
          1787 => x"53",
          1788 => x"fd",
          1789 => x"ca",
          1790 => x"9f",
          1791 => x"ff",
          1792 => x"11",
          1793 => x"70",
          1794 => x"18",
          1795 => x"76",
          1796 => x"53",
          1797 => x"91",
          1798 => x"80",
          1799 => x"83",
          1800 => x"b4",
          1801 => x"88",
          1802 => x"79",
          1803 => x"84",
          1804 => x"58",
          1805 => x"80",
          1806 => x"9f",
          1807 => x"80",
          1808 => x"88",
          1809 => x"08",
          1810 => x"51",
          1811 => x"91",
          1812 => x"80",
          1813 => x"10",
          1814 => x"74",
          1815 => x"51",
          1816 => x"91",
          1817 => x"83",
          1818 => x"58",
          1819 => x"87",
          1820 => x"08",
          1821 => x"51",
          1822 => x"91",
          1823 => x"9b",
          1824 => x"2b",
          1825 => x"74",
          1826 => x"51",
          1827 => x"91",
          1828 => x"f0",
          1829 => x"83",
          1830 => x"77",
          1831 => x"0c",
          1832 => x"04",
          1833 => x"7a",
          1834 => x"58",
          1835 => x"81",
          1836 => x"9e",
          1837 => x"17",
          1838 => x"96",
          1839 => x"53",
          1840 => x"81",
          1841 => x"79",
          1842 => x"72",
          1843 => x"38",
          1844 => x"72",
          1845 => x"b8",
          1846 => x"39",
          1847 => x"17",
          1848 => x"a4",
          1849 => x"53",
          1850 => x"fb",
          1851 => x"ca",
          1852 => x"91",
          1853 => x"81",
          1854 => x"83",
          1855 => x"b4",
          1856 => x"78",
          1857 => x"56",
          1858 => x"76",
          1859 => x"38",
          1860 => x"9f",
          1861 => x"33",
          1862 => x"07",
          1863 => x"74",
          1864 => x"83",
          1865 => x"89",
          1866 => x"08",
          1867 => x"51",
          1868 => x"91",
          1869 => x"59",
          1870 => x"08",
          1871 => x"74",
          1872 => x"16",
          1873 => x"84",
          1874 => x"76",
          1875 => x"88",
          1876 => x"81",
          1877 => x"8f",
          1878 => x"53",
          1879 => x"80",
          1880 => x"88",
          1881 => x"08",
          1882 => x"51",
          1883 => x"91",
          1884 => x"59",
          1885 => x"08",
          1886 => x"77",
          1887 => x"06",
          1888 => x"83",
          1889 => x"05",
          1890 => x"f7",
          1891 => x"39",
          1892 => x"a4",
          1893 => x"52",
          1894 => x"ef",
          1895 => x"88",
          1896 => x"ca",
          1897 => x"38",
          1898 => x"06",
          1899 => x"83",
          1900 => x"18",
          1901 => x"54",
          1902 => x"f6",
          1903 => x"ca",
          1904 => x"0a",
          1905 => x"52",
          1906 => x"83",
          1907 => x"83",
          1908 => x"91",
          1909 => x"8a",
          1910 => x"f8",
          1911 => x"7c",
          1912 => x"59",
          1913 => x"81",
          1914 => x"38",
          1915 => x"08",
          1916 => x"73",
          1917 => x"38",
          1918 => x"52",
          1919 => x"a4",
          1920 => x"88",
          1921 => x"ca",
          1922 => x"f2",
          1923 => x"82",
          1924 => x"39",
          1925 => x"e6",
          1926 => x"88",
          1927 => x"de",
          1928 => x"78",
          1929 => x"3f",
          1930 => x"08",
          1931 => x"88",
          1932 => x"80",
          1933 => x"ca",
          1934 => x"2e",
          1935 => x"ca",
          1936 => x"2e",
          1937 => x"53",
          1938 => x"51",
          1939 => x"91",
          1940 => x"c5",
          1941 => x"08",
          1942 => x"18",
          1943 => x"57",
          1944 => x"90",
          1945 => x"90",
          1946 => x"16",
          1947 => x"54",
          1948 => x"34",
          1949 => x"78",
          1950 => x"38",
          1951 => x"91",
          1952 => x"8a",
          1953 => x"f6",
          1954 => x"7e",
          1955 => x"5b",
          1956 => x"38",
          1957 => x"58",
          1958 => x"88",
          1959 => x"08",
          1960 => x"38",
          1961 => x"39",
          1962 => x"51",
          1963 => x"81",
          1964 => x"ca",
          1965 => x"82",
          1966 => x"ca",
          1967 => x"91",
          1968 => x"ff",
          1969 => x"38",
          1970 => x"91",
          1971 => x"26",
          1972 => x"79",
          1973 => x"08",
          1974 => x"73",
          1975 => x"b9",
          1976 => x"2e",
          1977 => x"80",
          1978 => x"1a",
          1979 => x"08",
          1980 => x"38",
          1981 => x"52",
          1982 => x"af",
          1983 => x"91",
          1984 => x"81",
          1985 => x"06",
          1986 => x"ca",
          1987 => x"91",
          1988 => x"09",
          1989 => x"72",
          1990 => x"70",
          1991 => x"ca",
          1992 => x"51",
          1993 => x"73",
          1994 => x"91",
          1995 => x"80",
          1996 => x"8c",
          1997 => x"81",
          1998 => x"38",
          1999 => x"08",
          2000 => x"73",
          2001 => x"75",
          2002 => x"77",
          2003 => x"56",
          2004 => x"76",
          2005 => x"82",
          2006 => x"26",
          2007 => x"75",
          2008 => x"f8",
          2009 => x"ca",
          2010 => x"2e",
          2011 => x"59",
          2012 => x"08",
          2013 => x"81",
          2014 => x"91",
          2015 => x"59",
          2016 => x"08",
          2017 => x"70",
          2018 => x"25",
          2019 => x"51",
          2020 => x"73",
          2021 => x"75",
          2022 => x"81",
          2023 => x"38",
          2024 => x"f5",
          2025 => x"75",
          2026 => x"f9",
          2027 => x"ca",
          2028 => x"ca",
          2029 => x"70",
          2030 => x"08",
          2031 => x"51",
          2032 => x"80",
          2033 => x"73",
          2034 => x"38",
          2035 => x"52",
          2036 => x"d0",
          2037 => x"88",
          2038 => x"a5",
          2039 => x"18",
          2040 => x"08",
          2041 => x"18",
          2042 => x"74",
          2043 => x"38",
          2044 => x"18",
          2045 => x"33",
          2046 => x"73",
          2047 => x"97",
          2048 => x"74",
          2049 => x"38",
          2050 => x"55",
          2051 => x"ca",
          2052 => x"85",
          2053 => x"75",
          2054 => x"ca",
          2055 => x"3d",
          2056 => x"3d",
          2057 => x"52",
          2058 => x"3f",
          2059 => x"08",
          2060 => x"91",
          2061 => x"80",
          2062 => x"52",
          2063 => x"c1",
          2064 => x"88",
          2065 => x"88",
          2066 => x"0c",
          2067 => x"53",
          2068 => x"15",
          2069 => x"f2",
          2070 => x"56",
          2071 => x"16",
          2072 => x"22",
          2073 => x"27",
          2074 => x"54",
          2075 => x"76",
          2076 => x"33",
          2077 => x"3f",
          2078 => x"08",
          2079 => x"38",
          2080 => x"76",
          2081 => x"70",
          2082 => x"9f",
          2083 => x"56",
          2084 => x"ca",
          2085 => x"3d",
          2086 => x"3d",
          2087 => x"71",
          2088 => x"57",
          2089 => x"0a",
          2090 => x"38",
          2091 => x"53",
          2092 => x"38",
          2093 => x"0c",
          2094 => x"54",
          2095 => x"75",
          2096 => x"73",
          2097 => x"a8",
          2098 => x"73",
          2099 => x"85",
          2100 => x"0b",
          2101 => x"5a",
          2102 => x"27",
          2103 => x"a8",
          2104 => x"18",
          2105 => x"39",
          2106 => x"70",
          2107 => x"58",
          2108 => x"b2",
          2109 => x"76",
          2110 => x"3f",
          2111 => x"08",
          2112 => x"88",
          2113 => x"bd",
          2114 => x"91",
          2115 => x"27",
          2116 => x"16",
          2117 => x"88",
          2118 => x"38",
          2119 => x"39",
          2120 => x"55",
          2121 => x"52",
          2122 => x"d5",
          2123 => x"88",
          2124 => x"0c",
          2125 => x"0c",
          2126 => x"53",
          2127 => x"80",
          2128 => x"85",
          2129 => x"94",
          2130 => x"2a",
          2131 => x"0c",
          2132 => x"06",
          2133 => x"9c",
          2134 => x"58",
          2135 => x"88",
          2136 => x"0d",
          2137 => x"0d",
          2138 => x"90",
          2139 => x"05",
          2140 => x"f0",
          2141 => x"27",
          2142 => x"0b",
          2143 => x"98",
          2144 => x"84",
          2145 => x"2e",
          2146 => x"76",
          2147 => x"58",
          2148 => x"38",
          2149 => x"15",
          2150 => x"08",
          2151 => x"38",
          2152 => x"88",
          2153 => x"53",
          2154 => x"81",
          2155 => x"c0",
          2156 => x"22",
          2157 => x"89",
          2158 => x"72",
          2159 => x"74",
          2160 => x"f3",
          2161 => x"ca",
          2162 => x"82",
          2163 => x"91",
          2164 => x"27",
          2165 => x"81",
          2166 => x"88",
          2167 => x"80",
          2168 => x"16",
          2169 => x"88",
          2170 => x"ca",
          2171 => x"38",
          2172 => x"0c",
          2173 => x"dd",
          2174 => x"08",
          2175 => x"f9",
          2176 => x"ca",
          2177 => x"87",
          2178 => x"88",
          2179 => x"80",
          2180 => x"55",
          2181 => x"08",
          2182 => x"38",
          2183 => x"ca",
          2184 => x"2e",
          2185 => x"ca",
          2186 => x"75",
          2187 => x"3f",
          2188 => x"08",
          2189 => x"94",
          2190 => x"52",
          2191 => x"c1",
          2192 => x"88",
          2193 => x"0c",
          2194 => x"0c",
          2195 => x"05",
          2196 => x"80",
          2197 => x"ca",
          2198 => x"3d",
          2199 => x"3d",
          2200 => x"71",
          2201 => x"57",
          2202 => x"51",
          2203 => x"91",
          2204 => x"54",
          2205 => x"08",
          2206 => x"91",
          2207 => x"56",
          2208 => x"52",
          2209 => x"83",
          2210 => x"88",
          2211 => x"ca",
          2212 => x"d2",
          2213 => x"88",
          2214 => x"08",
          2215 => x"54",
          2216 => x"e5",
          2217 => x"06",
          2218 => x"58",
          2219 => x"08",
          2220 => x"38",
          2221 => x"75",
          2222 => x"80",
          2223 => x"81",
          2224 => x"7a",
          2225 => x"06",
          2226 => x"39",
          2227 => x"08",
          2228 => x"76",
          2229 => x"3f",
          2230 => x"08",
          2231 => x"88",
          2232 => x"ff",
          2233 => x"84",
          2234 => x"06",
          2235 => x"54",
          2236 => x"88",
          2237 => x"0d",
          2238 => x"0d",
          2239 => x"52",
          2240 => x"3f",
          2241 => x"08",
          2242 => x"06",
          2243 => x"51",
          2244 => x"83",
          2245 => x"06",
          2246 => x"14",
          2247 => x"3f",
          2248 => x"08",
          2249 => x"07",
          2250 => x"ca",
          2251 => x"3d",
          2252 => x"3d",
          2253 => x"70",
          2254 => x"06",
          2255 => x"53",
          2256 => x"ed",
          2257 => x"33",
          2258 => x"83",
          2259 => x"06",
          2260 => x"90",
          2261 => x"15",
          2262 => x"3f",
          2263 => x"04",
          2264 => x"7b",
          2265 => x"84",
          2266 => x"58",
          2267 => x"80",
          2268 => x"38",
          2269 => x"52",
          2270 => x"8f",
          2271 => x"88",
          2272 => x"ca",
          2273 => x"f5",
          2274 => x"08",
          2275 => x"53",
          2276 => x"84",
          2277 => x"39",
          2278 => x"70",
          2279 => x"81",
          2280 => x"51",
          2281 => x"16",
          2282 => x"88",
          2283 => x"81",
          2284 => x"38",
          2285 => x"ae",
          2286 => x"81",
          2287 => x"54",
          2288 => x"2e",
          2289 => x"8f",
          2290 => x"91",
          2291 => x"76",
          2292 => x"54",
          2293 => x"09",
          2294 => x"38",
          2295 => x"7a",
          2296 => x"80",
          2297 => x"fa",
          2298 => x"ca",
          2299 => x"91",
          2300 => x"89",
          2301 => x"08",
          2302 => x"86",
          2303 => x"98",
          2304 => x"91",
          2305 => x"8b",
          2306 => x"fb",
          2307 => x"70",
          2308 => x"81",
          2309 => x"fc",
          2310 => x"ca",
          2311 => x"91",
          2312 => x"b4",
          2313 => x"08",
          2314 => x"ec",
          2315 => x"ca",
          2316 => x"91",
          2317 => x"a0",
          2318 => x"91",
          2319 => x"52",
          2320 => x"51",
          2321 => x"8b",
          2322 => x"52",
          2323 => x"51",
          2324 => x"81",
          2325 => x"34",
          2326 => x"88",
          2327 => x"0d",
          2328 => x"0d",
          2329 => x"98",
          2330 => x"70",
          2331 => x"ec",
          2332 => x"ca",
          2333 => x"38",
          2334 => x"53",
          2335 => x"81",
          2336 => x"34",
          2337 => x"04",
          2338 => x"78",
          2339 => x"80",
          2340 => x"34",
          2341 => x"80",
          2342 => x"38",
          2343 => x"18",
          2344 => x"9c",
          2345 => x"70",
          2346 => x"56",
          2347 => x"a0",
          2348 => x"71",
          2349 => x"81",
          2350 => x"81",
          2351 => x"89",
          2352 => x"06",
          2353 => x"73",
          2354 => x"55",
          2355 => x"55",
          2356 => x"81",
          2357 => x"81",
          2358 => x"74",
          2359 => x"75",
          2360 => x"52",
          2361 => x"13",
          2362 => x"08",
          2363 => x"33",
          2364 => x"9c",
          2365 => x"11",
          2366 => x"8a",
          2367 => x"88",
          2368 => x"96",
          2369 => x"e7",
          2370 => x"88",
          2371 => x"23",
          2372 => x"e7",
          2373 => x"ca",
          2374 => x"17",
          2375 => x"0d",
          2376 => x"0d",
          2377 => x"5e",
          2378 => x"70",
          2379 => x"55",
          2380 => x"83",
          2381 => x"73",
          2382 => x"91",
          2383 => x"2e",
          2384 => x"1d",
          2385 => x"0c",
          2386 => x"15",
          2387 => x"70",
          2388 => x"56",
          2389 => x"09",
          2390 => x"38",
          2391 => x"80",
          2392 => x"30",
          2393 => x"78",
          2394 => x"54",
          2395 => x"73",
          2396 => x"60",
          2397 => x"54",
          2398 => x"96",
          2399 => x"0b",
          2400 => x"80",
          2401 => x"f6",
          2402 => x"ca",
          2403 => x"85",
          2404 => x"3d",
          2405 => x"5c",
          2406 => x"53",
          2407 => x"51",
          2408 => x"80",
          2409 => x"88",
          2410 => x"5c",
          2411 => x"09",
          2412 => x"d4",
          2413 => x"70",
          2414 => x"71",
          2415 => x"30",
          2416 => x"73",
          2417 => x"51",
          2418 => x"57",
          2419 => x"38",
          2420 => x"75",
          2421 => x"17",
          2422 => x"75",
          2423 => x"30",
          2424 => x"51",
          2425 => x"80",
          2426 => x"38",
          2427 => x"87",
          2428 => x"26",
          2429 => x"77",
          2430 => x"a4",
          2431 => x"27",
          2432 => x"a0",
          2433 => x"39",
          2434 => x"33",
          2435 => x"57",
          2436 => x"27",
          2437 => x"75",
          2438 => x"30",
          2439 => x"32",
          2440 => x"80",
          2441 => x"25",
          2442 => x"56",
          2443 => x"80",
          2444 => x"84",
          2445 => x"58",
          2446 => x"70",
          2447 => x"55",
          2448 => x"09",
          2449 => x"38",
          2450 => x"80",
          2451 => x"30",
          2452 => x"77",
          2453 => x"54",
          2454 => x"81",
          2455 => x"ae",
          2456 => x"06",
          2457 => x"54",
          2458 => x"74",
          2459 => x"80",
          2460 => x"7b",
          2461 => x"30",
          2462 => x"70",
          2463 => x"25",
          2464 => x"07",
          2465 => x"51",
          2466 => x"a7",
          2467 => x"8b",
          2468 => x"39",
          2469 => x"54",
          2470 => x"8c",
          2471 => x"ff",
          2472 => x"94",
          2473 => x"54",
          2474 => x"e1",
          2475 => x"88",
          2476 => x"b2",
          2477 => x"70",
          2478 => x"71",
          2479 => x"54",
          2480 => x"91",
          2481 => x"80",
          2482 => x"38",
          2483 => x"76",
          2484 => x"df",
          2485 => x"54",
          2486 => x"81",
          2487 => x"55",
          2488 => x"34",
          2489 => x"52",
          2490 => x"51",
          2491 => x"91",
          2492 => x"bf",
          2493 => x"16",
          2494 => x"26",
          2495 => x"16",
          2496 => x"06",
          2497 => x"17",
          2498 => x"34",
          2499 => x"fd",
          2500 => x"19",
          2501 => x"80",
          2502 => x"79",
          2503 => x"81",
          2504 => x"81",
          2505 => x"85",
          2506 => x"54",
          2507 => x"8f",
          2508 => x"86",
          2509 => x"39",
          2510 => x"f3",
          2511 => x"73",
          2512 => x"80",
          2513 => x"52",
          2514 => x"ce",
          2515 => x"88",
          2516 => x"ca",
          2517 => x"d7",
          2518 => x"08",
          2519 => x"e6",
          2520 => x"ca",
          2521 => x"91",
          2522 => x"80",
          2523 => x"1b",
          2524 => x"55",
          2525 => x"2e",
          2526 => x"8b",
          2527 => x"06",
          2528 => x"1c",
          2529 => x"33",
          2530 => x"70",
          2531 => x"55",
          2532 => x"38",
          2533 => x"52",
          2534 => x"9f",
          2535 => x"88",
          2536 => x"8b",
          2537 => x"7a",
          2538 => x"3f",
          2539 => x"75",
          2540 => x"57",
          2541 => x"2e",
          2542 => x"84",
          2543 => x"06",
          2544 => x"75",
          2545 => x"81",
          2546 => x"2a",
          2547 => x"73",
          2548 => x"38",
          2549 => x"54",
          2550 => x"fb",
          2551 => x"80",
          2552 => x"34",
          2553 => x"c1",
          2554 => x"06",
          2555 => x"38",
          2556 => x"39",
          2557 => x"70",
          2558 => x"54",
          2559 => x"86",
          2560 => x"84",
          2561 => x"06",
          2562 => x"73",
          2563 => x"38",
          2564 => x"83",
          2565 => x"b4",
          2566 => x"51",
          2567 => x"91",
          2568 => x"88",
          2569 => x"ea",
          2570 => x"ca",
          2571 => x"3d",
          2572 => x"3d",
          2573 => x"ff",
          2574 => x"71",
          2575 => x"5c",
          2576 => x"80",
          2577 => x"38",
          2578 => x"05",
          2579 => x"a0",
          2580 => x"71",
          2581 => x"38",
          2582 => x"71",
          2583 => x"81",
          2584 => x"38",
          2585 => x"11",
          2586 => x"06",
          2587 => x"70",
          2588 => x"38",
          2589 => x"81",
          2590 => x"05",
          2591 => x"76",
          2592 => x"38",
          2593 => x"b9",
          2594 => x"77",
          2595 => x"57",
          2596 => x"05",
          2597 => x"70",
          2598 => x"33",
          2599 => x"53",
          2600 => x"99",
          2601 => x"e0",
          2602 => x"ff",
          2603 => x"ff",
          2604 => x"70",
          2605 => x"38",
          2606 => x"81",
          2607 => x"51",
          2608 => x"9f",
          2609 => x"72",
          2610 => x"81",
          2611 => x"70",
          2612 => x"72",
          2613 => x"32",
          2614 => x"72",
          2615 => x"73",
          2616 => x"53",
          2617 => x"70",
          2618 => x"38",
          2619 => x"19",
          2620 => x"75",
          2621 => x"38",
          2622 => x"83",
          2623 => x"74",
          2624 => x"59",
          2625 => x"39",
          2626 => x"33",
          2627 => x"ca",
          2628 => x"3d",
          2629 => x"3d",
          2630 => x"80",
          2631 => x"34",
          2632 => x"17",
          2633 => x"75",
          2634 => x"3f",
          2635 => x"ca",
          2636 => x"80",
          2637 => x"16",
          2638 => x"3f",
          2639 => x"08",
          2640 => x"06",
          2641 => x"73",
          2642 => x"2e",
          2643 => x"80",
          2644 => x"0b",
          2645 => x"56",
          2646 => x"e9",
          2647 => x"06",
          2648 => x"57",
          2649 => x"32",
          2650 => x"80",
          2651 => x"51",
          2652 => x"8a",
          2653 => x"e8",
          2654 => x"06",
          2655 => x"53",
          2656 => x"52",
          2657 => x"51",
          2658 => x"91",
          2659 => x"55",
          2660 => x"08",
          2661 => x"38",
          2662 => x"b8",
          2663 => x"86",
          2664 => x"97",
          2665 => x"88",
          2666 => x"ca",
          2667 => x"2e",
          2668 => x"55",
          2669 => x"88",
          2670 => x"0d",
          2671 => x"0d",
          2672 => x"05",
          2673 => x"33",
          2674 => x"75",
          2675 => x"fc",
          2676 => x"ca",
          2677 => x"8b",
          2678 => x"91",
          2679 => x"24",
          2680 => x"91",
          2681 => x"84",
          2682 => x"a4",
          2683 => x"55",
          2684 => x"73",
          2685 => x"e6",
          2686 => x"0c",
          2687 => x"06",
          2688 => x"57",
          2689 => x"ae",
          2690 => x"33",
          2691 => x"3f",
          2692 => x"08",
          2693 => x"70",
          2694 => x"55",
          2695 => x"76",
          2696 => x"b8",
          2697 => x"2a",
          2698 => x"51",
          2699 => x"72",
          2700 => x"86",
          2701 => x"74",
          2702 => x"15",
          2703 => x"81",
          2704 => x"d7",
          2705 => x"ca",
          2706 => x"ff",
          2707 => x"06",
          2708 => x"56",
          2709 => x"38",
          2710 => x"8f",
          2711 => x"2a",
          2712 => x"51",
          2713 => x"72",
          2714 => x"80",
          2715 => x"52",
          2716 => x"3f",
          2717 => x"08",
          2718 => x"57",
          2719 => x"09",
          2720 => x"e2",
          2721 => x"74",
          2722 => x"56",
          2723 => x"33",
          2724 => x"72",
          2725 => x"38",
          2726 => x"51",
          2727 => x"91",
          2728 => x"57",
          2729 => x"84",
          2730 => x"ff",
          2731 => x"56",
          2732 => x"25",
          2733 => x"0b",
          2734 => x"56",
          2735 => x"05",
          2736 => x"83",
          2737 => x"2e",
          2738 => x"52",
          2739 => x"c6",
          2740 => x"88",
          2741 => x"06",
          2742 => x"27",
          2743 => x"16",
          2744 => x"27",
          2745 => x"56",
          2746 => x"84",
          2747 => x"56",
          2748 => x"84",
          2749 => x"14",
          2750 => x"3f",
          2751 => x"08",
          2752 => x"06",
          2753 => x"80",
          2754 => x"06",
          2755 => x"80",
          2756 => x"db",
          2757 => x"ca",
          2758 => x"ff",
          2759 => x"77",
          2760 => x"d8",
          2761 => x"de",
          2762 => x"88",
          2763 => x"9c",
          2764 => x"c4",
          2765 => x"15",
          2766 => x"14",
          2767 => x"70",
          2768 => x"51",
          2769 => x"56",
          2770 => x"84",
          2771 => x"81",
          2772 => x"71",
          2773 => x"16",
          2774 => x"53",
          2775 => x"23",
          2776 => x"8b",
          2777 => x"73",
          2778 => x"80",
          2779 => x"8d",
          2780 => x"39",
          2781 => x"51",
          2782 => x"91",
          2783 => x"53",
          2784 => x"08",
          2785 => x"72",
          2786 => x"8d",
          2787 => x"ce",
          2788 => x"14",
          2789 => x"3f",
          2790 => x"08",
          2791 => x"06",
          2792 => x"38",
          2793 => x"51",
          2794 => x"91",
          2795 => x"55",
          2796 => x"51",
          2797 => x"91",
          2798 => x"83",
          2799 => x"53",
          2800 => x"80",
          2801 => x"38",
          2802 => x"78",
          2803 => x"2a",
          2804 => x"78",
          2805 => x"86",
          2806 => x"22",
          2807 => x"31",
          2808 => x"83",
          2809 => x"88",
          2810 => x"ca",
          2811 => x"2e",
          2812 => x"91",
          2813 => x"80",
          2814 => x"f5",
          2815 => x"83",
          2816 => x"ff",
          2817 => x"38",
          2818 => x"9f",
          2819 => x"38",
          2820 => x"39",
          2821 => x"80",
          2822 => x"38",
          2823 => x"98",
          2824 => x"a0",
          2825 => x"1c",
          2826 => x"0c",
          2827 => x"17",
          2828 => x"76",
          2829 => x"81",
          2830 => x"80",
          2831 => x"d9",
          2832 => x"ca",
          2833 => x"ff",
          2834 => x"8d",
          2835 => x"8e",
          2836 => x"8a",
          2837 => x"14",
          2838 => x"3f",
          2839 => x"08",
          2840 => x"74",
          2841 => x"a2",
          2842 => x"79",
          2843 => x"ee",
          2844 => x"a8",
          2845 => x"15",
          2846 => x"2e",
          2847 => x"10",
          2848 => x"2a",
          2849 => x"05",
          2850 => x"ff",
          2851 => x"53",
          2852 => x"9c",
          2853 => x"81",
          2854 => x"0b",
          2855 => x"ff",
          2856 => x"0c",
          2857 => x"84",
          2858 => x"83",
          2859 => x"06",
          2860 => x"80",
          2861 => x"d8",
          2862 => x"ca",
          2863 => x"ff",
          2864 => x"72",
          2865 => x"81",
          2866 => x"38",
          2867 => x"73",
          2868 => x"3f",
          2869 => x"08",
          2870 => x"91",
          2871 => x"84",
          2872 => x"b2",
          2873 => x"87",
          2874 => x"88",
          2875 => x"ff",
          2876 => x"82",
          2877 => x"09",
          2878 => x"c8",
          2879 => x"51",
          2880 => x"91",
          2881 => x"84",
          2882 => x"d2",
          2883 => x"06",
          2884 => x"98",
          2885 => x"ee",
          2886 => x"88",
          2887 => x"85",
          2888 => x"09",
          2889 => x"38",
          2890 => x"51",
          2891 => x"91",
          2892 => x"90",
          2893 => x"a0",
          2894 => x"ca",
          2895 => x"88",
          2896 => x"0c",
          2897 => x"91",
          2898 => x"81",
          2899 => x"91",
          2900 => x"72",
          2901 => x"80",
          2902 => x"0c",
          2903 => x"91",
          2904 => x"90",
          2905 => x"fb",
          2906 => x"54",
          2907 => x"80",
          2908 => x"73",
          2909 => x"80",
          2910 => x"72",
          2911 => x"80",
          2912 => x"86",
          2913 => x"15",
          2914 => x"71",
          2915 => x"81",
          2916 => x"81",
          2917 => x"d0",
          2918 => x"ca",
          2919 => x"06",
          2920 => x"38",
          2921 => x"54",
          2922 => x"80",
          2923 => x"71",
          2924 => x"91",
          2925 => x"87",
          2926 => x"fa",
          2927 => x"ab",
          2928 => x"58",
          2929 => x"05",
          2930 => x"e6",
          2931 => x"80",
          2932 => x"88",
          2933 => x"38",
          2934 => x"08",
          2935 => x"ca",
          2936 => x"08",
          2937 => x"80",
          2938 => x"80",
          2939 => x"54",
          2940 => x"84",
          2941 => x"34",
          2942 => x"75",
          2943 => x"2e",
          2944 => x"53",
          2945 => x"53",
          2946 => x"f7",
          2947 => x"ca",
          2948 => x"73",
          2949 => x"0c",
          2950 => x"04",
          2951 => x"67",
          2952 => x"80",
          2953 => x"59",
          2954 => x"78",
          2955 => x"c8",
          2956 => x"06",
          2957 => x"3d",
          2958 => x"99",
          2959 => x"52",
          2960 => x"3f",
          2961 => x"08",
          2962 => x"88",
          2963 => x"38",
          2964 => x"52",
          2965 => x"52",
          2966 => x"3f",
          2967 => x"08",
          2968 => x"88",
          2969 => x"02",
          2970 => x"33",
          2971 => x"55",
          2972 => x"25",
          2973 => x"55",
          2974 => x"54",
          2975 => x"81",
          2976 => x"80",
          2977 => x"74",
          2978 => x"81",
          2979 => x"75",
          2980 => x"3f",
          2981 => x"08",
          2982 => x"02",
          2983 => x"91",
          2984 => x"81",
          2985 => x"82",
          2986 => x"06",
          2987 => x"80",
          2988 => x"88",
          2989 => x"39",
          2990 => x"58",
          2991 => x"38",
          2992 => x"70",
          2993 => x"54",
          2994 => x"81",
          2995 => x"52",
          2996 => x"a5",
          2997 => x"88",
          2998 => x"88",
          2999 => x"62",
          3000 => x"d4",
          3001 => x"54",
          3002 => x"15",
          3003 => x"62",
          3004 => x"e8",
          3005 => x"52",
          3006 => x"51",
          3007 => x"7a",
          3008 => x"83",
          3009 => x"80",
          3010 => x"38",
          3011 => x"08",
          3012 => x"53",
          3013 => x"3d",
          3014 => x"dd",
          3015 => x"ca",
          3016 => x"91",
          3017 => x"82",
          3018 => x"39",
          3019 => x"38",
          3020 => x"33",
          3021 => x"70",
          3022 => x"55",
          3023 => x"2e",
          3024 => x"55",
          3025 => x"77",
          3026 => x"81",
          3027 => x"73",
          3028 => x"38",
          3029 => x"54",
          3030 => x"a0",
          3031 => x"82",
          3032 => x"52",
          3033 => x"a3",
          3034 => x"88",
          3035 => x"18",
          3036 => x"55",
          3037 => x"88",
          3038 => x"38",
          3039 => x"70",
          3040 => x"54",
          3041 => x"86",
          3042 => x"c0",
          3043 => x"b0",
          3044 => x"1b",
          3045 => x"1b",
          3046 => x"70",
          3047 => x"d9",
          3048 => x"88",
          3049 => x"88",
          3050 => x"0c",
          3051 => x"52",
          3052 => x"3f",
          3053 => x"08",
          3054 => x"08",
          3055 => x"77",
          3056 => x"86",
          3057 => x"1a",
          3058 => x"1a",
          3059 => x"91",
          3060 => x"0b",
          3061 => x"80",
          3062 => x"0c",
          3063 => x"70",
          3064 => x"54",
          3065 => x"81",
          3066 => x"ca",
          3067 => x"2e",
          3068 => x"91",
          3069 => x"94",
          3070 => x"17",
          3071 => x"2b",
          3072 => x"57",
          3073 => x"52",
          3074 => x"9f",
          3075 => x"88",
          3076 => x"ca",
          3077 => x"26",
          3078 => x"55",
          3079 => x"08",
          3080 => x"81",
          3081 => x"79",
          3082 => x"31",
          3083 => x"70",
          3084 => x"25",
          3085 => x"76",
          3086 => x"81",
          3087 => x"55",
          3088 => x"38",
          3089 => x"0c",
          3090 => x"75",
          3091 => x"54",
          3092 => x"a2",
          3093 => x"7a",
          3094 => x"3f",
          3095 => x"08",
          3096 => x"55",
          3097 => x"89",
          3098 => x"88",
          3099 => x"1a",
          3100 => x"80",
          3101 => x"54",
          3102 => x"88",
          3103 => x"0d",
          3104 => x"0d",
          3105 => x"64",
          3106 => x"59",
          3107 => x"90",
          3108 => x"52",
          3109 => x"cf",
          3110 => x"88",
          3111 => x"ca",
          3112 => x"38",
          3113 => x"55",
          3114 => x"86",
          3115 => x"82",
          3116 => x"19",
          3117 => x"55",
          3118 => x"80",
          3119 => x"38",
          3120 => x"0b",
          3121 => x"82",
          3122 => x"39",
          3123 => x"1a",
          3124 => x"82",
          3125 => x"19",
          3126 => x"08",
          3127 => x"7c",
          3128 => x"74",
          3129 => x"2e",
          3130 => x"94",
          3131 => x"83",
          3132 => x"56",
          3133 => x"38",
          3134 => x"22",
          3135 => x"89",
          3136 => x"55",
          3137 => x"75",
          3138 => x"19",
          3139 => x"39",
          3140 => x"52",
          3141 => x"93",
          3142 => x"88",
          3143 => x"75",
          3144 => x"38",
          3145 => x"ff",
          3146 => x"98",
          3147 => x"19",
          3148 => x"51",
          3149 => x"91",
          3150 => x"80",
          3151 => x"38",
          3152 => x"08",
          3153 => x"2a",
          3154 => x"80",
          3155 => x"38",
          3156 => x"8a",
          3157 => x"5c",
          3158 => x"27",
          3159 => x"7a",
          3160 => x"54",
          3161 => x"52",
          3162 => x"51",
          3163 => x"91",
          3164 => x"fe",
          3165 => x"83",
          3166 => x"56",
          3167 => x"9f",
          3168 => x"08",
          3169 => x"74",
          3170 => x"38",
          3171 => x"b4",
          3172 => x"16",
          3173 => x"89",
          3174 => x"51",
          3175 => x"77",
          3176 => x"b9",
          3177 => x"1a",
          3178 => x"08",
          3179 => x"84",
          3180 => x"57",
          3181 => x"27",
          3182 => x"56",
          3183 => x"52",
          3184 => x"c7",
          3185 => x"88",
          3186 => x"38",
          3187 => x"19",
          3188 => x"06",
          3189 => x"52",
          3190 => x"a2",
          3191 => x"31",
          3192 => x"7f",
          3193 => x"94",
          3194 => x"94",
          3195 => x"5c",
          3196 => x"80",
          3197 => x"ca",
          3198 => x"3d",
          3199 => x"3d",
          3200 => x"65",
          3201 => x"5d",
          3202 => x"0c",
          3203 => x"05",
          3204 => x"f6",
          3205 => x"ca",
          3206 => x"91",
          3207 => x"8a",
          3208 => x"33",
          3209 => x"2e",
          3210 => x"56",
          3211 => x"90",
          3212 => x"81",
          3213 => x"06",
          3214 => x"87",
          3215 => x"2e",
          3216 => x"95",
          3217 => x"91",
          3218 => x"56",
          3219 => x"81",
          3220 => x"34",
          3221 => x"8e",
          3222 => x"08",
          3223 => x"56",
          3224 => x"84",
          3225 => x"5c",
          3226 => x"82",
          3227 => x"18",
          3228 => x"ff",
          3229 => x"74",
          3230 => x"7e",
          3231 => x"ff",
          3232 => x"2a",
          3233 => x"7a",
          3234 => x"8c",
          3235 => x"08",
          3236 => x"38",
          3237 => x"39",
          3238 => x"52",
          3239 => x"e7",
          3240 => x"88",
          3241 => x"ca",
          3242 => x"2e",
          3243 => x"74",
          3244 => x"91",
          3245 => x"2e",
          3246 => x"74",
          3247 => x"88",
          3248 => x"38",
          3249 => x"0c",
          3250 => x"15",
          3251 => x"08",
          3252 => x"06",
          3253 => x"51",
          3254 => x"91",
          3255 => x"fe",
          3256 => x"18",
          3257 => x"51",
          3258 => x"91",
          3259 => x"80",
          3260 => x"38",
          3261 => x"08",
          3262 => x"2a",
          3263 => x"80",
          3264 => x"38",
          3265 => x"8a",
          3266 => x"5b",
          3267 => x"27",
          3268 => x"7b",
          3269 => x"54",
          3270 => x"52",
          3271 => x"51",
          3272 => x"91",
          3273 => x"fe",
          3274 => x"b0",
          3275 => x"31",
          3276 => x"79",
          3277 => x"84",
          3278 => x"16",
          3279 => x"89",
          3280 => x"52",
          3281 => x"cc",
          3282 => x"55",
          3283 => x"16",
          3284 => x"2b",
          3285 => x"39",
          3286 => x"94",
          3287 => x"93",
          3288 => x"cd",
          3289 => x"ca",
          3290 => x"e3",
          3291 => x"b0",
          3292 => x"76",
          3293 => x"94",
          3294 => x"ff",
          3295 => x"71",
          3296 => x"7b",
          3297 => x"38",
          3298 => x"18",
          3299 => x"51",
          3300 => x"91",
          3301 => x"fd",
          3302 => x"53",
          3303 => x"18",
          3304 => x"06",
          3305 => x"51",
          3306 => x"7e",
          3307 => x"83",
          3308 => x"76",
          3309 => x"17",
          3310 => x"1e",
          3311 => x"18",
          3312 => x"0c",
          3313 => x"58",
          3314 => x"74",
          3315 => x"38",
          3316 => x"8c",
          3317 => x"90",
          3318 => x"33",
          3319 => x"55",
          3320 => x"34",
          3321 => x"91",
          3322 => x"90",
          3323 => x"f8",
          3324 => x"8b",
          3325 => x"53",
          3326 => x"f2",
          3327 => x"ca",
          3328 => x"91",
          3329 => x"80",
          3330 => x"16",
          3331 => x"2a",
          3332 => x"51",
          3333 => x"80",
          3334 => x"38",
          3335 => x"52",
          3336 => x"e7",
          3337 => x"88",
          3338 => x"ca",
          3339 => x"d4",
          3340 => x"08",
          3341 => x"a0",
          3342 => x"73",
          3343 => x"88",
          3344 => x"74",
          3345 => x"51",
          3346 => x"8c",
          3347 => x"9c",
          3348 => x"fb",
          3349 => x"b2",
          3350 => x"15",
          3351 => x"3f",
          3352 => x"15",
          3353 => x"3f",
          3354 => x"0b",
          3355 => x"78",
          3356 => x"3f",
          3357 => x"08",
          3358 => x"81",
          3359 => x"57",
          3360 => x"34",
          3361 => x"88",
          3362 => x"0d",
          3363 => x"0d",
          3364 => x"54",
          3365 => x"91",
          3366 => x"53",
          3367 => x"08",
          3368 => x"3d",
          3369 => x"73",
          3370 => x"3f",
          3371 => x"08",
          3372 => x"88",
          3373 => x"91",
          3374 => x"74",
          3375 => x"ca",
          3376 => x"3d",
          3377 => x"3d",
          3378 => x"51",
          3379 => x"8b",
          3380 => x"91",
          3381 => x"24",
          3382 => x"ca",
          3383 => x"ca",
          3384 => x"52",
          3385 => x"88",
          3386 => x"0d",
          3387 => x"0d",
          3388 => x"3d",
          3389 => x"94",
          3390 => x"c1",
          3391 => x"88",
          3392 => x"ca",
          3393 => x"e0",
          3394 => x"63",
          3395 => x"d4",
          3396 => x"8d",
          3397 => x"88",
          3398 => x"ca",
          3399 => x"38",
          3400 => x"05",
          3401 => x"2b",
          3402 => x"80",
          3403 => x"76",
          3404 => x"0c",
          3405 => x"02",
          3406 => x"70",
          3407 => x"81",
          3408 => x"56",
          3409 => x"9e",
          3410 => x"53",
          3411 => x"db",
          3412 => x"ca",
          3413 => x"15",
          3414 => x"91",
          3415 => x"84",
          3416 => x"06",
          3417 => x"55",
          3418 => x"88",
          3419 => x"0d",
          3420 => x"0d",
          3421 => x"5b",
          3422 => x"80",
          3423 => x"ff",
          3424 => x"9f",
          3425 => x"b5",
          3426 => x"88",
          3427 => x"ca",
          3428 => x"fc",
          3429 => x"7a",
          3430 => x"08",
          3431 => x"64",
          3432 => x"2e",
          3433 => x"a0",
          3434 => x"70",
          3435 => x"ea",
          3436 => x"88",
          3437 => x"ca",
          3438 => x"d4",
          3439 => x"7b",
          3440 => x"3f",
          3441 => x"08",
          3442 => x"88",
          3443 => x"38",
          3444 => x"51",
          3445 => x"91",
          3446 => x"45",
          3447 => x"51",
          3448 => x"91",
          3449 => x"57",
          3450 => x"08",
          3451 => x"80",
          3452 => x"da",
          3453 => x"ca",
          3454 => x"91",
          3455 => x"a4",
          3456 => x"7b",
          3457 => x"3f",
          3458 => x"88",
          3459 => x"38",
          3460 => x"51",
          3461 => x"91",
          3462 => x"57",
          3463 => x"08",
          3464 => x"38",
          3465 => x"09",
          3466 => x"38",
          3467 => x"e0",
          3468 => x"dc",
          3469 => x"ff",
          3470 => x"74",
          3471 => x"3f",
          3472 => x"78",
          3473 => x"33",
          3474 => x"56",
          3475 => x"91",
          3476 => x"05",
          3477 => x"81",
          3478 => x"56",
          3479 => x"f5",
          3480 => x"54",
          3481 => x"81",
          3482 => x"80",
          3483 => x"78",
          3484 => x"55",
          3485 => x"11",
          3486 => x"18",
          3487 => x"58",
          3488 => x"34",
          3489 => x"ff",
          3490 => x"55",
          3491 => x"34",
          3492 => x"77",
          3493 => x"81",
          3494 => x"ff",
          3495 => x"55",
          3496 => x"34",
          3497 => x"ca",
          3498 => x"84",
          3499 => x"84",
          3500 => x"70",
          3501 => x"56",
          3502 => x"76",
          3503 => x"81",
          3504 => x"70",
          3505 => x"56",
          3506 => x"82",
          3507 => x"78",
          3508 => x"80",
          3509 => x"27",
          3510 => x"19",
          3511 => x"7a",
          3512 => x"5c",
          3513 => x"55",
          3514 => x"7a",
          3515 => x"5c",
          3516 => x"2e",
          3517 => x"85",
          3518 => x"94",
          3519 => x"81",
          3520 => x"73",
          3521 => x"81",
          3522 => x"7a",
          3523 => x"38",
          3524 => x"76",
          3525 => x"0c",
          3526 => x"04",
          3527 => x"7b",
          3528 => x"fc",
          3529 => x"53",
          3530 => x"bb",
          3531 => x"88",
          3532 => x"ca",
          3533 => x"fa",
          3534 => x"33",
          3535 => x"f2",
          3536 => x"08",
          3537 => x"27",
          3538 => x"15",
          3539 => x"2a",
          3540 => x"51",
          3541 => x"83",
          3542 => x"94",
          3543 => x"80",
          3544 => x"0c",
          3545 => x"2e",
          3546 => x"79",
          3547 => x"70",
          3548 => x"51",
          3549 => x"2e",
          3550 => x"52",
          3551 => x"ff",
          3552 => x"91",
          3553 => x"ff",
          3554 => x"70",
          3555 => x"ff",
          3556 => x"91",
          3557 => x"73",
          3558 => x"76",
          3559 => x"06",
          3560 => x"0c",
          3561 => x"98",
          3562 => x"58",
          3563 => x"39",
          3564 => x"54",
          3565 => x"73",
          3566 => x"cd",
          3567 => x"ca",
          3568 => x"91",
          3569 => x"81",
          3570 => x"38",
          3571 => x"08",
          3572 => x"9b",
          3573 => x"88",
          3574 => x"0c",
          3575 => x"0c",
          3576 => x"81",
          3577 => x"76",
          3578 => x"38",
          3579 => x"94",
          3580 => x"94",
          3581 => x"16",
          3582 => x"2a",
          3583 => x"51",
          3584 => x"72",
          3585 => x"38",
          3586 => x"51",
          3587 => x"91",
          3588 => x"54",
          3589 => x"08",
          3590 => x"ca",
          3591 => x"a7",
          3592 => x"74",
          3593 => x"3f",
          3594 => x"08",
          3595 => x"2e",
          3596 => x"74",
          3597 => x"79",
          3598 => x"14",
          3599 => x"38",
          3600 => x"0c",
          3601 => x"94",
          3602 => x"94",
          3603 => x"83",
          3604 => x"72",
          3605 => x"38",
          3606 => x"51",
          3607 => x"91",
          3608 => x"94",
          3609 => x"91",
          3610 => x"53",
          3611 => x"81",
          3612 => x"34",
          3613 => x"39",
          3614 => x"91",
          3615 => x"05",
          3616 => x"08",
          3617 => x"08",
          3618 => x"38",
          3619 => x"0c",
          3620 => x"80",
          3621 => x"72",
          3622 => x"73",
          3623 => x"53",
          3624 => x"8c",
          3625 => x"16",
          3626 => x"38",
          3627 => x"0c",
          3628 => x"91",
          3629 => x"8b",
          3630 => x"f9",
          3631 => x"56",
          3632 => x"80",
          3633 => x"38",
          3634 => x"3d",
          3635 => x"8a",
          3636 => x"51",
          3637 => x"91",
          3638 => x"55",
          3639 => x"08",
          3640 => x"77",
          3641 => x"52",
          3642 => x"b5",
          3643 => x"88",
          3644 => x"ca",
          3645 => x"c3",
          3646 => x"33",
          3647 => x"55",
          3648 => x"24",
          3649 => x"16",
          3650 => x"2a",
          3651 => x"51",
          3652 => x"80",
          3653 => x"9c",
          3654 => x"77",
          3655 => x"3f",
          3656 => x"08",
          3657 => x"77",
          3658 => x"22",
          3659 => x"74",
          3660 => x"ce",
          3661 => x"ca",
          3662 => x"74",
          3663 => x"81",
          3664 => x"85",
          3665 => x"74",
          3666 => x"38",
          3667 => x"74",
          3668 => x"ca",
          3669 => x"3d",
          3670 => x"3d",
          3671 => x"3d",
          3672 => x"70",
          3673 => x"ff",
          3674 => x"88",
          3675 => x"91",
          3676 => x"73",
          3677 => x"0d",
          3678 => x"0d",
          3679 => x"3d",
          3680 => x"71",
          3681 => x"e7",
          3682 => x"ca",
          3683 => x"91",
          3684 => x"80",
          3685 => x"93",
          3686 => x"88",
          3687 => x"51",
          3688 => x"91",
          3689 => x"53",
          3690 => x"91",
          3691 => x"52",
          3692 => x"ac",
          3693 => x"88",
          3694 => x"ca",
          3695 => x"2e",
          3696 => x"85",
          3697 => x"87",
          3698 => x"88",
          3699 => x"74",
          3700 => x"d5",
          3701 => x"52",
          3702 => x"89",
          3703 => x"88",
          3704 => x"70",
          3705 => x"07",
          3706 => x"91",
          3707 => x"06",
          3708 => x"54",
          3709 => x"88",
          3710 => x"0d",
          3711 => x"0d",
          3712 => x"53",
          3713 => x"53",
          3714 => x"56",
          3715 => x"91",
          3716 => x"55",
          3717 => x"08",
          3718 => x"52",
          3719 => x"81",
          3720 => x"88",
          3721 => x"ca",
          3722 => x"38",
          3723 => x"05",
          3724 => x"2b",
          3725 => x"80",
          3726 => x"86",
          3727 => x"76",
          3728 => x"38",
          3729 => x"51",
          3730 => x"74",
          3731 => x"0c",
          3732 => x"04",
          3733 => x"63",
          3734 => x"80",
          3735 => x"ec",
          3736 => x"3d",
          3737 => x"3f",
          3738 => x"08",
          3739 => x"88",
          3740 => x"38",
          3741 => x"73",
          3742 => x"08",
          3743 => x"13",
          3744 => x"58",
          3745 => x"26",
          3746 => x"7c",
          3747 => x"39",
          3748 => x"cc",
          3749 => x"81",
          3750 => x"ca",
          3751 => x"33",
          3752 => x"81",
          3753 => x"06",
          3754 => x"75",
          3755 => x"52",
          3756 => x"05",
          3757 => x"3f",
          3758 => x"08",
          3759 => x"38",
          3760 => x"08",
          3761 => x"38",
          3762 => x"08",
          3763 => x"ca",
          3764 => x"80",
          3765 => x"81",
          3766 => x"59",
          3767 => x"14",
          3768 => x"ca",
          3769 => x"39",
          3770 => x"91",
          3771 => x"57",
          3772 => x"38",
          3773 => x"18",
          3774 => x"ff",
          3775 => x"91",
          3776 => x"5b",
          3777 => x"08",
          3778 => x"7c",
          3779 => x"12",
          3780 => x"52",
          3781 => x"82",
          3782 => x"06",
          3783 => x"14",
          3784 => x"cb",
          3785 => x"88",
          3786 => x"ff",
          3787 => x"70",
          3788 => x"82",
          3789 => x"51",
          3790 => x"b4",
          3791 => x"bb",
          3792 => x"ca",
          3793 => x"0a",
          3794 => x"70",
          3795 => x"84",
          3796 => x"51",
          3797 => x"ff",
          3798 => x"56",
          3799 => x"38",
          3800 => x"7c",
          3801 => x"0c",
          3802 => x"81",
          3803 => x"74",
          3804 => x"7a",
          3805 => x"0c",
          3806 => x"04",
          3807 => x"79",
          3808 => x"05",
          3809 => x"57",
          3810 => x"91",
          3811 => x"56",
          3812 => x"08",
          3813 => x"91",
          3814 => x"75",
          3815 => x"90",
          3816 => x"81",
          3817 => x"06",
          3818 => x"87",
          3819 => x"2e",
          3820 => x"94",
          3821 => x"73",
          3822 => x"27",
          3823 => x"73",
          3824 => x"ca",
          3825 => x"88",
          3826 => x"76",
          3827 => x"3f",
          3828 => x"08",
          3829 => x"0c",
          3830 => x"39",
          3831 => x"52",
          3832 => x"bf",
          3833 => x"ca",
          3834 => x"2e",
          3835 => x"83",
          3836 => x"91",
          3837 => x"81",
          3838 => x"06",
          3839 => x"56",
          3840 => x"a0",
          3841 => x"91",
          3842 => x"98",
          3843 => x"94",
          3844 => x"08",
          3845 => x"88",
          3846 => x"51",
          3847 => x"91",
          3848 => x"56",
          3849 => x"8c",
          3850 => x"17",
          3851 => x"07",
          3852 => x"18",
          3853 => x"2e",
          3854 => x"91",
          3855 => x"55",
          3856 => x"88",
          3857 => x"0d",
          3858 => x"0d",
          3859 => x"3d",
          3860 => x"52",
          3861 => x"da",
          3862 => x"ca",
          3863 => x"91",
          3864 => x"81",
          3865 => x"45",
          3866 => x"52",
          3867 => x"52",
          3868 => x"3f",
          3869 => x"08",
          3870 => x"88",
          3871 => x"38",
          3872 => x"05",
          3873 => x"2a",
          3874 => x"51",
          3875 => x"55",
          3876 => x"38",
          3877 => x"54",
          3878 => x"81",
          3879 => x"80",
          3880 => x"70",
          3881 => x"54",
          3882 => x"81",
          3883 => x"52",
          3884 => x"c5",
          3885 => x"88",
          3886 => x"2a",
          3887 => x"51",
          3888 => x"80",
          3889 => x"38",
          3890 => x"ca",
          3891 => x"15",
          3892 => x"86",
          3893 => x"91",
          3894 => x"5c",
          3895 => x"3d",
          3896 => x"c7",
          3897 => x"ca",
          3898 => x"91",
          3899 => x"80",
          3900 => x"ca",
          3901 => x"73",
          3902 => x"3f",
          3903 => x"08",
          3904 => x"88",
          3905 => x"87",
          3906 => x"39",
          3907 => x"08",
          3908 => x"38",
          3909 => x"08",
          3910 => x"77",
          3911 => x"3f",
          3912 => x"08",
          3913 => x"08",
          3914 => x"ca",
          3915 => x"80",
          3916 => x"55",
          3917 => x"94",
          3918 => x"2e",
          3919 => x"53",
          3920 => x"51",
          3921 => x"91",
          3922 => x"55",
          3923 => x"78",
          3924 => x"fe",
          3925 => x"88",
          3926 => x"91",
          3927 => x"a0",
          3928 => x"e9",
          3929 => x"53",
          3930 => x"05",
          3931 => x"51",
          3932 => x"91",
          3933 => x"54",
          3934 => x"08",
          3935 => x"78",
          3936 => x"8e",
          3937 => x"58",
          3938 => x"91",
          3939 => x"54",
          3940 => x"08",
          3941 => x"54",
          3942 => x"91",
          3943 => x"84",
          3944 => x"06",
          3945 => x"02",
          3946 => x"33",
          3947 => x"81",
          3948 => x"86",
          3949 => x"f6",
          3950 => x"74",
          3951 => x"70",
          3952 => x"c3",
          3953 => x"88",
          3954 => x"56",
          3955 => x"08",
          3956 => x"54",
          3957 => x"08",
          3958 => x"81",
          3959 => x"82",
          3960 => x"88",
          3961 => x"09",
          3962 => x"38",
          3963 => x"b4",
          3964 => x"b0",
          3965 => x"88",
          3966 => x"51",
          3967 => x"91",
          3968 => x"54",
          3969 => x"08",
          3970 => x"8b",
          3971 => x"b4",
          3972 => x"b7",
          3973 => x"54",
          3974 => x"15",
          3975 => x"90",
          3976 => x"34",
          3977 => x"0a",
          3978 => x"19",
          3979 => x"9f",
          3980 => x"78",
          3981 => x"51",
          3982 => x"a0",
          3983 => x"11",
          3984 => x"05",
          3985 => x"b6",
          3986 => x"ae",
          3987 => x"15",
          3988 => x"78",
          3989 => x"53",
          3990 => x"3f",
          3991 => x"0b",
          3992 => x"77",
          3993 => x"3f",
          3994 => x"08",
          3995 => x"88",
          3996 => x"82",
          3997 => x"52",
          3998 => x"51",
          3999 => x"3f",
          4000 => x"52",
          4001 => x"aa",
          4002 => x"90",
          4003 => x"34",
          4004 => x"0b",
          4005 => x"78",
          4006 => x"b6",
          4007 => x"88",
          4008 => x"39",
          4009 => x"52",
          4010 => x"be",
          4011 => x"91",
          4012 => x"99",
          4013 => x"da",
          4014 => x"3d",
          4015 => x"d2",
          4016 => x"53",
          4017 => x"84",
          4018 => x"3d",
          4019 => x"3f",
          4020 => x"08",
          4021 => x"88",
          4022 => x"38",
          4023 => x"3d",
          4024 => x"3d",
          4025 => x"cc",
          4026 => x"ca",
          4027 => x"91",
          4028 => x"82",
          4029 => x"81",
          4030 => x"81",
          4031 => x"86",
          4032 => x"aa",
          4033 => x"a4",
          4034 => x"a8",
          4035 => x"05",
          4036 => x"ea",
          4037 => x"77",
          4038 => x"70",
          4039 => x"b4",
          4040 => x"3d",
          4041 => x"51",
          4042 => x"91",
          4043 => x"55",
          4044 => x"08",
          4045 => x"6f",
          4046 => x"06",
          4047 => x"a2",
          4048 => x"92",
          4049 => x"81",
          4050 => x"ca",
          4051 => x"2e",
          4052 => x"81",
          4053 => x"51",
          4054 => x"91",
          4055 => x"55",
          4056 => x"08",
          4057 => x"68",
          4058 => x"a8",
          4059 => x"05",
          4060 => x"51",
          4061 => x"3f",
          4062 => x"33",
          4063 => x"8b",
          4064 => x"84",
          4065 => x"06",
          4066 => x"73",
          4067 => x"a0",
          4068 => x"8b",
          4069 => x"54",
          4070 => x"15",
          4071 => x"33",
          4072 => x"70",
          4073 => x"55",
          4074 => x"2e",
          4075 => x"6e",
          4076 => x"df",
          4077 => x"78",
          4078 => x"3f",
          4079 => x"08",
          4080 => x"ff",
          4081 => x"82",
          4082 => x"88",
          4083 => x"80",
          4084 => x"ca",
          4085 => x"78",
          4086 => x"af",
          4087 => x"88",
          4088 => x"d4",
          4089 => x"55",
          4090 => x"08",
          4091 => x"81",
          4092 => x"73",
          4093 => x"81",
          4094 => x"63",
          4095 => x"76",
          4096 => x"3f",
          4097 => x"0b",
          4098 => x"87",
          4099 => x"88",
          4100 => x"77",
          4101 => x"3f",
          4102 => x"08",
          4103 => x"88",
          4104 => x"78",
          4105 => x"aa",
          4106 => x"88",
          4107 => x"91",
          4108 => x"a8",
          4109 => x"ed",
          4110 => x"80",
          4111 => x"02",
          4112 => x"df",
          4113 => x"57",
          4114 => x"3d",
          4115 => x"96",
          4116 => x"e9",
          4117 => x"88",
          4118 => x"ca",
          4119 => x"cf",
          4120 => x"65",
          4121 => x"d4",
          4122 => x"b5",
          4123 => x"88",
          4124 => x"ca",
          4125 => x"38",
          4126 => x"05",
          4127 => x"06",
          4128 => x"73",
          4129 => x"a7",
          4130 => x"09",
          4131 => x"71",
          4132 => x"06",
          4133 => x"55",
          4134 => x"15",
          4135 => x"81",
          4136 => x"34",
          4137 => x"b4",
          4138 => x"ca",
          4139 => x"74",
          4140 => x"0c",
          4141 => x"04",
          4142 => x"64",
          4143 => x"93",
          4144 => x"52",
          4145 => x"d1",
          4146 => x"ca",
          4147 => x"91",
          4148 => x"80",
          4149 => x"58",
          4150 => x"3d",
          4151 => x"c8",
          4152 => x"ca",
          4153 => x"91",
          4154 => x"b4",
          4155 => x"c7",
          4156 => x"a0",
          4157 => x"55",
          4158 => x"84",
          4159 => x"17",
          4160 => x"2b",
          4161 => x"96",
          4162 => x"b0",
          4163 => x"54",
          4164 => x"15",
          4165 => x"ff",
          4166 => x"91",
          4167 => x"55",
          4168 => x"88",
          4169 => x"0d",
          4170 => x"0d",
          4171 => x"5a",
          4172 => x"3d",
          4173 => x"99",
          4174 => x"81",
          4175 => x"88",
          4176 => x"88",
          4177 => x"91",
          4178 => x"07",
          4179 => x"55",
          4180 => x"2e",
          4181 => x"81",
          4182 => x"55",
          4183 => x"2e",
          4184 => x"7b",
          4185 => x"80",
          4186 => x"70",
          4187 => x"be",
          4188 => x"ca",
          4189 => x"91",
          4190 => x"80",
          4191 => x"52",
          4192 => x"dc",
          4193 => x"88",
          4194 => x"ca",
          4195 => x"38",
          4196 => x"08",
          4197 => x"08",
          4198 => x"56",
          4199 => x"19",
          4200 => x"59",
          4201 => x"74",
          4202 => x"56",
          4203 => x"ec",
          4204 => x"75",
          4205 => x"74",
          4206 => x"2e",
          4207 => x"16",
          4208 => x"33",
          4209 => x"73",
          4210 => x"38",
          4211 => x"84",
          4212 => x"06",
          4213 => x"7a",
          4214 => x"76",
          4215 => x"07",
          4216 => x"54",
          4217 => x"80",
          4218 => x"80",
          4219 => x"7b",
          4220 => x"53",
          4221 => x"93",
          4222 => x"88",
          4223 => x"ca",
          4224 => x"38",
          4225 => x"55",
          4226 => x"56",
          4227 => x"8b",
          4228 => x"56",
          4229 => x"83",
          4230 => x"75",
          4231 => x"51",
          4232 => x"3f",
          4233 => x"08",
          4234 => x"91",
          4235 => x"98",
          4236 => x"e6",
          4237 => x"53",
          4238 => x"b8",
          4239 => x"3d",
          4240 => x"3f",
          4241 => x"08",
          4242 => x"08",
          4243 => x"ca",
          4244 => x"98",
          4245 => x"a0",
          4246 => x"70",
          4247 => x"ae",
          4248 => x"6d",
          4249 => x"81",
          4250 => x"57",
          4251 => x"74",
          4252 => x"38",
          4253 => x"81",
          4254 => x"81",
          4255 => x"52",
          4256 => x"89",
          4257 => x"88",
          4258 => x"a5",
          4259 => x"33",
          4260 => x"54",
          4261 => x"3f",
          4262 => x"08",
          4263 => x"38",
          4264 => x"76",
          4265 => x"05",
          4266 => x"39",
          4267 => x"08",
          4268 => x"15",
          4269 => x"ff",
          4270 => x"73",
          4271 => x"38",
          4272 => x"83",
          4273 => x"56",
          4274 => x"75",
          4275 => x"91",
          4276 => x"33",
          4277 => x"2e",
          4278 => x"52",
          4279 => x"51",
          4280 => x"3f",
          4281 => x"08",
          4282 => x"ff",
          4283 => x"38",
          4284 => x"88",
          4285 => x"8a",
          4286 => x"38",
          4287 => x"ec",
          4288 => x"75",
          4289 => x"74",
          4290 => x"73",
          4291 => x"05",
          4292 => x"17",
          4293 => x"70",
          4294 => x"34",
          4295 => x"70",
          4296 => x"ff",
          4297 => x"55",
          4298 => x"26",
          4299 => x"8b",
          4300 => x"86",
          4301 => x"e5",
          4302 => x"38",
          4303 => x"99",
          4304 => x"05",
          4305 => x"70",
          4306 => x"73",
          4307 => x"81",
          4308 => x"ff",
          4309 => x"ed",
          4310 => x"80",
          4311 => x"91",
          4312 => x"55",
          4313 => x"3f",
          4314 => x"08",
          4315 => x"88",
          4316 => x"38",
          4317 => x"51",
          4318 => x"3f",
          4319 => x"08",
          4320 => x"88",
          4321 => x"76",
          4322 => x"67",
          4323 => x"34",
          4324 => x"91",
          4325 => x"84",
          4326 => x"06",
          4327 => x"80",
          4328 => x"2e",
          4329 => x"81",
          4330 => x"ff",
          4331 => x"91",
          4332 => x"54",
          4333 => x"08",
          4334 => x"53",
          4335 => x"08",
          4336 => x"ff",
          4337 => x"67",
          4338 => x"8b",
          4339 => x"53",
          4340 => x"51",
          4341 => x"3f",
          4342 => x"0b",
          4343 => x"79",
          4344 => x"ee",
          4345 => x"88",
          4346 => x"55",
          4347 => x"88",
          4348 => x"0d",
          4349 => x"0d",
          4350 => x"88",
          4351 => x"05",
          4352 => x"fc",
          4353 => x"54",
          4354 => x"d2",
          4355 => x"ca",
          4356 => x"91",
          4357 => x"82",
          4358 => x"1a",
          4359 => x"82",
          4360 => x"80",
          4361 => x"8c",
          4362 => x"78",
          4363 => x"1a",
          4364 => x"2a",
          4365 => x"51",
          4366 => x"90",
          4367 => x"82",
          4368 => x"58",
          4369 => x"81",
          4370 => x"39",
          4371 => x"22",
          4372 => x"70",
          4373 => x"56",
          4374 => x"82",
          4375 => x"14",
          4376 => x"30",
          4377 => x"9f",
          4378 => x"88",
          4379 => x"19",
          4380 => x"5a",
          4381 => x"81",
          4382 => x"38",
          4383 => x"77",
          4384 => x"82",
          4385 => x"56",
          4386 => x"74",
          4387 => x"ff",
          4388 => x"81",
          4389 => x"55",
          4390 => x"75",
          4391 => x"82",
          4392 => x"88",
          4393 => x"ff",
          4394 => x"ca",
          4395 => x"2e",
          4396 => x"91",
          4397 => x"8e",
          4398 => x"56",
          4399 => x"09",
          4400 => x"38",
          4401 => x"59",
          4402 => x"77",
          4403 => x"06",
          4404 => x"87",
          4405 => x"39",
          4406 => x"ba",
          4407 => x"55",
          4408 => x"2e",
          4409 => x"15",
          4410 => x"2e",
          4411 => x"83",
          4412 => x"75",
          4413 => x"7e",
          4414 => x"a8",
          4415 => x"88",
          4416 => x"ca",
          4417 => x"ce",
          4418 => x"16",
          4419 => x"56",
          4420 => x"38",
          4421 => x"19",
          4422 => x"8c",
          4423 => x"7d",
          4424 => x"38",
          4425 => x"0c",
          4426 => x"0c",
          4427 => x"80",
          4428 => x"73",
          4429 => x"98",
          4430 => x"05",
          4431 => x"57",
          4432 => x"26",
          4433 => x"7b",
          4434 => x"0c",
          4435 => x"81",
          4436 => x"84",
          4437 => x"54",
          4438 => x"88",
          4439 => x"0d",
          4440 => x"0d",
          4441 => x"88",
          4442 => x"05",
          4443 => x"54",
          4444 => x"c5",
          4445 => x"56",
          4446 => x"ca",
          4447 => x"8b",
          4448 => x"ca",
          4449 => x"29",
          4450 => x"05",
          4451 => x"55",
          4452 => x"84",
          4453 => x"34",
          4454 => x"08",
          4455 => x"5f",
          4456 => x"51",
          4457 => x"3f",
          4458 => x"08",
          4459 => x"70",
          4460 => x"57",
          4461 => x"8b",
          4462 => x"82",
          4463 => x"06",
          4464 => x"56",
          4465 => x"38",
          4466 => x"05",
          4467 => x"7e",
          4468 => x"f0",
          4469 => x"88",
          4470 => x"67",
          4471 => x"2e",
          4472 => x"82",
          4473 => x"8b",
          4474 => x"75",
          4475 => x"80",
          4476 => x"81",
          4477 => x"2e",
          4478 => x"80",
          4479 => x"38",
          4480 => x"0a",
          4481 => x"ff",
          4482 => x"55",
          4483 => x"86",
          4484 => x"8a",
          4485 => x"89",
          4486 => x"2a",
          4487 => x"77",
          4488 => x"59",
          4489 => x"81",
          4490 => x"70",
          4491 => x"07",
          4492 => x"56",
          4493 => x"38",
          4494 => x"05",
          4495 => x"7e",
          4496 => x"80",
          4497 => x"91",
          4498 => x"8a",
          4499 => x"83",
          4500 => x"06",
          4501 => x"08",
          4502 => x"74",
          4503 => x"41",
          4504 => x"56",
          4505 => x"8a",
          4506 => x"61",
          4507 => x"55",
          4508 => x"27",
          4509 => x"93",
          4510 => x"80",
          4511 => x"38",
          4512 => x"70",
          4513 => x"43",
          4514 => x"95",
          4515 => x"06",
          4516 => x"2e",
          4517 => x"77",
          4518 => x"74",
          4519 => x"83",
          4520 => x"06",
          4521 => x"82",
          4522 => x"2e",
          4523 => x"78",
          4524 => x"2e",
          4525 => x"80",
          4526 => x"ae",
          4527 => x"2a",
          4528 => x"91",
          4529 => x"56",
          4530 => x"2e",
          4531 => x"77",
          4532 => x"91",
          4533 => x"79",
          4534 => x"70",
          4535 => x"5a",
          4536 => x"86",
          4537 => x"27",
          4538 => x"52",
          4539 => x"fc",
          4540 => x"ca",
          4541 => x"29",
          4542 => x"70",
          4543 => x"55",
          4544 => x"0b",
          4545 => x"08",
          4546 => x"05",
          4547 => x"ff",
          4548 => x"27",
          4549 => x"88",
          4550 => x"ae",
          4551 => x"2a",
          4552 => x"91",
          4553 => x"56",
          4554 => x"2e",
          4555 => x"77",
          4556 => x"91",
          4557 => x"79",
          4558 => x"70",
          4559 => x"5a",
          4560 => x"86",
          4561 => x"27",
          4562 => x"52",
          4563 => x"fc",
          4564 => x"ca",
          4565 => x"84",
          4566 => x"ca",
          4567 => x"f5",
          4568 => x"81",
          4569 => x"88",
          4570 => x"ca",
          4571 => x"71",
          4572 => x"83",
          4573 => x"5e",
          4574 => x"89",
          4575 => x"5c",
          4576 => x"1c",
          4577 => x"05",
          4578 => x"ff",
          4579 => x"70",
          4580 => x"31",
          4581 => x"57",
          4582 => x"83",
          4583 => x"06",
          4584 => x"1c",
          4585 => x"5c",
          4586 => x"1d",
          4587 => x"29",
          4588 => x"31",
          4589 => x"55",
          4590 => x"87",
          4591 => x"7c",
          4592 => x"7a",
          4593 => x"31",
          4594 => x"fb",
          4595 => x"ca",
          4596 => x"7d",
          4597 => x"81",
          4598 => x"91",
          4599 => x"83",
          4600 => x"80",
          4601 => x"87",
          4602 => x"81",
          4603 => x"fd",
          4604 => x"f8",
          4605 => x"2e",
          4606 => x"80",
          4607 => x"ff",
          4608 => x"ca",
          4609 => x"a0",
          4610 => x"38",
          4611 => x"74",
          4612 => x"86",
          4613 => x"fd",
          4614 => x"81",
          4615 => x"80",
          4616 => x"83",
          4617 => x"39",
          4618 => x"08",
          4619 => x"92",
          4620 => x"b8",
          4621 => x"59",
          4622 => x"27",
          4623 => x"86",
          4624 => x"55",
          4625 => x"09",
          4626 => x"38",
          4627 => x"f5",
          4628 => x"38",
          4629 => x"55",
          4630 => x"86",
          4631 => x"80",
          4632 => x"7a",
          4633 => x"b9",
          4634 => x"91",
          4635 => x"7a",
          4636 => x"8a",
          4637 => x"52",
          4638 => x"ff",
          4639 => x"79",
          4640 => x"7b",
          4641 => x"06",
          4642 => x"51",
          4643 => x"3f",
          4644 => x"1c",
          4645 => x"32",
          4646 => x"96",
          4647 => x"06",
          4648 => x"91",
          4649 => x"a1",
          4650 => x"55",
          4651 => x"ff",
          4652 => x"74",
          4653 => x"06",
          4654 => x"51",
          4655 => x"3f",
          4656 => x"52",
          4657 => x"ff",
          4658 => x"f8",
          4659 => x"34",
          4660 => x"1b",
          4661 => x"d9",
          4662 => x"52",
          4663 => x"ff",
          4664 => x"60",
          4665 => x"51",
          4666 => x"3f",
          4667 => x"09",
          4668 => x"cb",
          4669 => x"b2",
          4670 => x"c3",
          4671 => x"a0",
          4672 => x"52",
          4673 => x"ff",
          4674 => x"82",
          4675 => x"51",
          4676 => x"3f",
          4677 => x"1b",
          4678 => x"95",
          4679 => x"b2",
          4680 => x"a0",
          4681 => x"80",
          4682 => x"1c",
          4683 => x"80",
          4684 => x"93",
          4685 => x"dc",
          4686 => x"1b",
          4687 => x"82",
          4688 => x"52",
          4689 => x"ff",
          4690 => x"7c",
          4691 => x"06",
          4692 => x"51",
          4693 => x"3f",
          4694 => x"a4",
          4695 => x"0b",
          4696 => x"93",
          4697 => x"f0",
          4698 => x"51",
          4699 => x"3f",
          4700 => x"52",
          4701 => x"70",
          4702 => x"9f",
          4703 => x"54",
          4704 => x"52",
          4705 => x"9b",
          4706 => x"56",
          4707 => x"08",
          4708 => x"7d",
          4709 => x"81",
          4710 => x"38",
          4711 => x"86",
          4712 => x"52",
          4713 => x"9b",
          4714 => x"80",
          4715 => x"7a",
          4716 => x"ed",
          4717 => x"85",
          4718 => x"7a",
          4719 => x"8f",
          4720 => x"85",
          4721 => x"83",
          4722 => x"ff",
          4723 => x"ff",
          4724 => x"e8",
          4725 => x"9e",
          4726 => x"52",
          4727 => x"51",
          4728 => x"3f",
          4729 => x"52",
          4730 => x"9e",
          4731 => x"54",
          4732 => x"53",
          4733 => x"51",
          4734 => x"3f",
          4735 => x"16",
          4736 => x"7e",
          4737 => x"d8",
          4738 => x"80",
          4739 => x"ff",
          4740 => x"7f",
          4741 => x"7d",
          4742 => x"81",
          4743 => x"f8",
          4744 => x"ff",
          4745 => x"ff",
          4746 => x"51",
          4747 => x"3f",
          4748 => x"88",
          4749 => x"39",
          4750 => x"f8",
          4751 => x"2e",
          4752 => x"55",
          4753 => x"51",
          4754 => x"3f",
          4755 => x"57",
          4756 => x"83",
          4757 => x"76",
          4758 => x"7a",
          4759 => x"ff",
          4760 => x"91",
          4761 => x"82",
          4762 => x"80",
          4763 => x"88",
          4764 => x"51",
          4765 => x"3f",
          4766 => x"78",
          4767 => x"74",
          4768 => x"18",
          4769 => x"2e",
          4770 => x"79",
          4771 => x"2e",
          4772 => x"55",
          4773 => x"62",
          4774 => x"74",
          4775 => x"75",
          4776 => x"7e",
          4777 => x"b8",
          4778 => x"88",
          4779 => x"38",
          4780 => x"78",
          4781 => x"74",
          4782 => x"56",
          4783 => x"93",
          4784 => x"66",
          4785 => x"26",
          4786 => x"56",
          4787 => x"83",
          4788 => x"64",
          4789 => x"77",
          4790 => x"84",
          4791 => x"52",
          4792 => x"9d",
          4793 => x"d4",
          4794 => x"51",
          4795 => x"3f",
          4796 => x"55",
          4797 => x"81",
          4798 => x"34",
          4799 => x"16",
          4800 => x"16",
          4801 => x"16",
          4802 => x"05",
          4803 => x"c1",
          4804 => x"fe",
          4805 => x"fe",
          4806 => x"34",
          4807 => x"08",
          4808 => x"07",
          4809 => x"16",
          4810 => x"88",
          4811 => x"34",
          4812 => x"c6",
          4813 => x"9c",
          4814 => x"52",
          4815 => x"51",
          4816 => x"3f",
          4817 => x"53",
          4818 => x"51",
          4819 => x"3f",
          4820 => x"ca",
          4821 => x"38",
          4822 => x"52",
          4823 => x"99",
          4824 => x"56",
          4825 => x"08",
          4826 => x"39",
          4827 => x"39",
          4828 => x"39",
          4829 => x"08",
          4830 => x"ca",
          4831 => x"3d",
          4832 => x"3d",
          4833 => x"71",
          4834 => x"8e",
          4835 => x"29",
          4836 => x"05",
          4837 => x"04",
          4838 => x"51",
          4839 => x"91",
          4840 => x"80",
          4841 => x"bb",
          4842 => x"f2",
          4843 => x"8c",
          4844 => x"39",
          4845 => x"51",
          4846 => x"91",
          4847 => x"80",
          4848 => x"bc",
          4849 => x"d6",
          4850 => x"d0",
          4851 => x"39",
          4852 => x"51",
          4853 => x"91",
          4854 => x"80",
          4855 => x"bd",
          4856 => x"39",
          4857 => x"51",
          4858 => x"bd",
          4859 => x"39",
          4860 => x"51",
          4861 => x"be",
          4862 => x"39",
          4863 => x"51",
          4864 => x"be",
          4865 => x"39",
          4866 => x"51",
          4867 => x"be",
          4868 => x"39",
          4869 => x"51",
          4870 => x"bf",
          4871 => x"87",
          4872 => x"3d",
          4873 => x"3d",
          4874 => x"56",
          4875 => x"e7",
          4876 => x"74",
          4877 => x"e8",
          4878 => x"39",
          4879 => x"74",
          4880 => x"a3",
          4881 => x"88",
          4882 => x"51",
          4883 => x"3f",
          4884 => x"08",
          4885 => x"75",
          4886 => x"a0",
          4887 => x"a0",
          4888 => x"0d",
          4889 => x"0d",
          4890 => x"02",
          4891 => x"c7",
          4892 => x"73",
          4893 => x"5d",
          4894 => x"5c",
          4895 => x"91",
          4896 => x"ff",
          4897 => x"91",
          4898 => x"ff",
          4899 => x"80",
          4900 => x"27",
          4901 => x"79",
          4902 => x"38",
          4903 => x"a7",
          4904 => x"39",
          4905 => x"72",
          4906 => x"38",
          4907 => x"91",
          4908 => x"ff",
          4909 => x"89",
          4910 => x"dc",
          4911 => x"dc",
          4912 => x"55",
          4913 => x"74",
          4914 => x"78",
          4915 => x"72",
          4916 => x"bf",
          4917 => x"8c",
          4918 => x"39",
          4919 => x"51",
          4920 => x"3f",
          4921 => x"a1",
          4922 => x"53",
          4923 => x"8e",
          4924 => x"52",
          4925 => x"51",
          4926 => x"3f",
          4927 => x"bf",
          4928 => x"86",
          4929 => x"15",
          4930 => x"fe",
          4931 => x"ff",
          4932 => x"bf",
          4933 => x"86",
          4934 => x"55",
          4935 => x"aa",
          4936 => x"70",
          4937 => x"26",
          4938 => x"9f",
          4939 => x"38",
          4940 => x"8b",
          4941 => x"fe",
          4942 => x"73",
          4943 => x"a0",
          4944 => x"d7",
          4945 => x"55",
          4946 => x"bf",
          4947 => x"85",
          4948 => x"16",
          4949 => x"56",
          4950 => x"3f",
          4951 => x"08",
          4952 => x"98",
          4953 => x"74",
          4954 => x"81",
          4955 => x"fe",
          4956 => x"91",
          4957 => x"98",
          4958 => x"2c",
          4959 => x"70",
          4960 => x"07",
          4961 => x"56",
          4962 => x"74",
          4963 => x"38",
          4964 => x"74",
          4965 => x"81",
          4966 => x"80",
          4967 => x"7a",
          4968 => x"76",
          4969 => x"38",
          4970 => x"91",
          4971 => x"8d",
          4972 => x"ec",
          4973 => x"02",
          4974 => x"e3",
          4975 => x"72",
          4976 => x"07",
          4977 => x"87",
          4978 => x"07",
          4979 => x"5a",
          4980 => x"57",
          4981 => x"38",
          4982 => x"52",
          4983 => x"52",
          4984 => x"3f",
          4985 => x"08",
          4986 => x"88",
          4987 => x"91",
          4988 => x"87",
          4989 => x"0c",
          4990 => x"08",
          4991 => x"d4",
          4992 => x"80",
          4993 => x"76",
          4994 => x"3f",
          4995 => x"08",
          4996 => x"88",
          4997 => x"7a",
          4998 => x"2e",
          4999 => x"19",
          5000 => x"59",
          5001 => x"3d",
          5002 => x"cc",
          5003 => x"30",
          5004 => x"80",
          5005 => x"79",
          5006 => x"38",
          5007 => x"90",
          5008 => x"f8",
          5009 => x"98",
          5010 => x"78",
          5011 => x"3f",
          5012 => x"91",
          5013 => x"96",
          5014 => x"f9",
          5015 => x"02",
          5016 => x"05",
          5017 => x"ff",
          5018 => x"7a",
          5019 => x"fe",
          5020 => x"ca",
          5021 => x"38",
          5022 => x"88",
          5023 => x"2e",
          5024 => x"39",
          5025 => x"54",
          5026 => x"53",
          5027 => x"51",
          5028 => x"ca",
          5029 => x"83",
          5030 => x"76",
          5031 => x"0c",
          5032 => x"04",
          5033 => x"02",
          5034 => x"91",
          5035 => x"91",
          5036 => x"55",
          5037 => x"3f",
          5038 => x"22",
          5039 => x"e2",
          5040 => x"94",
          5041 => x"a0",
          5042 => x"89",
          5043 => x"c0",
          5044 => x"88",
          5045 => x"80",
          5046 => x"fe",
          5047 => x"86",
          5048 => x"fe",
          5049 => x"c0",
          5050 => x"53",
          5051 => x"3f",
          5052 => x"f6",
          5053 => x"c0",
          5054 => x"f8",
          5055 => x"51",
          5056 => x"3f",
          5057 => x"70",
          5058 => x"52",
          5059 => x"95",
          5060 => x"fe",
          5061 => x"91",
          5062 => x"fe",
          5063 => x"80",
          5064 => x"dd",
          5065 => x"2a",
          5066 => x"51",
          5067 => x"2e",
          5068 => x"51",
          5069 => x"3f",
          5070 => x"51",
          5071 => x"3f",
          5072 => x"f5",
          5073 => x"83",
          5074 => x"06",
          5075 => x"80",
          5076 => x"81",
          5077 => x"a9",
          5078 => x"84",
          5079 => x"a1",
          5080 => x"fe",
          5081 => x"72",
          5082 => x"81",
          5083 => x"71",
          5084 => x"38",
          5085 => x"f5",
          5086 => x"c1",
          5087 => x"f7",
          5088 => x"51",
          5089 => x"3f",
          5090 => x"70",
          5091 => x"52",
          5092 => x"95",
          5093 => x"fe",
          5094 => x"91",
          5095 => x"fe",
          5096 => x"80",
          5097 => x"d9",
          5098 => x"2a",
          5099 => x"51",
          5100 => x"2e",
          5101 => x"51",
          5102 => x"3f",
          5103 => x"51",
          5104 => x"3f",
          5105 => x"f4",
          5106 => x"87",
          5107 => x"06",
          5108 => x"80",
          5109 => x"81",
          5110 => x"a5",
          5111 => x"d4",
          5112 => x"9d",
          5113 => x"fe",
          5114 => x"72",
          5115 => x"81",
          5116 => x"71",
          5117 => x"38",
          5118 => x"f4",
          5119 => x"c1",
          5120 => x"f5",
          5121 => x"51",
          5122 => x"3f",
          5123 => x"3f",
          5124 => x"04",
          5125 => x"78",
          5126 => x"55",
          5127 => x"80",
          5128 => x"38",
          5129 => x"77",
          5130 => x"33",
          5131 => x"39",
          5132 => x"80",
          5133 => x"81",
          5134 => x"57",
          5135 => x"2e",
          5136 => x"53",
          5137 => x"84",
          5138 => x"38",
          5139 => x"06",
          5140 => x"2e",
          5141 => x"88",
          5142 => x"70",
          5143 => x"34",
          5144 => x"90",
          5145 => x"a8",
          5146 => x"53",
          5147 => x"55",
          5148 => x"3f",
          5149 => x"08",
          5150 => x"15",
          5151 => x"81",
          5152 => x"38",
          5153 => x"81",
          5154 => x"53",
          5155 => x"d2",
          5156 => x"72",
          5157 => x"0c",
          5158 => x"04",
          5159 => x"80",
          5160 => x"e1",
          5161 => x"5c",
          5162 => x"51",
          5163 => x"3f",
          5164 => x"08",
          5165 => x"59",
          5166 => x"09",
          5167 => x"38",
          5168 => x"52",
          5169 => x"52",
          5170 => x"ca",
          5171 => x"78",
          5172 => x"b8",
          5173 => x"e3",
          5174 => x"88",
          5175 => x"88",
          5176 => x"ac",
          5177 => x"39",
          5178 => x"5c",
          5179 => x"51",
          5180 => x"3f",
          5181 => x"46",
          5182 => x"53",
          5183 => x"51",
          5184 => x"3f",
          5185 => x"64",
          5186 => x"ce",
          5187 => x"fe",
          5188 => x"fd",
          5189 => x"ca",
          5190 => x"2b",
          5191 => x"51",
          5192 => x"c2",
          5193 => x"38",
          5194 => x"24",
          5195 => x"78",
          5196 => x"ef",
          5197 => x"24",
          5198 => x"84",
          5199 => x"38",
          5200 => x"90",
          5201 => x"2e",
          5202 => x"78",
          5203 => x"a9",
          5204 => x"39",
          5205 => x"82",
          5206 => x"ab",
          5207 => x"38",
          5208 => x"78",
          5209 => x"f2",
          5210 => x"24",
          5211 => x"bc",
          5212 => x"38",
          5213 => x"84",
          5214 => x"c8",
          5215 => x"c0",
          5216 => x"38",
          5217 => x"2e",
          5218 => x"8e",
          5219 => x"80",
          5220 => x"a5",
          5221 => x"f8",
          5222 => x"78",
          5223 => x"8c",
          5224 => x"80",
          5225 => x"38",
          5226 => x"2e",
          5227 => x"78",
          5228 => x"8c",
          5229 => x"8c",
          5230 => x"d4",
          5231 => x"38",
          5232 => x"2e",
          5233 => x"8d",
          5234 => x"81",
          5235 => x"e0",
          5236 => x"83",
          5237 => x"78",
          5238 => x"8d",
          5239 => x"81",
          5240 => x"bd",
          5241 => x"39",
          5242 => x"2e",
          5243 => x"78",
          5244 => x"fd",
          5245 => x"cc",
          5246 => x"fe",
          5247 => x"fe",
          5248 => x"ff",
          5249 => x"91",
          5250 => x"88",
          5251 => x"e8",
          5252 => x"39",
          5253 => x"f0",
          5254 => x"f8",
          5255 => x"83",
          5256 => x"ca",
          5257 => x"2e",
          5258 => x"63",
          5259 => x"80",
          5260 => x"cb",
          5261 => x"02",
          5262 => x"33",
          5263 => x"b7",
          5264 => x"88",
          5265 => x"06",
          5266 => x"38",
          5267 => x"51",
          5268 => x"3f",
          5269 => x"94",
          5270 => x"88",
          5271 => x"39",
          5272 => x"f4",
          5273 => x"f8",
          5274 => x"83",
          5275 => x"ca",
          5276 => x"2e",
          5277 => x"80",
          5278 => x"02",
          5279 => x"33",
          5280 => x"c0",
          5281 => x"88",
          5282 => x"c3",
          5283 => x"8a",
          5284 => x"fe",
          5285 => x"fe",
          5286 => x"ff",
          5287 => x"91",
          5288 => x"80",
          5289 => x"63",
          5290 => x"c0",
          5291 => x"fe",
          5292 => x"fe",
          5293 => x"ff",
          5294 => x"91",
          5295 => x"86",
          5296 => x"88",
          5297 => x"53",
          5298 => x"52",
          5299 => x"80",
          5300 => x"80",
          5301 => x"53",
          5302 => x"84",
          5303 => x"cb",
          5304 => x"ff",
          5305 => x"91",
          5306 => x"81",
          5307 => x"c2",
          5308 => x"fa",
          5309 => x"5c",
          5310 => x"b7",
          5311 => x"05",
          5312 => x"ae",
          5313 => x"88",
          5314 => x"fe",
          5315 => x"5b",
          5316 => x"3f",
          5317 => x"ca",
          5318 => x"7a",
          5319 => x"3f",
          5320 => x"b7",
          5321 => x"05",
          5322 => x"86",
          5323 => x"88",
          5324 => x"fe",
          5325 => x"5b",
          5326 => x"3f",
          5327 => x"08",
          5328 => x"f8",
          5329 => x"fe",
          5330 => x"91",
          5331 => x"b8",
          5332 => x"05",
          5333 => x"ea",
          5334 => x"c6",
          5335 => x"ca",
          5336 => x"56",
          5337 => x"ca",
          5338 => x"ff",
          5339 => x"53",
          5340 => x"51",
          5341 => x"91",
          5342 => x"80",
          5343 => x"38",
          5344 => x"08",
          5345 => x"3f",
          5346 => x"b7",
          5347 => x"11",
          5348 => x"05",
          5349 => x"dd",
          5350 => x"88",
          5351 => x"fa",
          5352 => x"3d",
          5353 => x"53",
          5354 => x"51",
          5355 => x"3f",
          5356 => x"08",
          5357 => x"b4",
          5358 => x"fe",
          5359 => x"fe",
          5360 => x"ff",
          5361 => x"91",
          5362 => x"86",
          5363 => x"88",
          5364 => x"c3",
          5365 => x"f8",
          5366 => x"63",
          5367 => x"7b",
          5368 => x"38",
          5369 => x"7a",
          5370 => x"5c",
          5371 => x"26",
          5372 => x"e1",
          5373 => x"fe",
          5374 => x"fe",
          5375 => x"fe",
          5376 => x"91",
          5377 => x"80",
          5378 => x"38",
          5379 => x"f0",
          5380 => x"f8",
          5381 => x"ff",
          5382 => x"ca",
          5383 => x"2e",
          5384 => x"b7",
          5385 => x"11",
          5386 => x"05",
          5387 => x"c5",
          5388 => x"88",
          5389 => x"f9",
          5390 => x"c3",
          5391 => x"f7",
          5392 => x"5a",
          5393 => x"81",
          5394 => x"59",
          5395 => x"05",
          5396 => x"34",
          5397 => x"42",
          5398 => x"3d",
          5399 => x"53",
          5400 => x"51",
          5401 => x"3f",
          5402 => x"08",
          5403 => x"fc",
          5404 => x"fe",
          5405 => x"fe",
          5406 => x"fe",
          5407 => x"91",
          5408 => x"80",
          5409 => x"38",
          5410 => x"ec",
          5411 => x"f8",
          5412 => x"fe",
          5413 => x"ca",
          5414 => x"2e",
          5415 => x"91",
          5416 => x"fe",
          5417 => x"63",
          5418 => x"27",
          5419 => x"70",
          5420 => x"41",
          5421 => x"7f",
          5422 => x"78",
          5423 => x"79",
          5424 => x"52",
          5425 => x"51",
          5426 => x"3f",
          5427 => x"81",
          5428 => x"d5",
          5429 => x"f4",
          5430 => x"39",
          5431 => x"f4",
          5432 => x"f8",
          5433 => x"fe",
          5434 => x"ca",
          5435 => x"c4",
          5436 => x"91",
          5437 => x"80",
          5438 => x"91",
          5439 => x"44",
          5440 => x"c7",
          5441 => x"78",
          5442 => x"38",
          5443 => x"08",
          5444 => x"91",
          5445 => x"59",
          5446 => x"91",
          5447 => x"59",
          5448 => x"88",
          5449 => x"f4",
          5450 => x"39",
          5451 => x"08",
          5452 => x"44",
          5453 => x"f0",
          5454 => x"f8",
          5455 => x"fd",
          5456 => x"ca",
          5457 => x"c3",
          5458 => x"91",
          5459 => x"80",
          5460 => x"91",
          5461 => x"43",
          5462 => x"c7",
          5463 => x"78",
          5464 => x"38",
          5465 => x"08",
          5466 => x"91",
          5467 => x"59",
          5468 => x"91",
          5469 => x"59",
          5470 => x"88",
          5471 => x"f8",
          5472 => x"39",
          5473 => x"08",
          5474 => x"b7",
          5475 => x"11",
          5476 => x"05",
          5477 => x"dd",
          5478 => x"88",
          5479 => x"9b",
          5480 => x"5b",
          5481 => x"2e",
          5482 => x"59",
          5483 => x"8d",
          5484 => x"2e",
          5485 => x"a0",
          5486 => x"88",
          5487 => x"f0",
          5488 => x"d8",
          5489 => x"63",
          5490 => x"62",
          5491 => x"ed",
          5492 => x"c4",
          5493 => x"bd",
          5494 => x"fe",
          5495 => x"fe",
          5496 => x"fe",
          5497 => x"91",
          5498 => x"80",
          5499 => x"38",
          5500 => x"f0",
          5501 => x"f8",
          5502 => x"fb",
          5503 => x"ca",
          5504 => x"2e",
          5505 => x"59",
          5506 => x"05",
          5507 => x"63",
          5508 => x"b7",
          5509 => x"11",
          5510 => x"05",
          5511 => x"d5",
          5512 => x"88",
          5513 => x"f5",
          5514 => x"70",
          5515 => x"91",
          5516 => x"fe",
          5517 => x"80",
          5518 => x"51",
          5519 => x"3f",
          5520 => x"33",
          5521 => x"2e",
          5522 => x"9f",
          5523 => x"38",
          5524 => x"f0",
          5525 => x"f8",
          5526 => x"fb",
          5527 => x"ca",
          5528 => x"2e",
          5529 => x"59",
          5530 => x"05",
          5531 => x"63",
          5532 => x"ff",
          5533 => x"c4",
          5534 => x"f3",
          5535 => x"aa",
          5536 => x"fe",
          5537 => x"fe",
          5538 => x"fe",
          5539 => x"91",
          5540 => x"80",
          5541 => x"38",
          5542 => x"e4",
          5543 => x"f8",
          5544 => x"fc",
          5545 => x"ca",
          5546 => x"2e",
          5547 => x"59",
          5548 => x"22",
          5549 => x"05",
          5550 => x"41",
          5551 => x"e4",
          5552 => x"f8",
          5553 => x"fc",
          5554 => x"ca",
          5555 => x"38",
          5556 => x"60",
          5557 => x"52",
          5558 => x"51",
          5559 => x"3f",
          5560 => x"79",
          5561 => x"f2",
          5562 => x"79",
          5563 => x"ae",
          5564 => x"38",
          5565 => x"87",
          5566 => x"05",
          5567 => x"b7",
          5568 => x"11",
          5569 => x"05",
          5570 => x"db",
          5571 => x"88",
          5572 => x"92",
          5573 => x"02",
          5574 => x"79",
          5575 => x"5b",
          5576 => x"ff",
          5577 => x"c4",
          5578 => x"f1",
          5579 => x"a3",
          5580 => x"fe",
          5581 => x"fe",
          5582 => x"fe",
          5583 => x"91",
          5584 => x"80",
          5585 => x"38",
          5586 => x"e4",
          5587 => x"f8",
          5588 => x"fb",
          5589 => x"ca",
          5590 => x"2e",
          5591 => x"60",
          5592 => x"60",
          5593 => x"b7",
          5594 => x"11",
          5595 => x"05",
          5596 => x"f3",
          5597 => x"88",
          5598 => x"f2",
          5599 => x"70",
          5600 => x"91",
          5601 => x"fe",
          5602 => x"80",
          5603 => x"51",
          5604 => x"3f",
          5605 => x"33",
          5606 => x"2e",
          5607 => x"9f",
          5608 => x"38",
          5609 => x"e4",
          5610 => x"f8",
          5611 => x"fa",
          5612 => x"ca",
          5613 => x"2e",
          5614 => x"53",
          5615 => x"c4",
          5616 => x"f6",
          5617 => x"60",
          5618 => x"60",
          5619 => x"ff",
          5620 => x"c4",
          5621 => x"f0",
          5622 => x"a2",
          5623 => x"b8",
          5624 => x"b8",
          5625 => x"fe",
          5626 => x"f1",
          5627 => x"c4",
          5628 => x"f0",
          5629 => x"51",
          5630 => x"3f",
          5631 => x"84",
          5632 => x"87",
          5633 => x"0c",
          5634 => x"0b",
          5635 => x"94",
          5636 => x"e8",
          5637 => x"84",
          5638 => x"39",
          5639 => x"51",
          5640 => x"3f",
          5641 => x"0b",
          5642 => x"84",
          5643 => x"83",
          5644 => x"94",
          5645 => x"b4",
          5646 => x"fe",
          5647 => x"fe",
          5648 => x"fe",
          5649 => x"91",
          5650 => x"80",
          5651 => x"38",
          5652 => x"c5",
          5653 => x"f5",
          5654 => x"59",
          5655 => x"3d",
          5656 => x"53",
          5657 => x"51",
          5658 => x"3f",
          5659 => x"08",
          5660 => x"f8",
          5661 => x"91",
          5662 => x"fe",
          5663 => x"63",
          5664 => x"91",
          5665 => x"5e",
          5666 => x"08",
          5667 => x"dc",
          5668 => x"88",
          5669 => x"c5",
          5670 => x"f4",
          5671 => x"cc",
          5672 => x"e4",
          5673 => x"f4",
          5674 => x"d4",
          5675 => x"39",
          5676 => x"51",
          5677 => x"3f",
          5678 => x"a0",
          5679 => x"b0",
          5680 => x"39",
          5681 => x"51",
          5682 => x"2e",
          5683 => x"7b",
          5684 => x"d2",
          5685 => x"2e",
          5686 => x"b7",
          5687 => x"05",
          5688 => x"ce",
          5689 => x"94",
          5690 => x"88",
          5691 => x"c6",
          5692 => x"53",
          5693 => x"52",
          5694 => x"52",
          5695 => x"96",
          5696 => x"e4",
          5697 => x"bc",
          5698 => x"64",
          5699 => x"81",
          5700 => x"54",
          5701 => x"53",
          5702 => x"52",
          5703 => x"bb",
          5704 => x"88",
          5705 => x"81",
          5706 => x"32",
          5707 => x"8a",
          5708 => x"2e",
          5709 => x"ef",
          5710 => x"c6",
          5711 => x"f3",
          5712 => x"a8",
          5713 => x"0d",
          5714 => x"ca",
          5715 => x"94",
          5716 => x"ca",
          5717 => x"97",
          5718 => x"ca",
          5719 => x"e5",
          5720 => x"ec",
          5721 => x"c6",
          5722 => x"e3",
          5723 => x"c6",
          5724 => x"ed",
          5725 => x"9d",
          5726 => x"eb",
          5727 => x"51",
          5728 => x"ee",
          5729 => x"04",
          5730 => x"3e",
          5731 => x"44",
          5732 => x"4a",
          5733 => x"50",
          5734 => x"56",
          5735 => x"14",
          5736 => x"98",
          5737 => x"9f",
          5738 => x"a6",
          5739 => x"ad",
          5740 => x"b4",
          5741 => x"bb",
          5742 => x"c2",
          5743 => x"c9",
          5744 => x"d0",
          5745 => x"d7",
          5746 => x"de",
          5747 => x"e4",
          5748 => x"ea",
          5749 => x"f0",
          5750 => x"f6",
          5751 => x"fc",
          5752 => x"02",
          5753 => x"08",
          5754 => x"0e",
          5755 => x"25",
          5756 => x"64",
          5757 => x"3a",
          5758 => x"25",
          5759 => x"64",
          5760 => x"00",
          5761 => x"20",
          5762 => x"66",
          5763 => x"72",
          5764 => x"6f",
          5765 => x"00",
          5766 => x"72",
          5767 => x"53",
          5768 => x"63",
          5769 => x"69",
          5770 => x"00",
          5771 => x"65",
          5772 => x"65",
          5773 => x"6d",
          5774 => x"6d",
          5775 => x"65",
          5776 => x"00",
          5777 => x"20",
          5778 => x"4e",
          5779 => x"41",
          5780 => x"53",
          5781 => x"74",
          5782 => x"38",
          5783 => x"53",
          5784 => x"3d",
          5785 => x"58",
          5786 => x"00",
          5787 => x"20",
          5788 => x"4d",
          5789 => x"74",
          5790 => x"3d",
          5791 => x"58",
          5792 => x"69",
          5793 => x"25",
          5794 => x"29",
          5795 => x"00",
          5796 => x"20",
          5797 => x"20",
          5798 => x"61",
          5799 => x"25",
          5800 => x"2c",
          5801 => x"7a",
          5802 => x"30",
          5803 => x"2e",
          5804 => x"00",
          5805 => x"20",
          5806 => x"54",
          5807 => x"00",
          5808 => x"20",
          5809 => x"0a",
          5810 => x"00",
          5811 => x"20",
          5812 => x"0a",
          5813 => x"00",
          5814 => x"20",
          5815 => x"43",
          5816 => x"20",
          5817 => x"76",
          5818 => x"73",
          5819 => x"32",
          5820 => x"0a",
          5821 => x"00",
          5822 => x"20",
          5823 => x"45",
          5824 => x"50",
          5825 => x"4f",
          5826 => x"4f",
          5827 => x"52",
          5828 => x"00",
          5829 => x"20",
          5830 => x"45",
          5831 => x"28",
          5832 => x"65",
          5833 => x"25",
          5834 => x"29",
          5835 => x"00",
          5836 => x"72",
          5837 => x"65",
          5838 => x"00",
          5839 => x"20",
          5840 => x"20",
          5841 => x"65",
          5842 => x"65",
          5843 => x"72",
          5844 => x"64",
          5845 => x"73",
          5846 => x"25",
          5847 => x"0a",
          5848 => x"00",
          5849 => x"20",
          5850 => x"20",
          5851 => x"6f",
          5852 => x"53",
          5853 => x"74",
          5854 => x"64",
          5855 => x"73",
          5856 => x"25",
          5857 => x"0a",
          5858 => x"00",
          5859 => x"20",
          5860 => x"63",
          5861 => x"74",
          5862 => x"20",
          5863 => x"72",
          5864 => x"20",
          5865 => x"20",
          5866 => x"25",
          5867 => x"0a",
          5868 => x"00",
          5869 => x"20",
          5870 => x"20",
          5871 => x"20",
          5872 => x"20",
          5873 => x"20",
          5874 => x"20",
          5875 => x"20",
          5876 => x"25",
          5877 => x"0a",
          5878 => x"00",
          5879 => x"20",
          5880 => x"74",
          5881 => x"43",
          5882 => x"6b",
          5883 => x"65",
          5884 => x"20",
          5885 => x"20",
          5886 => x"25",
          5887 => x"0a",
          5888 => x"00",
          5889 => x"6c",
          5890 => x"00",
          5891 => x"69",
          5892 => x"00",
          5893 => x"78",
          5894 => x"00",
          5895 => x"00",
          5896 => x"6d",
          5897 => x"00",
          5898 => x"6e",
          5899 => x"00",
          5900 => x"00",
          5901 => x"2c",
          5902 => x"3d",
          5903 => x"5d",
          5904 => x"00",
          5905 => x"00",
          5906 => x"33",
          5907 => x"00",
          5908 => x"4d",
          5909 => x"53",
          5910 => x"00",
          5911 => x"4e",
          5912 => x"20",
          5913 => x"46",
          5914 => x"32",
          5915 => x"00",
          5916 => x"4e",
          5917 => x"20",
          5918 => x"46",
          5919 => x"20",
          5920 => x"00",
          5921 => x"30",
          5922 => x"00",
          5923 => x"00",
          5924 => x"00",
          5925 => x"41",
          5926 => x"80",
          5927 => x"49",
          5928 => x"8f",
          5929 => x"4f",
          5930 => x"55",
          5931 => x"9b",
          5932 => x"9f",
          5933 => x"55",
          5934 => x"a7",
          5935 => x"ab",
          5936 => x"af",
          5937 => x"b3",
          5938 => x"b7",
          5939 => x"bb",
          5940 => x"bf",
          5941 => x"c3",
          5942 => x"c7",
          5943 => x"cb",
          5944 => x"cf",
          5945 => x"d3",
          5946 => x"d7",
          5947 => x"db",
          5948 => x"df",
          5949 => x"e3",
          5950 => x"e7",
          5951 => x"eb",
          5952 => x"ef",
          5953 => x"f3",
          5954 => x"f7",
          5955 => x"fb",
          5956 => x"ff",
          5957 => x"3b",
          5958 => x"2f",
          5959 => x"3a",
          5960 => x"7c",
          5961 => x"00",
          5962 => x"04",
          5963 => x"40",
          5964 => x"00",
          5965 => x"00",
          5966 => x"02",
          5967 => x"08",
          5968 => x"20",
          5969 => x"00",
          5970 => x"69",
          5971 => x"00",
          5972 => x"63",
          5973 => x"00",
          5974 => x"69",
          5975 => x"00",
          5976 => x"61",
          5977 => x"00",
          5978 => x"65",
          5979 => x"00",
          5980 => x"65",
          5981 => x"00",
          5982 => x"70",
          5983 => x"00",
          5984 => x"66",
          5985 => x"00",
          5986 => x"6d",
          5987 => x"00",
          5988 => x"00",
          5989 => x"00",
          5990 => x"00",
          5991 => x"00",
          5992 => x"00",
          5993 => x"00",
          5994 => x"00",
          5995 => x"6c",
          5996 => x"00",
          5997 => x"00",
          5998 => x"74",
          5999 => x"00",
          6000 => x"65",
          6001 => x"00",
          6002 => x"6f",
          6003 => x"00",
          6004 => x"74",
          6005 => x"00",
          6006 => x"6b",
          6007 => x"72",
          6008 => x"00",
          6009 => x"65",
          6010 => x"6c",
          6011 => x"72",
          6012 => x"0a",
          6013 => x"00",
          6014 => x"6b",
          6015 => x"74",
          6016 => x"61",
          6017 => x"0a",
          6018 => x"00",
          6019 => x"66",
          6020 => x"20",
          6021 => x"6e",
          6022 => x"00",
          6023 => x"70",
          6024 => x"20",
          6025 => x"6e",
          6026 => x"00",
          6027 => x"61",
          6028 => x"20",
          6029 => x"65",
          6030 => x"65",
          6031 => x"00",
          6032 => x"65",
          6033 => x"64",
          6034 => x"65",
          6035 => x"00",
          6036 => x"65",
          6037 => x"72",
          6038 => x"79",
          6039 => x"69",
          6040 => x"2e",
          6041 => x"00",
          6042 => x"65",
          6043 => x"6e",
          6044 => x"20",
          6045 => x"61",
          6046 => x"2e",
          6047 => x"00",
          6048 => x"69",
          6049 => x"72",
          6050 => x"20",
          6051 => x"74",
          6052 => x"65",
          6053 => x"00",
          6054 => x"76",
          6055 => x"75",
          6056 => x"72",
          6057 => x"20",
          6058 => x"61",
          6059 => x"2e",
          6060 => x"00",
          6061 => x"6b",
          6062 => x"74",
          6063 => x"61",
          6064 => x"64",
          6065 => x"00",
          6066 => x"63",
          6067 => x"61",
          6068 => x"6c",
          6069 => x"69",
          6070 => x"79",
          6071 => x"6d",
          6072 => x"75",
          6073 => x"6f",
          6074 => x"69",
          6075 => x"0a",
          6076 => x"00",
          6077 => x"6d",
          6078 => x"61",
          6079 => x"74",
          6080 => x"0a",
          6081 => x"00",
          6082 => x"65",
          6083 => x"2c",
          6084 => x"65",
          6085 => x"69",
          6086 => x"63",
          6087 => x"65",
          6088 => x"64",
          6089 => x"00",
          6090 => x"65",
          6091 => x"20",
          6092 => x"6b",
          6093 => x"0a",
          6094 => x"00",
          6095 => x"75",
          6096 => x"63",
          6097 => x"74",
          6098 => x"6d",
          6099 => x"2e",
          6100 => x"00",
          6101 => x"20",
          6102 => x"79",
          6103 => x"65",
          6104 => x"69",
          6105 => x"2e",
          6106 => x"00",
          6107 => x"61",
          6108 => x"65",
          6109 => x"69",
          6110 => x"72",
          6111 => x"74",
          6112 => x"00",
          6113 => x"63",
          6114 => x"2e",
          6115 => x"00",
          6116 => x"6e",
          6117 => x"20",
          6118 => x"6f",
          6119 => x"00",
          6120 => x"75",
          6121 => x"74",
          6122 => x"25",
          6123 => x"74",
          6124 => x"75",
          6125 => x"74",
          6126 => x"73",
          6127 => x"0a",
          6128 => x"00",
          6129 => x"58",
          6130 => x"00",
          6131 => x"00",
          6132 => x"58",
          6133 => x"00",
          6134 => x"20",
          6135 => x"20",
          6136 => x"00",
          6137 => x"58",
          6138 => x"00",
          6139 => x"00",
          6140 => x"00",
          6141 => x"00",
          6142 => x"64",
          6143 => x"00",
          6144 => x"54",
          6145 => x"00",
          6146 => x"20",
          6147 => x"28",
          6148 => x"00",
          6149 => x"30",
          6150 => x"30",
          6151 => x"00",
          6152 => x"33",
          6153 => x"00",
          6154 => x"55",
          6155 => x"65",
          6156 => x"30",
          6157 => x"20",
          6158 => x"25",
          6159 => x"2a",
          6160 => x"00",
          6161 => x"54",
          6162 => x"6e",
          6163 => x"72",
          6164 => x"20",
          6165 => x"64",
          6166 => x"0a",
          6167 => x"00",
          6168 => x"65",
          6169 => x"6e",
          6170 => x"72",
          6171 => x"0a",
          6172 => x"00",
          6173 => x"20",
          6174 => x"65",
          6175 => x"70",
          6176 => x"00",
          6177 => x"54",
          6178 => x"44",
          6179 => x"74",
          6180 => x"75",
          6181 => x"00",
          6182 => x"54",
          6183 => x"52",
          6184 => x"74",
          6185 => x"75",
          6186 => x"00",
          6187 => x"54",
          6188 => x"58",
          6189 => x"74",
          6190 => x"75",
          6191 => x"00",
          6192 => x"54",
          6193 => x"58",
          6194 => x"74",
          6195 => x"75",
          6196 => x"00",
          6197 => x"54",
          6198 => x"58",
          6199 => x"74",
          6200 => x"75",
          6201 => x"00",
          6202 => x"54",
          6203 => x"58",
          6204 => x"74",
          6205 => x"75",
          6206 => x"00",
          6207 => x"74",
          6208 => x"20",
          6209 => x"74",
          6210 => x"72",
          6211 => x"0a",
          6212 => x"00",
          6213 => x"62",
          6214 => x"67",
          6215 => x"6d",
          6216 => x"2e",
          6217 => x"00",
          6218 => x"00",
          6219 => x"6c",
          6220 => x"74",
          6221 => x"6e",
          6222 => x"61",
          6223 => x"65",
          6224 => x"20",
          6225 => x"64",
          6226 => x"20",
          6227 => x"61",
          6228 => x"69",
          6229 => x"20",
          6230 => x"75",
          6231 => x"79",
          6232 => x"00",
          6233 => x"00",
          6234 => x"20",
          6235 => x"6b",
          6236 => x"21",
          6237 => x"00",
          6238 => x"74",
          6239 => x"69",
          6240 => x"2e",
          6241 => x"00",
          6242 => x"6c",
          6243 => x"74",
          6244 => x"6e",
          6245 => x"61",
          6246 => x"65",
          6247 => x"00",
          6248 => x"25",
          6249 => x"00",
          6250 => x"00",
          6251 => x"61",
          6252 => x"67",
          6253 => x"00",
          6254 => x"79",
          6255 => x"2e",
          6256 => x"00",
          6257 => x"70",
          6258 => x"6e",
          6259 => x"2e",
          6260 => x"00",
          6261 => x"6c",
          6262 => x"30",
          6263 => x"2d",
          6264 => x"38",
          6265 => x"25",
          6266 => x"29",
          6267 => x"00",
          6268 => x"70",
          6269 => x"6d",
          6270 => x"0a",
          6271 => x"00",
          6272 => x"6d",
          6273 => x"74",
          6274 => x"00",
          6275 => x"58",
          6276 => x"32",
          6277 => x"00",
          6278 => x"0a",
          6279 => x"00",
          6280 => x"58",
          6281 => x"34",
          6282 => x"00",
          6283 => x"58",
          6284 => x"38",
          6285 => x"00",
          6286 => x"61",
          6287 => x"6e",
          6288 => x"6e",
          6289 => x"72",
          6290 => x"73",
          6291 => x"00",
          6292 => x"62",
          6293 => x"67",
          6294 => x"74",
          6295 => x"75",
          6296 => x"0a",
          6297 => x"00",
          6298 => x"61",
          6299 => x"64",
          6300 => x"72",
          6301 => x"69",
          6302 => x"00",
          6303 => x"62",
          6304 => x"67",
          6305 => x"72",
          6306 => x"69",
          6307 => x"00",
          6308 => x"63",
          6309 => x"6e",
          6310 => x"6f",
          6311 => x"40",
          6312 => x"38",
          6313 => x"2e",
          6314 => x"00",
          6315 => x"6c",
          6316 => x"20",
          6317 => x"65",
          6318 => x"25",
          6319 => x"20",
          6320 => x"0a",
          6321 => x"00",
          6322 => x"6c",
          6323 => x"74",
          6324 => x"65",
          6325 => x"6f",
          6326 => x"28",
          6327 => x"2e",
          6328 => x"00",
          6329 => x"74",
          6330 => x"69",
          6331 => x"61",
          6332 => x"69",
          6333 => x"69",
          6334 => x"2e",
          6335 => x"00",
          6336 => x"64",
          6337 => x"62",
          6338 => x"69",
          6339 => x"2e",
          6340 => x"00",
          6341 => x"00",
          6342 => x"00",
          6343 => x"5c",
          6344 => x"25",
          6345 => x"73",
          6346 => x"00",
          6347 => x"20",
          6348 => x"6d",
          6349 => x"2e",
          6350 => x"00",
          6351 => x"6e",
          6352 => x"2e",
          6353 => x"00",
          6354 => x"62",
          6355 => x"67",
          6356 => x"74",
          6357 => x"75",
          6358 => x"2e",
          6359 => x"00",
          6360 => x"00",
          6361 => x"00",
          6362 => x"ff",
          6363 => x"00",
          6364 => x"ff",
          6365 => x"00",
          6366 => x"ff",
          6367 => x"00",
          6368 => x"00",
          6369 => x"00",
          6370 => x"00",
          6371 => x"00",
          6372 => x"01",
          6373 => x"01",
          6374 => x"01",
          6375 => x"00",
          6376 => x"00",
          6377 => x"00",
          6378 => x"48",
          6379 => x"00",
          6380 => x"00",
          6381 => x"00",
          6382 => x"50",
          6383 => x"00",
          6384 => x"00",
          6385 => x"00",
          6386 => x"58",
          6387 => x"00",
          6388 => x"00",
          6389 => x"00",
          6390 => x"60",
          6391 => x"00",
          6392 => x"00",
          6393 => x"00",
          6394 => x"68",
          6395 => x"00",
          6396 => x"00",
          6397 => x"00",
          6398 => x"70",
          6399 => x"00",
          6400 => x"00",
          6401 => x"00",
          6402 => x"78",
          6403 => x"00",
          6404 => x"00",
          6405 => x"00",
          6406 => x"80",
          6407 => x"00",
          6408 => x"00",
          6409 => x"00",
          6410 => x"88",
          6411 => x"00",
          6412 => x"00",
          6413 => x"00",
          6414 => x"90",
          6415 => x"00",
          6416 => x"00",
          6417 => x"00",
          6418 => x"94",
          6419 => x"00",
          6420 => x"00",
          6421 => x"00",
          6422 => x"98",
          6423 => x"00",
          6424 => x"00",
          6425 => x"00",
          6426 => x"9c",
          6427 => x"00",
          6428 => x"00",
          6429 => x"00",
          6430 => x"a0",
          6431 => x"00",
          6432 => x"00",
          6433 => x"00",
          6434 => x"a4",
          6435 => x"00",
          6436 => x"00",
          6437 => x"00",
          6438 => x"a8",
          6439 => x"00",
          6440 => x"00",
          6441 => x"00",
          6442 => x"ac",
          6443 => x"00",
          6444 => x"00",
          6445 => x"00",
          6446 => x"b4",
          6447 => x"00",
          6448 => x"00",
          6449 => x"00",
          6450 => x"b8",
          6451 => x"00",
          6452 => x"00",
          6453 => x"00",
          6454 => x"c0",
          6455 => x"00",
          6456 => x"00",
          6457 => x"00",
          6458 => x"c8",
          6459 => x"00",
          6460 => x"00",
          6461 => x"00",
          6462 => x"d0",
          6463 => x"00",
          6464 => x"00",
          6465 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"90",
             1 => x"0b",
             2 => x"c6",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"90",
             9 => x"0b",
            10 => x"85",
            11 => x"90",
            12 => x"0b",
            13 => x"a7",
            14 => x"90",
            15 => x"0b",
            16 => x"c9",
            17 => x"90",
            18 => x"0b",
            19 => x"eb",
            20 => x"90",
            21 => x"0b",
            22 => x"8d",
            23 => x"90",
            24 => x"0b",
            25 => x"af",
            26 => x"90",
            27 => x"0b",
            28 => x"d1",
            29 => x"90",
            30 => x"0b",
            31 => x"f3",
            32 => x"90",
            33 => x"0b",
            34 => x"95",
            35 => x"90",
            36 => x"0b",
            37 => x"b7",
            38 => x"90",
            39 => x"0b",
            40 => x"d9",
            41 => x"90",
            42 => x"0b",
            43 => x"fb",
            44 => x"90",
            45 => x"0b",
            46 => x"9d",
            47 => x"90",
            48 => x"0b",
            49 => x"bf",
            50 => x"90",
            51 => x"0b",
            52 => x"e1",
            53 => x"90",
            54 => x"0b",
            55 => x"83",
            56 => x"90",
            57 => x"0b",
            58 => x"a5",
            59 => x"90",
            60 => x"0b",
            61 => x"c7",
            62 => x"90",
            63 => x"0b",
            64 => x"e9",
            65 => x"90",
            66 => x"0b",
            67 => x"8b",
            68 => x"90",
            69 => x"0b",
            70 => x"ad",
            71 => x"90",
            72 => x"0b",
            73 => x"cf",
            74 => x"90",
            75 => x"0b",
            76 => x"f1",
            77 => x"90",
            78 => x"0b",
            79 => x"93",
            80 => x"90",
            81 => x"0b",
            82 => x"b5",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"84",
           129 => x"ca",
           130 => x"95",
           131 => x"ca",
           132 => x"c0",
           133 => x"91",
           134 => x"90",
           135 => x"91",
           136 => x"88",
           137 => x"04",
           138 => x"0c",
           139 => x"2d",
           140 => x"08",
           141 => x"90",
           142 => x"94",
           143 => x"9c",
           144 => x"94",
           145 => x"80",
           146 => x"ca",
           147 => x"a6",
           148 => x"ca",
           149 => x"c0",
           150 => x"91",
           151 => x"90",
           152 => x"91",
           153 => x"88",
           154 => x"04",
           155 => x"0c",
           156 => x"2d",
           157 => x"08",
           158 => x"90",
           159 => x"94",
           160 => x"f5",
           161 => x"94",
           162 => x"80",
           163 => x"ca",
           164 => x"a9",
           165 => x"ca",
           166 => x"c0",
           167 => x"91",
           168 => x"90",
           169 => x"91",
           170 => x"88",
           171 => x"04",
           172 => x"0c",
           173 => x"2d",
           174 => x"08",
           175 => x"90",
           176 => x"94",
           177 => x"ba",
           178 => x"94",
           179 => x"80",
           180 => x"ca",
           181 => x"97",
           182 => x"ca",
           183 => x"c0",
           184 => x"91",
           185 => x"90",
           186 => x"91",
           187 => x"88",
           188 => x"04",
           189 => x"0c",
           190 => x"2d",
           191 => x"08",
           192 => x"90",
           193 => x"94",
           194 => x"be",
           195 => x"94",
           196 => x"80",
           197 => x"ca",
           198 => x"92",
           199 => x"ca",
           200 => x"c0",
           201 => x"91",
           202 => x"90",
           203 => x"91",
           204 => x"88",
           205 => x"04",
           206 => x"0c",
           207 => x"2d",
           208 => x"08",
           209 => x"90",
           210 => x"94",
           211 => x"81",
           212 => x"94",
           213 => x"80",
           214 => x"ca",
           215 => x"e3",
           216 => x"ca",
           217 => x"c0",
           218 => x"91",
           219 => x"90",
           220 => x"91",
           221 => x"88",
           222 => x"04",
           223 => x"0c",
           224 => x"2d",
           225 => x"08",
           226 => x"90",
           227 => x"94",
           228 => x"ef",
           229 => x"94",
           230 => x"80",
           231 => x"ca",
           232 => x"f1",
           233 => x"ca",
           234 => x"c0",
           235 => x"91",
           236 => x"90",
           237 => x"91",
           238 => x"88",
           239 => x"04",
           240 => x"0c",
           241 => x"2d",
           242 => x"08",
           243 => x"90",
           244 => x"94",
           245 => x"e3",
           246 => x"94",
           247 => x"80",
           248 => x"ca",
           249 => x"f8",
           250 => x"ca",
           251 => x"c0",
           252 => x"91",
           253 => x"90",
           254 => x"91",
           255 => x"88",
           256 => x"04",
           257 => x"0c",
           258 => x"2d",
           259 => x"08",
           260 => x"90",
           261 => x"94",
           262 => x"b7",
           263 => x"94",
           264 => x"80",
           265 => x"ca",
           266 => x"81",
           267 => x"ca",
           268 => x"c0",
           269 => x"91",
           270 => x"90",
           271 => x"91",
           272 => x"88",
           273 => x"04",
           274 => x"0c",
           275 => x"2d",
           276 => x"08",
           277 => x"90",
           278 => x"94",
           279 => x"f1",
           280 => x"94",
           281 => x"80",
           282 => x"ca",
           283 => x"f4",
           284 => x"ca",
           285 => x"c0",
           286 => x"91",
           287 => x"91",
           288 => x"91",
           289 => x"88",
           290 => x"04",
           291 => x"0c",
           292 => x"2d",
           293 => x"08",
           294 => x"90",
           295 => x"94",
           296 => x"f5",
           297 => x"94",
           298 => x"80",
           299 => x"ca",
           300 => x"db",
           301 => x"ca",
           302 => x"c0",
           303 => x"91",
           304 => x"91",
           305 => x"91",
           306 => x"88",
           307 => x"04",
           308 => x"0c",
           309 => x"2d",
           310 => x"08",
           311 => x"90",
           312 => x"94",
           313 => x"e0",
           314 => x"94",
           315 => x"80",
           316 => x"ca",
           317 => x"b0",
           318 => x"ca",
           319 => x"c0",
           320 => x"91",
           321 => x"90",
           322 => x"91",
           323 => x"88",
           324 => x"04",
           325 => x"0c",
           326 => x"2d",
           327 => x"08",
           328 => x"90",
           329 => x"94",
           330 => x"81",
           331 => x"94",
           332 => x"80",
           333 => x"ca",
           334 => x"97",
           335 => x"ca",
           336 => x"c0",
           337 => x"91",
           338 => x"91",
           339 => x"8e",
           340 => x"70",
           341 => x"0c",
           342 => x"8a",
           343 => x"84",
           344 => x"b2",
           345 => x"04",
           346 => x"08",
           347 => x"94",
           348 => x"0d",
           349 => x"ca",
           350 => x"05",
           351 => x"ca",
           352 => x"05",
           353 => x"c5",
           354 => x"88",
           355 => x"ca",
           356 => x"85",
           357 => x"ca",
           358 => x"91",
           359 => x"02",
           360 => x"0c",
           361 => x"81",
           362 => x"94",
           363 => x"08",
           364 => x"94",
           365 => x"08",
           366 => x"91",
           367 => x"70",
           368 => x"0c",
           369 => x"0d",
           370 => x"0c",
           371 => x"94",
           372 => x"ca",
           373 => x"3d",
           374 => x"91",
           375 => x"fc",
           376 => x"0b",
           377 => x"08",
           378 => x"91",
           379 => x"8c",
           380 => x"ca",
           381 => x"05",
           382 => x"38",
           383 => x"08",
           384 => x"80",
           385 => x"80",
           386 => x"94",
           387 => x"08",
           388 => x"91",
           389 => x"8c",
           390 => x"91",
           391 => x"8c",
           392 => x"ca",
           393 => x"05",
           394 => x"ca",
           395 => x"05",
           396 => x"39",
           397 => x"08",
           398 => x"80",
           399 => x"38",
           400 => x"08",
           401 => x"91",
           402 => x"88",
           403 => x"ad",
           404 => x"94",
           405 => x"08",
           406 => x"08",
           407 => x"31",
           408 => x"08",
           409 => x"91",
           410 => x"f8",
           411 => x"ca",
           412 => x"05",
           413 => x"ca",
           414 => x"05",
           415 => x"94",
           416 => x"08",
           417 => x"ca",
           418 => x"05",
           419 => x"94",
           420 => x"08",
           421 => x"ca",
           422 => x"05",
           423 => x"39",
           424 => x"08",
           425 => x"80",
           426 => x"91",
           427 => x"88",
           428 => x"91",
           429 => x"f4",
           430 => x"91",
           431 => x"94",
           432 => x"08",
           433 => x"94",
           434 => x"0c",
           435 => x"94",
           436 => x"08",
           437 => x"0c",
           438 => x"91",
           439 => x"04",
           440 => x"76",
           441 => x"8c",
           442 => x"33",
           443 => x"55",
           444 => x"8a",
           445 => x"06",
           446 => x"2e",
           447 => x"12",
           448 => x"2e",
           449 => x"73",
           450 => x"55",
           451 => x"52",
           452 => x"09",
           453 => x"38",
           454 => x"88",
           455 => x"0d",
           456 => x"88",
           457 => x"70",
           458 => x"07",
           459 => x"8f",
           460 => x"38",
           461 => x"84",
           462 => x"72",
           463 => x"05",
           464 => x"71",
           465 => x"53",
           466 => x"70",
           467 => x"0c",
           468 => x"71",
           469 => x"38",
           470 => x"90",
           471 => x"70",
           472 => x"0c",
           473 => x"71",
           474 => x"38",
           475 => x"8e",
           476 => x"0d",
           477 => x"72",
           478 => x"53",
           479 => x"93",
           480 => x"73",
           481 => x"54",
           482 => x"2e",
           483 => x"73",
           484 => x"71",
           485 => x"ff",
           486 => x"70",
           487 => x"38",
           488 => x"70",
           489 => x"81",
           490 => x"81",
           491 => x"71",
           492 => x"ff",
           493 => x"54",
           494 => x"38",
           495 => x"73",
           496 => x"75",
           497 => x"71",
           498 => x"ca",
           499 => x"52",
           500 => x"04",
           501 => x"f7",
           502 => x"14",
           503 => x"84",
           504 => x"06",
           505 => x"70",
           506 => x"14",
           507 => x"08",
           508 => x"71",
           509 => x"dc",
           510 => x"54",
           511 => x"39",
           512 => x"ca",
           513 => x"3d",
           514 => x"3d",
           515 => x"83",
           516 => x"2b",
           517 => x"3f",
           518 => x"08",
           519 => x"72",
           520 => x"54",
           521 => x"25",
           522 => x"91",
           523 => x"84",
           524 => x"fb",
           525 => x"70",
           526 => x"53",
           527 => x"2e",
           528 => x"71",
           529 => x"a0",
           530 => x"06",
           531 => x"12",
           532 => x"71",
           533 => x"81",
           534 => x"73",
           535 => x"ff",
           536 => x"55",
           537 => x"83",
           538 => x"70",
           539 => x"38",
           540 => x"73",
           541 => x"51",
           542 => x"09",
           543 => x"38",
           544 => x"81",
           545 => x"72",
           546 => x"51",
           547 => x"88",
           548 => x"0d",
           549 => x"0d",
           550 => x"08",
           551 => x"38",
           552 => x"05",
           553 => x"98",
           554 => x"ca",
           555 => x"38",
           556 => x"39",
           557 => x"91",
           558 => x"86",
           559 => x"fc",
           560 => x"82",
           561 => x"05",
           562 => x"52",
           563 => x"81",
           564 => x"13",
           565 => x"51",
           566 => x"9e",
           567 => x"38",
           568 => x"51",
           569 => x"97",
           570 => x"38",
           571 => x"51",
           572 => x"bb",
           573 => x"38",
           574 => x"51",
           575 => x"bb",
           576 => x"38",
           577 => x"55",
           578 => x"87",
           579 => x"d9",
           580 => x"22",
           581 => x"73",
           582 => x"80",
           583 => x"0b",
           584 => x"9c",
           585 => x"87",
           586 => x"0c",
           587 => x"87",
           588 => x"0c",
           589 => x"87",
           590 => x"0c",
           591 => x"87",
           592 => x"0c",
           593 => x"87",
           594 => x"0c",
           595 => x"87",
           596 => x"0c",
           597 => x"98",
           598 => x"87",
           599 => x"0c",
           600 => x"c0",
           601 => x"80",
           602 => x"ca",
           603 => x"3d",
           604 => x"3d",
           605 => x"87",
           606 => x"5d",
           607 => x"87",
           608 => x"08",
           609 => x"23",
           610 => x"b8",
           611 => x"82",
           612 => x"c0",
           613 => x"5a",
           614 => x"34",
           615 => x"b0",
           616 => x"84",
           617 => x"c0",
           618 => x"5a",
           619 => x"34",
           620 => x"a8",
           621 => x"86",
           622 => x"c0",
           623 => x"5c",
           624 => x"23",
           625 => x"a0",
           626 => x"8a",
           627 => x"7d",
           628 => x"ff",
           629 => x"7b",
           630 => x"06",
           631 => x"33",
           632 => x"33",
           633 => x"33",
           634 => x"33",
           635 => x"33",
           636 => x"ff",
           637 => x"91",
           638 => x"92",
           639 => x"3d",
           640 => x"3d",
           641 => x"05",
           642 => x"70",
           643 => x"52",
           644 => x"0b",
           645 => x"34",
           646 => x"04",
           647 => x"77",
           648 => x"c6",
           649 => x"81",
           650 => x"55",
           651 => x"94",
           652 => x"80",
           653 => x"87",
           654 => x"51",
           655 => x"96",
           656 => x"06",
           657 => x"70",
           658 => x"38",
           659 => x"70",
           660 => x"51",
           661 => x"72",
           662 => x"81",
           663 => x"70",
           664 => x"38",
           665 => x"70",
           666 => x"51",
           667 => x"38",
           668 => x"06",
           669 => x"94",
           670 => x"80",
           671 => x"87",
           672 => x"52",
           673 => x"75",
           674 => x"0c",
           675 => x"04",
           676 => x"02",
           677 => x"0b",
           678 => x"e0",
           679 => x"ff",
           680 => x"56",
           681 => x"84",
           682 => x"2e",
           683 => x"c0",
           684 => x"70",
           685 => x"2a",
           686 => x"53",
           687 => x"80",
           688 => x"71",
           689 => x"81",
           690 => x"70",
           691 => x"81",
           692 => x"06",
           693 => x"80",
           694 => x"71",
           695 => x"81",
           696 => x"70",
           697 => x"73",
           698 => x"51",
           699 => x"80",
           700 => x"2e",
           701 => x"c0",
           702 => x"75",
           703 => x"3d",
           704 => x"3d",
           705 => x"80",
           706 => x"81",
           707 => x"53",
           708 => x"2e",
           709 => x"71",
           710 => x"81",
           711 => x"91",
           712 => x"70",
           713 => x"59",
           714 => x"87",
           715 => x"51",
           716 => x"86",
           717 => x"94",
           718 => x"08",
           719 => x"70",
           720 => x"54",
           721 => x"2e",
           722 => x"91",
           723 => x"06",
           724 => x"d7",
           725 => x"32",
           726 => x"51",
           727 => x"2e",
           728 => x"93",
           729 => x"06",
           730 => x"ff",
           731 => x"81",
           732 => x"87",
           733 => x"52",
           734 => x"86",
           735 => x"94",
           736 => x"72",
           737 => x"74",
           738 => x"ff",
           739 => x"57",
           740 => x"38",
           741 => x"88",
           742 => x"0d",
           743 => x"0d",
           744 => x"c6",
           745 => x"81",
           746 => x"52",
           747 => x"84",
           748 => x"2e",
           749 => x"c0",
           750 => x"70",
           751 => x"2a",
           752 => x"51",
           753 => x"80",
           754 => x"71",
           755 => x"51",
           756 => x"80",
           757 => x"2e",
           758 => x"c0",
           759 => x"71",
           760 => x"ff",
           761 => x"88",
           762 => x"3d",
           763 => x"3d",
           764 => x"91",
           765 => x"70",
           766 => x"52",
           767 => x"94",
           768 => x"80",
           769 => x"87",
           770 => x"52",
           771 => x"82",
           772 => x"06",
           773 => x"ff",
           774 => x"2e",
           775 => x"81",
           776 => x"87",
           777 => x"52",
           778 => x"86",
           779 => x"94",
           780 => x"08",
           781 => x"70",
           782 => x"53",
           783 => x"ca",
           784 => x"3d",
           785 => x"3d",
           786 => x"9e",
           787 => x"9c",
           788 => x"51",
           789 => x"2e",
           790 => x"87",
           791 => x"08",
           792 => x"0c",
           793 => x"a0",
           794 => x"e8",
           795 => x"9e",
           796 => x"c6",
           797 => x"c0",
           798 => x"91",
           799 => x"87",
           800 => x"08",
           801 => x"0c",
           802 => x"98",
           803 => x"f8",
           804 => x"9e",
           805 => x"c6",
           806 => x"c0",
           807 => x"91",
           808 => x"87",
           809 => x"08",
           810 => x"0c",
           811 => x"80",
           812 => x"91",
           813 => x"87",
           814 => x"08",
           815 => x"0c",
           816 => x"c7",
           817 => x"0b",
           818 => x"88",
           819 => x"80",
           820 => x"52",
           821 => x"83",
           822 => x"71",
           823 => x"34",
           824 => x"c0",
           825 => x"70",
           826 => x"06",
           827 => x"70",
           828 => x"38",
           829 => x"91",
           830 => x"80",
           831 => x"9e",
           832 => x"80",
           833 => x"51",
           834 => x"80",
           835 => x"81",
           836 => x"c7",
           837 => x"0b",
           838 => x"88",
           839 => x"80",
           840 => x"52",
           841 => x"83",
           842 => x"71",
           843 => x"34",
           844 => x"c0",
           845 => x"70",
           846 => x"51",
           847 => x"80",
           848 => x"81",
           849 => x"c7",
           850 => x"0b",
           851 => x"88",
           852 => x"80",
           853 => x"52",
           854 => x"83",
           855 => x"71",
           856 => x"34",
           857 => x"c0",
           858 => x"70",
           859 => x"51",
           860 => x"80",
           861 => x"81",
           862 => x"c7",
           863 => x"0b",
           864 => x"88",
           865 => x"80",
           866 => x"52",
           867 => x"83",
           868 => x"71",
           869 => x"34",
           870 => x"88",
           871 => x"e0",
           872 => x"2c",
           873 => x"70",
           874 => x"34",
           875 => x"c0",
           876 => x"70",
           877 => x"52",
           878 => x"2e",
           879 => x"52",
           880 => x"9a",
           881 => x"87",
           882 => x"08",
           883 => x"51",
           884 => x"80",
           885 => x"81",
           886 => x"c7",
           887 => x"c0",
           888 => x"70",
           889 => x"51",
           890 => x"9c",
           891 => x"0d",
           892 => x"0d",
           893 => x"51",
           894 => x"91",
           895 => x"54",
           896 => x"88",
           897 => x"98",
           898 => x"3f",
           899 => x"51",
           900 => x"91",
           901 => x"54",
           902 => x"92",
           903 => x"e8",
           904 => x"c6",
           905 => x"91",
           906 => x"89",
           907 => x"c7",
           908 => x"73",
           909 => x"38",
           910 => x"08",
           911 => x"ec",
           912 => x"b4",
           913 => x"b9",
           914 => x"93",
           915 => x"8b",
           916 => x"94",
           917 => x"80",
           918 => x"91",
           919 => x"53",
           920 => x"08",
           921 => x"90",
           922 => x"3f",
           923 => x"33",
           924 => x"2e",
           925 => x"b5",
           926 => x"a1",
           927 => x"96",
           928 => x"80",
           929 => x"91",
           930 => x"83",
           931 => x"c7",
           932 => x"73",
           933 => x"38",
           934 => x"51",
           935 => x"91",
           936 => x"54",
           937 => x"8d",
           938 => x"99",
           939 => x"b5",
           940 => x"cd",
           941 => x"9a",
           942 => x"80",
           943 => x"91",
           944 => x"82",
           945 => x"c7",
           946 => x"73",
           947 => x"38",
           948 => x"33",
           949 => x"94",
           950 => x"3f",
           951 => x"51",
           952 => x"91",
           953 => x"52",
           954 => x"51",
           955 => x"91",
           956 => x"52",
           957 => x"51",
           958 => x"91",
           959 => x"52",
           960 => x"51",
           961 => x"91",
           962 => x"52",
           963 => x"51",
           964 => x"91",
           965 => x"52",
           966 => x"51",
           967 => x"85",
           968 => x"fe",
           969 => x"92",
           970 => x"05",
           971 => x"26",
           972 => x"84",
           973 => x"91",
           974 => x"52",
           975 => x"91",
           976 => x"9d",
           977 => x"8c",
           978 => x"91",
           979 => x"91",
           980 => x"9c",
           981 => x"91",
           982 => x"85",
           983 => x"a8",
           984 => x"3f",
           985 => x"04",
           986 => x"0c",
           987 => x"87",
           988 => x"0c",
           989 => x"0d",
           990 => x"84",
           991 => x"52",
           992 => x"70",
           993 => x"91",
           994 => x"72",
           995 => x"0d",
           996 => x"0d",
           997 => x"84",
           998 => x"c7",
           999 => x"80",
          1000 => x"09",
          1001 => x"a0",
          1002 => x"91",
          1003 => x"73",
          1004 => x"3d",
          1005 => x"c7",
          1006 => x"c0",
          1007 => x"04",
          1008 => x"02",
          1009 => x"53",
          1010 => x"09",
          1011 => x"38",
          1012 => x"3f",
          1013 => x"08",
          1014 => x"2e",
          1015 => x"72",
          1016 => x"a0",
          1017 => x"91",
          1018 => x"8f",
          1019 => x"98",
          1020 => x"80",
          1021 => x"72",
          1022 => x"84",
          1023 => x"fe",
          1024 => x"97",
          1025 => x"ca",
          1026 => x"91",
          1027 => x"54",
          1028 => x"3f",
          1029 => x"98",
          1030 => x"0d",
          1031 => x"0d",
          1032 => x"33",
          1033 => x"06",
          1034 => x"80",
          1035 => x"72",
          1036 => x"51",
          1037 => x"ff",
          1038 => x"39",
          1039 => x"04",
          1040 => x"77",
          1041 => x"08",
          1042 => x"98",
          1043 => x"73",
          1044 => x"ff",
          1045 => x"71",
          1046 => x"38",
          1047 => x"06",
          1048 => x"54",
          1049 => x"e7",
          1050 => x"ca",
          1051 => x"3d",
          1052 => x"3d",
          1053 => x"59",
          1054 => x"81",
          1055 => x"56",
          1056 => x"84",
          1057 => x"a5",
          1058 => x"06",
          1059 => x"80",
          1060 => x"81",
          1061 => x"58",
          1062 => x"b0",
          1063 => x"06",
          1064 => x"5a",
          1065 => x"ad",
          1066 => x"06",
          1067 => x"5a",
          1068 => x"05",
          1069 => x"75",
          1070 => x"81",
          1071 => x"77",
          1072 => x"08",
          1073 => x"05",
          1074 => x"5d",
          1075 => x"39",
          1076 => x"72",
          1077 => x"38",
          1078 => x"7b",
          1079 => x"05",
          1080 => x"70",
          1081 => x"33",
          1082 => x"39",
          1083 => x"32",
          1084 => x"72",
          1085 => x"78",
          1086 => x"70",
          1087 => x"07",
          1088 => x"07",
          1089 => x"51",
          1090 => x"80",
          1091 => x"79",
          1092 => x"70",
          1093 => x"33",
          1094 => x"80",
          1095 => x"38",
          1096 => x"e0",
          1097 => x"38",
          1098 => x"81",
          1099 => x"53",
          1100 => x"2e",
          1101 => x"73",
          1102 => x"a2",
          1103 => x"c3",
          1104 => x"38",
          1105 => x"24",
          1106 => x"80",
          1107 => x"8c",
          1108 => x"39",
          1109 => x"2e",
          1110 => x"81",
          1111 => x"80",
          1112 => x"80",
          1113 => x"d5",
          1114 => x"73",
          1115 => x"8e",
          1116 => x"39",
          1117 => x"2e",
          1118 => x"80",
          1119 => x"84",
          1120 => x"56",
          1121 => x"74",
          1122 => x"72",
          1123 => x"38",
          1124 => x"15",
          1125 => x"54",
          1126 => x"38",
          1127 => x"56",
          1128 => x"81",
          1129 => x"72",
          1130 => x"38",
          1131 => x"90",
          1132 => x"06",
          1133 => x"2e",
          1134 => x"51",
          1135 => x"74",
          1136 => x"53",
          1137 => x"fd",
          1138 => x"51",
          1139 => x"ef",
          1140 => x"19",
          1141 => x"53",
          1142 => x"39",
          1143 => x"39",
          1144 => x"39",
          1145 => x"39",
          1146 => x"39",
          1147 => x"d0",
          1148 => x"39",
          1149 => x"70",
          1150 => x"53",
          1151 => x"88",
          1152 => x"19",
          1153 => x"39",
          1154 => x"54",
          1155 => x"74",
          1156 => x"70",
          1157 => x"07",
          1158 => x"55",
          1159 => x"80",
          1160 => x"72",
          1161 => x"38",
          1162 => x"90",
          1163 => x"80",
          1164 => x"5e",
          1165 => x"74",
          1166 => x"3f",
          1167 => x"08",
          1168 => x"7c",
          1169 => x"54",
          1170 => x"91",
          1171 => x"55",
          1172 => x"92",
          1173 => x"53",
          1174 => x"2e",
          1175 => x"14",
          1176 => x"ff",
          1177 => x"14",
          1178 => x"70",
          1179 => x"34",
          1180 => x"30",
          1181 => x"9f",
          1182 => x"57",
          1183 => x"85",
          1184 => x"b1",
          1185 => x"2a",
          1186 => x"51",
          1187 => x"2e",
          1188 => x"3d",
          1189 => x"05",
          1190 => x"34",
          1191 => x"76",
          1192 => x"54",
          1193 => x"72",
          1194 => x"54",
          1195 => x"70",
          1196 => x"56",
          1197 => x"81",
          1198 => x"7b",
          1199 => x"73",
          1200 => x"3f",
          1201 => x"53",
          1202 => x"74",
          1203 => x"53",
          1204 => x"eb",
          1205 => x"77",
          1206 => x"53",
          1207 => x"14",
          1208 => x"54",
          1209 => x"3f",
          1210 => x"74",
          1211 => x"53",
          1212 => x"fb",
          1213 => x"51",
          1214 => x"ef",
          1215 => x"0d",
          1216 => x"0d",
          1217 => x"70",
          1218 => x"08",
          1219 => x"51",
          1220 => x"85",
          1221 => x"fe",
          1222 => x"91",
          1223 => x"85",
          1224 => x"52",
          1225 => x"ca",
          1226 => x"a0",
          1227 => x"73",
          1228 => x"91",
          1229 => x"84",
          1230 => x"fd",
          1231 => x"ca",
          1232 => x"91",
          1233 => x"87",
          1234 => x"53",
          1235 => x"fa",
          1236 => x"91",
          1237 => x"85",
          1238 => x"fb",
          1239 => x"79",
          1240 => x"08",
          1241 => x"57",
          1242 => x"71",
          1243 => x"e0",
          1244 => x"9c",
          1245 => x"2d",
          1246 => x"08",
          1247 => x"53",
          1248 => x"80",
          1249 => x"8d",
          1250 => x"72",
          1251 => x"30",
          1252 => x"51",
          1253 => x"80",
          1254 => x"71",
          1255 => x"38",
          1256 => x"97",
          1257 => x"25",
          1258 => x"16",
          1259 => x"25",
          1260 => x"14",
          1261 => x"34",
          1262 => x"72",
          1263 => x"3f",
          1264 => x"73",
          1265 => x"72",
          1266 => x"f7",
          1267 => x"53",
          1268 => x"88",
          1269 => x"0d",
          1270 => x"0d",
          1271 => x"08",
          1272 => x"9c",
          1273 => x"76",
          1274 => x"ef",
          1275 => x"ca",
          1276 => x"3d",
          1277 => x"3d",
          1278 => x"5a",
          1279 => x"7a",
          1280 => x"08",
          1281 => x"53",
          1282 => x"09",
          1283 => x"38",
          1284 => x"0c",
          1285 => x"ad",
          1286 => x"06",
          1287 => x"76",
          1288 => x"0c",
          1289 => x"33",
          1290 => x"73",
          1291 => x"81",
          1292 => x"38",
          1293 => x"05",
          1294 => x"08",
          1295 => x"53",
          1296 => x"2e",
          1297 => x"57",
          1298 => x"2e",
          1299 => x"39",
          1300 => x"13",
          1301 => x"08",
          1302 => x"53",
          1303 => x"55",
          1304 => x"80",
          1305 => x"14",
          1306 => x"88",
          1307 => x"27",
          1308 => x"eb",
          1309 => x"53",
          1310 => x"89",
          1311 => x"38",
          1312 => x"55",
          1313 => x"8a",
          1314 => x"a0",
          1315 => x"c2",
          1316 => x"74",
          1317 => x"e0",
          1318 => x"ff",
          1319 => x"d0",
          1320 => x"ff",
          1321 => x"90",
          1322 => x"38",
          1323 => x"81",
          1324 => x"53",
          1325 => x"ca",
          1326 => x"27",
          1327 => x"77",
          1328 => x"08",
          1329 => x"0c",
          1330 => x"33",
          1331 => x"ff",
          1332 => x"80",
          1333 => x"74",
          1334 => x"79",
          1335 => x"74",
          1336 => x"0c",
          1337 => x"04",
          1338 => x"7a",
          1339 => x"80",
          1340 => x"58",
          1341 => x"33",
          1342 => x"a0",
          1343 => x"06",
          1344 => x"13",
          1345 => x"39",
          1346 => x"09",
          1347 => x"38",
          1348 => x"11",
          1349 => x"08",
          1350 => x"54",
          1351 => x"2e",
          1352 => x"80",
          1353 => x"08",
          1354 => x"0c",
          1355 => x"33",
          1356 => x"80",
          1357 => x"38",
          1358 => x"80",
          1359 => x"38",
          1360 => x"57",
          1361 => x"0c",
          1362 => x"33",
          1363 => x"39",
          1364 => x"74",
          1365 => x"38",
          1366 => x"80",
          1367 => x"89",
          1368 => x"38",
          1369 => x"d0",
          1370 => x"55",
          1371 => x"80",
          1372 => x"39",
          1373 => x"d9",
          1374 => x"80",
          1375 => x"27",
          1376 => x"80",
          1377 => x"89",
          1378 => x"70",
          1379 => x"55",
          1380 => x"70",
          1381 => x"55",
          1382 => x"27",
          1383 => x"14",
          1384 => x"06",
          1385 => x"74",
          1386 => x"73",
          1387 => x"38",
          1388 => x"14",
          1389 => x"05",
          1390 => x"08",
          1391 => x"54",
          1392 => x"39",
          1393 => x"84",
          1394 => x"55",
          1395 => x"81",
          1396 => x"ca",
          1397 => x"3d",
          1398 => x"3d",
          1399 => x"05",
          1400 => x"52",
          1401 => x"87",
          1402 => x"a4",
          1403 => x"71",
          1404 => x"0c",
          1405 => x"04",
          1406 => x"02",
          1407 => x"02",
          1408 => x"05",
          1409 => x"83",
          1410 => x"26",
          1411 => x"72",
          1412 => x"c0",
          1413 => x"53",
          1414 => x"74",
          1415 => x"38",
          1416 => x"73",
          1417 => x"c0",
          1418 => x"51",
          1419 => x"85",
          1420 => x"98",
          1421 => x"52",
          1422 => x"82",
          1423 => x"70",
          1424 => x"38",
          1425 => x"8c",
          1426 => x"ec",
          1427 => x"fc",
          1428 => x"52",
          1429 => x"87",
          1430 => x"08",
          1431 => x"2e",
          1432 => x"91",
          1433 => x"34",
          1434 => x"13",
          1435 => x"91",
          1436 => x"86",
          1437 => x"f3",
          1438 => x"62",
          1439 => x"05",
          1440 => x"57",
          1441 => x"83",
          1442 => x"fe",
          1443 => x"ca",
          1444 => x"06",
          1445 => x"71",
          1446 => x"71",
          1447 => x"2b",
          1448 => x"80",
          1449 => x"92",
          1450 => x"c0",
          1451 => x"41",
          1452 => x"5a",
          1453 => x"87",
          1454 => x"0c",
          1455 => x"84",
          1456 => x"08",
          1457 => x"70",
          1458 => x"53",
          1459 => x"2e",
          1460 => x"08",
          1461 => x"70",
          1462 => x"34",
          1463 => x"80",
          1464 => x"53",
          1465 => x"2e",
          1466 => x"53",
          1467 => x"26",
          1468 => x"80",
          1469 => x"87",
          1470 => x"08",
          1471 => x"38",
          1472 => x"8c",
          1473 => x"80",
          1474 => x"78",
          1475 => x"99",
          1476 => x"0c",
          1477 => x"8c",
          1478 => x"08",
          1479 => x"51",
          1480 => x"38",
          1481 => x"8d",
          1482 => x"17",
          1483 => x"81",
          1484 => x"53",
          1485 => x"2e",
          1486 => x"fc",
          1487 => x"52",
          1488 => x"7d",
          1489 => x"ed",
          1490 => x"80",
          1491 => x"71",
          1492 => x"38",
          1493 => x"53",
          1494 => x"88",
          1495 => x"0d",
          1496 => x"0d",
          1497 => x"02",
          1498 => x"05",
          1499 => x"58",
          1500 => x"80",
          1501 => x"fc",
          1502 => x"ca",
          1503 => x"06",
          1504 => x"71",
          1505 => x"81",
          1506 => x"38",
          1507 => x"2b",
          1508 => x"80",
          1509 => x"92",
          1510 => x"c0",
          1511 => x"40",
          1512 => x"5a",
          1513 => x"c0",
          1514 => x"76",
          1515 => x"76",
          1516 => x"75",
          1517 => x"2a",
          1518 => x"51",
          1519 => x"80",
          1520 => x"7a",
          1521 => x"5c",
          1522 => x"81",
          1523 => x"81",
          1524 => x"06",
          1525 => x"80",
          1526 => x"87",
          1527 => x"08",
          1528 => x"38",
          1529 => x"8c",
          1530 => x"80",
          1531 => x"77",
          1532 => x"99",
          1533 => x"0c",
          1534 => x"8c",
          1535 => x"08",
          1536 => x"51",
          1537 => x"38",
          1538 => x"8d",
          1539 => x"70",
          1540 => x"84",
          1541 => x"5b",
          1542 => x"2e",
          1543 => x"fc",
          1544 => x"52",
          1545 => x"7d",
          1546 => x"f8",
          1547 => x"80",
          1548 => x"71",
          1549 => x"38",
          1550 => x"53",
          1551 => x"88",
          1552 => x"0d",
          1553 => x"0d",
          1554 => x"05",
          1555 => x"02",
          1556 => x"05",
          1557 => x"54",
          1558 => x"fe",
          1559 => x"88",
          1560 => x"53",
          1561 => x"80",
          1562 => x"0b",
          1563 => x"8c",
          1564 => x"71",
          1565 => x"dc",
          1566 => x"24",
          1567 => x"84",
          1568 => x"92",
          1569 => x"54",
          1570 => x"8d",
          1571 => x"39",
          1572 => x"80",
          1573 => x"cb",
          1574 => x"70",
          1575 => x"81",
          1576 => x"52",
          1577 => x"8a",
          1578 => x"98",
          1579 => x"71",
          1580 => x"c0",
          1581 => x"52",
          1582 => x"81",
          1583 => x"c0",
          1584 => x"53",
          1585 => x"82",
          1586 => x"71",
          1587 => x"39",
          1588 => x"39",
          1589 => x"77",
          1590 => x"81",
          1591 => x"72",
          1592 => x"84",
          1593 => x"73",
          1594 => x"0c",
          1595 => x"04",
          1596 => x"74",
          1597 => x"71",
          1598 => x"2b",
          1599 => x"88",
          1600 => x"84",
          1601 => x"fd",
          1602 => x"83",
          1603 => x"12",
          1604 => x"2b",
          1605 => x"07",
          1606 => x"70",
          1607 => x"2b",
          1608 => x"07",
          1609 => x"0c",
          1610 => x"56",
          1611 => x"3d",
          1612 => x"3d",
          1613 => x"84",
          1614 => x"22",
          1615 => x"72",
          1616 => x"54",
          1617 => x"2a",
          1618 => x"34",
          1619 => x"04",
          1620 => x"73",
          1621 => x"70",
          1622 => x"05",
          1623 => x"88",
          1624 => x"72",
          1625 => x"54",
          1626 => x"2a",
          1627 => x"70",
          1628 => x"34",
          1629 => x"51",
          1630 => x"83",
          1631 => x"fe",
          1632 => x"75",
          1633 => x"51",
          1634 => x"92",
          1635 => x"81",
          1636 => x"73",
          1637 => x"55",
          1638 => x"51",
          1639 => x"3d",
          1640 => x"3d",
          1641 => x"76",
          1642 => x"72",
          1643 => x"05",
          1644 => x"11",
          1645 => x"38",
          1646 => x"04",
          1647 => x"78",
          1648 => x"56",
          1649 => x"81",
          1650 => x"74",
          1651 => x"56",
          1652 => x"31",
          1653 => x"52",
          1654 => x"80",
          1655 => x"71",
          1656 => x"38",
          1657 => x"88",
          1658 => x"0d",
          1659 => x"0d",
          1660 => x"51",
          1661 => x"73",
          1662 => x"81",
          1663 => x"33",
          1664 => x"38",
          1665 => x"ca",
          1666 => x"3d",
          1667 => x"0b",
          1668 => x"0c",
          1669 => x"91",
          1670 => x"04",
          1671 => x"7b",
          1672 => x"83",
          1673 => x"5a",
          1674 => x"80",
          1675 => x"54",
          1676 => x"53",
          1677 => x"53",
          1678 => x"52",
          1679 => x"3f",
          1680 => x"08",
          1681 => x"81",
          1682 => x"91",
          1683 => x"83",
          1684 => x"16",
          1685 => x"18",
          1686 => x"18",
          1687 => x"58",
          1688 => x"9f",
          1689 => x"33",
          1690 => x"2e",
          1691 => x"93",
          1692 => x"76",
          1693 => x"52",
          1694 => x"51",
          1695 => x"83",
          1696 => x"79",
          1697 => x"0c",
          1698 => x"04",
          1699 => x"78",
          1700 => x"80",
          1701 => x"17",
          1702 => x"38",
          1703 => x"fc",
          1704 => x"88",
          1705 => x"ca",
          1706 => x"38",
          1707 => x"53",
          1708 => x"81",
          1709 => x"f7",
          1710 => x"ca",
          1711 => x"2e",
          1712 => x"55",
          1713 => x"b0",
          1714 => x"91",
          1715 => x"88",
          1716 => x"f8",
          1717 => x"70",
          1718 => x"c0",
          1719 => x"88",
          1720 => x"ca",
          1721 => x"91",
          1722 => x"55",
          1723 => x"09",
          1724 => x"f0",
          1725 => x"33",
          1726 => x"2e",
          1727 => x"80",
          1728 => x"80",
          1729 => x"88",
          1730 => x"17",
          1731 => x"fd",
          1732 => x"d4",
          1733 => x"b2",
          1734 => x"96",
          1735 => x"85",
          1736 => x"75",
          1737 => x"3f",
          1738 => x"e4",
          1739 => x"98",
          1740 => x"9c",
          1741 => x"08",
          1742 => x"17",
          1743 => x"3f",
          1744 => x"52",
          1745 => x"51",
          1746 => x"a0",
          1747 => x"05",
          1748 => x"0c",
          1749 => x"75",
          1750 => x"33",
          1751 => x"3f",
          1752 => x"34",
          1753 => x"52",
          1754 => x"51",
          1755 => x"91",
          1756 => x"80",
          1757 => x"81",
          1758 => x"ca",
          1759 => x"3d",
          1760 => x"3d",
          1761 => x"1a",
          1762 => x"fe",
          1763 => x"54",
          1764 => x"73",
          1765 => x"8a",
          1766 => x"71",
          1767 => x"08",
          1768 => x"75",
          1769 => x"0c",
          1770 => x"04",
          1771 => x"7a",
          1772 => x"56",
          1773 => x"77",
          1774 => x"38",
          1775 => x"08",
          1776 => x"38",
          1777 => x"54",
          1778 => x"2e",
          1779 => x"72",
          1780 => x"38",
          1781 => x"8d",
          1782 => x"39",
          1783 => x"81",
          1784 => x"b6",
          1785 => x"2a",
          1786 => x"2a",
          1787 => x"05",
          1788 => x"55",
          1789 => x"91",
          1790 => x"81",
          1791 => x"83",
          1792 => x"b4",
          1793 => x"17",
          1794 => x"a4",
          1795 => x"55",
          1796 => x"57",
          1797 => x"3f",
          1798 => x"08",
          1799 => x"74",
          1800 => x"14",
          1801 => x"70",
          1802 => x"07",
          1803 => x"71",
          1804 => x"52",
          1805 => x"72",
          1806 => x"75",
          1807 => x"58",
          1808 => x"76",
          1809 => x"15",
          1810 => x"73",
          1811 => x"3f",
          1812 => x"08",
          1813 => x"76",
          1814 => x"06",
          1815 => x"05",
          1816 => x"3f",
          1817 => x"08",
          1818 => x"06",
          1819 => x"76",
          1820 => x"15",
          1821 => x"73",
          1822 => x"3f",
          1823 => x"08",
          1824 => x"82",
          1825 => x"06",
          1826 => x"05",
          1827 => x"3f",
          1828 => x"08",
          1829 => x"58",
          1830 => x"58",
          1831 => x"88",
          1832 => x"0d",
          1833 => x"0d",
          1834 => x"5a",
          1835 => x"59",
          1836 => x"82",
          1837 => x"98",
          1838 => x"82",
          1839 => x"33",
          1840 => x"2e",
          1841 => x"72",
          1842 => x"38",
          1843 => x"8d",
          1844 => x"39",
          1845 => x"81",
          1846 => x"f7",
          1847 => x"2a",
          1848 => x"2a",
          1849 => x"05",
          1850 => x"55",
          1851 => x"91",
          1852 => x"59",
          1853 => x"08",
          1854 => x"74",
          1855 => x"16",
          1856 => x"16",
          1857 => x"59",
          1858 => x"53",
          1859 => x"8f",
          1860 => x"2b",
          1861 => x"74",
          1862 => x"71",
          1863 => x"72",
          1864 => x"0b",
          1865 => x"74",
          1866 => x"17",
          1867 => x"75",
          1868 => x"3f",
          1869 => x"08",
          1870 => x"88",
          1871 => x"38",
          1872 => x"06",
          1873 => x"78",
          1874 => x"54",
          1875 => x"77",
          1876 => x"33",
          1877 => x"71",
          1878 => x"51",
          1879 => x"34",
          1880 => x"76",
          1881 => x"17",
          1882 => x"75",
          1883 => x"3f",
          1884 => x"08",
          1885 => x"88",
          1886 => x"38",
          1887 => x"ff",
          1888 => x"10",
          1889 => x"76",
          1890 => x"51",
          1891 => x"be",
          1892 => x"2a",
          1893 => x"05",
          1894 => x"f9",
          1895 => x"ca",
          1896 => x"91",
          1897 => x"ab",
          1898 => x"0a",
          1899 => x"2b",
          1900 => x"70",
          1901 => x"70",
          1902 => x"54",
          1903 => x"91",
          1904 => x"8f",
          1905 => x"07",
          1906 => x"f7",
          1907 => x"0b",
          1908 => x"78",
          1909 => x"0c",
          1910 => x"04",
          1911 => x"7a",
          1912 => x"08",
          1913 => x"59",
          1914 => x"a4",
          1915 => x"17",
          1916 => x"38",
          1917 => x"aa",
          1918 => x"73",
          1919 => x"fd",
          1920 => x"ca",
          1921 => x"91",
          1922 => x"80",
          1923 => x"39",
          1924 => x"eb",
          1925 => x"80",
          1926 => x"ca",
          1927 => x"80",
          1928 => x"52",
          1929 => x"84",
          1930 => x"88",
          1931 => x"ca",
          1932 => x"2e",
          1933 => x"91",
          1934 => x"81",
          1935 => x"91",
          1936 => x"ff",
          1937 => x"80",
          1938 => x"75",
          1939 => x"3f",
          1940 => x"08",
          1941 => x"16",
          1942 => x"90",
          1943 => x"55",
          1944 => x"27",
          1945 => x"15",
          1946 => x"84",
          1947 => x"07",
          1948 => x"17",
          1949 => x"76",
          1950 => x"a6",
          1951 => x"73",
          1952 => x"0c",
          1953 => x"04",
          1954 => x"7c",
          1955 => x"59",
          1956 => x"95",
          1957 => x"08",
          1958 => x"2e",
          1959 => x"17",
          1960 => x"b2",
          1961 => x"ae",
          1962 => x"7a",
          1963 => x"3f",
          1964 => x"91",
          1965 => x"27",
          1966 => x"91",
          1967 => x"55",
          1968 => x"08",
          1969 => x"d2",
          1970 => x"08",
          1971 => x"08",
          1972 => x"38",
          1973 => x"17",
          1974 => x"54",
          1975 => x"82",
          1976 => x"7a",
          1977 => x"06",
          1978 => x"81",
          1979 => x"17",
          1980 => x"83",
          1981 => x"75",
          1982 => x"f9",
          1983 => x"59",
          1984 => x"08",
          1985 => x"81",
          1986 => x"91",
          1987 => x"59",
          1988 => x"08",
          1989 => x"70",
          1990 => x"25",
          1991 => x"91",
          1992 => x"54",
          1993 => x"55",
          1994 => x"38",
          1995 => x"08",
          1996 => x"38",
          1997 => x"54",
          1998 => x"90",
          1999 => x"18",
          2000 => x"38",
          2001 => x"39",
          2002 => x"38",
          2003 => x"16",
          2004 => x"08",
          2005 => x"38",
          2006 => x"78",
          2007 => x"38",
          2008 => x"51",
          2009 => x"91",
          2010 => x"80",
          2011 => x"80",
          2012 => x"88",
          2013 => x"09",
          2014 => x"38",
          2015 => x"08",
          2016 => x"88",
          2017 => x"30",
          2018 => x"80",
          2019 => x"07",
          2020 => x"55",
          2021 => x"38",
          2022 => x"09",
          2023 => x"ae",
          2024 => x"80",
          2025 => x"53",
          2026 => x"51",
          2027 => x"91",
          2028 => x"91",
          2029 => x"30",
          2030 => x"88",
          2031 => x"25",
          2032 => x"79",
          2033 => x"38",
          2034 => x"8f",
          2035 => x"79",
          2036 => x"f9",
          2037 => x"ca",
          2038 => x"74",
          2039 => x"8c",
          2040 => x"17",
          2041 => x"90",
          2042 => x"54",
          2043 => x"86",
          2044 => x"90",
          2045 => x"17",
          2046 => x"54",
          2047 => x"34",
          2048 => x"56",
          2049 => x"90",
          2050 => x"80",
          2051 => x"91",
          2052 => x"55",
          2053 => x"56",
          2054 => x"91",
          2055 => x"8c",
          2056 => x"f8",
          2057 => x"70",
          2058 => x"f0",
          2059 => x"88",
          2060 => x"56",
          2061 => x"08",
          2062 => x"7b",
          2063 => x"f6",
          2064 => x"ca",
          2065 => x"ca",
          2066 => x"17",
          2067 => x"80",
          2068 => x"b4",
          2069 => x"57",
          2070 => x"77",
          2071 => x"81",
          2072 => x"15",
          2073 => x"78",
          2074 => x"81",
          2075 => x"53",
          2076 => x"15",
          2077 => x"e9",
          2078 => x"88",
          2079 => x"df",
          2080 => x"22",
          2081 => x"30",
          2082 => x"70",
          2083 => x"51",
          2084 => x"91",
          2085 => x"8a",
          2086 => x"f8",
          2087 => x"7c",
          2088 => x"56",
          2089 => x"80",
          2090 => x"f1",
          2091 => x"06",
          2092 => x"e9",
          2093 => x"18",
          2094 => x"08",
          2095 => x"38",
          2096 => x"82",
          2097 => x"38",
          2098 => x"54",
          2099 => x"74",
          2100 => x"82",
          2101 => x"22",
          2102 => x"79",
          2103 => x"38",
          2104 => x"98",
          2105 => x"cd",
          2106 => x"22",
          2107 => x"54",
          2108 => x"26",
          2109 => x"52",
          2110 => x"b0",
          2111 => x"88",
          2112 => x"ca",
          2113 => x"2e",
          2114 => x"0b",
          2115 => x"08",
          2116 => x"98",
          2117 => x"ca",
          2118 => x"85",
          2119 => x"bd",
          2120 => x"31",
          2121 => x"73",
          2122 => x"f4",
          2123 => x"ca",
          2124 => x"18",
          2125 => x"18",
          2126 => x"08",
          2127 => x"72",
          2128 => x"38",
          2129 => x"58",
          2130 => x"89",
          2131 => x"18",
          2132 => x"ff",
          2133 => x"05",
          2134 => x"80",
          2135 => x"ca",
          2136 => x"3d",
          2137 => x"3d",
          2138 => x"08",
          2139 => x"a0",
          2140 => x"54",
          2141 => x"77",
          2142 => x"80",
          2143 => x"0c",
          2144 => x"53",
          2145 => x"80",
          2146 => x"38",
          2147 => x"06",
          2148 => x"b5",
          2149 => x"98",
          2150 => x"14",
          2151 => x"92",
          2152 => x"2a",
          2153 => x"56",
          2154 => x"26",
          2155 => x"80",
          2156 => x"16",
          2157 => x"77",
          2158 => x"53",
          2159 => x"38",
          2160 => x"51",
          2161 => x"91",
          2162 => x"53",
          2163 => x"0b",
          2164 => x"08",
          2165 => x"38",
          2166 => x"ca",
          2167 => x"2e",
          2168 => x"98",
          2169 => x"ca",
          2170 => x"80",
          2171 => x"8a",
          2172 => x"15",
          2173 => x"80",
          2174 => x"14",
          2175 => x"51",
          2176 => x"91",
          2177 => x"53",
          2178 => x"ca",
          2179 => x"2e",
          2180 => x"82",
          2181 => x"88",
          2182 => x"ba",
          2183 => x"91",
          2184 => x"ff",
          2185 => x"91",
          2186 => x"52",
          2187 => x"f3",
          2188 => x"88",
          2189 => x"72",
          2190 => x"72",
          2191 => x"f2",
          2192 => x"ca",
          2193 => x"15",
          2194 => x"15",
          2195 => x"b4",
          2196 => x"0c",
          2197 => x"91",
          2198 => x"8a",
          2199 => x"f7",
          2200 => x"7d",
          2201 => x"5b",
          2202 => x"76",
          2203 => x"3f",
          2204 => x"08",
          2205 => x"88",
          2206 => x"38",
          2207 => x"08",
          2208 => x"08",
          2209 => x"f0",
          2210 => x"ca",
          2211 => x"91",
          2212 => x"80",
          2213 => x"ca",
          2214 => x"18",
          2215 => x"51",
          2216 => x"81",
          2217 => x"81",
          2218 => x"81",
          2219 => x"88",
          2220 => x"83",
          2221 => x"77",
          2222 => x"72",
          2223 => x"38",
          2224 => x"75",
          2225 => x"81",
          2226 => x"a5",
          2227 => x"88",
          2228 => x"52",
          2229 => x"8e",
          2230 => x"88",
          2231 => x"ca",
          2232 => x"2e",
          2233 => x"73",
          2234 => x"81",
          2235 => x"87",
          2236 => x"ca",
          2237 => x"3d",
          2238 => x"3d",
          2239 => x"11",
          2240 => x"ec",
          2241 => x"88",
          2242 => x"ff",
          2243 => x"33",
          2244 => x"71",
          2245 => x"81",
          2246 => x"94",
          2247 => x"d0",
          2248 => x"88",
          2249 => x"73",
          2250 => x"91",
          2251 => x"85",
          2252 => x"fc",
          2253 => x"79",
          2254 => x"ff",
          2255 => x"12",
          2256 => x"eb",
          2257 => x"70",
          2258 => x"72",
          2259 => x"81",
          2260 => x"73",
          2261 => x"94",
          2262 => x"d6",
          2263 => x"0d",
          2264 => x"0d",
          2265 => x"55",
          2266 => x"5a",
          2267 => x"08",
          2268 => x"8a",
          2269 => x"08",
          2270 => x"ee",
          2271 => x"ca",
          2272 => x"91",
          2273 => x"80",
          2274 => x"15",
          2275 => x"55",
          2276 => x"38",
          2277 => x"e6",
          2278 => x"33",
          2279 => x"70",
          2280 => x"58",
          2281 => x"86",
          2282 => x"ca",
          2283 => x"73",
          2284 => x"83",
          2285 => x"73",
          2286 => x"38",
          2287 => x"06",
          2288 => x"80",
          2289 => x"75",
          2290 => x"38",
          2291 => x"08",
          2292 => x"54",
          2293 => x"2e",
          2294 => x"83",
          2295 => x"73",
          2296 => x"38",
          2297 => x"51",
          2298 => x"91",
          2299 => x"58",
          2300 => x"08",
          2301 => x"15",
          2302 => x"38",
          2303 => x"0b",
          2304 => x"77",
          2305 => x"0c",
          2306 => x"04",
          2307 => x"77",
          2308 => x"54",
          2309 => x"51",
          2310 => x"91",
          2311 => x"55",
          2312 => x"08",
          2313 => x"14",
          2314 => x"51",
          2315 => x"91",
          2316 => x"55",
          2317 => x"08",
          2318 => x"53",
          2319 => x"08",
          2320 => x"08",
          2321 => x"3f",
          2322 => x"14",
          2323 => x"08",
          2324 => x"3f",
          2325 => x"17",
          2326 => x"ca",
          2327 => x"3d",
          2328 => x"3d",
          2329 => x"08",
          2330 => x"54",
          2331 => x"53",
          2332 => x"91",
          2333 => x"8d",
          2334 => x"08",
          2335 => x"34",
          2336 => x"15",
          2337 => x"0d",
          2338 => x"0d",
          2339 => x"57",
          2340 => x"17",
          2341 => x"08",
          2342 => x"82",
          2343 => x"89",
          2344 => x"55",
          2345 => x"14",
          2346 => x"16",
          2347 => x"71",
          2348 => x"38",
          2349 => x"09",
          2350 => x"38",
          2351 => x"73",
          2352 => x"81",
          2353 => x"ae",
          2354 => x"05",
          2355 => x"15",
          2356 => x"70",
          2357 => x"34",
          2358 => x"8a",
          2359 => x"38",
          2360 => x"05",
          2361 => x"81",
          2362 => x"17",
          2363 => x"12",
          2364 => x"34",
          2365 => x"9c",
          2366 => x"e8",
          2367 => x"ca",
          2368 => x"0c",
          2369 => x"e7",
          2370 => x"ca",
          2371 => x"17",
          2372 => x"51",
          2373 => x"91",
          2374 => x"84",
          2375 => x"3d",
          2376 => x"3d",
          2377 => x"08",
          2378 => x"61",
          2379 => x"55",
          2380 => x"2e",
          2381 => x"55",
          2382 => x"2e",
          2383 => x"80",
          2384 => x"94",
          2385 => x"1c",
          2386 => x"81",
          2387 => x"61",
          2388 => x"56",
          2389 => x"2e",
          2390 => x"83",
          2391 => x"73",
          2392 => x"70",
          2393 => x"25",
          2394 => x"51",
          2395 => x"38",
          2396 => x"0c",
          2397 => x"51",
          2398 => x"26",
          2399 => x"80",
          2400 => x"34",
          2401 => x"51",
          2402 => x"91",
          2403 => x"55",
          2404 => x"91",
          2405 => x"1d",
          2406 => x"8b",
          2407 => x"79",
          2408 => x"3f",
          2409 => x"57",
          2410 => x"55",
          2411 => x"2e",
          2412 => x"80",
          2413 => x"18",
          2414 => x"1a",
          2415 => x"70",
          2416 => x"2a",
          2417 => x"07",
          2418 => x"5a",
          2419 => x"8c",
          2420 => x"54",
          2421 => x"81",
          2422 => x"39",
          2423 => x"70",
          2424 => x"2a",
          2425 => x"75",
          2426 => x"8c",
          2427 => x"2e",
          2428 => x"a0",
          2429 => x"38",
          2430 => x"0c",
          2431 => x"76",
          2432 => x"38",
          2433 => x"b8",
          2434 => x"70",
          2435 => x"5a",
          2436 => x"76",
          2437 => x"38",
          2438 => x"70",
          2439 => x"dc",
          2440 => x"72",
          2441 => x"80",
          2442 => x"51",
          2443 => x"73",
          2444 => x"38",
          2445 => x"18",
          2446 => x"1a",
          2447 => x"55",
          2448 => x"2e",
          2449 => x"83",
          2450 => x"73",
          2451 => x"70",
          2452 => x"25",
          2453 => x"51",
          2454 => x"38",
          2455 => x"75",
          2456 => x"81",
          2457 => x"81",
          2458 => x"27",
          2459 => x"73",
          2460 => x"38",
          2461 => x"70",
          2462 => x"32",
          2463 => x"80",
          2464 => x"2a",
          2465 => x"56",
          2466 => x"81",
          2467 => x"57",
          2468 => x"f5",
          2469 => x"2b",
          2470 => x"25",
          2471 => x"80",
          2472 => x"b9",
          2473 => x"57",
          2474 => x"e6",
          2475 => x"ca",
          2476 => x"2e",
          2477 => x"18",
          2478 => x"1a",
          2479 => x"56",
          2480 => x"3f",
          2481 => x"08",
          2482 => x"e8",
          2483 => x"54",
          2484 => x"80",
          2485 => x"17",
          2486 => x"34",
          2487 => x"11",
          2488 => x"74",
          2489 => x"75",
          2490 => x"b4",
          2491 => x"3f",
          2492 => x"08",
          2493 => x"9f",
          2494 => x"99",
          2495 => x"e0",
          2496 => x"ff",
          2497 => x"79",
          2498 => x"74",
          2499 => x"57",
          2500 => x"77",
          2501 => x"76",
          2502 => x"38",
          2503 => x"73",
          2504 => x"09",
          2505 => x"38",
          2506 => x"84",
          2507 => x"27",
          2508 => x"39",
          2509 => x"f2",
          2510 => x"80",
          2511 => x"54",
          2512 => x"34",
          2513 => x"58",
          2514 => x"f2",
          2515 => x"ca",
          2516 => x"91",
          2517 => x"80",
          2518 => x"1b",
          2519 => x"51",
          2520 => x"91",
          2521 => x"56",
          2522 => x"08",
          2523 => x"9c",
          2524 => x"33",
          2525 => x"80",
          2526 => x"38",
          2527 => x"bf",
          2528 => x"86",
          2529 => x"15",
          2530 => x"2a",
          2531 => x"51",
          2532 => x"92",
          2533 => x"79",
          2534 => x"e4",
          2535 => x"ca",
          2536 => x"2e",
          2537 => x"52",
          2538 => x"ba",
          2539 => x"39",
          2540 => x"33",
          2541 => x"80",
          2542 => x"74",
          2543 => x"81",
          2544 => x"38",
          2545 => x"70",
          2546 => x"82",
          2547 => x"54",
          2548 => x"96",
          2549 => x"06",
          2550 => x"2e",
          2551 => x"ff",
          2552 => x"1c",
          2553 => x"80",
          2554 => x"81",
          2555 => x"ba",
          2556 => x"b6",
          2557 => x"2a",
          2558 => x"51",
          2559 => x"38",
          2560 => x"70",
          2561 => x"81",
          2562 => x"55",
          2563 => x"e1",
          2564 => x"08",
          2565 => x"1d",
          2566 => x"7c",
          2567 => x"3f",
          2568 => x"08",
          2569 => x"fa",
          2570 => x"91",
          2571 => x"8f",
          2572 => x"f6",
          2573 => x"5b",
          2574 => x"70",
          2575 => x"59",
          2576 => x"73",
          2577 => x"c6",
          2578 => x"81",
          2579 => x"70",
          2580 => x"52",
          2581 => x"8d",
          2582 => x"38",
          2583 => x"09",
          2584 => x"a5",
          2585 => x"d0",
          2586 => x"ff",
          2587 => x"53",
          2588 => x"91",
          2589 => x"73",
          2590 => x"d0",
          2591 => x"71",
          2592 => x"f7",
          2593 => x"91",
          2594 => x"55",
          2595 => x"55",
          2596 => x"81",
          2597 => x"74",
          2598 => x"56",
          2599 => x"12",
          2600 => x"70",
          2601 => x"38",
          2602 => x"81",
          2603 => x"51",
          2604 => x"51",
          2605 => x"89",
          2606 => x"70",
          2607 => x"53",
          2608 => x"70",
          2609 => x"51",
          2610 => x"09",
          2611 => x"38",
          2612 => x"38",
          2613 => x"77",
          2614 => x"70",
          2615 => x"2a",
          2616 => x"07",
          2617 => x"51",
          2618 => x"8f",
          2619 => x"84",
          2620 => x"83",
          2621 => x"94",
          2622 => x"74",
          2623 => x"38",
          2624 => x"0c",
          2625 => x"86",
          2626 => x"b8",
          2627 => x"91",
          2628 => x"8c",
          2629 => x"fa",
          2630 => x"56",
          2631 => x"17",
          2632 => x"b0",
          2633 => x"52",
          2634 => x"e0",
          2635 => x"91",
          2636 => x"81",
          2637 => x"b2",
          2638 => x"b4",
          2639 => x"88",
          2640 => x"ff",
          2641 => x"55",
          2642 => x"d5",
          2643 => x"06",
          2644 => x"80",
          2645 => x"33",
          2646 => x"81",
          2647 => x"81",
          2648 => x"81",
          2649 => x"eb",
          2650 => x"70",
          2651 => x"07",
          2652 => x"73",
          2653 => x"81",
          2654 => x"81",
          2655 => x"83",
          2656 => x"c4",
          2657 => x"16",
          2658 => x"3f",
          2659 => x"08",
          2660 => x"88",
          2661 => x"9d",
          2662 => x"91",
          2663 => x"81",
          2664 => x"e0",
          2665 => x"ca",
          2666 => x"91",
          2667 => x"80",
          2668 => x"82",
          2669 => x"ca",
          2670 => x"3d",
          2671 => x"3d",
          2672 => x"84",
          2673 => x"05",
          2674 => x"80",
          2675 => x"51",
          2676 => x"91",
          2677 => x"58",
          2678 => x"0b",
          2679 => x"08",
          2680 => x"38",
          2681 => x"08",
          2682 => x"ca",
          2683 => x"08",
          2684 => x"56",
          2685 => x"86",
          2686 => x"75",
          2687 => x"fe",
          2688 => x"54",
          2689 => x"2e",
          2690 => x"14",
          2691 => x"ca",
          2692 => x"88",
          2693 => x"06",
          2694 => x"54",
          2695 => x"38",
          2696 => x"86",
          2697 => x"82",
          2698 => x"06",
          2699 => x"56",
          2700 => x"38",
          2701 => x"80",
          2702 => x"81",
          2703 => x"52",
          2704 => x"51",
          2705 => x"91",
          2706 => x"81",
          2707 => x"81",
          2708 => x"83",
          2709 => x"87",
          2710 => x"2e",
          2711 => x"82",
          2712 => x"06",
          2713 => x"56",
          2714 => x"38",
          2715 => x"74",
          2716 => x"a3",
          2717 => x"88",
          2718 => x"06",
          2719 => x"2e",
          2720 => x"80",
          2721 => x"3d",
          2722 => x"83",
          2723 => x"15",
          2724 => x"53",
          2725 => x"8d",
          2726 => x"15",
          2727 => x"3f",
          2728 => x"08",
          2729 => x"70",
          2730 => x"0c",
          2731 => x"16",
          2732 => x"80",
          2733 => x"80",
          2734 => x"54",
          2735 => x"84",
          2736 => x"5b",
          2737 => x"80",
          2738 => x"7a",
          2739 => x"fc",
          2740 => x"ca",
          2741 => x"ff",
          2742 => x"77",
          2743 => x"81",
          2744 => x"76",
          2745 => x"81",
          2746 => x"2e",
          2747 => x"8d",
          2748 => x"26",
          2749 => x"bf",
          2750 => x"f4",
          2751 => x"88",
          2752 => x"ff",
          2753 => x"84",
          2754 => x"81",
          2755 => x"38",
          2756 => x"51",
          2757 => x"91",
          2758 => x"83",
          2759 => x"58",
          2760 => x"80",
          2761 => x"db",
          2762 => x"ca",
          2763 => x"77",
          2764 => x"80",
          2765 => x"82",
          2766 => x"c4",
          2767 => x"11",
          2768 => x"06",
          2769 => x"8d",
          2770 => x"26",
          2771 => x"74",
          2772 => x"78",
          2773 => x"c1",
          2774 => x"59",
          2775 => x"15",
          2776 => x"2e",
          2777 => x"13",
          2778 => x"72",
          2779 => x"38",
          2780 => x"eb",
          2781 => x"14",
          2782 => x"3f",
          2783 => x"08",
          2784 => x"88",
          2785 => x"23",
          2786 => x"57",
          2787 => x"83",
          2788 => x"c7",
          2789 => x"d8",
          2790 => x"88",
          2791 => x"ff",
          2792 => x"8d",
          2793 => x"14",
          2794 => x"3f",
          2795 => x"08",
          2796 => x"14",
          2797 => x"3f",
          2798 => x"08",
          2799 => x"06",
          2800 => x"72",
          2801 => x"97",
          2802 => x"22",
          2803 => x"84",
          2804 => x"5a",
          2805 => x"83",
          2806 => x"14",
          2807 => x"79",
          2808 => x"b3",
          2809 => x"ca",
          2810 => x"91",
          2811 => x"80",
          2812 => x"38",
          2813 => x"08",
          2814 => x"ff",
          2815 => x"38",
          2816 => x"83",
          2817 => x"83",
          2818 => x"74",
          2819 => x"85",
          2820 => x"89",
          2821 => x"76",
          2822 => x"c3",
          2823 => x"70",
          2824 => x"7b",
          2825 => x"73",
          2826 => x"17",
          2827 => x"ac",
          2828 => x"55",
          2829 => x"09",
          2830 => x"38",
          2831 => x"51",
          2832 => x"91",
          2833 => x"83",
          2834 => x"53",
          2835 => x"82",
          2836 => x"82",
          2837 => x"e0",
          2838 => x"ab",
          2839 => x"88",
          2840 => x"0c",
          2841 => x"53",
          2842 => x"56",
          2843 => x"81",
          2844 => x"13",
          2845 => x"74",
          2846 => x"82",
          2847 => x"74",
          2848 => x"81",
          2849 => x"06",
          2850 => x"83",
          2851 => x"2a",
          2852 => x"72",
          2853 => x"26",
          2854 => x"ff",
          2855 => x"0c",
          2856 => x"15",
          2857 => x"0b",
          2858 => x"76",
          2859 => x"81",
          2860 => x"38",
          2861 => x"51",
          2862 => x"91",
          2863 => x"83",
          2864 => x"53",
          2865 => x"09",
          2866 => x"f9",
          2867 => x"52",
          2868 => x"b8",
          2869 => x"88",
          2870 => x"38",
          2871 => x"08",
          2872 => x"84",
          2873 => x"d8",
          2874 => x"ca",
          2875 => x"ff",
          2876 => x"72",
          2877 => x"2e",
          2878 => x"80",
          2879 => x"14",
          2880 => x"3f",
          2881 => x"08",
          2882 => x"a4",
          2883 => x"81",
          2884 => x"84",
          2885 => x"d7",
          2886 => x"ca",
          2887 => x"8a",
          2888 => x"2e",
          2889 => x"9d",
          2890 => x"14",
          2891 => x"3f",
          2892 => x"08",
          2893 => x"84",
          2894 => x"d7",
          2895 => x"ca",
          2896 => x"15",
          2897 => x"34",
          2898 => x"22",
          2899 => x"72",
          2900 => x"23",
          2901 => x"23",
          2902 => x"15",
          2903 => x"75",
          2904 => x"0c",
          2905 => x"04",
          2906 => x"77",
          2907 => x"73",
          2908 => x"38",
          2909 => x"72",
          2910 => x"38",
          2911 => x"71",
          2912 => x"38",
          2913 => x"84",
          2914 => x"52",
          2915 => x"09",
          2916 => x"38",
          2917 => x"51",
          2918 => x"91",
          2919 => x"81",
          2920 => x"88",
          2921 => x"08",
          2922 => x"39",
          2923 => x"73",
          2924 => x"74",
          2925 => x"0c",
          2926 => x"04",
          2927 => x"02",
          2928 => x"7a",
          2929 => x"fc",
          2930 => x"f4",
          2931 => x"54",
          2932 => x"ca",
          2933 => x"bc",
          2934 => x"88",
          2935 => x"91",
          2936 => x"70",
          2937 => x"73",
          2938 => x"38",
          2939 => x"78",
          2940 => x"2e",
          2941 => x"74",
          2942 => x"0c",
          2943 => x"80",
          2944 => x"80",
          2945 => x"70",
          2946 => x"51",
          2947 => x"91",
          2948 => x"54",
          2949 => x"88",
          2950 => x"0d",
          2951 => x"0d",
          2952 => x"05",
          2953 => x"33",
          2954 => x"54",
          2955 => x"84",
          2956 => x"bf",
          2957 => x"98",
          2958 => x"53",
          2959 => x"05",
          2960 => x"fa",
          2961 => x"88",
          2962 => x"ca",
          2963 => x"a4",
          2964 => x"68",
          2965 => x"70",
          2966 => x"c6",
          2967 => x"88",
          2968 => x"ca",
          2969 => x"38",
          2970 => x"05",
          2971 => x"2b",
          2972 => x"80",
          2973 => x"86",
          2974 => x"06",
          2975 => x"2e",
          2976 => x"74",
          2977 => x"38",
          2978 => x"09",
          2979 => x"38",
          2980 => x"f8",
          2981 => x"88",
          2982 => x"39",
          2983 => x"33",
          2984 => x"73",
          2985 => x"77",
          2986 => x"81",
          2987 => x"73",
          2988 => x"38",
          2989 => x"bc",
          2990 => x"07",
          2991 => x"b4",
          2992 => x"2a",
          2993 => x"51",
          2994 => x"2e",
          2995 => x"62",
          2996 => x"e8",
          2997 => x"ca",
          2998 => x"82",
          2999 => x"52",
          3000 => x"51",
          3001 => x"62",
          3002 => x"8b",
          3003 => x"53",
          3004 => x"51",
          3005 => x"80",
          3006 => x"05",
          3007 => x"3f",
          3008 => x"0b",
          3009 => x"75",
          3010 => x"f1",
          3011 => x"11",
          3012 => x"80",
          3013 => x"97",
          3014 => x"51",
          3015 => x"91",
          3016 => x"55",
          3017 => x"08",
          3018 => x"b7",
          3019 => x"c4",
          3020 => x"05",
          3021 => x"2a",
          3022 => x"51",
          3023 => x"80",
          3024 => x"84",
          3025 => x"39",
          3026 => x"70",
          3027 => x"54",
          3028 => x"a9",
          3029 => x"06",
          3030 => x"2e",
          3031 => x"55",
          3032 => x"73",
          3033 => x"d6",
          3034 => x"ca",
          3035 => x"ff",
          3036 => x"0c",
          3037 => x"ca",
          3038 => x"f8",
          3039 => x"2a",
          3040 => x"51",
          3041 => x"2e",
          3042 => x"80",
          3043 => x"7a",
          3044 => x"a0",
          3045 => x"a4",
          3046 => x"53",
          3047 => x"e6",
          3048 => x"ca",
          3049 => x"ca",
          3050 => x"1b",
          3051 => x"05",
          3052 => x"d3",
          3053 => x"88",
          3054 => x"88",
          3055 => x"0c",
          3056 => x"56",
          3057 => x"84",
          3058 => x"90",
          3059 => x"0b",
          3060 => x"80",
          3061 => x"0c",
          3062 => x"1a",
          3063 => x"2a",
          3064 => x"51",
          3065 => x"2e",
          3066 => x"91",
          3067 => x"80",
          3068 => x"38",
          3069 => x"08",
          3070 => x"8a",
          3071 => x"89",
          3072 => x"59",
          3073 => x"76",
          3074 => x"d7",
          3075 => x"ca",
          3076 => x"91",
          3077 => x"81",
          3078 => x"82",
          3079 => x"88",
          3080 => x"09",
          3081 => x"38",
          3082 => x"78",
          3083 => x"30",
          3084 => x"80",
          3085 => x"77",
          3086 => x"38",
          3087 => x"06",
          3088 => x"c3",
          3089 => x"1a",
          3090 => x"38",
          3091 => x"06",
          3092 => x"2e",
          3093 => x"52",
          3094 => x"a6",
          3095 => x"88",
          3096 => x"82",
          3097 => x"75",
          3098 => x"ca",
          3099 => x"9c",
          3100 => x"39",
          3101 => x"74",
          3102 => x"ca",
          3103 => x"3d",
          3104 => x"3d",
          3105 => x"65",
          3106 => x"5d",
          3107 => x"0c",
          3108 => x"05",
          3109 => x"f9",
          3110 => x"ca",
          3111 => x"91",
          3112 => x"8a",
          3113 => x"33",
          3114 => x"2e",
          3115 => x"56",
          3116 => x"90",
          3117 => x"06",
          3118 => x"74",
          3119 => x"b6",
          3120 => x"82",
          3121 => x"34",
          3122 => x"aa",
          3123 => x"91",
          3124 => x"56",
          3125 => x"8c",
          3126 => x"1a",
          3127 => x"74",
          3128 => x"38",
          3129 => x"80",
          3130 => x"38",
          3131 => x"70",
          3132 => x"56",
          3133 => x"b2",
          3134 => x"11",
          3135 => x"77",
          3136 => x"5b",
          3137 => x"38",
          3138 => x"88",
          3139 => x"8f",
          3140 => x"08",
          3141 => x"d5",
          3142 => x"ca",
          3143 => x"81",
          3144 => x"9f",
          3145 => x"2e",
          3146 => x"74",
          3147 => x"98",
          3148 => x"7e",
          3149 => x"3f",
          3150 => x"08",
          3151 => x"83",
          3152 => x"88",
          3153 => x"89",
          3154 => x"77",
          3155 => x"d6",
          3156 => x"7f",
          3157 => x"58",
          3158 => x"75",
          3159 => x"75",
          3160 => x"77",
          3161 => x"7c",
          3162 => x"33",
          3163 => x"3f",
          3164 => x"08",
          3165 => x"7e",
          3166 => x"56",
          3167 => x"2e",
          3168 => x"16",
          3169 => x"55",
          3170 => x"94",
          3171 => x"53",
          3172 => x"b0",
          3173 => x"31",
          3174 => x"05",
          3175 => x"3f",
          3176 => x"56",
          3177 => x"9c",
          3178 => x"19",
          3179 => x"06",
          3180 => x"31",
          3181 => x"76",
          3182 => x"7b",
          3183 => x"08",
          3184 => x"d1",
          3185 => x"ca",
          3186 => x"81",
          3187 => x"94",
          3188 => x"ff",
          3189 => x"05",
          3190 => x"cf",
          3191 => x"76",
          3192 => x"17",
          3193 => x"1e",
          3194 => x"18",
          3195 => x"5e",
          3196 => x"39",
          3197 => x"91",
          3198 => x"90",
          3199 => x"f2",
          3200 => x"63",
          3201 => x"40",
          3202 => x"7e",
          3203 => x"fc",
          3204 => x"51",
          3205 => x"91",
          3206 => x"55",
          3207 => x"08",
          3208 => x"18",
          3209 => x"80",
          3210 => x"74",
          3211 => x"39",
          3212 => x"70",
          3213 => x"81",
          3214 => x"56",
          3215 => x"80",
          3216 => x"38",
          3217 => x"0b",
          3218 => x"82",
          3219 => x"39",
          3220 => x"19",
          3221 => x"83",
          3222 => x"18",
          3223 => x"56",
          3224 => x"27",
          3225 => x"09",
          3226 => x"2e",
          3227 => x"94",
          3228 => x"83",
          3229 => x"56",
          3230 => x"38",
          3231 => x"22",
          3232 => x"89",
          3233 => x"55",
          3234 => x"75",
          3235 => x"18",
          3236 => x"9c",
          3237 => x"85",
          3238 => x"08",
          3239 => x"d7",
          3240 => x"ca",
          3241 => x"91",
          3242 => x"80",
          3243 => x"38",
          3244 => x"ff",
          3245 => x"ff",
          3246 => x"38",
          3247 => x"0c",
          3248 => x"85",
          3249 => x"19",
          3250 => x"b0",
          3251 => x"19",
          3252 => x"81",
          3253 => x"74",
          3254 => x"3f",
          3255 => x"08",
          3256 => x"98",
          3257 => x"7e",
          3258 => x"3f",
          3259 => x"08",
          3260 => x"d2",
          3261 => x"88",
          3262 => x"89",
          3263 => x"78",
          3264 => x"d5",
          3265 => x"7f",
          3266 => x"58",
          3267 => x"75",
          3268 => x"75",
          3269 => x"78",
          3270 => x"7c",
          3271 => x"33",
          3272 => x"3f",
          3273 => x"08",
          3274 => x"7e",
          3275 => x"78",
          3276 => x"74",
          3277 => x"38",
          3278 => x"b0",
          3279 => x"31",
          3280 => x"05",
          3281 => x"51",
          3282 => x"7e",
          3283 => x"83",
          3284 => x"89",
          3285 => x"db",
          3286 => x"08",
          3287 => x"26",
          3288 => x"51",
          3289 => x"91",
          3290 => x"fd",
          3291 => x"77",
          3292 => x"55",
          3293 => x"0c",
          3294 => x"83",
          3295 => x"80",
          3296 => x"55",
          3297 => x"83",
          3298 => x"9c",
          3299 => x"7e",
          3300 => x"3f",
          3301 => x"08",
          3302 => x"75",
          3303 => x"94",
          3304 => x"ff",
          3305 => x"05",
          3306 => x"3f",
          3307 => x"0b",
          3308 => x"7b",
          3309 => x"08",
          3310 => x"76",
          3311 => x"08",
          3312 => x"1c",
          3313 => x"08",
          3314 => x"5c",
          3315 => x"83",
          3316 => x"74",
          3317 => x"fd",
          3318 => x"18",
          3319 => x"07",
          3320 => x"19",
          3321 => x"75",
          3322 => x"0c",
          3323 => x"04",
          3324 => x"7a",
          3325 => x"05",
          3326 => x"56",
          3327 => x"91",
          3328 => x"57",
          3329 => x"08",
          3330 => x"90",
          3331 => x"86",
          3332 => x"06",
          3333 => x"73",
          3334 => x"e9",
          3335 => x"08",
          3336 => x"cc",
          3337 => x"ca",
          3338 => x"91",
          3339 => x"80",
          3340 => x"16",
          3341 => x"33",
          3342 => x"55",
          3343 => x"34",
          3344 => x"53",
          3345 => x"08",
          3346 => x"3f",
          3347 => x"52",
          3348 => x"c9",
          3349 => x"88",
          3350 => x"96",
          3351 => x"f0",
          3352 => x"92",
          3353 => x"ca",
          3354 => x"81",
          3355 => x"34",
          3356 => x"df",
          3357 => x"88",
          3358 => x"33",
          3359 => x"55",
          3360 => x"17",
          3361 => x"ca",
          3362 => x"3d",
          3363 => x"3d",
          3364 => x"52",
          3365 => x"3f",
          3366 => x"08",
          3367 => x"88",
          3368 => x"86",
          3369 => x"52",
          3370 => x"bc",
          3371 => x"88",
          3372 => x"ca",
          3373 => x"38",
          3374 => x"08",
          3375 => x"91",
          3376 => x"86",
          3377 => x"ff",
          3378 => x"3d",
          3379 => x"3f",
          3380 => x"0b",
          3381 => x"08",
          3382 => x"91",
          3383 => x"91",
          3384 => x"80",
          3385 => x"ca",
          3386 => x"3d",
          3387 => x"3d",
          3388 => x"93",
          3389 => x"52",
          3390 => x"e9",
          3391 => x"ca",
          3392 => x"91",
          3393 => x"80",
          3394 => x"58",
          3395 => x"3d",
          3396 => x"e0",
          3397 => x"ca",
          3398 => x"91",
          3399 => x"bc",
          3400 => x"c7",
          3401 => x"98",
          3402 => x"73",
          3403 => x"38",
          3404 => x"12",
          3405 => x"39",
          3406 => x"33",
          3407 => x"70",
          3408 => x"55",
          3409 => x"2e",
          3410 => x"7f",
          3411 => x"54",
          3412 => x"91",
          3413 => x"94",
          3414 => x"39",
          3415 => x"08",
          3416 => x"81",
          3417 => x"85",
          3418 => x"ca",
          3419 => x"3d",
          3420 => x"3d",
          3421 => x"5b",
          3422 => x"34",
          3423 => x"3d",
          3424 => x"52",
          3425 => x"e8",
          3426 => x"ca",
          3427 => x"91",
          3428 => x"82",
          3429 => x"43",
          3430 => x"11",
          3431 => x"58",
          3432 => x"80",
          3433 => x"38",
          3434 => x"3d",
          3435 => x"d5",
          3436 => x"ca",
          3437 => x"91",
          3438 => x"82",
          3439 => x"52",
          3440 => x"c8",
          3441 => x"88",
          3442 => x"ca",
          3443 => x"c1",
          3444 => x"7b",
          3445 => x"3f",
          3446 => x"08",
          3447 => x"74",
          3448 => x"3f",
          3449 => x"08",
          3450 => x"88",
          3451 => x"38",
          3452 => x"51",
          3453 => x"91",
          3454 => x"57",
          3455 => x"08",
          3456 => x"52",
          3457 => x"f2",
          3458 => x"ca",
          3459 => x"a6",
          3460 => x"74",
          3461 => x"3f",
          3462 => x"08",
          3463 => x"88",
          3464 => x"cc",
          3465 => x"2e",
          3466 => x"86",
          3467 => x"81",
          3468 => x"81",
          3469 => x"3d",
          3470 => x"52",
          3471 => x"c9",
          3472 => x"3d",
          3473 => x"11",
          3474 => x"5a",
          3475 => x"2e",
          3476 => x"b9",
          3477 => x"16",
          3478 => x"33",
          3479 => x"73",
          3480 => x"16",
          3481 => x"26",
          3482 => x"75",
          3483 => x"38",
          3484 => x"05",
          3485 => x"6f",
          3486 => x"ff",
          3487 => x"55",
          3488 => x"74",
          3489 => x"38",
          3490 => x"11",
          3491 => x"74",
          3492 => x"39",
          3493 => x"09",
          3494 => x"38",
          3495 => x"11",
          3496 => x"74",
          3497 => x"91",
          3498 => x"70",
          3499 => x"b9",
          3500 => x"08",
          3501 => x"5c",
          3502 => x"73",
          3503 => x"38",
          3504 => x"1a",
          3505 => x"55",
          3506 => x"38",
          3507 => x"73",
          3508 => x"38",
          3509 => x"76",
          3510 => x"74",
          3511 => x"33",
          3512 => x"05",
          3513 => x"15",
          3514 => x"ba",
          3515 => x"05",
          3516 => x"ff",
          3517 => x"06",
          3518 => x"57",
          3519 => x"18",
          3520 => x"54",
          3521 => x"70",
          3522 => x"34",
          3523 => x"ee",
          3524 => x"34",
          3525 => x"88",
          3526 => x"0d",
          3527 => x"0d",
          3528 => x"3d",
          3529 => x"71",
          3530 => x"ec",
          3531 => x"ca",
          3532 => x"91",
          3533 => x"82",
          3534 => x"15",
          3535 => x"82",
          3536 => x"15",
          3537 => x"76",
          3538 => x"90",
          3539 => x"81",
          3540 => x"06",
          3541 => x"72",
          3542 => x"56",
          3543 => x"54",
          3544 => x"17",
          3545 => x"78",
          3546 => x"38",
          3547 => x"22",
          3548 => x"59",
          3549 => x"78",
          3550 => x"76",
          3551 => x"51",
          3552 => x"3f",
          3553 => x"08",
          3554 => x"54",
          3555 => x"53",
          3556 => x"3f",
          3557 => x"08",
          3558 => x"38",
          3559 => x"75",
          3560 => x"18",
          3561 => x"31",
          3562 => x"57",
          3563 => x"b1",
          3564 => x"08",
          3565 => x"38",
          3566 => x"51",
          3567 => x"91",
          3568 => x"54",
          3569 => x"08",
          3570 => x"9a",
          3571 => x"88",
          3572 => x"81",
          3573 => x"ca",
          3574 => x"16",
          3575 => x"16",
          3576 => x"2e",
          3577 => x"76",
          3578 => x"dc",
          3579 => x"31",
          3580 => x"18",
          3581 => x"90",
          3582 => x"81",
          3583 => x"06",
          3584 => x"56",
          3585 => x"9a",
          3586 => x"74",
          3587 => x"3f",
          3588 => x"08",
          3589 => x"88",
          3590 => x"91",
          3591 => x"56",
          3592 => x"52",
          3593 => x"84",
          3594 => x"88",
          3595 => x"ff",
          3596 => x"81",
          3597 => x"38",
          3598 => x"98",
          3599 => x"a6",
          3600 => x"16",
          3601 => x"39",
          3602 => x"16",
          3603 => x"75",
          3604 => x"53",
          3605 => x"aa",
          3606 => x"79",
          3607 => x"3f",
          3608 => x"08",
          3609 => x"0b",
          3610 => x"82",
          3611 => x"39",
          3612 => x"16",
          3613 => x"bb",
          3614 => x"2a",
          3615 => x"08",
          3616 => x"15",
          3617 => x"15",
          3618 => x"90",
          3619 => x"16",
          3620 => x"33",
          3621 => x"53",
          3622 => x"34",
          3623 => x"06",
          3624 => x"2e",
          3625 => x"9c",
          3626 => x"85",
          3627 => x"16",
          3628 => x"72",
          3629 => x"0c",
          3630 => x"04",
          3631 => x"79",
          3632 => x"75",
          3633 => x"8a",
          3634 => x"89",
          3635 => x"52",
          3636 => x"05",
          3637 => x"3f",
          3638 => x"08",
          3639 => x"88",
          3640 => x"38",
          3641 => x"7a",
          3642 => x"d8",
          3643 => x"ca",
          3644 => x"91",
          3645 => x"80",
          3646 => x"16",
          3647 => x"2b",
          3648 => x"74",
          3649 => x"86",
          3650 => x"84",
          3651 => x"06",
          3652 => x"73",
          3653 => x"38",
          3654 => x"52",
          3655 => x"da",
          3656 => x"88",
          3657 => x"0c",
          3658 => x"14",
          3659 => x"23",
          3660 => x"51",
          3661 => x"91",
          3662 => x"55",
          3663 => x"09",
          3664 => x"38",
          3665 => x"39",
          3666 => x"84",
          3667 => x"0c",
          3668 => x"91",
          3669 => x"89",
          3670 => x"fc",
          3671 => x"87",
          3672 => x"53",
          3673 => x"e7",
          3674 => x"ca",
          3675 => x"38",
          3676 => x"08",
          3677 => x"3d",
          3678 => x"3d",
          3679 => x"89",
          3680 => x"54",
          3681 => x"54",
          3682 => x"91",
          3683 => x"53",
          3684 => x"08",
          3685 => x"74",
          3686 => x"ca",
          3687 => x"73",
          3688 => x"3f",
          3689 => x"08",
          3690 => x"39",
          3691 => x"08",
          3692 => x"d3",
          3693 => x"ca",
          3694 => x"91",
          3695 => x"84",
          3696 => x"06",
          3697 => x"53",
          3698 => x"ca",
          3699 => x"38",
          3700 => x"51",
          3701 => x"72",
          3702 => x"cf",
          3703 => x"ca",
          3704 => x"32",
          3705 => x"72",
          3706 => x"70",
          3707 => x"08",
          3708 => x"54",
          3709 => x"ca",
          3710 => x"3d",
          3711 => x"3d",
          3712 => x"80",
          3713 => x"70",
          3714 => x"52",
          3715 => x"3f",
          3716 => x"08",
          3717 => x"88",
          3718 => x"64",
          3719 => x"d6",
          3720 => x"ca",
          3721 => x"91",
          3722 => x"a0",
          3723 => x"cb",
          3724 => x"98",
          3725 => x"73",
          3726 => x"38",
          3727 => x"39",
          3728 => x"88",
          3729 => x"75",
          3730 => x"3f",
          3731 => x"88",
          3732 => x"0d",
          3733 => x"0d",
          3734 => x"5c",
          3735 => x"3d",
          3736 => x"93",
          3737 => x"d6",
          3738 => x"88",
          3739 => x"ca",
          3740 => x"80",
          3741 => x"0c",
          3742 => x"11",
          3743 => x"90",
          3744 => x"56",
          3745 => x"74",
          3746 => x"75",
          3747 => x"e4",
          3748 => x"81",
          3749 => x"5b",
          3750 => x"91",
          3751 => x"75",
          3752 => x"73",
          3753 => x"81",
          3754 => x"82",
          3755 => x"76",
          3756 => x"f0",
          3757 => x"f4",
          3758 => x"88",
          3759 => x"d1",
          3760 => x"88",
          3761 => x"ce",
          3762 => x"88",
          3763 => x"91",
          3764 => x"07",
          3765 => x"05",
          3766 => x"53",
          3767 => x"98",
          3768 => x"26",
          3769 => x"f9",
          3770 => x"08",
          3771 => x"08",
          3772 => x"98",
          3773 => x"81",
          3774 => x"58",
          3775 => x"3f",
          3776 => x"08",
          3777 => x"88",
          3778 => x"38",
          3779 => x"77",
          3780 => x"5d",
          3781 => x"74",
          3782 => x"81",
          3783 => x"b4",
          3784 => x"bb",
          3785 => x"ca",
          3786 => x"ff",
          3787 => x"30",
          3788 => x"1b",
          3789 => x"5b",
          3790 => x"39",
          3791 => x"ff",
          3792 => x"91",
          3793 => x"f0",
          3794 => x"30",
          3795 => x"1b",
          3796 => x"5b",
          3797 => x"83",
          3798 => x"58",
          3799 => x"92",
          3800 => x"0c",
          3801 => x"12",
          3802 => x"33",
          3803 => x"54",
          3804 => x"34",
          3805 => x"88",
          3806 => x"0d",
          3807 => x"0d",
          3808 => x"fc",
          3809 => x"52",
          3810 => x"3f",
          3811 => x"08",
          3812 => x"88",
          3813 => x"38",
          3814 => x"56",
          3815 => x"38",
          3816 => x"70",
          3817 => x"81",
          3818 => x"55",
          3819 => x"80",
          3820 => x"38",
          3821 => x"54",
          3822 => x"08",
          3823 => x"38",
          3824 => x"91",
          3825 => x"53",
          3826 => x"52",
          3827 => x"8c",
          3828 => x"88",
          3829 => x"19",
          3830 => x"c9",
          3831 => x"08",
          3832 => x"ff",
          3833 => x"91",
          3834 => x"ff",
          3835 => x"06",
          3836 => x"56",
          3837 => x"08",
          3838 => x"81",
          3839 => x"82",
          3840 => x"75",
          3841 => x"54",
          3842 => x"08",
          3843 => x"27",
          3844 => x"17",
          3845 => x"ca",
          3846 => x"76",
          3847 => x"3f",
          3848 => x"08",
          3849 => x"08",
          3850 => x"90",
          3851 => x"c0",
          3852 => x"90",
          3853 => x"80",
          3854 => x"75",
          3855 => x"75",
          3856 => x"ca",
          3857 => x"3d",
          3858 => x"3d",
          3859 => x"a0",
          3860 => x"05",
          3861 => x"51",
          3862 => x"91",
          3863 => x"55",
          3864 => x"08",
          3865 => x"78",
          3866 => x"08",
          3867 => x"70",
          3868 => x"ae",
          3869 => x"88",
          3870 => x"ca",
          3871 => x"db",
          3872 => x"fb",
          3873 => x"85",
          3874 => x"06",
          3875 => x"86",
          3876 => x"c7",
          3877 => x"2b",
          3878 => x"24",
          3879 => x"02",
          3880 => x"33",
          3881 => x"58",
          3882 => x"76",
          3883 => x"6b",
          3884 => x"cc",
          3885 => x"ca",
          3886 => x"84",
          3887 => x"06",
          3888 => x"73",
          3889 => x"d4",
          3890 => x"91",
          3891 => x"94",
          3892 => x"81",
          3893 => x"5a",
          3894 => x"08",
          3895 => x"8a",
          3896 => x"54",
          3897 => x"91",
          3898 => x"55",
          3899 => x"08",
          3900 => x"91",
          3901 => x"52",
          3902 => x"e5",
          3903 => x"88",
          3904 => x"ca",
          3905 => x"38",
          3906 => x"cf",
          3907 => x"88",
          3908 => x"88",
          3909 => x"88",
          3910 => x"38",
          3911 => x"c2",
          3912 => x"88",
          3913 => x"88",
          3914 => x"91",
          3915 => x"07",
          3916 => x"55",
          3917 => x"2e",
          3918 => x"80",
          3919 => x"80",
          3920 => x"77",
          3921 => x"3f",
          3922 => x"08",
          3923 => x"38",
          3924 => x"ba",
          3925 => x"ca",
          3926 => x"74",
          3927 => x"0c",
          3928 => x"04",
          3929 => x"82",
          3930 => x"c0",
          3931 => x"3d",
          3932 => x"3f",
          3933 => x"08",
          3934 => x"88",
          3935 => x"38",
          3936 => x"52",
          3937 => x"52",
          3938 => x"3f",
          3939 => x"08",
          3940 => x"88",
          3941 => x"88",
          3942 => x"39",
          3943 => x"08",
          3944 => x"81",
          3945 => x"38",
          3946 => x"05",
          3947 => x"2a",
          3948 => x"55",
          3949 => x"81",
          3950 => x"5a",
          3951 => x"3d",
          3952 => x"c1",
          3953 => x"ca",
          3954 => x"55",
          3955 => x"88",
          3956 => x"87",
          3957 => x"88",
          3958 => x"09",
          3959 => x"38",
          3960 => x"ca",
          3961 => x"2e",
          3962 => x"86",
          3963 => x"81",
          3964 => x"81",
          3965 => x"ca",
          3966 => x"78",
          3967 => x"3f",
          3968 => x"08",
          3969 => x"88",
          3970 => x"38",
          3971 => x"52",
          3972 => x"ff",
          3973 => x"78",
          3974 => x"b4",
          3975 => x"54",
          3976 => x"15",
          3977 => x"b2",
          3978 => x"ca",
          3979 => x"b6",
          3980 => x"53",
          3981 => x"53",
          3982 => x"3f",
          3983 => x"b4",
          3984 => x"d4",
          3985 => x"b6",
          3986 => x"54",
          3987 => x"d5",
          3988 => x"53",
          3989 => x"11",
          3990 => x"d7",
          3991 => x"81",
          3992 => x"34",
          3993 => x"a4",
          3994 => x"88",
          3995 => x"ca",
          3996 => x"38",
          3997 => x"0a",
          3998 => x"05",
          3999 => x"d0",
          4000 => x"64",
          4001 => x"c9",
          4002 => x"54",
          4003 => x"15",
          4004 => x"81",
          4005 => x"34",
          4006 => x"b8",
          4007 => x"ca",
          4008 => x"8b",
          4009 => x"75",
          4010 => x"ff",
          4011 => x"73",
          4012 => x"0c",
          4013 => x"04",
          4014 => x"a9",
          4015 => x"51",
          4016 => x"82",
          4017 => x"ff",
          4018 => x"a9",
          4019 => x"ee",
          4020 => x"88",
          4021 => x"ca",
          4022 => x"d3",
          4023 => x"a9",
          4024 => x"9d",
          4025 => x"58",
          4026 => x"91",
          4027 => x"55",
          4028 => x"08",
          4029 => x"02",
          4030 => x"33",
          4031 => x"54",
          4032 => x"82",
          4033 => x"53",
          4034 => x"52",
          4035 => x"88",
          4036 => x"b4",
          4037 => x"53",
          4038 => x"3d",
          4039 => x"ff",
          4040 => x"aa",
          4041 => x"73",
          4042 => x"3f",
          4043 => x"08",
          4044 => x"88",
          4045 => x"63",
          4046 => x"81",
          4047 => x"65",
          4048 => x"2e",
          4049 => x"55",
          4050 => x"91",
          4051 => x"84",
          4052 => x"06",
          4053 => x"73",
          4054 => x"3f",
          4055 => x"08",
          4056 => x"88",
          4057 => x"38",
          4058 => x"53",
          4059 => x"95",
          4060 => x"16",
          4061 => x"87",
          4062 => x"05",
          4063 => x"34",
          4064 => x"70",
          4065 => x"81",
          4066 => x"55",
          4067 => x"74",
          4068 => x"73",
          4069 => x"78",
          4070 => x"83",
          4071 => x"16",
          4072 => x"2a",
          4073 => x"51",
          4074 => x"80",
          4075 => x"38",
          4076 => x"80",
          4077 => x"52",
          4078 => x"be",
          4079 => x"88",
          4080 => x"51",
          4081 => x"3f",
          4082 => x"ca",
          4083 => x"2e",
          4084 => x"91",
          4085 => x"52",
          4086 => x"b5",
          4087 => x"ca",
          4088 => x"80",
          4089 => x"58",
          4090 => x"88",
          4091 => x"38",
          4092 => x"54",
          4093 => x"09",
          4094 => x"38",
          4095 => x"52",
          4096 => x"af",
          4097 => x"81",
          4098 => x"34",
          4099 => x"ca",
          4100 => x"38",
          4101 => x"ca",
          4102 => x"88",
          4103 => x"ca",
          4104 => x"38",
          4105 => x"b5",
          4106 => x"ca",
          4107 => x"74",
          4108 => x"0c",
          4109 => x"04",
          4110 => x"02",
          4111 => x"33",
          4112 => x"80",
          4113 => x"57",
          4114 => x"95",
          4115 => x"52",
          4116 => x"d2",
          4117 => x"ca",
          4118 => x"91",
          4119 => x"80",
          4120 => x"5a",
          4121 => x"3d",
          4122 => x"c9",
          4123 => x"ca",
          4124 => x"91",
          4125 => x"b8",
          4126 => x"cf",
          4127 => x"a0",
          4128 => x"55",
          4129 => x"75",
          4130 => x"71",
          4131 => x"33",
          4132 => x"74",
          4133 => x"57",
          4134 => x"8b",
          4135 => x"54",
          4136 => x"15",
          4137 => x"ff",
          4138 => x"91",
          4139 => x"55",
          4140 => x"88",
          4141 => x"0d",
          4142 => x"0d",
          4143 => x"53",
          4144 => x"05",
          4145 => x"51",
          4146 => x"91",
          4147 => x"55",
          4148 => x"08",
          4149 => x"76",
          4150 => x"93",
          4151 => x"51",
          4152 => x"91",
          4153 => x"55",
          4154 => x"08",
          4155 => x"80",
          4156 => x"81",
          4157 => x"86",
          4158 => x"38",
          4159 => x"86",
          4160 => x"90",
          4161 => x"54",
          4162 => x"ff",
          4163 => x"76",
          4164 => x"83",
          4165 => x"51",
          4166 => x"3f",
          4167 => x"08",
          4168 => x"ca",
          4169 => x"3d",
          4170 => x"3d",
          4171 => x"5c",
          4172 => x"98",
          4173 => x"52",
          4174 => x"d1",
          4175 => x"ca",
          4176 => x"ca",
          4177 => x"70",
          4178 => x"08",
          4179 => x"51",
          4180 => x"80",
          4181 => x"38",
          4182 => x"06",
          4183 => x"80",
          4184 => x"38",
          4185 => x"5f",
          4186 => x"3d",
          4187 => x"ff",
          4188 => x"91",
          4189 => x"57",
          4190 => x"08",
          4191 => x"74",
          4192 => x"c3",
          4193 => x"ca",
          4194 => x"91",
          4195 => x"bf",
          4196 => x"88",
          4197 => x"88",
          4198 => x"59",
          4199 => x"81",
          4200 => x"56",
          4201 => x"33",
          4202 => x"16",
          4203 => x"27",
          4204 => x"56",
          4205 => x"80",
          4206 => x"80",
          4207 => x"ff",
          4208 => x"70",
          4209 => x"56",
          4210 => x"e8",
          4211 => x"76",
          4212 => x"81",
          4213 => x"80",
          4214 => x"57",
          4215 => x"78",
          4216 => x"51",
          4217 => x"2e",
          4218 => x"73",
          4219 => x"38",
          4220 => x"08",
          4221 => x"b1",
          4222 => x"ca",
          4223 => x"91",
          4224 => x"a7",
          4225 => x"33",
          4226 => x"c3",
          4227 => x"2e",
          4228 => x"e4",
          4229 => x"2e",
          4230 => x"56",
          4231 => x"05",
          4232 => x"e3",
          4233 => x"88",
          4234 => x"76",
          4235 => x"0c",
          4236 => x"04",
          4237 => x"82",
          4238 => x"ff",
          4239 => x"9d",
          4240 => x"fa",
          4241 => x"88",
          4242 => x"88",
          4243 => x"91",
          4244 => x"83",
          4245 => x"53",
          4246 => x"3d",
          4247 => x"ff",
          4248 => x"73",
          4249 => x"70",
          4250 => x"52",
          4251 => x"9f",
          4252 => x"bc",
          4253 => x"74",
          4254 => x"6d",
          4255 => x"70",
          4256 => x"af",
          4257 => x"ca",
          4258 => x"2e",
          4259 => x"70",
          4260 => x"57",
          4261 => x"fd",
          4262 => x"88",
          4263 => x"8d",
          4264 => x"2b",
          4265 => x"81",
          4266 => x"86",
          4267 => x"88",
          4268 => x"9f",
          4269 => x"ff",
          4270 => x"54",
          4271 => x"8a",
          4272 => x"70",
          4273 => x"06",
          4274 => x"ff",
          4275 => x"38",
          4276 => x"15",
          4277 => x"80",
          4278 => x"74",
          4279 => x"94",
          4280 => x"89",
          4281 => x"88",
          4282 => x"81",
          4283 => x"88",
          4284 => x"26",
          4285 => x"39",
          4286 => x"86",
          4287 => x"81",
          4288 => x"ff",
          4289 => x"38",
          4290 => x"54",
          4291 => x"81",
          4292 => x"81",
          4293 => x"78",
          4294 => x"5a",
          4295 => x"6d",
          4296 => x"81",
          4297 => x"57",
          4298 => x"9f",
          4299 => x"38",
          4300 => x"54",
          4301 => x"81",
          4302 => x"b1",
          4303 => x"2e",
          4304 => x"a7",
          4305 => x"15",
          4306 => x"54",
          4307 => x"09",
          4308 => x"38",
          4309 => x"76",
          4310 => x"41",
          4311 => x"52",
          4312 => x"52",
          4313 => x"b3",
          4314 => x"88",
          4315 => x"ca",
          4316 => x"f7",
          4317 => x"74",
          4318 => x"e5",
          4319 => x"88",
          4320 => x"ca",
          4321 => x"38",
          4322 => x"38",
          4323 => x"74",
          4324 => x"39",
          4325 => x"08",
          4326 => x"81",
          4327 => x"38",
          4328 => x"74",
          4329 => x"38",
          4330 => x"51",
          4331 => x"3f",
          4332 => x"08",
          4333 => x"88",
          4334 => x"a0",
          4335 => x"88",
          4336 => x"51",
          4337 => x"3f",
          4338 => x"0b",
          4339 => x"8b",
          4340 => x"67",
          4341 => x"a7",
          4342 => x"81",
          4343 => x"34",
          4344 => x"ad",
          4345 => x"ca",
          4346 => x"73",
          4347 => x"ca",
          4348 => x"3d",
          4349 => x"3d",
          4350 => x"02",
          4351 => x"cb",
          4352 => x"3d",
          4353 => x"72",
          4354 => x"5a",
          4355 => x"91",
          4356 => x"58",
          4357 => x"08",
          4358 => x"91",
          4359 => x"77",
          4360 => x"7c",
          4361 => x"38",
          4362 => x"59",
          4363 => x"90",
          4364 => x"81",
          4365 => x"06",
          4366 => x"73",
          4367 => x"54",
          4368 => x"82",
          4369 => x"39",
          4370 => x"8b",
          4371 => x"11",
          4372 => x"2b",
          4373 => x"54",
          4374 => x"ff",
          4375 => x"ff",
          4376 => x"70",
          4377 => x"07",
          4378 => x"ca",
          4379 => x"8c",
          4380 => x"40",
          4381 => x"55",
          4382 => x"88",
          4383 => x"08",
          4384 => x"38",
          4385 => x"77",
          4386 => x"56",
          4387 => x"51",
          4388 => x"3f",
          4389 => x"55",
          4390 => x"08",
          4391 => x"38",
          4392 => x"ca",
          4393 => x"2e",
          4394 => x"91",
          4395 => x"ff",
          4396 => x"38",
          4397 => x"08",
          4398 => x"16",
          4399 => x"2e",
          4400 => x"87",
          4401 => x"74",
          4402 => x"74",
          4403 => x"81",
          4404 => x"38",
          4405 => x"ff",
          4406 => x"2e",
          4407 => x"7b",
          4408 => x"80",
          4409 => x"81",
          4410 => x"81",
          4411 => x"06",
          4412 => x"56",
          4413 => x"52",
          4414 => x"af",
          4415 => x"ca",
          4416 => x"91",
          4417 => x"80",
          4418 => x"81",
          4419 => x"56",
          4420 => x"d3",
          4421 => x"ff",
          4422 => x"7c",
          4423 => x"55",
          4424 => x"b3",
          4425 => x"1b",
          4426 => x"1b",
          4427 => x"33",
          4428 => x"54",
          4429 => x"34",
          4430 => x"fe",
          4431 => x"08",
          4432 => x"74",
          4433 => x"75",
          4434 => x"16",
          4435 => x"33",
          4436 => x"73",
          4437 => x"77",
          4438 => x"ca",
          4439 => x"3d",
          4440 => x"3d",
          4441 => x"02",
          4442 => x"eb",
          4443 => x"3d",
          4444 => x"59",
          4445 => x"8b",
          4446 => x"91",
          4447 => x"24",
          4448 => x"91",
          4449 => x"84",
          4450 => x"a4",
          4451 => x"51",
          4452 => x"2e",
          4453 => x"75",
          4454 => x"88",
          4455 => x"06",
          4456 => x"7e",
          4457 => x"d0",
          4458 => x"88",
          4459 => x"06",
          4460 => x"56",
          4461 => x"74",
          4462 => x"76",
          4463 => x"81",
          4464 => x"8a",
          4465 => x"b2",
          4466 => x"fc",
          4467 => x"52",
          4468 => x"a4",
          4469 => x"ca",
          4470 => x"38",
          4471 => x"80",
          4472 => x"74",
          4473 => x"26",
          4474 => x"15",
          4475 => x"74",
          4476 => x"38",
          4477 => x"80",
          4478 => x"84",
          4479 => x"92",
          4480 => x"80",
          4481 => x"38",
          4482 => x"06",
          4483 => x"2e",
          4484 => x"56",
          4485 => x"78",
          4486 => x"89",
          4487 => x"2b",
          4488 => x"43",
          4489 => x"38",
          4490 => x"30",
          4491 => x"77",
          4492 => x"91",
          4493 => x"c2",
          4494 => x"f8",
          4495 => x"52",
          4496 => x"a4",
          4497 => x"56",
          4498 => x"08",
          4499 => x"77",
          4500 => x"77",
          4501 => x"88",
          4502 => x"45",
          4503 => x"bf",
          4504 => x"8e",
          4505 => x"26",
          4506 => x"74",
          4507 => x"48",
          4508 => x"75",
          4509 => x"38",
          4510 => x"81",
          4511 => x"fa",
          4512 => x"2a",
          4513 => x"56",
          4514 => x"2e",
          4515 => x"87",
          4516 => x"82",
          4517 => x"38",
          4518 => x"55",
          4519 => x"83",
          4520 => x"81",
          4521 => x"56",
          4522 => x"80",
          4523 => x"38",
          4524 => x"83",
          4525 => x"06",
          4526 => x"78",
          4527 => x"91",
          4528 => x"0b",
          4529 => x"22",
          4530 => x"80",
          4531 => x"74",
          4532 => x"38",
          4533 => x"56",
          4534 => x"17",
          4535 => x"57",
          4536 => x"2e",
          4537 => x"75",
          4538 => x"79",
          4539 => x"fe",
          4540 => x"91",
          4541 => x"84",
          4542 => x"05",
          4543 => x"5e",
          4544 => x"80",
          4545 => x"88",
          4546 => x"8a",
          4547 => x"fd",
          4548 => x"75",
          4549 => x"38",
          4550 => x"78",
          4551 => x"8c",
          4552 => x"0b",
          4553 => x"22",
          4554 => x"80",
          4555 => x"74",
          4556 => x"38",
          4557 => x"56",
          4558 => x"17",
          4559 => x"57",
          4560 => x"2e",
          4561 => x"75",
          4562 => x"79",
          4563 => x"fe",
          4564 => x"91",
          4565 => x"10",
          4566 => x"91",
          4567 => x"9f",
          4568 => x"38",
          4569 => x"ca",
          4570 => x"91",
          4571 => x"05",
          4572 => x"2a",
          4573 => x"56",
          4574 => x"17",
          4575 => x"81",
          4576 => x"60",
          4577 => x"65",
          4578 => x"12",
          4579 => x"30",
          4580 => x"74",
          4581 => x"59",
          4582 => x"7d",
          4583 => x"81",
          4584 => x"76",
          4585 => x"41",
          4586 => x"76",
          4587 => x"90",
          4588 => x"62",
          4589 => x"51",
          4590 => x"26",
          4591 => x"75",
          4592 => x"31",
          4593 => x"65",
          4594 => x"fe",
          4595 => x"91",
          4596 => x"58",
          4597 => x"09",
          4598 => x"38",
          4599 => x"08",
          4600 => x"26",
          4601 => x"78",
          4602 => x"79",
          4603 => x"78",
          4604 => x"86",
          4605 => x"82",
          4606 => x"06",
          4607 => x"83",
          4608 => x"91",
          4609 => x"27",
          4610 => x"8f",
          4611 => x"55",
          4612 => x"26",
          4613 => x"59",
          4614 => x"62",
          4615 => x"74",
          4616 => x"38",
          4617 => x"88",
          4618 => x"88",
          4619 => x"26",
          4620 => x"86",
          4621 => x"1a",
          4622 => x"79",
          4623 => x"38",
          4624 => x"80",
          4625 => x"2e",
          4626 => x"83",
          4627 => x"9f",
          4628 => x"8b",
          4629 => x"06",
          4630 => x"74",
          4631 => x"84",
          4632 => x"52",
          4633 => x"a2",
          4634 => x"53",
          4635 => x"52",
          4636 => x"a2",
          4637 => x"80",
          4638 => x"51",
          4639 => x"3f",
          4640 => x"34",
          4641 => x"ff",
          4642 => x"1b",
          4643 => x"a2",
          4644 => x"90",
          4645 => x"83",
          4646 => x"70",
          4647 => x"80",
          4648 => x"55",
          4649 => x"ff",
          4650 => x"66",
          4651 => x"ff",
          4652 => x"38",
          4653 => x"ff",
          4654 => x"1b",
          4655 => x"f2",
          4656 => x"74",
          4657 => x"51",
          4658 => x"3f",
          4659 => x"1c",
          4660 => x"98",
          4661 => x"a0",
          4662 => x"ff",
          4663 => x"51",
          4664 => x"3f",
          4665 => x"1b",
          4666 => x"e4",
          4667 => x"2e",
          4668 => x"80",
          4669 => x"88",
          4670 => x"80",
          4671 => x"ff",
          4672 => x"7c",
          4673 => x"51",
          4674 => x"3f",
          4675 => x"1b",
          4676 => x"bc",
          4677 => x"b0",
          4678 => x"a0",
          4679 => x"52",
          4680 => x"ff",
          4681 => x"ff",
          4682 => x"c0",
          4683 => x"0b",
          4684 => x"34",
          4685 => x"b8",
          4686 => x"c7",
          4687 => x"39",
          4688 => x"0a",
          4689 => x"51",
          4690 => x"3f",
          4691 => x"ff",
          4692 => x"1b",
          4693 => x"da",
          4694 => x"0b",
          4695 => x"a9",
          4696 => x"34",
          4697 => x"b8",
          4698 => x"1b",
          4699 => x"8f",
          4700 => x"d5",
          4701 => x"1b",
          4702 => x"ff",
          4703 => x"81",
          4704 => x"7a",
          4705 => x"ff",
          4706 => x"81",
          4707 => x"88",
          4708 => x"38",
          4709 => x"09",
          4710 => x"ee",
          4711 => x"60",
          4712 => x"7a",
          4713 => x"ff",
          4714 => x"84",
          4715 => x"52",
          4716 => x"9f",
          4717 => x"8b",
          4718 => x"52",
          4719 => x"9f",
          4720 => x"8a",
          4721 => x"52",
          4722 => x"51",
          4723 => x"3f",
          4724 => x"83",
          4725 => x"ff",
          4726 => x"82",
          4727 => x"1b",
          4728 => x"ec",
          4729 => x"d5",
          4730 => x"ff",
          4731 => x"75",
          4732 => x"05",
          4733 => x"7e",
          4734 => x"e5",
          4735 => x"60",
          4736 => x"52",
          4737 => x"9a",
          4738 => x"53",
          4739 => x"51",
          4740 => x"3f",
          4741 => x"58",
          4742 => x"09",
          4743 => x"38",
          4744 => x"51",
          4745 => x"3f",
          4746 => x"1b",
          4747 => x"a0",
          4748 => x"52",
          4749 => x"91",
          4750 => x"ff",
          4751 => x"81",
          4752 => x"f8",
          4753 => x"7a",
          4754 => x"84",
          4755 => x"61",
          4756 => x"26",
          4757 => x"57",
          4758 => x"53",
          4759 => x"51",
          4760 => x"3f",
          4761 => x"08",
          4762 => x"84",
          4763 => x"ca",
          4764 => x"7a",
          4765 => x"aa",
          4766 => x"75",
          4767 => x"56",
          4768 => x"81",
          4769 => x"80",
          4770 => x"38",
          4771 => x"83",
          4772 => x"63",
          4773 => x"74",
          4774 => x"38",
          4775 => x"54",
          4776 => x"52",
          4777 => x"99",
          4778 => x"ca",
          4779 => x"c1",
          4780 => x"75",
          4781 => x"56",
          4782 => x"8c",
          4783 => x"2e",
          4784 => x"56",
          4785 => x"ff",
          4786 => x"84",
          4787 => x"2e",
          4788 => x"56",
          4789 => x"58",
          4790 => x"38",
          4791 => x"77",
          4792 => x"ff",
          4793 => x"82",
          4794 => x"78",
          4795 => x"c2",
          4796 => x"1b",
          4797 => x"34",
          4798 => x"16",
          4799 => x"82",
          4800 => x"83",
          4801 => x"84",
          4802 => x"67",
          4803 => x"fd",
          4804 => x"51",
          4805 => x"3f",
          4806 => x"16",
          4807 => x"88",
          4808 => x"bf",
          4809 => x"86",
          4810 => x"ca",
          4811 => x"16",
          4812 => x"83",
          4813 => x"ff",
          4814 => x"66",
          4815 => x"1b",
          4816 => x"8c",
          4817 => x"77",
          4818 => x"7e",
          4819 => x"91",
          4820 => x"91",
          4821 => x"a2",
          4822 => x"80",
          4823 => x"ff",
          4824 => x"81",
          4825 => x"88",
          4826 => x"89",
          4827 => x"8a",
          4828 => x"86",
          4829 => x"88",
          4830 => x"91",
          4831 => x"99",
          4832 => x"ff",
          4833 => x"52",
          4834 => x"81",
          4835 => x"84",
          4836 => x"9c",
          4837 => x"08",
          4838 => x"d8",
          4839 => x"39",
          4840 => x"51",
          4841 => x"91",
          4842 => x"80",
          4843 => x"bc",
          4844 => x"eb",
          4845 => x"9c",
          4846 => x"39",
          4847 => x"51",
          4848 => x"91",
          4849 => x"80",
          4850 => x"bc",
          4851 => x"cf",
          4852 => x"e8",
          4853 => x"39",
          4854 => x"51",
          4855 => x"91",
          4856 => x"bb",
          4857 => x"b4",
          4858 => x"91",
          4859 => x"af",
          4860 => x"f4",
          4861 => x"91",
          4862 => x"a3",
          4863 => x"a8",
          4864 => x"91",
          4865 => x"97",
          4866 => x"d4",
          4867 => x"91",
          4868 => x"8b",
          4869 => x"84",
          4870 => x"91",
          4871 => x"ff",
          4872 => x"83",
          4873 => x"fb",
          4874 => x"79",
          4875 => x"87",
          4876 => x"38",
          4877 => x"87",
          4878 => x"91",
          4879 => x"52",
          4880 => x"f2",
          4881 => x"ca",
          4882 => x"75",
          4883 => x"98",
          4884 => x"88",
          4885 => x"53",
          4886 => x"bf",
          4887 => x"8d",
          4888 => x"3d",
          4889 => x"3d",
          4890 => x"61",
          4891 => x"80",
          4892 => x"73",
          4893 => x"5f",
          4894 => x"5c",
          4895 => x"52",
          4896 => x"51",
          4897 => x"3f",
          4898 => x"51",
          4899 => x"3f",
          4900 => x"77",
          4901 => x"38",
          4902 => x"89",
          4903 => x"2e",
          4904 => x"c6",
          4905 => x"53",
          4906 => x"8e",
          4907 => x"52",
          4908 => x"51",
          4909 => x"3f",
          4910 => x"bf",
          4911 => x"86",
          4912 => x"15",
          4913 => x"39",
          4914 => x"72",
          4915 => x"38",
          4916 => x"91",
          4917 => x"ff",
          4918 => x"89",
          4919 => x"d8",
          4920 => x"b9",
          4921 => x"55",
          4922 => x"16",
          4923 => x"27",
          4924 => x"33",
          4925 => x"e4",
          4926 => x"85",
          4927 => x"91",
          4928 => x"ff",
          4929 => x"81",
          4930 => x"51",
          4931 => x"3f",
          4932 => x"91",
          4933 => x"ff",
          4934 => x"80",
          4935 => x"27",
          4936 => x"16",
          4937 => x"72",
          4938 => x"53",
          4939 => x"90",
          4940 => x"2e",
          4941 => x"80",
          4942 => x"38",
          4943 => x"39",
          4944 => x"f9",
          4945 => x"15",
          4946 => x"91",
          4947 => x"ff",
          4948 => x"76",
          4949 => x"5a",
          4950 => x"92",
          4951 => x"88",
          4952 => x"70",
          4953 => x"55",
          4954 => x"09",
          4955 => x"38",
          4956 => x"3f",
          4957 => x"08",
          4958 => x"98",
          4959 => x"32",
          4960 => x"72",
          4961 => x"51",
          4962 => x"55",
          4963 => x"8c",
          4964 => x"38",
          4965 => x"09",
          4966 => x"38",
          4967 => x"39",
          4968 => x"72",
          4969 => x"d6",
          4970 => x"72",
          4971 => x"0c",
          4972 => x"04",
          4973 => x"66",
          4974 => x"80",
          4975 => x"69",
          4976 => x"74",
          4977 => x"70",
          4978 => x"27",
          4979 => x"58",
          4980 => x"93",
          4981 => x"fb",
          4982 => x"75",
          4983 => x"70",
          4984 => x"b9",
          4985 => x"88",
          4986 => x"ca",
          4987 => x"38",
          4988 => x"08",
          4989 => x"88",
          4990 => x"88",
          4991 => x"3d",
          4992 => x"84",
          4993 => x"52",
          4994 => x"f6",
          4995 => x"88",
          4996 => x"ca",
          4997 => x"38",
          4998 => x"80",
          4999 => x"74",
          5000 => x"59",
          5001 => x"96",
          5002 => x"51",
          5003 => x"75",
          5004 => x"07",
          5005 => x"55",
          5006 => x"95",
          5007 => x"2e",
          5008 => x"bf",
          5009 => x"c0",
          5010 => x"52",
          5011 => x"d7",
          5012 => x"76",
          5013 => x"0c",
          5014 => x"04",
          5015 => x"7b",
          5016 => x"b3",
          5017 => x"58",
          5018 => x"53",
          5019 => x"51",
          5020 => x"91",
          5021 => x"a4",
          5022 => x"2e",
          5023 => x"81",
          5024 => x"98",
          5025 => x"7f",
          5026 => x"88",
          5027 => x"7d",
          5028 => x"91",
          5029 => x"57",
          5030 => x"04",
          5031 => x"88",
          5032 => x"0d",
          5033 => x"0d",
          5034 => x"33",
          5035 => x"53",
          5036 => x"52",
          5037 => x"c9",
          5038 => x"88",
          5039 => x"80",
          5040 => x"c0",
          5041 => x"c0",
          5042 => x"c7",
          5043 => x"91",
          5044 => x"ff",
          5045 => x"74",
          5046 => x"38",
          5047 => x"3f",
          5048 => x"04",
          5049 => x"87",
          5050 => x"08",
          5051 => x"fd",
          5052 => x"fe",
          5053 => x"91",
          5054 => x"fe",
          5055 => x"80",
          5056 => x"fe",
          5057 => x"2a",
          5058 => x"51",
          5059 => x"2e",
          5060 => x"51",
          5061 => x"3f",
          5062 => x"51",
          5063 => x"3f",
          5064 => x"f5",
          5065 => x"82",
          5066 => x"06",
          5067 => x"80",
          5068 => x"81",
          5069 => x"ca",
          5070 => x"f4",
          5071 => x"c2",
          5072 => x"fe",
          5073 => x"72",
          5074 => x"81",
          5075 => x"71",
          5076 => x"38",
          5077 => x"f5",
          5078 => x"c1",
          5079 => x"f7",
          5080 => x"51",
          5081 => x"3f",
          5082 => x"70",
          5083 => x"52",
          5084 => x"95",
          5085 => x"fe",
          5086 => x"91",
          5087 => x"fe",
          5088 => x"80",
          5089 => x"fa",
          5090 => x"2a",
          5091 => x"51",
          5092 => x"2e",
          5093 => x"51",
          5094 => x"3f",
          5095 => x"51",
          5096 => x"3f",
          5097 => x"f4",
          5098 => x"86",
          5099 => x"06",
          5100 => x"80",
          5101 => x"81",
          5102 => x"c6",
          5103 => x"c0",
          5104 => x"be",
          5105 => x"fe",
          5106 => x"72",
          5107 => x"81",
          5108 => x"71",
          5109 => x"38",
          5110 => x"f4",
          5111 => x"c1",
          5112 => x"f6",
          5113 => x"51",
          5114 => x"3f",
          5115 => x"70",
          5116 => x"52",
          5117 => x"95",
          5118 => x"fe",
          5119 => x"91",
          5120 => x"fe",
          5121 => x"80",
          5122 => x"f6",
          5123 => x"a6",
          5124 => x"0d",
          5125 => x"0d",
          5126 => x"70",
          5127 => x"73",
          5128 => x"f0",
          5129 => x"73",
          5130 => x"15",
          5131 => x"e4",
          5132 => x"54",
          5133 => x"70",
          5134 => x"57",
          5135 => x"a0",
          5136 => x"81",
          5137 => x"2e",
          5138 => x"e5",
          5139 => x"ff",
          5140 => x"a0",
          5141 => x"06",
          5142 => x"74",
          5143 => x"56",
          5144 => x"75",
          5145 => x"c7",
          5146 => x"08",
          5147 => x"52",
          5148 => x"fd",
          5149 => x"88",
          5150 => x"84",
          5151 => x"72",
          5152 => x"a3",
          5153 => x"70",
          5154 => x"57",
          5155 => x"27",
          5156 => x"53",
          5157 => x"88",
          5158 => x"0d",
          5159 => x"0d",
          5160 => x"91",
          5161 => x"5e",
          5162 => x"7b",
          5163 => x"c8",
          5164 => x"88",
          5165 => x"06",
          5166 => x"2e",
          5167 => x"a2",
          5168 => x"a8",
          5169 => x"70",
          5170 => x"84",
          5171 => x"53",
          5172 => x"cb",
          5173 => x"b9",
          5174 => x"ca",
          5175 => x"2e",
          5176 => x"c2",
          5177 => x"d7",
          5178 => x"5e",
          5179 => x"e4",
          5180 => x"a9",
          5181 => x"70",
          5182 => x"f8",
          5183 => x"79",
          5184 => x"dc",
          5185 => x"52",
          5186 => x"84",
          5187 => x"3d",
          5188 => x"51",
          5189 => x"91",
          5190 => x"90",
          5191 => x"2c",
          5192 => x"80",
          5193 => x"da",
          5194 => x"c2",
          5195 => x"38",
          5196 => x"83",
          5197 => x"b0",
          5198 => x"78",
          5199 => x"a1",
          5200 => x"24",
          5201 => x"80",
          5202 => x"38",
          5203 => x"81",
          5204 => x"f1",
          5205 => x"2e",
          5206 => x"78",
          5207 => x"9c",
          5208 => x"39",
          5209 => x"85",
          5210 => x"bf",
          5211 => x"78",
          5212 => x"98",
          5213 => x"2e",
          5214 => x"8e",
          5215 => x"80",
          5216 => x"d9",
          5217 => x"c1",
          5218 => x"38",
          5219 => x"78",
          5220 => x"8d",
          5221 => x"80",
          5222 => x"38",
          5223 => x"2e",
          5224 => x"78",
          5225 => x"92",
          5226 => x"c3",
          5227 => x"38",
          5228 => x"2e",
          5229 => x"8e",
          5230 => x"80",
          5231 => x"c0",
          5232 => x"d5",
          5233 => x"38",
          5234 => x"78",
          5235 => x"8d",
          5236 => x"81",
          5237 => x"38",
          5238 => x"2e",
          5239 => x"78",
          5240 => x"8d",
          5241 => x"dd",
          5242 => x"85",
          5243 => x"38",
          5244 => x"2e",
          5245 => x"8d",
          5246 => x"3d",
          5247 => x"53",
          5248 => x"51",
          5249 => x"3f",
          5250 => x"08",
          5251 => x"c2",
          5252 => x"ab",
          5253 => x"fe",
          5254 => x"fe",
          5255 => x"ff",
          5256 => x"91",
          5257 => x"80",
          5258 => x"81",
          5259 => x"38",
          5260 => x"80",
          5261 => x"52",
          5262 => x"05",
          5263 => x"87",
          5264 => x"ca",
          5265 => x"ff",
          5266 => x"8e",
          5267 => x"f8",
          5268 => x"c9",
          5269 => x"fd",
          5270 => x"c3",
          5271 => x"b6",
          5272 => x"fe",
          5273 => x"fe",
          5274 => x"ff",
          5275 => x"91",
          5276 => x"80",
          5277 => x"38",
          5278 => x"52",
          5279 => x"05",
          5280 => x"8b",
          5281 => x"ca",
          5282 => x"91",
          5283 => x"8c",
          5284 => x"3d",
          5285 => x"53",
          5286 => x"51",
          5287 => x"3f",
          5288 => x"08",
          5289 => x"38",
          5290 => x"fc",
          5291 => x"3d",
          5292 => x"53",
          5293 => x"51",
          5294 => x"3f",
          5295 => x"08",
          5296 => x"ca",
          5297 => x"63",
          5298 => x"a8",
          5299 => x"ff",
          5300 => x"02",
          5301 => x"33",
          5302 => x"63",
          5303 => x"91",
          5304 => x"51",
          5305 => x"3f",
          5306 => x"08",
          5307 => x"91",
          5308 => x"fe",
          5309 => x"81",
          5310 => x"39",
          5311 => x"f8",
          5312 => x"ea",
          5313 => x"ca",
          5314 => x"3d",
          5315 => x"52",
          5316 => x"81",
          5317 => x"91",
          5318 => x"52",
          5319 => x"94",
          5320 => x"39",
          5321 => x"f8",
          5322 => x"ea",
          5323 => x"ca",
          5324 => x"3d",
          5325 => x"52",
          5326 => x"d9",
          5327 => x"88",
          5328 => x"fe",
          5329 => x"5a",
          5330 => x"3f",
          5331 => x"08",
          5332 => x"f8",
          5333 => x"fe",
          5334 => x"91",
          5335 => x"91",
          5336 => x"80",
          5337 => x"91",
          5338 => x"81",
          5339 => x"78",
          5340 => x"7a",
          5341 => x"3f",
          5342 => x"08",
          5343 => x"ed",
          5344 => x"88",
          5345 => x"fb",
          5346 => x"39",
          5347 => x"f4",
          5348 => x"f8",
          5349 => x"80",
          5350 => x"ca",
          5351 => x"2e",
          5352 => x"b7",
          5353 => x"11",
          5354 => x"05",
          5355 => x"c6",
          5356 => x"88",
          5357 => x"fa",
          5358 => x"3d",
          5359 => x"53",
          5360 => x"51",
          5361 => x"3f",
          5362 => x"08",
          5363 => x"ca",
          5364 => x"91",
          5365 => x"fe",
          5366 => x"63",
          5367 => x"79",
          5368 => x"f2",
          5369 => x"78",
          5370 => x"05",
          5371 => x"7a",
          5372 => x"81",
          5373 => x"3d",
          5374 => x"53",
          5375 => x"51",
          5376 => x"3f",
          5377 => x"08",
          5378 => x"e1",
          5379 => x"fe",
          5380 => x"fe",
          5381 => x"fe",
          5382 => x"91",
          5383 => x"80",
          5384 => x"38",
          5385 => x"ec",
          5386 => x"f8",
          5387 => x"ff",
          5388 => x"ca",
          5389 => x"2e",
          5390 => x"91",
          5391 => x"fe",
          5392 => x"63",
          5393 => x"27",
          5394 => x"61",
          5395 => x"81",
          5396 => x"79",
          5397 => x"05",
          5398 => x"b7",
          5399 => x"11",
          5400 => x"05",
          5401 => x"8e",
          5402 => x"88",
          5403 => x"f8",
          5404 => x"3d",
          5405 => x"53",
          5406 => x"51",
          5407 => x"3f",
          5408 => x"08",
          5409 => x"e5",
          5410 => x"fe",
          5411 => x"fe",
          5412 => x"fe",
          5413 => x"91",
          5414 => x"80",
          5415 => x"38",
          5416 => x"51",
          5417 => x"3f",
          5418 => x"63",
          5419 => x"61",
          5420 => x"33",
          5421 => x"78",
          5422 => x"38",
          5423 => x"54",
          5424 => x"79",
          5425 => x"d4",
          5426 => x"b5",
          5427 => x"62",
          5428 => x"5a",
          5429 => x"c2",
          5430 => x"ba",
          5431 => x"fe",
          5432 => x"fe",
          5433 => x"fe",
          5434 => x"91",
          5435 => x"80",
          5436 => x"c7",
          5437 => x"78",
          5438 => x"38",
          5439 => x"08",
          5440 => x"91",
          5441 => x"59",
          5442 => x"88",
          5443 => x"ec",
          5444 => x"39",
          5445 => x"33",
          5446 => x"38",
          5447 => x"33",
          5448 => x"2e",
          5449 => x"c6",
          5450 => x"89",
          5451 => x"84",
          5452 => x"05",
          5453 => x"fe",
          5454 => x"fe",
          5455 => x"fe",
          5456 => x"91",
          5457 => x"80",
          5458 => x"c7",
          5459 => x"78",
          5460 => x"38",
          5461 => x"08",
          5462 => x"91",
          5463 => x"59",
          5464 => x"88",
          5465 => x"f0",
          5466 => x"39",
          5467 => x"33",
          5468 => x"38",
          5469 => x"33",
          5470 => x"2e",
          5471 => x"c6",
          5472 => x"88",
          5473 => x"84",
          5474 => x"43",
          5475 => x"ec",
          5476 => x"f8",
          5477 => x"fc",
          5478 => x"ca",
          5479 => x"2e",
          5480 => x"62",
          5481 => x"88",
          5482 => x"81",
          5483 => x"2e",
          5484 => x"80",
          5485 => x"79",
          5486 => x"38",
          5487 => x"c3",
          5488 => x"f4",
          5489 => x"55",
          5490 => x"53",
          5491 => x"51",
          5492 => x"91",
          5493 => x"84",
          5494 => x"3d",
          5495 => x"53",
          5496 => x"51",
          5497 => x"3f",
          5498 => x"08",
          5499 => x"fd",
          5500 => x"fe",
          5501 => x"fe",
          5502 => x"fe",
          5503 => x"91",
          5504 => x"80",
          5505 => x"63",
          5506 => x"cb",
          5507 => x"34",
          5508 => x"44",
          5509 => x"f0",
          5510 => x"f8",
          5511 => x"fb",
          5512 => x"ca",
          5513 => x"38",
          5514 => x"63",
          5515 => x"52",
          5516 => x"51",
          5517 => x"3f",
          5518 => x"79",
          5519 => x"9b",
          5520 => x"79",
          5521 => x"ae",
          5522 => x"38",
          5523 => x"a0",
          5524 => x"fe",
          5525 => x"fe",
          5526 => x"fe",
          5527 => x"91",
          5528 => x"80",
          5529 => x"63",
          5530 => x"cb",
          5531 => x"34",
          5532 => x"44",
          5533 => x"91",
          5534 => x"fe",
          5535 => x"ff",
          5536 => x"3d",
          5537 => x"53",
          5538 => x"51",
          5539 => x"3f",
          5540 => x"08",
          5541 => x"d5",
          5542 => x"fe",
          5543 => x"fe",
          5544 => x"fe",
          5545 => x"91",
          5546 => x"80",
          5547 => x"60",
          5548 => x"05",
          5549 => x"82",
          5550 => x"78",
          5551 => x"fe",
          5552 => x"fe",
          5553 => x"fe",
          5554 => x"91",
          5555 => x"df",
          5556 => x"39",
          5557 => x"54",
          5558 => x"a0",
          5559 => x"a1",
          5560 => x"52",
          5561 => x"f8",
          5562 => x"45",
          5563 => x"78",
          5564 => x"f9",
          5565 => x"26",
          5566 => x"84",
          5567 => x"39",
          5568 => x"e4",
          5569 => x"f8",
          5570 => x"fb",
          5571 => x"ca",
          5572 => x"2e",
          5573 => x"59",
          5574 => x"22",
          5575 => x"05",
          5576 => x"41",
          5577 => x"91",
          5578 => x"fe",
          5579 => x"ff",
          5580 => x"3d",
          5581 => x"53",
          5582 => x"51",
          5583 => x"3f",
          5584 => x"08",
          5585 => x"a5",
          5586 => x"fe",
          5587 => x"fe",
          5588 => x"fe",
          5589 => x"91",
          5590 => x"80",
          5591 => x"60",
          5592 => x"59",
          5593 => x"41",
          5594 => x"e4",
          5595 => x"f8",
          5596 => x"fa",
          5597 => x"ca",
          5598 => x"38",
          5599 => x"60",
          5600 => x"52",
          5601 => x"51",
          5602 => x"3f",
          5603 => x"79",
          5604 => x"c7",
          5605 => x"79",
          5606 => x"ae",
          5607 => x"38",
          5608 => x"a8",
          5609 => x"fe",
          5610 => x"fe",
          5611 => x"fe",
          5612 => x"91",
          5613 => x"80",
          5614 => x"7f",
          5615 => x"91",
          5616 => x"fe",
          5617 => x"60",
          5618 => x"59",
          5619 => x"41",
          5620 => x"91",
          5621 => x"fe",
          5622 => x"ff",
          5623 => x"c4",
          5624 => x"f0",
          5625 => x"51",
          5626 => x"3f",
          5627 => x"91",
          5628 => x"fe",
          5629 => x"a2",
          5630 => x"f9",
          5631 => x"39",
          5632 => x"0b",
          5633 => x"84",
          5634 => x"81",
          5635 => x"94",
          5636 => x"c4",
          5637 => x"f0",
          5638 => x"d1",
          5639 => x"fc",
          5640 => x"f9",
          5641 => x"83",
          5642 => x"94",
          5643 => x"80",
          5644 => x"c0",
          5645 => x"f1",
          5646 => x"3d",
          5647 => x"53",
          5648 => x"51",
          5649 => x"3f",
          5650 => x"08",
          5651 => x"9d",
          5652 => x"91",
          5653 => x"fe",
          5654 => x"63",
          5655 => x"b7",
          5656 => x"11",
          5657 => x"05",
          5658 => x"8a",
          5659 => x"88",
          5660 => x"f0",
          5661 => x"52",
          5662 => x"51",
          5663 => x"3f",
          5664 => x"2d",
          5665 => x"08",
          5666 => x"88",
          5667 => x"f0",
          5668 => x"ca",
          5669 => x"91",
          5670 => x"fe",
          5671 => x"f0",
          5672 => x"c5",
          5673 => x"ee",
          5674 => x"ce",
          5675 => x"bd",
          5676 => x"80",
          5677 => x"e5",
          5678 => x"ff",
          5679 => x"ea",
          5680 => x"a9",
          5681 => x"33",
          5682 => x"80",
          5683 => x"38",
          5684 => x"80",
          5685 => x"80",
          5686 => x"38",
          5687 => x"f8",
          5688 => x"de",
          5689 => x"c6",
          5690 => x"ca",
          5691 => x"91",
          5692 => x"80",
          5693 => x"9c",
          5694 => x"70",
          5695 => x"f4",
          5696 => x"c6",
          5697 => x"ca",
          5698 => x"56",
          5699 => x"46",
          5700 => x"80",
          5701 => x"0a",
          5702 => x"0a",
          5703 => x"ea",
          5704 => x"ca",
          5705 => x"7c",
          5706 => x"81",
          5707 => x"78",
          5708 => x"ff",
          5709 => x"06",
          5710 => x"91",
          5711 => x"fe",
          5712 => x"ef",
          5713 => x"3d",
          5714 => x"91",
          5715 => x"90",
          5716 => x"91",
          5717 => x"90",
          5718 => x"91",
          5719 => x"fe",
          5720 => x"fe",
          5721 => x"91",
          5722 => x"fe",
          5723 => x"91",
          5724 => x"fe",
          5725 => x"91",
          5726 => x"fe",
          5727 => x"81",
          5728 => x"3f",
          5729 => x"80",
          5730 => x"0f",
          5731 => x"0f",
          5732 => x"0f",
          5733 => x"0f",
          5734 => x"0f",
          5735 => x"4c",
          5736 => x"4b",
          5737 => x"4b",
          5738 => x"4b",
          5739 => x"4b",
          5740 => x"4b",
          5741 => x"4b",
          5742 => x"4b",
          5743 => x"4b",
          5744 => x"4b",
          5745 => x"4b",
          5746 => x"4b",
          5747 => x"4b",
          5748 => x"4b",
          5749 => x"4b",
          5750 => x"4b",
          5751 => x"4b",
          5752 => x"4c",
          5753 => x"4c",
          5754 => x"4c",
          5755 => x"2f",
          5756 => x"25",
          5757 => x"64",
          5758 => x"3a",
          5759 => x"25",
          5760 => x"0a",
          5761 => x"43",
          5762 => x"6e",
          5763 => x"75",
          5764 => x"69",
          5765 => x"00",
          5766 => x"66",
          5767 => x"20",
          5768 => x"20",
          5769 => x"66",
          5770 => x"00",
          5771 => x"44",
          5772 => x"63",
          5773 => x"69",
          5774 => x"65",
          5775 => x"74",
          5776 => x"0a",
          5777 => x"20",
          5778 => x"53",
          5779 => x"52",
          5780 => x"28",
          5781 => x"72",
          5782 => x"30",
          5783 => x"20",
          5784 => x"65",
          5785 => x"38",
          5786 => x"0a",
          5787 => x"20",
          5788 => x"41",
          5789 => x"53",
          5790 => x"74",
          5791 => x"38",
          5792 => x"53",
          5793 => x"3d",
          5794 => x"58",
          5795 => x"00",
          5796 => x"20",
          5797 => x"4d",
          5798 => x"74",
          5799 => x"3d",
          5800 => x"58",
          5801 => x"69",
          5802 => x"25",
          5803 => x"29",
          5804 => x"00",
          5805 => x"20",
          5806 => x"43",
          5807 => x"00",
          5808 => x"20",
          5809 => x"32",
          5810 => x"00",
          5811 => x"20",
          5812 => x"49",
          5813 => x"00",
          5814 => x"20",
          5815 => x"20",
          5816 => x"64",
          5817 => x"65",
          5818 => x"65",
          5819 => x"30",
          5820 => x"2e",
          5821 => x"00",
          5822 => x"20",
          5823 => x"54",
          5824 => x"55",
          5825 => x"43",
          5826 => x"52",
          5827 => x"45",
          5828 => x"00",
          5829 => x"20",
          5830 => x"4d",
          5831 => x"20",
          5832 => x"6d",
          5833 => x"3d",
          5834 => x"58",
          5835 => x"00",
          5836 => x"64",
          5837 => x"73",
          5838 => x"0a",
          5839 => x"20",
          5840 => x"55",
          5841 => x"73",
          5842 => x"56",
          5843 => x"6f",
          5844 => x"64",
          5845 => x"73",
          5846 => x"20",
          5847 => x"58",
          5848 => x"00",
          5849 => x"20",
          5850 => x"55",
          5851 => x"6d",
          5852 => x"20",
          5853 => x"72",
          5854 => x"64",
          5855 => x"73",
          5856 => x"20",
          5857 => x"58",
          5858 => x"00",
          5859 => x"20",
          5860 => x"61",
          5861 => x"53",
          5862 => x"74",
          5863 => x"64",
          5864 => x"73",
          5865 => x"20",
          5866 => x"20",
          5867 => x"58",
          5868 => x"00",
          5869 => x"20",
          5870 => x"55",
          5871 => x"20",
          5872 => x"20",
          5873 => x"20",
          5874 => x"20",
          5875 => x"20",
          5876 => x"20",
          5877 => x"58",
          5878 => x"00",
          5879 => x"20",
          5880 => x"73",
          5881 => x"20",
          5882 => x"63",
          5883 => x"72",
          5884 => x"20",
          5885 => x"20",
          5886 => x"20",
          5887 => x"58",
          5888 => x"00",
          5889 => x"61",
          5890 => x"00",
          5891 => x"64",
          5892 => x"00",
          5893 => x"65",
          5894 => x"00",
          5895 => x"4f",
          5896 => x"4f",
          5897 => x"00",
          5898 => x"6b",
          5899 => x"6e",
          5900 => x"00",
          5901 => x"2b",
          5902 => x"3c",
          5903 => x"5b",
          5904 => x"00",
          5905 => x"54",
          5906 => x"54",
          5907 => x"00",
          5908 => x"90",
          5909 => x"4f",
          5910 => x"30",
          5911 => x"20",
          5912 => x"45",
          5913 => x"20",
          5914 => x"33",
          5915 => x"20",
          5916 => x"20",
          5917 => x"45",
          5918 => x"20",
          5919 => x"20",
          5920 => x"20",
          5921 => x"5c",
          5922 => x"00",
          5923 => x"00",
          5924 => x"00",
          5925 => x"45",
          5926 => x"8f",
          5927 => x"45",
          5928 => x"8e",
          5929 => x"92",
          5930 => x"55",
          5931 => x"9a",
          5932 => x"9e",
          5933 => x"4f",
          5934 => x"a6",
          5935 => x"aa",
          5936 => x"ae",
          5937 => x"b2",
          5938 => x"b6",
          5939 => x"ba",
          5940 => x"be",
          5941 => x"c2",
          5942 => x"c6",
          5943 => x"ca",
          5944 => x"ce",
          5945 => x"d2",
          5946 => x"d6",
          5947 => x"da",
          5948 => x"de",
          5949 => x"e2",
          5950 => x"e6",
          5951 => x"ea",
          5952 => x"ee",
          5953 => x"f2",
          5954 => x"f6",
          5955 => x"fa",
          5956 => x"fe",
          5957 => x"2c",
          5958 => x"5d",
          5959 => x"2a",
          5960 => x"3f",
          5961 => x"00",
          5962 => x"00",
          5963 => x"00",
          5964 => x"02",
          5965 => x"00",
          5966 => x"00",
          5967 => x"00",
          5968 => x"00",
          5969 => x"00",
          5970 => x"6e",
          5971 => x"00",
          5972 => x"6f",
          5973 => x"00",
          5974 => x"6e",
          5975 => x"00",
          5976 => x"6f",
          5977 => x"00",
          5978 => x"78",
          5979 => x"00",
          5980 => x"6c",
          5981 => x"00",
          5982 => x"6f",
          5983 => x"00",
          5984 => x"69",
          5985 => x"00",
          5986 => x"75",
          5987 => x"00",
          5988 => x"62",
          5989 => x"68",
          5990 => x"77",
          5991 => x"64",
          5992 => x"65",
          5993 => x"64",
          5994 => x"65",
          5995 => x"6c",
          5996 => x"00",
          5997 => x"70",
          5998 => x"73",
          5999 => x"74",
          6000 => x"73",
          6001 => x"00",
          6002 => x"66",
          6003 => x"00",
          6004 => x"73",
          6005 => x"00",
          6006 => x"73",
          6007 => x"72",
          6008 => x"0a",
          6009 => x"74",
          6010 => x"61",
          6011 => x"72",
          6012 => x"2e",
          6013 => x"00",
          6014 => x"73",
          6015 => x"6f",
          6016 => x"65",
          6017 => x"2e",
          6018 => x"00",
          6019 => x"20",
          6020 => x"65",
          6021 => x"75",
          6022 => x"0a",
          6023 => x"20",
          6024 => x"68",
          6025 => x"75",
          6026 => x"0a",
          6027 => x"76",
          6028 => x"64",
          6029 => x"6c",
          6030 => x"6d",
          6031 => x"00",
          6032 => x"63",
          6033 => x"20",
          6034 => x"69",
          6035 => x"0a",
          6036 => x"6c",
          6037 => x"6c",
          6038 => x"64",
          6039 => x"78",
          6040 => x"73",
          6041 => x"00",
          6042 => x"6c",
          6043 => x"61",
          6044 => x"65",
          6045 => x"76",
          6046 => x"64",
          6047 => x"00",
          6048 => x"20",
          6049 => x"77",
          6050 => x"65",
          6051 => x"6f",
          6052 => x"74",
          6053 => x"0a",
          6054 => x"69",
          6055 => x"6e",
          6056 => x"65",
          6057 => x"73",
          6058 => x"76",
          6059 => x"64",
          6060 => x"00",
          6061 => x"73",
          6062 => x"6f",
          6063 => x"6e",
          6064 => x"65",
          6065 => x"00",
          6066 => x"20",
          6067 => x"70",
          6068 => x"62",
          6069 => x"66",
          6070 => x"73",
          6071 => x"65",
          6072 => x"6f",
          6073 => x"20",
          6074 => x"64",
          6075 => x"2e",
          6076 => x"00",
          6077 => x"72",
          6078 => x"20",
          6079 => x"72",
          6080 => x"2e",
          6081 => x"00",
          6082 => x"6d",
          6083 => x"74",
          6084 => x"70",
          6085 => x"74",
          6086 => x"20",
          6087 => x"63",
          6088 => x"65",
          6089 => x"00",
          6090 => x"6c",
          6091 => x"73",
          6092 => x"63",
          6093 => x"2e",
          6094 => x"00",
          6095 => x"73",
          6096 => x"69",
          6097 => x"6e",
          6098 => x"65",
          6099 => x"79",
          6100 => x"00",
          6101 => x"6f",
          6102 => x"6e",
          6103 => x"70",
          6104 => x"66",
          6105 => x"73",
          6106 => x"00",
          6107 => x"72",
          6108 => x"74",
          6109 => x"20",
          6110 => x"6f",
          6111 => x"63",
          6112 => x"00",
          6113 => x"63",
          6114 => x"73",
          6115 => x"00",
          6116 => x"6b",
          6117 => x"6e",
          6118 => x"72",
          6119 => x"0a",
          6120 => x"6c",
          6121 => x"79",
          6122 => x"20",
          6123 => x"61",
          6124 => x"6c",
          6125 => x"79",
          6126 => x"2f",
          6127 => x"2e",
          6128 => x"00",
          6129 => x"38",
          6130 => x"00",
          6131 => x"20",
          6132 => x"34",
          6133 => x"00",
          6134 => x"20",
          6135 => x"20",
          6136 => x"00",
          6137 => x"32",
          6138 => x"00",
          6139 => x"00",
          6140 => x"00",
          6141 => x"0a",
          6142 => x"61",
          6143 => x"00",
          6144 => x"55",
          6145 => x"00",
          6146 => x"2a",
          6147 => x"20",
          6148 => x"00",
          6149 => x"2f",
          6150 => x"32",
          6151 => x"00",
          6152 => x"2e",
          6153 => x"00",
          6154 => x"50",
          6155 => x"72",
          6156 => x"25",
          6157 => x"29",
          6158 => x"20",
          6159 => x"2a",
          6160 => x"00",
          6161 => x"55",
          6162 => x"49",
          6163 => x"72",
          6164 => x"74",
          6165 => x"6e",
          6166 => x"72",
          6167 => x"00",
          6168 => x"6d",
          6169 => x"69",
          6170 => x"72",
          6171 => x"74",
          6172 => x"00",
          6173 => x"32",
          6174 => x"74",
          6175 => x"75",
          6176 => x"00",
          6177 => x"43",
          6178 => x"52",
          6179 => x"6e",
          6180 => x"72",
          6181 => x"0a",
          6182 => x"43",
          6183 => x"57",
          6184 => x"6e",
          6185 => x"72",
          6186 => x"0a",
          6187 => x"52",
          6188 => x"52",
          6189 => x"6e",
          6190 => x"72",
          6191 => x"0a",
          6192 => x"52",
          6193 => x"54",
          6194 => x"6e",
          6195 => x"72",
          6196 => x"0a",
          6197 => x"52",
          6198 => x"52",
          6199 => x"6e",
          6200 => x"72",
          6201 => x"0a",
          6202 => x"52",
          6203 => x"54",
          6204 => x"6e",
          6205 => x"72",
          6206 => x"0a",
          6207 => x"74",
          6208 => x"67",
          6209 => x"20",
          6210 => x"65",
          6211 => x"2e",
          6212 => x"00",
          6213 => x"61",
          6214 => x"6e",
          6215 => x"69",
          6216 => x"2e",
          6217 => x"00",
          6218 => x"00",
          6219 => x"69",
          6220 => x"20",
          6221 => x"69",
          6222 => x"69",
          6223 => x"73",
          6224 => x"64",
          6225 => x"72",
          6226 => x"2c",
          6227 => x"65",
          6228 => x"20",
          6229 => x"74",
          6230 => x"6e",
          6231 => x"6c",
          6232 => x"00",
          6233 => x"00",
          6234 => x"64",
          6235 => x"73",
          6236 => x"64",
          6237 => x"00",
          6238 => x"69",
          6239 => x"6c",
          6240 => x"64",
          6241 => x"00",
          6242 => x"69",
          6243 => x"20",
          6244 => x"69",
          6245 => x"69",
          6246 => x"73",
          6247 => x"00",
          6248 => x"3d",
          6249 => x"00",
          6250 => x"3a",
          6251 => x"65",
          6252 => x"6e",
          6253 => x"2e",
          6254 => x"70",
          6255 => x"67",
          6256 => x"00",
          6257 => x"6d",
          6258 => x"69",
          6259 => x"2e",
          6260 => x"00",
          6261 => x"38",
          6262 => x"25",
          6263 => x"29",
          6264 => x"30",
          6265 => x"28",
          6266 => x"78",
          6267 => x"00",
          6268 => x"6d",
          6269 => x"65",
          6270 => x"79",
          6271 => x"00",
          6272 => x"6f",
          6273 => x"65",
          6274 => x"0a",
          6275 => x"38",
          6276 => x"30",
          6277 => x"00",
          6278 => x"3f",
          6279 => x"00",
          6280 => x"38",
          6281 => x"30",
          6282 => x"00",
          6283 => x"38",
          6284 => x"30",
          6285 => x"00",
          6286 => x"73",
          6287 => x"69",
          6288 => x"69",
          6289 => x"72",
          6290 => x"74",
          6291 => x"00",
          6292 => x"61",
          6293 => x"6e",
          6294 => x"6e",
          6295 => x"72",
          6296 => x"73",
          6297 => x"00",
          6298 => x"73",
          6299 => x"65",
          6300 => x"61",
          6301 => x"66",
          6302 => x"0a",
          6303 => x"61",
          6304 => x"6e",
          6305 => x"61",
          6306 => x"66",
          6307 => x"0a",
          6308 => x"65",
          6309 => x"69",
          6310 => x"63",
          6311 => x"20",
          6312 => x"30",
          6313 => x"2e",
          6314 => x"00",
          6315 => x"6c",
          6316 => x"67",
          6317 => x"64",
          6318 => x"20",
          6319 => x"78",
          6320 => x"2e",
          6321 => x"00",
          6322 => x"6c",
          6323 => x"65",
          6324 => x"6e",
          6325 => x"63",
          6326 => x"20",
          6327 => x"29",
          6328 => x"00",
          6329 => x"73",
          6330 => x"74",
          6331 => x"20",
          6332 => x"6c",
          6333 => x"74",
          6334 => x"2e",
          6335 => x"00",
          6336 => x"6c",
          6337 => x"65",
          6338 => x"74",
          6339 => x"2e",
          6340 => x"00",
          6341 => x"55",
          6342 => x"6e",
          6343 => x"3a",
          6344 => x"5c",
          6345 => x"25",
          6346 => x"00",
          6347 => x"64",
          6348 => x"6d",
          6349 => x"64",
          6350 => x"00",
          6351 => x"6e",
          6352 => x"67",
          6353 => x"0a",
          6354 => x"61",
          6355 => x"6e",
          6356 => x"6e",
          6357 => x"72",
          6358 => x"73",
          6359 => x"0a",
          6360 => x"00",
          6361 => x"00",
          6362 => x"7f",
          6363 => x"00",
          6364 => x"7f",
          6365 => x"00",
          6366 => x"7f",
          6367 => x"00",
          6368 => x"00",
          6369 => x"78",
          6370 => x"00",
          6371 => x"e1",
          6372 => x"01",
          6373 => x"01",
          6374 => x"01",
          6375 => x"00",
          6376 => x"00",
          6377 => x"00",
          6378 => x"5d",
          6379 => x"01",
          6380 => x"00",
          6381 => x"00",
          6382 => x"5d",
          6383 => x"01",
          6384 => x"00",
          6385 => x"00",
          6386 => x"5d",
          6387 => x"03",
          6388 => x"00",
          6389 => x"00",
          6390 => x"5d",
          6391 => x"03",
          6392 => x"00",
          6393 => x"00",
          6394 => x"5d",
          6395 => x"03",
          6396 => x"00",
          6397 => x"00",
          6398 => x"5d",
          6399 => x"04",
          6400 => x"00",
          6401 => x"00",
          6402 => x"5d",
          6403 => x"04",
          6404 => x"00",
          6405 => x"00",
          6406 => x"5d",
          6407 => x"04",
          6408 => x"00",
          6409 => x"00",
          6410 => x"5d",
          6411 => x"04",
          6412 => x"00",
          6413 => x"00",
          6414 => x"5d",
          6415 => x"04",
          6416 => x"00",
          6417 => x"00",
          6418 => x"5d",
          6419 => x"04",
          6420 => x"00",
          6421 => x"00",
          6422 => x"5d",
          6423 => x"04",
          6424 => x"00",
          6425 => x"00",
          6426 => x"5d",
          6427 => x"05",
          6428 => x"00",
          6429 => x"00",
          6430 => x"5d",
          6431 => x"05",
          6432 => x"00",
          6433 => x"00",
          6434 => x"5d",
          6435 => x"05",
          6436 => x"00",
          6437 => x"00",
          6438 => x"5d",
          6439 => x"05",
          6440 => x"00",
          6441 => x"00",
          6442 => x"5d",
          6443 => x"07",
          6444 => x"00",
          6445 => x"00",
          6446 => x"5d",
          6447 => x"07",
          6448 => x"00",
          6449 => x"00",
          6450 => x"5d",
          6451 => x"08",
          6452 => x"00",
          6453 => x"00",
          6454 => x"5d",
          6455 => x"08",
          6456 => x"00",
          6457 => x"00",
          6458 => x"5d",
          6459 => x"08",
          6460 => x"00",
          6461 => x"00",
          6462 => x"5d",
          6463 => x"08",
          6464 => x"00",
          6465 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"8a",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"84",
            11 => x"0b",
            12 => x"04",
            13 => x"84",
            14 => x"0b",
            15 => x"04",
            16 => x"84",
            17 => x"0b",
            18 => x"04",
            19 => x"84",
            20 => x"0b",
            21 => x"04",
            22 => x"85",
            23 => x"0b",
            24 => x"04",
            25 => x"85",
            26 => x"0b",
            27 => x"04",
            28 => x"85",
            29 => x"0b",
            30 => x"04",
            31 => x"85",
            32 => x"0b",
            33 => x"04",
            34 => x"86",
            35 => x"0b",
            36 => x"04",
            37 => x"86",
            38 => x"0b",
            39 => x"04",
            40 => x"86",
            41 => x"0b",
            42 => x"04",
            43 => x"86",
            44 => x"0b",
            45 => x"04",
            46 => x"87",
            47 => x"0b",
            48 => x"04",
            49 => x"87",
            50 => x"0b",
            51 => x"04",
            52 => x"87",
            53 => x"0b",
            54 => x"04",
            55 => x"88",
            56 => x"0b",
            57 => x"04",
            58 => x"88",
            59 => x"0b",
            60 => x"04",
            61 => x"88",
            62 => x"0b",
            63 => x"04",
            64 => x"88",
            65 => x"0b",
            66 => x"04",
            67 => x"89",
            68 => x"0b",
            69 => x"04",
            70 => x"89",
            71 => x"0b",
            72 => x"04",
            73 => x"89",
            74 => x"0b",
            75 => x"04",
            76 => x"89",
            77 => x"0b",
            78 => x"04",
            79 => x"8a",
            80 => x"0b",
            81 => x"04",
            82 => x"8a",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"90",
           129 => x"91",
           130 => x"90",
           131 => x"91",
           132 => x"88",
           133 => x"04",
           134 => x"0c",
           135 => x"2d",
           136 => x"08",
           137 => x"90",
           138 => x"94",
           139 => x"fe",
           140 => x"94",
           141 => x"80",
           142 => x"ca",
           143 => x"a0",
           144 => x"ca",
           145 => x"c0",
           146 => x"91",
           147 => x"90",
           148 => x"91",
           149 => x"88",
           150 => x"04",
           151 => x"0c",
           152 => x"2d",
           153 => x"08",
           154 => x"90",
           155 => x"94",
           156 => x"bf",
           157 => x"94",
           158 => x"80",
           159 => x"ca",
           160 => x"a7",
           161 => x"ca",
           162 => x"c0",
           163 => x"91",
           164 => x"90",
           165 => x"91",
           166 => x"88",
           167 => x"04",
           168 => x"0c",
           169 => x"2d",
           170 => x"08",
           171 => x"90",
           172 => x"94",
           173 => x"96",
           174 => x"94",
           175 => x"80",
           176 => x"ca",
           177 => x"a6",
           178 => x"ca",
           179 => x"c0",
           180 => x"91",
           181 => x"90",
           182 => x"91",
           183 => x"88",
           184 => x"04",
           185 => x"0c",
           186 => x"2d",
           187 => x"08",
           188 => x"90",
           189 => x"94",
           190 => x"89",
           191 => x"94",
           192 => x"80",
           193 => x"ca",
           194 => x"91",
           195 => x"ca",
           196 => x"c0",
           197 => x"91",
           198 => x"90",
           199 => x"91",
           200 => x"88",
           201 => x"04",
           202 => x"0c",
           203 => x"2d",
           204 => x"08",
           205 => x"90",
           206 => x"94",
           207 => x"8d",
           208 => x"94",
           209 => x"80",
           210 => x"ca",
           211 => x"e1",
           212 => x"ca",
           213 => x"c0",
           214 => x"91",
           215 => x"90",
           216 => x"91",
           217 => x"88",
           218 => x"04",
           219 => x"0c",
           220 => x"2d",
           221 => x"08",
           222 => x"90",
           223 => x"94",
           224 => x"fc",
           225 => x"94",
           226 => x"80",
           227 => x"ca",
           228 => x"e7",
           229 => x"ca",
           230 => x"c0",
           231 => x"91",
           232 => x"90",
           233 => x"91",
           234 => x"88",
           235 => x"04",
           236 => x"0c",
           237 => x"2d",
           238 => x"08",
           239 => x"90",
           240 => x"94",
           241 => x"f9",
           242 => x"94",
           243 => x"80",
           244 => x"ca",
           245 => x"fa",
           246 => x"ca",
           247 => x"c0",
           248 => x"91",
           249 => x"90",
           250 => x"91",
           251 => x"88",
           252 => x"04",
           253 => x"0c",
           254 => x"2d",
           255 => x"08",
           256 => x"90",
           257 => x"94",
           258 => x"fd",
           259 => x"94",
           260 => x"80",
           261 => x"ca",
           262 => x"80",
           263 => x"ca",
           264 => x"c0",
           265 => x"91",
           266 => x"91",
           267 => x"91",
           268 => x"88",
           269 => x"04",
           270 => x"0c",
           271 => x"2d",
           272 => x"08",
           273 => x"90",
           274 => x"94",
           275 => x"c6",
           276 => x"94",
           277 => x"80",
           278 => x"ca",
           279 => x"ea",
           280 => x"ca",
           281 => x"c0",
           282 => x"91",
           283 => x"90",
           284 => x"91",
           285 => x"88",
           286 => x"04",
           287 => x"0c",
           288 => x"2d",
           289 => x"08",
           290 => x"90",
           291 => x"94",
           292 => x"b3",
           293 => x"94",
           294 => x"80",
           295 => x"ca",
           296 => x"87",
           297 => x"ca",
           298 => x"c0",
           299 => x"91",
           300 => x"90",
           301 => x"91",
           302 => x"88",
           303 => x"04",
           304 => x"0c",
           305 => x"2d",
           306 => x"08",
           307 => x"90",
           308 => x"94",
           309 => x"f6",
           310 => x"94",
           311 => x"80",
           312 => x"ca",
           313 => x"ae",
           314 => x"ca",
           315 => x"c0",
           316 => x"91",
           317 => x"90",
           318 => x"91",
           319 => x"88",
           320 => x"04",
           321 => x"0c",
           322 => x"2d",
           323 => x"08",
           324 => x"90",
           325 => x"94",
           326 => x"94",
           327 => x"94",
           328 => x"80",
           329 => x"ca",
           330 => x"94",
           331 => x"ca",
           332 => x"c0",
           333 => x"91",
           334 => x"91",
           335 => x"91",
           336 => x"88",
           337 => x"04",
           338 => x"70",
           339 => x"27",
           340 => x"71",
           341 => x"53",
           342 => x"90",
           343 => x"90",
           344 => x"91",
           345 => x"3c",
           346 => x"94",
           347 => x"ca",
           348 => x"3d",
           349 => x"91",
           350 => x"8c",
           351 => x"91",
           352 => x"88",
           353 => x"80",
           354 => x"ca",
           355 => x"91",
           356 => x"54",
           357 => x"91",
           358 => x"04",
           359 => x"08",
           360 => x"94",
           361 => x"0d",
           362 => x"ca",
           363 => x"05",
           364 => x"ca",
           365 => x"05",
           366 => x"3f",
           367 => x"08",
           368 => x"88",
           369 => x"3d",
           370 => x"94",
           371 => x"ca",
           372 => x"91",
           373 => x"fd",
           374 => x"0b",
           375 => x"08",
           376 => x"80",
           377 => x"94",
           378 => x"0c",
           379 => x"08",
           380 => x"91",
           381 => x"88",
           382 => x"b9",
           383 => x"94",
           384 => x"08",
           385 => x"38",
           386 => x"ca",
           387 => x"05",
           388 => x"38",
           389 => x"08",
           390 => x"10",
           391 => x"08",
           392 => x"91",
           393 => x"fc",
           394 => x"91",
           395 => x"fc",
           396 => x"b8",
           397 => x"94",
           398 => x"08",
           399 => x"e1",
           400 => x"94",
           401 => x"08",
           402 => x"08",
           403 => x"26",
           404 => x"ca",
           405 => x"05",
           406 => x"94",
           407 => x"08",
           408 => x"94",
           409 => x"0c",
           410 => x"08",
           411 => x"91",
           412 => x"fc",
           413 => x"91",
           414 => x"f8",
           415 => x"ca",
           416 => x"05",
           417 => x"91",
           418 => x"fc",
           419 => x"ca",
           420 => x"05",
           421 => x"91",
           422 => x"8c",
           423 => x"95",
           424 => x"94",
           425 => x"08",
           426 => x"38",
           427 => x"08",
           428 => x"70",
           429 => x"08",
           430 => x"51",
           431 => x"ca",
           432 => x"05",
           433 => x"ca",
           434 => x"05",
           435 => x"ca",
           436 => x"05",
           437 => x"88",
           438 => x"0d",
           439 => x"0c",
           440 => x"0d",
           441 => x"02",
           442 => x"05",
           443 => x"53",
           444 => x"27",
           445 => x"83",
           446 => x"80",
           447 => x"ff",
           448 => x"ff",
           449 => x"73",
           450 => x"05",
           451 => x"12",
           452 => x"2e",
           453 => x"ef",
           454 => x"ca",
           455 => x"3d",
           456 => x"74",
           457 => x"07",
           458 => x"2b",
           459 => x"51",
           460 => x"a5",
           461 => x"70",
           462 => x"0c",
           463 => x"84",
           464 => x"72",
           465 => x"05",
           466 => x"71",
           467 => x"53",
           468 => x"52",
           469 => x"dd",
           470 => x"27",
           471 => x"71",
           472 => x"53",
           473 => x"52",
           474 => x"f2",
           475 => x"ff",
           476 => x"3d",
           477 => x"70",
           478 => x"06",
           479 => x"70",
           480 => x"73",
           481 => x"56",
           482 => x"08",
           483 => x"38",
           484 => x"52",
           485 => x"81",
           486 => x"54",
           487 => x"9d",
           488 => x"55",
           489 => x"09",
           490 => x"38",
           491 => x"14",
           492 => x"81",
           493 => x"56",
           494 => x"e5",
           495 => x"55",
           496 => x"06",
           497 => x"06",
           498 => x"91",
           499 => x"52",
           500 => x"0d",
           501 => x"70",
           502 => x"ff",
           503 => x"f8",
           504 => x"80",
           505 => x"51",
           506 => x"84",
           507 => x"71",
           508 => x"54",
           509 => x"2e",
           510 => x"75",
           511 => x"94",
           512 => x"91",
           513 => x"87",
           514 => x"fe",
           515 => x"52",
           516 => x"88",
           517 => x"86",
           518 => x"88",
           519 => x"06",
           520 => x"14",
           521 => x"80",
           522 => x"71",
           523 => x"0c",
           524 => x"04",
           525 => x"77",
           526 => x"53",
           527 => x"80",
           528 => x"38",
           529 => x"70",
           530 => x"81",
           531 => x"81",
           532 => x"39",
           533 => x"39",
           534 => x"80",
           535 => x"81",
           536 => x"55",
           537 => x"2e",
           538 => x"55",
           539 => x"84",
           540 => x"38",
           541 => x"06",
           542 => x"2e",
           543 => x"88",
           544 => x"70",
           545 => x"34",
           546 => x"71",
           547 => x"ca",
           548 => x"3d",
           549 => x"3d",
           550 => x"72",
           551 => x"91",
           552 => x"fc",
           553 => x"51",
           554 => x"91",
           555 => x"85",
           556 => x"83",
           557 => x"72",
           558 => x"0c",
           559 => x"04",
           560 => x"76",
           561 => x"ff",
           562 => x"81",
           563 => x"26",
           564 => x"83",
           565 => x"05",
           566 => x"70",
           567 => x"8a",
           568 => x"33",
           569 => x"70",
           570 => x"fe",
           571 => x"33",
           572 => x"70",
           573 => x"f2",
           574 => x"33",
           575 => x"70",
           576 => x"e6",
           577 => x"22",
           578 => x"74",
           579 => x"80",
           580 => x"13",
           581 => x"52",
           582 => x"26",
           583 => x"81",
           584 => x"98",
           585 => x"22",
           586 => x"bc",
           587 => x"33",
           588 => x"b8",
           589 => x"33",
           590 => x"b4",
           591 => x"33",
           592 => x"b0",
           593 => x"33",
           594 => x"ac",
           595 => x"33",
           596 => x"a8",
           597 => x"c0",
           598 => x"73",
           599 => x"a0",
           600 => x"87",
           601 => x"0c",
           602 => x"91",
           603 => x"86",
           604 => x"f3",
           605 => x"5b",
           606 => x"9c",
           607 => x"0c",
           608 => x"bc",
           609 => x"7b",
           610 => x"98",
           611 => x"79",
           612 => x"87",
           613 => x"08",
           614 => x"1c",
           615 => x"98",
           616 => x"79",
           617 => x"87",
           618 => x"08",
           619 => x"1c",
           620 => x"98",
           621 => x"79",
           622 => x"87",
           623 => x"08",
           624 => x"1c",
           625 => x"98",
           626 => x"79",
           627 => x"80",
           628 => x"83",
           629 => x"59",
           630 => x"ff",
           631 => x"1b",
           632 => x"1b",
           633 => x"1b",
           634 => x"1b",
           635 => x"1b",
           636 => x"83",
           637 => x"52",
           638 => x"51",
           639 => x"8f",
           640 => x"ff",
           641 => x"8f",
           642 => x"30",
           643 => x"51",
           644 => x"0b",
           645 => x"e0",
           646 => x"0d",
           647 => x"0d",
           648 => x"91",
           649 => x"70",
           650 => x"57",
           651 => x"c0",
           652 => x"74",
           653 => x"38",
           654 => x"94",
           655 => x"70",
           656 => x"81",
           657 => x"52",
           658 => x"8c",
           659 => x"2a",
           660 => x"51",
           661 => x"38",
           662 => x"70",
           663 => x"51",
           664 => x"8d",
           665 => x"2a",
           666 => x"51",
           667 => x"be",
           668 => x"ff",
           669 => x"c0",
           670 => x"70",
           671 => x"38",
           672 => x"90",
           673 => x"0c",
           674 => x"88",
           675 => x"0d",
           676 => x"0d",
           677 => x"33",
           678 => x"c6",
           679 => x"81",
           680 => x"55",
           681 => x"94",
           682 => x"80",
           683 => x"87",
           684 => x"51",
           685 => x"96",
           686 => x"06",
           687 => x"70",
           688 => x"38",
           689 => x"70",
           690 => x"51",
           691 => x"72",
           692 => x"81",
           693 => x"70",
           694 => x"38",
           695 => x"70",
           696 => x"51",
           697 => x"38",
           698 => x"06",
           699 => x"94",
           700 => x"80",
           701 => x"87",
           702 => x"52",
           703 => x"87",
           704 => x"f9",
           705 => x"54",
           706 => x"70",
           707 => x"53",
           708 => x"77",
           709 => x"38",
           710 => x"06",
           711 => x"0b",
           712 => x"33",
           713 => x"06",
           714 => x"58",
           715 => x"84",
           716 => x"2e",
           717 => x"c0",
           718 => x"70",
           719 => x"2a",
           720 => x"53",
           721 => x"80",
           722 => x"71",
           723 => x"81",
           724 => x"70",
           725 => x"81",
           726 => x"06",
           727 => x"80",
           728 => x"71",
           729 => x"81",
           730 => x"70",
           731 => x"74",
           732 => x"51",
           733 => x"80",
           734 => x"2e",
           735 => x"c0",
           736 => x"77",
           737 => x"17",
           738 => x"81",
           739 => x"53",
           740 => x"84",
           741 => x"ca",
           742 => x"3d",
           743 => x"3d",
           744 => x"91",
           745 => x"70",
           746 => x"54",
           747 => x"94",
           748 => x"80",
           749 => x"87",
           750 => x"51",
           751 => x"82",
           752 => x"06",
           753 => x"70",
           754 => x"38",
           755 => x"06",
           756 => x"94",
           757 => x"80",
           758 => x"87",
           759 => x"52",
           760 => x"81",
           761 => x"ca",
           762 => x"84",
           763 => x"fe",
           764 => x"0b",
           765 => x"33",
           766 => x"06",
           767 => x"c0",
           768 => x"70",
           769 => x"38",
           770 => x"94",
           771 => x"70",
           772 => x"81",
           773 => x"51",
           774 => x"80",
           775 => x"72",
           776 => x"51",
           777 => x"80",
           778 => x"2e",
           779 => x"c0",
           780 => x"71",
           781 => x"2b",
           782 => x"51",
           783 => x"91",
           784 => x"84",
           785 => x"ff",
           786 => x"c0",
           787 => x"70",
           788 => x"06",
           789 => x"80",
           790 => x"38",
           791 => x"9c",
           792 => x"e4",
           793 => x"9e",
           794 => x"c6",
           795 => x"c0",
           796 => x"91",
           797 => x"87",
           798 => x"08",
           799 => x"0c",
           800 => x"94",
           801 => x"f4",
           802 => x"9e",
           803 => x"c6",
           804 => x"c0",
           805 => x"91",
           806 => x"87",
           807 => x"08",
           808 => x"0c",
           809 => x"ac",
           810 => x"84",
           811 => x"9e",
           812 => x"70",
           813 => x"23",
           814 => x"84",
           815 => x"8c",
           816 => x"91",
           817 => x"80",
           818 => x"9e",
           819 => x"a0",
           820 => x"52",
           821 => x"2e",
           822 => x"52",
           823 => x"91",
           824 => x"87",
           825 => x"08",
           826 => x"80",
           827 => x"52",
           828 => x"83",
           829 => x"71",
           830 => x"34",
           831 => x"c0",
           832 => x"70",
           833 => x"06",
           834 => x"70",
           835 => x"38",
           836 => x"91",
           837 => x"80",
           838 => x"9e",
           839 => x"90",
           840 => x"52",
           841 => x"2e",
           842 => x"52",
           843 => x"94",
           844 => x"87",
           845 => x"08",
           846 => x"06",
           847 => x"70",
           848 => x"38",
           849 => x"91",
           850 => x"80",
           851 => x"9e",
           852 => x"84",
           853 => x"52",
           854 => x"2e",
           855 => x"52",
           856 => x"96",
           857 => x"87",
           858 => x"08",
           859 => x"06",
           860 => x"70",
           861 => x"38",
           862 => x"91",
           863 => x"80",
           864 => x"9e",
           865 => x"81",
           866 => x"52",
           867 => x"2e",
           868 => x"52",
           869 => x"98",
           870 => x"9e",
           871 => x"80",
           872 => x"86",
           873 => x"51",
           874 => x"99",
           875 => x"87",
           876 => x"08",
           877 => x"51",
           878 => x"80",
           879 => x"81",
           880 => x"c7",
           881 => x"0b",
           882 => x"88",
           883 => x"06",
           884 => x"70",
           885 => x"38",
           886 => x"91",
           887 => x"87",
           888 => x"08",
           889 => x"51",
           890 => x"c7",
           891 => x"3d",
           892 => x"3d",
           893 => x"84",
           894 => x"3f",
           895 => x"33",
           896 => x"2e",
           897 => x"b4",
           898 => x"92",
           899 => x"ac",
           900 => x"3f",
           901 => x"33",
           902 => x"2e",
           903 => x"c6",
           904 => x"91",
           905 => x"52",
           906 => x"51",
           907 => x"91",
           908 => x"54",
           909 => x"92",
           910 => x"f0",
           911 => x"c6",
           912 => x"91",
           913 => x"89",
           914 => x"c7",
           915 => x"73",
           916 => x"c7",
           917 => x"73",
           918 => x"38",
           919 => x"08",
           920 => x"f4",
           921 => x"b5",
           922 => x"96",
           923 => x"95",
           924 => x"80",
           925 => x"91",
           926 => x"83",
           927 => x"c7",
           928 => x"73",
           929 => x"38",
           930 => x"51",
           931 => x"91",
           932 => x"54",
           933 => x"88",
           934 => x"cc",
           935 => x"3f",
           936 => x"33",
           937 => x"2e",
           938 => x"c7",
           939 => x"91",
           940 => x"88",
           941 => x"c7",
           942 => x"73",
           943 => x"38",
           944 => x"51",
           945 => x"91",
           946 => x"54",
           947 => x"8d",
           948 => x"9c",
           949 => x"b6",
           950 => x"a6",
           951 => x"b0",
           952 => x"3f",
           953 => x"08",
           954 => x"bc",
           955 => x"3f",
           956 => x"08",
           957 => x"e4",
           958 => x"3f",
           959 => x"08",
           960 => x"8c",
           961 => x"3f",
           962 => x"22",
           963 => x"b4",
           964 => x"3f",
           965 => x"08",
           966 => x"dc",
           967 => x"3f",
           968 => x"04",
           969 => x"02",
           970 => x"ff",
           971 => x"84",
           972 => x"71",
           973 => x"0b",
           974 => x"05",
           975 => x"04",
           976 => x"51",
           977 => x"b8",
           978 => x"39",
           979 => x"51",
           980 => x"b8",
           981 => x"39",
           982 => x"51",
           983 => x"b8",
           984 => x"9f",
           985 => x"0d",
           986 => x"80",
           987 => x"0b",
           988 => x"84",
           989 => x"3d",
           990 => x"96",
           991 => x"52",
           992 => x"0c",
           993 => x"70",
           994 => x"0c",
           995 => x"3d",
           996 => x"3d",
           997 => x"96",
           998 => x"91",
           999 => x"52",
          1000 => x"73",
          1001 => x"c7",
          1002 => x"70",
          1003 => x"0c",
          1004 => x"83",
          1005 => x"91",
          1006 => x"87",
          1007 => x"0c",
          1008 => x"0d",
          1009 => x"33",
          1010 => x"2e",
          1011 => x"85",
          1012 => x"ed",
          1013 => x"a0",
          1014 => x"80",
          1015 => x"72",
          1016 => x"ca",
          1017 => x"05",
          1018 => x"0c",
          1019 => x"ca",
          1020 => x"71",
          1021 => x"38",
          1022 => x"2d",
          1023 => x"04",
          1024 => x"02",
          1025 => x"91",
          1026 => x"76",
          1027 => x"0c",
          1028 => x"ad",
          1029 => x"ca",
          1030 => x"3d",
          1031 => x"3d",
          1032 => x"73",
          1033 => x"ff",
          1034 => x"71",
          1035 => x"38",
          1036 => x"06",
          1037 => x"54",
          1038 => x"e7",
          1039 => x"0d",
          1040 => x"0d",
          1041 => x"98",
          1042 => x"ca",
          1043 => x"54",
          1044 => x"81",
          1045 => x"53",
          1046 => x"8e",
          1047 => x"ff",
          1048 => x"14",
          1049 => x"3f",
          1050 => x"91",
          1051 => x"86",
          1052 => x"ec",
          1053 => x"68",
          1054 => x"70",
          1055 => x"33",
          1056 => x"2e",
          1057 => x"75",
          1058 => x"81",
          1059 => x"38",
          1060 => x"70",
          1061 => x"33",
          1062 => x"75",
          1063 => x"81",
          1064 => x"81",
          1065 => x"75",
          1066 => x"81",
          1067 => x"82",
          1068 => x"81",
          1069 => x"56",
          1070 => x"09",
          1071 => x"38",
          1072 => x"71",
          1073 => x"81",
          1074 => x"59",
          1075 => x"9d",
          1076 => x"53",
          1077 => x"95",
          1078 => x"29",
          1079 => x"76",
          1080 => x"79",
          1081 => x"5b",
          1082 => x"e5",
          1083 => x"ec",
          1084 => x"70",
          1085 => x"25",
          1086 => x"32",
          1087 => x"72",
          1088 => x"73",
          1089 => x"58",
          1090 => x"73",
          1091 => x"38",
          1092 => x"79",
          1093 => x"5b",
          1094 => x"75",
          1095 => x"de",
          1096 => x"80",
          1097 => x"89",
          1098 => x"70",
          1099 => x"55",
          1100 => x"cf",
          1101 => x"38",
          1102 => x"24",
          1103 => x"80",
          1104 => x"8e",
          1105 => x"c3",
          1106 => x"73",
          1107 => x"81",
          1108 => x"99",
          1109 => x"c4",
          1110 => x"38",
          1111 => x"73",
          1112 => x"81",
          1113 => x"80",
          1114 => x"38",
          1115 => x"2e",
          1116 => x"f9",
          1117 => x"d8",
          1118 => x"38",
          1119 => x"77",
          1120 => x"08",
          1121 => x"80",
          1122 => x"55",
          1123 => x"8d",
          1124 => x"70",
          1125 => x"51",
          1126 => x"f5",
          1127 => x"2a",
          1128 => x"74",
          1129 => x"53",
          1130 => x"8f",
          1131 => x"fc",
          1132 => x"81",
          1133 => x"80",
          1134 => x"73",
          1135 => x"3f",
          1136 => x"56",
          1137 => x"27",
          1138 => x"a0",
          1139 => x"3f",
          1140 => x"84",
          1141 => x"33",
          1142 => x"93",
          1143 => x"95",
          1144 => x"91",
          1145 => x"8d",
          1146 => x"89",
          1147 => x"fb",
          1148 => x"86",
          1149 => x"2a",
          1150 => x"51",
          1151 => x"2e",
          1152 => x"84",
          1153 => x"86",
          1154 => x"78",
          1155 => x"08",
          1156 => x"32",
          1157 => x"72",
          1158 => x"51",
          1159 => x"74",
          1160 => x"38",
          1161 => x"88",
          1162 => x"7a",
          1163 => x"55",
          1164 => x"3d",
          1165 => x"52",
          1166 => x"e0",
          1167 => x"88",
          1168 => x"06",
          1169 => x"52",
          1170 => x"3f",
          1171 => x"08",
          1172 => x"27",
          1173 => x"14",
          1174 => x"f8",
          1175 => x"87",
          1176 => x"81",
          1177 => x"b0",
          1178 => x"7d",
          1179 => x"5f",
          1180 => x"75",
          1181 => x"07",
          1182 => x"54",
          1183 => x"26",
          1184 => x"ff",
          1185 => x"84",
          1186 => x"06",
          1187 => x"80",
          1188 => x"96",
          1189 => x"e0",
          1190 => x"73",
          1191 => x"57",
          1192 => x"06",
          1193 => x"54",
          1194 => x"a0",
          1195 => x"2a",
          1196 => x"54",
          1197 => x"38",
          1198 => x"76",
          1199 => x"38",
          1200 => x"fd",
          1201 => x"06",
          1202 => x"38",
          1203 => x"56",
          1204 => x"26",
          1205 => x"3d",
          1206 => x"05",
          1207 => x"ff",
          1208 => x"53",
          1209 => x"d9",
          1210 => x"38",
          1211 => x"56",
          1212 => x"27",
          1213 => x"a0",
          1214 => x"3f",
          1215 => x"3d",
          1216 => x"3d",
          1217 => x"70",
          1218 => x"52",
          1219 => x"73",
          1220 => x"3f",
          1221 => x"04",
          1222 => x"74",
          1223 => x"0c",
          1224 => x"05",
          1225 => x"fa",
          1226 => x"ca",
          1227 => x"80",
          1228 => x"0b",
          1229 => x"0c",
          1230 => x"04",
          1231 => x"91",
          1232 => x"76",
          1233 => x"0c",
          1234 => x"05",
          1235 => x"53",
          1236 => x"72",
          1237 => x"0c",
          1238 => x"04",
          1239 => x"77",
          1240 => x"9c",
          1241 => x"54",
          1242 => x"54",
          1243 => x"80",
          1244 => x"ca",
          1245 => x"71",
          1246 => x"88",
          1247 => x"06",
          1248 => x"2e",
          1249 => x"72",
          1250 => x"38",
          1251 => x"70",
          1252 => x"25",
          1253 => x"73",
          1254 => x"38",
          1255 => x"86",
          1256 => x"54",
          1257 => x"73",
          1258 => x"ff",
          1259 => x"72",
          1260 => x"74",
          1261 => x"72",
          1262 => x"54",
          1263 => x"81",
          1264 => x"39",
          1265 => x"80",
          1266 => x"51",
          1267 => x"81",
          1268 => x"ca",
          1269 => x"3d",
          1270 => x"3d",
          1271 => x"9c",
          1272 => x"ca",
          1273 => x"53",
          1274 => x"fe",
          1275 => x"91",
          1276 => x"84",
          1277 => x"f8",
          1278 => x"7c",
          1279 => x"70",
          1280 => x"75",
          1281 => x"55",
          1282 => x"2e",
          1283 => x"87",
          1284 => x"76",
          1285 => x"73",
          1286 => x"81",
          1287 => x"81",
          1288 => x"77",
          1289 => x"70",
          1290 => x"58",
          1291 => x"09",
          1292 => x"c2",
          1293 => x"81",
          1294 => x"75",
          1295 => x"55",
          1296 => x"e2",
          1297 => x"90",
          1298 => x"f8",
          1299 => x"8f",
          1300 => x"81",
          1301 => x"75",
          1302 => x"55",
          1303 => x"81",
          1304 => x"27",
          1305 => x"d0",
          1306 => x"55",
          1307 => x"73",
          1308 => x"80",
          1309 => x"14",
          1310 => x"72",
          1311 => x"e0",
          1312 => x"80",
          1313 => x"39",
          1314 => x"55",
          1315 => x"80",
          1316 => x"e0",
          1317 => x"38",
          1318 => x"81",
          1319 => x"53",
          1320 => x"81",
          1321 => x"53",
          1322 => x"8e",
          1323 => x"70",
          1324 => x"55",
          1325 => x"27",
          1326 => x"77",
          1327 => x"74",
          1328 => x"76",
          1329 => x"77",
          1330 => x"70",
          1331 => x"55",
          1332 => x"77",
          1333 => x"38",
          1334 => x"74",
          1335 => x"55",
          1336 => x"88",
          1337 => x"0d",
          1338 => x"0d",
          1339 => x"56",
          1340 => x"0c",
          1341 => x"70",
          1342 => x"73",
          1343 => x"81",
          1344 => x"81",
          1345 => x"ed",
          1346 => x"2e",
          1347 => x"8e",
          1348 => x"08",
          1349 => x"76",
          1350 => x"56",
          1351 => x"b0",
          1352 => x"06",
          1353 => x"75",
          1354 => x"76",
          1355 => x"70",
          1356 => x"73",
          1357 => x"8b",
          1358 => x"73",
          1359 => x"85",
          1360 => x"82",
          1361 => x"76",
          1362 => x"70",
          1363 => x"ac",
          1364 => x"a0",
          1365 => x"fa",
          1366 => x"53",
          1367 => x"57",
          1368 => x"98",
          1369 => x"39",
          1370 => x"80",
          1371 => x"26",
          1372 => x"86",
          1373 => x"80",
          1374 => x"57",
          1375 => x"74",
          1376 => x"38",
          1377 => x"27",
          1378 => x"14",
          1379 => x"06",
          1380 => x"14",
          1381 => x"06",
          1382 => x"74",
          1383 => x"f9",
          1384 => x"ff",
          1385 => x"89",
          1386 => x"38",
          1387 => x"c5",
          1388 => x"29",
          1389 => x"81",
          1390 => x"76",
          1391 => x"56",
          1392 => x"ba",
          1393 => x"2e",
          1394 => x"30",
          1395 => x"0c",
          1396 => x"91",
          1397 => x"8a",
          1398 => x"ff",
          1399 => x"8f",
          1400 => x"81",
          1401 => x"26",
          1402 => x"c7",
          1403 => x"52",
          1404 => x"88",
          1405 => x"0d",
          1406 => x"0d",
          1407 => x"33",
          1408 => x"9f",
          1409 => x"53",
          1410 => x"81",
          1411 => x"38",
          1412 => x"87",
          1413 => x"11",
          1414 => x"54",
          1415 => x"84",
          1416 => x"54",
          1417 => x"87",
          1418 => x"11",
          1419 => x"0c",
          1420 => x"c0",
          1421 => x"70",
          1422 => x"70",
          1423 => x"51",
          1424 => x"8a",
          1425 => x"98",
          1426 => x"70",
          1427 => x"08",
          1428 => x"06",
          1429 => x"38",
          1430 => x"8c",
          1431 => x"80",
          1432 => x"71",
          1433 => x"14",
          1434 => x"a4",
          1435 => x"70",
          1436 => x"0c",
          1437 => x"04",
          1438 => x"60",
          1439 => x"8c",
          1440 => x"33",
          1441 => x"5b",
          1442 => x"5a",
          1443 => x"91",
          1444 => x"81",
          1445 => x"52",
          1446 => x"38",
          1447 => x"84",
          1448 => x"92",
          1449 => x"c0",
          1450 => x"87",
          1451 => x"13",
          1452 => x"57",
          1453 => x"0b",
          1454 => x"8c",
          1455 => x"0c",
          1456 => x"75",
          1457 => x"2a",
          1458 => x"51",
          1459 => x"80",
          1460 => x"7b",
          1461 => x"7b",
          1462 => x"5d",
          1463 => x"59",
          1464 => x"06",
          1465 => x"73",
          1466 => x"81",
          1467 => x"ff",
          1468 => x"72",
          1469 => x"38",
          1470 => x"8c",
          1471 => x"c3",
          1472 => x"98",
          1473 => x"71",
          1474 => x"38",
          1475 => x"2e",
          1476 => x"76",
          1477 => x"92",
          1478 => x"72",
          1479 => x"06",
          1480 => x"f7",
          1481 => x"5a",
          1482 => x"80",
          1483 => x"70",
          1484 => x"5a",
          1485 => x"80",
          1486 => x"73",
          1487 => x"06",
          1488 => x"38",
          1489 => x"fe",
          1490 => x"fc",
          1491 => x"52",
          1492 => x"83",
          1493 => x"71",
          1494 => x"ca",
          1495 => x"3d",
          1496 => x"3d",
          1497 => x"64",
          1498 => x"bf",
          1499 => x"40",
          1500 => x"59",
          1501 => x"58",
          1502 => x"91",
          1503 => x"81",
          1504 => x"52",
          1505 => x"09",
          1506 => x"b1",
          1507 => x"84",
          1508 => x"92",
          1509 => x"c0",
          1510 => x"87",
          1511 => x"13",
          1512 => x"56",
          1513 => x"87",
          1514 => x"0c",
          1515 => x"82",
          1516 => x"58",
          1517 => x"84",
          1518 => x"06",
          1519 => x"71",
          1520 => x"38",
          1521 => x"05",
          1522 => x"0c",
          1523 => x"73",
          1524 => x"81",
          1525 => x"71",
          1526 => x"38",
          1527 => x"8c",
          1528 => x"d0",
          1529 => x"98",
          1530 => x"71",
          1531 => x"38",
          1532 => x"2e",
          1533 => x"76",
          1534 => x"92",
          1535 => x"72",
          1536 => x"06",
          1537 => x"f7",
          1538 => x"59",
          1539 => x"1a",
          1540 => x"06",
          1541 => x"59",
          1542 => x"80",
          1543 => x"73",
          1544 => x"06",
          1545 => x"38",
          1546 => x"fe",
          1547 => x"fc",
          1548 => x"52",
          1549 => x"83",
          1550 => x"71",
          1551 => x"ca",
          1552 => x"3d",
          1553 => x"3d",
          1554 => x"84",
          1555 => x"33",
          1556 => x"b7",
          1557 => x"54",
          1558 => x"fa",
          1559 => x"ca",
          1560 => x"06",
          1561 => x"72",
          1562 => x"85",
          1563 => x"98",
          1564 => x"56",
          1565 => x"80",
          1566 => x"76",
          1567 => x"74",
          1568 => x"c0",
          1569 => x"54",
          1570 => x"2e",
          1571 => x"d4",
          1572 => x"2e",
          1573 => x"80",
          1574 => x"08",
          1575 => x"70",
          1576 => x"51",
          1577 => x"2e",
          1578 => x"c0",
          1579 => x"52",
          1580 => x"87",
          1581 => x"08",
          1582 => x"38",
          1583 => x"87",
          1584 => x"14",
          1585 => x"70",
          1586 => x"52",
          1587 => x"96",
          1588 => x"92",
          1589 => x"0a",
          1590 => x"39",
          1591 => x"0c",
          1592 => x"39",
          1593 => x"54",
          1594 => x"88",
          1595 => x"0d",
          1596 => x"0d",
          1597 => x"33",
          1598 => x"88",
          1599 => x"ca",
          1600 => x"51",
          1601 => x"04",
          1602 => x"75",
          1603 => x"82",
          1604 => x"90",
          1605 => x"2b",
          1606 => x"33",
          1607 => x"88",
          1608 => x"71",
          1609 => x"88",
          1610 => x"54",
          1611 => x"85",
          1612 => x"ff",
          1613 => x"02",
          1614 => x"05",
          1615 => x"70",
          1616 => x"05",
          1617 => x"88",
          1618 => x"72",
          1619 => x"0d",
          1620 => x"0d",
          1621 => x"52",
          1622 => x"81",
          1623 => x"70",
          1624 => x"70",
          1625 => x"05",
          1626 => x"88",
          1627 => x"72",
          1628 => x"54",
          1629 => x"2a",
          1630 => x"34",
          1631 => x"04",
          1632 => x"76",
          1633 => x"54",
          1634 => x"2e",
          1635 => x"70",
          1636 => x"33",
          1637 => x"05",
          1638 => x"11",
          1639 => x"84",
          1640 => x"fe",
          1641 => x"77",
          1642 => x"53",
          1643 => x"81",
          1644 => x"ff",
          1645 => x"f4",
          1646 => x"0d",
          1647 => x"0d",
          1648 => x"56",
          1649 => x"70",
          1650 => x"33",
          1651 => x"05",
          1652 => x"71",
          1653 => x"56",
          1654 => x"72",
          1655 => x"38",
          1656 => x"e2",
          1657 => x"ca",
          1658 => x"3d",
          1659 => x"3d",
          1660 => x"54",
          1661 => x"71",
          1662 => x"38",
          1663 => x"70",
          1664 => x"f3",
          1665 => x"91",
          1666 => x"84",
          1667 => x"80",
          1668 => x"88",
          1669 => x"0b",
          1670 => x"0c",
          1671 => x"0d",
          1672 => x"0b",
          1673 => x"56",
          1674 => x"2e",
          1675 => x"81",
          1676 => x"08",
          1677 => x"70",
          1678 => x"33",
          1679 => x"a2",
          1680 => x"88",
          1681 => x"09",
          1682 => x"38",
          1683 => x"08",
          1684 => x"b0",
          1685 => x"a4",
          1686 => x"9c",
          1687 => x"56",
          1688 => x"27",
          1689 => x"16",
          1690 => x"82",
          1691 => x"06",
          1692 => x"54",
          1693 => x"78",
          1694 => x"33",
          1695 => x"3f",
          1696 => x"5a",
          1697 => x"88",
          1698 => x"0d",
          1699 => x"0d",
          1700 => x"56",
          1701 => x"b0",
          1702 => x"af",
          1703 => x"fe",
          1704 => x"ca",
          1705 => x"91",
          1706 => x"9f",
          1707 => x"74",
          1708 => x"52",
          1709 => x"51",
          1710 => x"91",
          1711 => x"80",
          1712 => x"ff",
          1713 => x"74",
          1714 => x"76",
          1715 => x"0c",
          1716 => x"04",
          1717 => x"7a",
          1718 => x"fe",
          1719 => x"ca",
          1720 => x"91",
          1721 => x"81",
          1722 => x"33",
          1723 => x"2e",
          1724 => x"80",
          1725 => x"17",
          1726 => x"81",
          1727 => x"06",
          1728 => x"84",
          1729 => x"ca",
          1730 => x"b4",
          1731 => x"56",
          1732 => x"82",
          1733 => x"84",
          1734 => x"fc",
          1735 => x"8b",
          1736 => x"52",
          1737 => x"a9",
          1738 => x"85",
          1739 => x"84",
          1740 => x"fc",
          1741 => x"17",
          1742 => x"9c",
          1743 => x"91",
          1744 => x"08",
          1745 => x"17",
          1746 => x"3f",
          1747 => x"81",
          1748 => x"19",
          1749 => x"53",
          1750 => x"17",
          1751 => x"82",
          1752 => x"18",
          1753 => x"80",
          1754 => x"33",
          1755 => x"3f",
          1756 => x"08",
          1757 => x"38",
          1758 => x"91",
          1759 => x"8a",
          1760 => x"fb",
          1761 => x"fe",
          1762 => x"08",
          1763 => x"56",
          1764 => x"74",
          1765 => x"38",
          1766 => x"75",
          1767 => x"16",
          1768 => x"53",
          1769 => x"88",
          1770 => x"0d",
          1771 => x"0d",
          1772 => x"08",
          1773 => x"81",
          1774 => x"df",
          1775 => x"15",
          1776 => x"d7",
          1777 => x"33",
          1778 => x"82",
          1779 => x"38",
          1780 => x"89",
          1781 => x"2e",
          1782 => x"bf",
          1783 => x"2e",
          1784 => x"81",
          1785 => x"81",
          1786 => x"89",
          1787 => x"08",
          1788 => x"52",
          1789 => x"3f",
          1790 => x"08",
          1791 => x"74",
          1792 => x"14",
          1793 => x"81",
          1794 => x"2a",
          1795 => x"05",
          1796 => x"57",
          1797 => x"f5",
          1798 => x"88",
          1799 => x"38",
          1800 => x"06",
          1801 => x"33",
          1802 => x"78",
          1803 => x"06",
          1804 => x"5c",
          1805 => x"53",
          1806 => x"38",
          1807 => x"06",
          1808 => x"39",
          1809 => x"a4",
          1810 => x"52",
          1811 => x"bd",
          1812 => x"88",
          1813 => x"38",
          1814 => x"fe",
          1815 => x"b4",
          1816 => x"8d",
          1817 => x"88",
          1818 => x"ff",
          1819 => x"39",
          1820 => x"a4",
          1821 => x"52",
          1822 => x"91",
          1823 => x"88",
          1824 => x"76",
          1825 => x"fc",
          1826 => x"b4",
          1827 => x"f8",
          1828 => x"88",
          1829 => x"06",
          1830 => x"81",
          1831 => x"ca",
          1832 => x"3d",
          1833 => x"3d",
          1834 => x"7e",
          1835 => x"82",
          1836 => x"27",
          1837 => x"76",
          1838 => x"27",
          1839 => x"75",
          1840 => x"79",
          1841 => x"38",
          1842 => x"89",
          1843 => x"2e",
          1844 => x"80",
          1845 => x"2e",
          1846 => x"81",
          1847 => x"81",
          1848 => x"89",
          1849 => x"08",
          1850 => x"52",
          1851 => x"3f",
          1852 => x"08",
          1853 => x"88",
          1854 => x"38",
          1855 => x"06",
          1856 => x"81",
          1857 => x"06",
          1858 => x"77",
          1859 => x"2e",
          1860 => x"84",
          1861 => x"06",
          1862 => x"06",
          1863 => x"53",
          1864 => x"81",
          1865 => x"34",
          1866 => x"a4",
          1867 => x"52",
          1868 => x"d9",
          1869 => x"88",
          1870 => x"ca",
          1871 => x"94",
          1872 => x"ff",
          1873 => x"05",
          1874 => x"54",
          1875 => x"38",
          1876 => x"74",
          1877 => x"06",
          1878 => x"07",
          1879 => x"74",
          1880 => x"39",
          1881 => x"a4",
          1882 => x"52",
          1883 => x"9d",
          1884 => x"88",
          1885 => x"ca",
          1886 => x"d8",
          1887 => x"ff",
          1888 => x"76",
          1889 => x"06",
          1890 => x"05",
          1891 => x"3f",
          1892 => x"87",
          1893 => x"08",
          1894 => x"51",
          1895 => x"91",
          1896 => x"59",
          1897 => x"08",
          1898 => x"f0",
          1899 => x"82",
          1900 => x"06",
          1901 => x"05",
          1902 => x"54",
          1903 => x"3f",
          1904 => x"08",
          1905 => x"74",
          1906 => x"51",
          1907 => x"81",
          1908 => x"34",
          1909 => x"88",
          1910 => x"0d",
          1911 => x"0d",
          1912 => x"72",
          1913 => x"56",
          1914 => x"27",
          1915 => x"98",
          1916 => x"9d",
          1917 => x"2e",
          1918 => x"53",
          1919 => x"51",
          1920 => x"91",
          1921 => x"54",
          1922 => x"08",
          1923 => x"93",
          1924 => x"80",
          1925 => x"54",
          1926 => x"91",
          1927 => x"54",
          1928 => x"74",
          1929 => x"fb",
          1930 => x"ca",
          1931 => x"91",
          1932 => x"80",
          1933 => x"38",
          1934 => x"08",
          1935 => x"38",
          1936 => x"08",
          1937 => x"38",
          1938 => x"52",
          1939 => x"d6",
          1940 => x"88",
          1941 => x"98",
          1942 => x"11",
          1943 => x"57",
          1944 => x"74",
          1945 => x"81",
          1946 => x"0c",
          1947 => x"81",
          1948 => x"84",
          1949 => x"55",
          1950 => x"ff",
          1951 => x"54",
          1952 => x"88",
          1953 => x"0d",
          1954 => x"0d",
          1955 => x"08",
          1956 => x"79",
          1957 => x"17",
          1958 => x"80",
          1959 => x"98",
          1960 => x"26",
          1961 => x"58",
          1962 => x"52",
          1963 => x"fd",
          1964 => x"74",
          1965 => x"08",
          1966 => x"38",
          1967 => x"08",
          1968 => x"88",
          1969 => x"82",
          1970 => x"17",
          1971 => x"88",
          1972 => x"c7",
          1973 => x"90",
          1974 => x"56",
          1975 => x"2e",
          1976 => x"77",
          1977 => x"81",
          1978 => x"38",
          1979 => x"98",
          1980 => x"26",
          1981 => x"56",
          1982 => x"51",
          1983 => x"80",
          1984 => x"88",
          1985 => x"09",
          1986 => x"38",
          1987 => x"08",
          1988 => x"88",
          1989 => x"30",
          1990 => x"80",
          1991 => x"07",
          1992 => x"08",
          1993 => x"55",
          1994 => x"ef",
          1995 => x"88",
          1996 => x"95",
          1997 => x"08",
          1998 => x"27",
          1999 => x"98",
          2000 => x"89",
          2001 => x"85",
          2002 => x"db",
          2003 => x"81",
          2004 => x"17",
          2005 => x"89",
          2006 => x"75",
          2007 => x"ac",
          2008 => x"7a",
          2009 => x"3f",
          2010 => x"08",
          2011 => x"38",
          2012 => x"ca",
          2013 => x"2e",
          2014 => x"86",
          2015 => x"88",
          2016 => x"ca",
          2017 => x"70",
          2018 => x"07",
          2019 => x"7c",
          2020 => x"55",
          2021 => x"f8",
          2022 => x"2e",
          2023 => x"ff",
          2024 => x"55",
          2025 => x"ff",
          2026 => x"76",
          2027 => x"3f",
          2028 => x"08",
          2029 => x"08",
          2030 => x"ca",
          2031 => x"80",
          2032 => x"55",
          2033 => x"94",
          2034 => x"2e",
          2035 => x"53",
          2036 => x"51",
          2037 => x"91",
          2038 => x"55",
          2039 => x"75",
          2040 => x"98",
          2041 => x"05",
          2042 => x"56",
          2043 => x"26",
          2044 => x"15",
          2045 => x"84",
          2046 => x"07",
          2047 => x"18",
          2048 => x"ff",
          2049 => x"2e",
          2050 => x"39",
          2051 => x"39",
          2052 => x"08",
          2053 => x"81",
          2054 => x"74",
          2055 => x"0c",
          2056 => x"04",
          2057 => x"7a",
          2058 => x"f3",
          2059 => x"ca",
          2060 => x"81",
          2061 => x"88",
          2062 => x"38",
          2063 => x"51",
          2064 => x"91",
          2065 => x"91",
          2066 => x"b0",
          2067 => x"84",
          2068 => x"52",
          2069 => x"52",
          2070 => x"3f",
          2071 => x"39",
          2072 => x"8a",
          2073 => x"75",
          2074 => x"38",
          2075 => x"19",
          2076 => x"81",
          2077 => x"ed",
          2078 => x"ca",
          2079 => x"2e",
          2080 => x"15",
          2081 => x"70",
          2082 => x"07",
          2083 => x"53",
          2084 => x"75",
          2085 => x"0c",
          2086 => x"04",
          2087 => x"7a",
          2088 => x"58",
          2089 => x"f0",
          2090 => x"80",
          2091 => x"9f",
          2092 => x"80",
          2093 => x"90",
          2094 => x"17",
          2095 => x"aa",
          2096 => x"53",
          2097 => x"88",
          2098 => x"08",
          2099 => x"38",
          2100 => x"53",
          2101 => x"17",
          2102 => x"72",
          2103 => x"fe",
          2104 => x"08",
          2105 => x"80",
          2106 => x"16",
          2107 => x"2b",
          2108 => x"75",
          2109 => x"73",
          2110 => x"f5",
          2111 => x"ca",
          2112 => x"91",
          2113 => x"ff",
          2114 => x"81",
          2115 => x"88",
          2116 => x"38",
          2117 => x"91",
          2118 => x"26",
          2119 => x"58",
          2120 => x"73",
          2121 => x"39",
          2122 => x"51",
          2123 => x"91",
          2124 => x"98",
          2125 => x"94",
          2126 => x"17",
          2127 => x"58",
          2128 => x"9a",
          2129 => x"81",
          2130 => x"74",
          2131 => x"98",
          2132 => x"83",
          2133 => x"b4",
          2134 => x"0c",
          2135 => x"91",
          2136 => x"8a",
          2137 => x"f8",
          2138 => x"70",
          2139 => x"08",
          2140 => x"57",
          2141 => x"0a",
          2142 => x"38",
          2143 => x"15",
          2144 => x"08",
          2145 => x"72",
          2146 => x"cb",
          2147 => x"ff",
          2148 => x"81",
          2149 => x"13",
          2150 => x"94",
          2151 => x"74",
          2152 => x"85",
          2153 => x"22",
          2154 => x"73",
          2155 => x"38",
          2156 => x"8a",
          2157 => x"05",
          2158 => x"06",
          2159 => x"8a",
          2160 => x"73",
          2161 => x"3f",
          2162 => x"08",
          2163 => x"81",
          2164 => x"88",
          2165 => x"ff",
          2166 => x"91",
          2167 => x"ff",
          2168 => x"38",
          2169 => x"91",
          2170 => x"26",
          2171 => x"7b",
          2172 => x"98",
          2173 => x"55",
          2174 => x"94",
          2175 => x"73",
          2176 => x"3f",
          2177 => x"08",
          2178 => x"91",
          2179 => x"80",
          2180 => x"38",
          2181 => x"ca",
          2182 => x"2e",
          2183 => x"55",
          2184 => x"08",
          2185 => x"38",
          2186 => x"08",
          2187 => x"fb",
          2188 => x"ca",
          2189 => x"38",
          2190 => x"0c",
          2191 => x"51",
          2192 => x"91",
          2193 => x"98",
          2194 => x"90",
          2195 => x"16",
          2196 => x"15",
          2197 => x"74",
          2198 => x"0c",
          2199 => x"04",
          2200 => x"7b",
          2201 => x"5b",
          2202 => x"52",
          2203 => x"ac",
          2204 => x"88",
          2205 => x"ca",
          2206 => x"ec",
          2207 => x"88",
          2208 => x"17",
          2209 => x"51",
          2210 => x"91",
          2211 => x"54",
          2212 => x"08",
          2213 => x"91",
          2214 => x"9c",
          2215 => x"33",
          2216 => x"72",
          2217 => x"09",
          2218 => x"38",
          2219 => x"ca",
          2220 => x"72",
          2221 => x"55",
          2222 => x"53",
          2223 => x"8e",
          2224 => x"56",
          2225 => x"09",
          2226 => x"38",
          2227 => x"ca",
          2228 => x"81",
          2229 => x"fd",
          2230 => x"ca",
          2231 => x"91",
          2232 => x"80",
          2233 => x"38",
          2234 => x"09",
          2235 => x"38",
          2236 => x"91",
          2237 => x"8b",
          2238 => x"fd",
          2239 => x"9a",
          2240 => x"eb",
          2241 => x"ca",
          2242 => x"ff",
          2243 => x"70",
          2244 => x"53",
          2245 => x"09",
          2246 => x"38",
          2247 => x"eb",
          2248 => x"ca",
          2249 => x"2b",
          2250 => x"72",
          2251 => x"0c",
          2252 => x"04",
          2253 => x"77",
          2254 => x"ff",
          2255 => x"9a",
          2256 => x"55",
          2257 => x"76",
          2258 => x"53",
          2259 => x"09",
          2260 => x"38",
          2261 => x"52",
          2262 => x"eb",
          2263 => x"3d",
          2264 => x"3d",
          2265 => x"5b",
          2266 => x"08",
          2267 => x"15",
          2268 => x"81",
          2269 => x"15",
          2270 => x"51",
          2271 => x"91",
          2272 => x"58",
          2273 => x"08",
          2274 => x"9c",
          2275 => x"33",
          2276 => x"86",
          2277 => x"80",
          2278 => x"13",
          2279 => x"06",
          2280 => x"06",
          2281 => x"72",
          2282 => x"91",
          2283 => x"53",
          2284 => x"2e",
          2285 => x"53",
          2286 => x"a9",
          2287 => x"74",
          2288 => x"72",
          2289 => x"38",
          2290 => x"99",
          2291 => x"88",
          2292 => x"06",
          2293 => x"88",
          2294 => x"06",
          2295 => x"54",
          2296 => x"a0",
          2297 => x"74",
          2298 => x"3f",
          2299 => x"08",
          2300 => x"88",
          2301 => x"98",
          2302 => x"fa",
          2303 => x"80",
          2304 => x"0c",
          2305 => x"88",
          2306 => x"0d",
          2307 => x"0d",
          2308 => x"57",
          2309 => x"73",
          2310 => x"3f",
          2311 => x"08",
          2312 => x"88",
          2313 => x"98",
          2314 => x"75",
          2315 => x"3f",
          2316 => x"08",
          2317 => x"88",
          2318 => x"a0",
          2319 => x"88",
          2320 => x"14",
          2321 => x"db",
          2322 => x"a0",
          2323 => x"14",
          2324 => x"ac",
          2325 => x"83",
          2326 => x"91",
          2327 => x"87",
          2328 => x"fd",
          2329 => x"70",
          2330 => x"08",
          2331 => x"55",
          2332 => x"3f",
          2333 => x"08",
          2334 => x"13",
          2335 => x"73",
          2336 => x"83",
          2337 => x"3d",
          2338 => x"3d",
          2339 => x"57",
          2340 => x"89",
          2341 => x"17",
          2342 => x"81",
          2343 => x"70",
          2344 => x"55",
          2345 => x"08",
          2346 => x"81",
          2347 => x"52",
          2348 => x"a8",
          2349 => x"2e",
          2350 => x"84",
          2351 => x"52",
          2352 => x"09",
          2353 => x"38",
          2354 => x"81",
          2355 => x"81",
          2356 => x"73",
          2357 => x"55",
          2358 => x"55",
          2359 => x"c5",
          2360 => x"88",
          2361 => x"0b",
          2362 => x"9c",
          2363 => x"8b",
          2364 => x"17",
          2365 => x"08",
          2366 => x"52",
          2367 => x"91",
          2368 => x"76",
          2369 => x"51",
          2370 => x"91",
          2371 => x"86",
          2372 => x"12",
          2373 => x"3f",
          2374 => x"08",
          2375 => x"88",
          2376 => x"f3",
          2377 => x"70",
          2378 => x"80",
          2379 => x"51",
          2380 => x"af",
          2381 => x"81",
          2382 => x"dc",
          2383 => x"74",
          2384 => x"38",
          2385 => x"88",
          2386 => x"39",
          2387 => x"80",
          2388 => x"56",
          2389 => x"af",
          2390 => x"06",
          2391 => x"56",
          2392 => x"32",
          2393 => x"80",
          2394 => x"51",
          2395 => x"dc",
          2396 => x"1c",
          2397 => x"33",
          2398 => x"9f",
          2399 => x"ff",
          2400 => x"1c",
          2401 => x"7a",
          2402 => x"3f",
          2403 => x"08",
          2404 => x"39",
          2405 => x"a0",
          2406 => x"5e",
          2407 => x"52",
          2408 => x"ff",
          2409 => x"59",
          2410 => x"33",
          2411 => x"ae",
          2412 => x"06",
          2413 => x"78",
          2414 => x"81",
          2415 => x"32",
          2416 => x"9f",
          2417 => x"26",
          2418 => x"53",
          2419 => x"73",
          2420 => x"17",
          2421 => x"34",
          2422 => x"db",
          2423 => x"32",
          2424 => x"9f",
          2425 => x"54",
          2426 => x"2e",
          2427 => x"80",
          2428 => x"75",
          2429 => x"bd",
          2430 => x"7e",
          2431 => x"a0",
          2432 => x"bd",
          2433 => x"82",
          2434 => x"18",
          2435 => x"1a",
          2436 => x"a0",
          2437 => x"fc",
          2438 => x"32",
          2439 => x"80",
          2440 => x"30",
          2441 => x"71",
          2442 => x"51",
          2443 => x"55",
          2444 => x"ac",
          2445 => x"81",
          2446 => x"78",
          2447 => x"51",
          2448 => x"af",
          2449 => x"06",
          2450 => x"55",
          2451 => x"32",
          2452 => x"80",
          2453 => x"51",
          2454 => x"db",
          2455 => x"39",
          2456 => x"09",
          2457 => x"38",
          2458 => x"7c",
          2459 => x"54",
          2460 => x"a2",
          2461 => x"32",
          2462 => x"ae",
          2463 => x"72",
          2464 => x"9f",
          2465 => x"51",
          2466 => x"74",
          2467 => x"88",
          2468 => x"fe",
          2469 => x"98",
          2470 => x"80",
          2471 => x"75",
          2472 => x"91",
          2473 => x"33",
          2474 => x"51",
          2475 => x"91",
          2476 => x"80",
          2477 => x"78",
          2478 => x"81",
          2479 => x"5a",
          2480 => x"d2",
          2481 => x"88",
          2482 => x"80",
          2483 => x"1c",
          2484 => x"27",
          2485 => x"79",
          2486 => x"74",
          2487 => x"7a",
          2488 => x"74",
          2489 => x"39",
          2490 => x"b8",
          2491 => x"fe",
          2492 => x"88",
          2493 => x"ff",
          2494 => x"73",
          2495 => x"38",
          2496 => x"81",
          2497 => x"54",
          2498 => x"75",
          2499 => x"17",
          2500 => x"39",
          2501 => x"0c",
          2502 => x"99",
          2503 => x"54",
          2504 => x"2e",
          2505 => x"84",
          2506 => x"34",
          2507 => x"76",
          2508 => x"8b",
          2509 => x"81",
          2510 => x"56",
          2511 => x"80",
          2512 => x"1b",
          2513 => x"08",
          2514 => x"51",
          2515 => x"91",
          2516 => x"56",
          2517 => x"08",
          2518 => x"98",
          2519 => x"76",
          2520 => x"3f",
          2521 => x"08",
          2522 => x"88",
          2523 => x"38",
          2524 => x"70",
          2525 => x"73",
          2526 => x"be",
          2527 => x"33",
          2528 => x"73",
          2529 => x"8b",
          2530 => x"83",
          2531 => x"06",
          2532 => x"73",
          2533 => x"53",
          2534 => x"51",
          2535 => x"91",
          2536 => x"80",
          2537 => x"75",
          2538 => x"f3",
          2539 => x"9f",
          2540 => x"1c",
          2541 => x"74",
          2542 => x"38",
          2543 => x"09",
          2544 => x"e7",
          2545 => x"2a",
          2546 => x"77",
          2547 => x"51",
          2548 => x"2e",
          2549 => x"81",
          2550 => x"80",
          2551 => x"38",
          2552 => x"ab",
          2553 => x"55",
          2554 => x"75",
          2555 => x"73",
          2556 => x"55",
          2557 => x"82",
          2558 => x"06",
          2559 => x"ab",
          2560 => x"33",
          2561 => x"70",
          2562 => x"55",
          2563 => x"2e",
          2564 => x"1b",
          2565 => x"06",
          2566 => x"52",
          2567 => x"db",
          2568 => x"88",
          2569 => x"0c",
          2570 => x"74",
          2571 => x"0c",
          2572 => x"04",
          2573 => x"7c",
          2574 => x"08",
          2575 => x"55",
          2576 => x"59",
          2577 => x"81",
          2578 => x"70",
          2579 => x"33",
          2580 => x"52",
          2581 => x"2e",
          2582 => x"ee",
          2583 => x"2e",
          2584 => x"81",
          2585 => x"33",
          2586 => x"81",
          2587 => x"52",
          2588 => x"26",
          2589 => x"14",
          2590 => x"06",
          2591 => x"52",
          2592 => x"80",
          2593 => x"0b",
          2594 => x"59",
          2595 => x"7a",
          2596 => x"70",
          2597 => x"33",
          2598 => x"05",
          2599 => x"9f",
          2600 => x"53",
          2601 => x"89",
          2602 => x"70",
          2603 => x"54",
          2604 => x"12",
          2605 => x"26",
          2606 => x"12",
          2607 => x"06",
          2608 => x"30",
          2609 => x"51",
          2610 => x"2e",
          2611 => x"85",
          2612 => x"be",
          2613 => x"74",
          2614 => x"30",
          2615 => x"9f",
          2616 => x"2a",
          2617 => x"54",
          2618 => x"2e",
          2619 => x"15",
          2620 => x"55",
          2621 => x"ff",
          2622 => x"39",
          2623 => x"86",
          2624 => x"7c",
          2625 => x"51",
          2626 => x"ca",
          2627 => x"70",
          2628 => x"0c",
          2629 => x"04",
          2630 => x"78",
          2631 => x"83",
          2632 => x"0b",
          2633 => x"79",
          2634 => x"e2",
          2635 => x"55",
          2636 => x"08",
          2637 => x"84",
          2638 => x"df",
          2639 => x"ca",
          2640 => x"ff",
          2641 => x"83",
          2642 => x"d4",
          2643 => x"81",
          2644 => x"38",
          2645 => x"17",
          2646 => x"74",
          2647 => x"09",
          2648 => x"38",
          2649 => x"81",
          2650 => x"30",
          2651 => x"79",
          2652 => x"54",
          2653 => x"74",
          2654 => x"09",
          2655 => x"38",
          2656 => x"b8",
          2657 => x"ea",
          2658 => x"b1",
          2659 => x"88",
          2660 => x"ca",
          2661 => x"2e",
          2662 => x"53",
          2663 => x"52",
          2664 => x"51",
          2665 => x"91",
          2666 => x"55",
          2667 => x"08",
          2668 => x"38",
          2669 => x"91",
          2670 => x"88",
          2671 => x"f2",
          2672 => x"02",
          2673 => x"cb",
          2674 => x"55",
          2675 => x"60",
          2676 => x"3f",
          2677 => x"08",
          2678 => x"80",
          2679 => x"88",
          2680 => x"fc",
          2681 => x"88",
          2682 => x"91",
          2683 => x"70",
          2684 => x"8c",
          2685 => x"2e",
          2686 => x"73",
          2687 => x"81",
          2688 => x"33",
          2689 => x"80",
          2690 => x"81",
          2691 => x"d7",
          2692 => x"ca",
          2693 => x"ff",
          2694 => x"06",
          2695 => x"98",
          2696 => x"2e",
          2697 => x"74",
          2698 => x"81",
          2699 => x"8a",
          2700 => x"ac",
          2701 => x"39",
          2702 => x"77",
          2703 => x"81",
          2704 => x"33",
          2705 => x"3f",
          2706 => x"08",
          2707 => x"70",
          2708 => x"55",
          2709 => x"86",
          2710 => x"80",
          2711 => x"74",
          2712 => x"81",
          2713 => x"8a",
          2714 => x"f4",
          2715 => x"53",
          2716 => x"fd",
          2717 => x"ca",
          2718 => x"ff",
          2719 => x"82",
          2720 => x"06",
          2721 => x"8c",
          2722 => x"58",
          2723 => x"f6",
          2724 => x"58",
          2725 => x"2e",
          2726 => x"fa",
          2727 => x"e8",
          2728 => x"88",
          2729 => x"78",
          2730 => x"5a",
          2731 => x"90",
          2732 => x"75",
          2733 => x"38",
          2734 => x"3d",
          2735 => x"70",
          2736 => x"08",
          2737 => x"7a",
          2738 => x"38",
          2739 => x"51",
          2740 => x"91",
          2741 => x"81",
          2742 => x"81",
          2743 => x"38",
          2744 => x"83",
          2745 => x"38",
          2746 => x"84",
          2747 => x"38",
          2748 => x"81",
          2749 => x"38",
          2750 => x"db",
          2751 => x"ca",
          2752 => x"ff",
          2753 => x"72",
          2754 => x"09",
          2755 => x"d0",
          2756 => x"14",
          2757 => x"3f",
          2758 => x"08",
          2759 => x"06",
          2760 => x"38",
          2761 => x"51",
          2762 => x"91",
          2763 => x"58",
          2764 => x"0c",
          2765 => x"33",
          2766 => x"80",
          2767 => x"ff",
          2768 => x"ff",
          2769 => x"55",
          2770 => x"81",
          2771 => x"38",
          2772 => x"06",
          2773 => x"80",
          2774 => x"52",
          2775 => x"8a",
          2776 => x"80",
          2777 => x"ff",
          2778 => x"53",
          2779 => x"86",
          2780 => x"83",
          2781 => x"c5",
          2782 => x"f5",
          2783 => x"88",
          2784 => x"ca",
          2785 => x"15",
          2786 => x"06",
          2787 => x"76",
          2788 => x"80",
          2789 => x"da",
          2790 => x"ca",
          2791 => x"ff",
          2792 => x"74",
          2793 => x"d4",
          2794 => x"dc",
          2795 => x"88",
          2796 => x"c2",
          2797 => x"b9",
          2798 => x"88",
          2799 => x"ff",
          2800 => x"56",
          2801 => x"83",
          2802 => x"14",
          2803 => x"71",
          2804 => x"5a",
          2805 => x"26",
          2806 => x"8a",
          2807 => x"74",
          2808 => x"ff",
          2809 => x"91",
          2810 => x"55",
          2811 => x"08",
          2812 => x"ec",
          2813 => x"88",
          2814 => x"ff",
          2815 => x"83",
          2816 => x"74",
          2817 => x"26",
          2818 => x"57",
          2819 => x"26",
          2820 => x"57",
          2821 => x"56",
          2822 => x"82",
          2823 => x"15",
          2824 => x"0c",
          2825 => x"0c",
          2826 => x"a4",
          2827 => x"1d",
          2828 => x"54",
          2829 => x"2e",
          2830 => x"af",
          2831 => x"14",
          2832 => x"3f",
          2833 => x"08",
          2834 => x"06",
          2835 => x"72",
          2836 => x"79",
          2837 => x"80",
          2838 => x"d9",
          2839 => x"ca",
          2840 => x"15",
          2841 => x"2b",
          2842 => x"8d",
          2843 => x"2e",
          2844 => x"77",
          2845 => x"0c",
          2846 => x"76",
          2847 => x"38",
          2848 => x"70",
          2849 => x"81",
          2850 => x"53",
          2851 => x"89",
          2852 => x"56",
          2853 => x"08",
          2854 => x"38",
          2855 => x"15",
          2856 => x"8c",
          2857 => x"80",
          2858 => x"34",
          2859 => x"09",
          2860 => x"92",
          2861 => x"14",
          2862 => x"3f",
          2863 => x"08",
          2864 => x"06",
          2865 => x"2e",
          2866 => x"80",
          2867 => x"1b",
          2868 => x"db",
          2869 => x"ca",
          2870 => x"ea",
          2871 => x"88",
          2872 => x"34",
          2873 => x"51",
          2874 => x"91",
          2875 => x"83",
          2876 => x"53",
          2877 => x"d5",
          2878 => x"06",
          2879 => x"b4",
          2880 => x"84",
          2881 => x"88",
          2882 => x"85",
          2883 => x"09",
          2884 => x"38",
          2885 => x"51",
          2886 => x"91",
          2887 => x"86",
          2888 => x"f2",
          2889 => x"06",
          2890 => x"9c",
          2891 => x"d8",
          2892 => x"88",
          2893 => x"0c",
          2894 => x"51",
          2895 => x"91",
          2896 => x"8c",
          2897 => x"74",
          2898 => x"b4",
          2899 => x"53",
          2900 => x"b4",
          2901 => x"15",
          2902 => x"94",
          2903 => x"56",
          2904 => x"88",
          2905 => x"0d",
          2906 => x"0d",
          2907 => x"55",
          2908 => x"b9",
          2909 => x"53",
          2910 => x"b1",
          2911 => x"52",
          2912 => x"a9",
          2913 => x"22",
          2914 => x"57",
          2915 => x"2e",
          2916 => x"99",
          2917 => x"33",
          2918 => x"3f",
          2919 => x"08",
          2920 => x"71",
          2921 => x"74",
          2922 => x"83",
          2923 => x"78",
          2924 => x"52",
          2925 => x"88",
          2926 => x"0d",
          2927 => x"0d",
          2928 => x"33",
          2929 => x"3d",
          2930 => x"56",
          2931 => x"8b",
          2932 => x"91",
          2933 => x"24",
          2934 => x"ca",
          2935 => x"29",
          2936 => x"05",
          2937 => x"55",
          2938 => x"84",
          2939 => x"34",
          2940 => x"80",
          2941 => x"80",
          2942 => x"75",
          2943 => x"75",
          2944 => x"38",
          2945 => x"3d",
          2946 => x"05",
          2947 => x"3f",
          2948 => x"08",
          2949 => x"ca",
          2950 => x"3d",
          2951 => x"3d",
          2952 => x"84",
          2953 => x"05",
          2954 => x"89",
          2955 => x"2e",
          2956 => x"77",
          2957 => x"54",
          2958 => x"05",
          2959 => x"84",
          2960 => x"f6",
          2961 => x"ca",
          2962 => x"91",
          2963 => x"84",
          2964 => x"5c",
          2965 => x"3d",
          2966 => x"ed",
          2967 => x"ca",
          2968 => x"91",
          2969 => x"92",
          2970 => x"d7",
          2971 => x"98",
          2972 => x"73",
          2973 => x"38",
          2974 => x"9c",
          2975 => x"80",
          2976 => x"38",
          2977 => x"95",
          2978 => x"2e",
          2979 => x"aa",
          2980 => x"ea",
          2981 => x"ca",
          2982 => x"9e",
          2983 => x"05",
          2984 => x"54",
          2985 => x"38",
          2986 => x"70",
          2987 => x"54",
          2988 => x"8e",
          2989 => x"83",
          2990 => x"88",
          2991 => x"83",
          2992 => x"83",
          2993 => x"06",
          2994 => x"80",
          2995 => x"38",
          2996 => x"51",
          2997 => x"91",
          2998 => x"56",
          2999 => x"0a",
          3000 => x"05",
          3001 => x"3f",
          3002 => x"0b",
          3003 => x"80",
          3004 => x"7a",
          3005 => x"3f",
          3006 => x"9c",
          3007 => x"d1",
          3008 => x"81",
          3009 => x"34",
          3010 => x"80",
          3011 => x"b0",
          3012 => x"54",
          3013 => x"52",
          3014 => x"05",
          3015 => x"3f",
          3016 => x"08",
          3017 => x"88",
          3018 => x"38",
          3019 => x"82",
          3020 => x"b2",
          3021 => x"84",
          3022 => x"06",
          3023 => x"73",
          3024 => x"38",
          3025 => x"ad",
          3026 => x"2a",
          3027 => x"51",
          3028 => x"2e",
          3029 => x"81",
          3030 => x"80",
          3031 => x"87",
          3032 => x"39",
          3033 => x"51",
          3034 => x"91",
          3035 => x"7b",
          3036 => x"12",
          3037 => x"91",
          3038 => x"81",
          3039 => x"83",
          3040 => x"06",
          3041 => x"80",
          3042 => x"77",
          3043 => x"58",
          3044 => x"08",
          3045 => x"63",
          3046 => x"63",
          3047 => x"57",
          3048 => x"91",
          3049 => x"91",
          3050 => x"88",
          3051 => x"9c",
          3052 => x"d2",
          3053 => x"ca",
          3054 => x"ca",
          3055 => x"1b",
          3056 => x"0c",
          3057 => x"22",
          3058 => x"77",
          3059 => x"80",
          3060 => x"34",
          3061 => x"1a",
          3062 => x"94",
          3063 => x"85",
          3064 => x"06",
          3065 => x"80",
          3066 => x"38",
          3067 => x"08",
          3068 => x"84",
          3069 => x"88",
          3070 => x"0c",
          3071 => x"70",
          3072 => x"52",
          3073 => x"39",
          3074 => x"51",
          3075 => x"91",
          3076 => x"57",
          3077 => x"08",
          3078 => x"38",
          3079 => x"ca",
          3080 => x"2e",
          3081 => x"83",
          3082 => x"75",
          3083 => x"74",
          3084 => x"07",
          3085 => x"54",
          3086 => x"8a",
          3087 => x"75",
          3088 => x"73",
          3089 => x"98",
          3090 => x"a9",
          3091 => x"ff",
          3092 => x"80",
          3093 => x"76",
          3094 => x"d6",
          3095 => x"ca",
          3096 => x"38",
          3097 => x"39",
          3098 => x"91",
          3099 => x"05",
          3100 => x"84",
          3101 => x"0c",
          3102 => x"91",
          3103 => x"97",
          3104 => x"f2",
          3105 => x"63",
          3106 => x"40",
          3107 => x"7e",
          3108 => x"fc",
          3109 => x"51",
          3110 => x"91",
          3111 => x"55",
          3112 => x"08",
          3113 => x"19",
          3114 => x"80",
          3115 => x"74",
          3116 => x"39",
          3117 => x"81",
          3118 => x"56",
          3119 => x"82",
          3120 => x"39",
          3121 => x"1a",
          3122 => x"82",
          3123 => x"0b",
          3124 => x"81",
          3125 => x"39",
          3126 => x"94",
          3127 => x"55",
          3128 => x"83",
          3129 => x"7b",
          3130 => x"89",
          3131 => x"08",
          3132 => x"06",
          3133 => x"81",
          3134 => x"8a",
          3135 => x"05",
          3136 => x"06",
          3137 => x"a8",
          3138 => x"38",
          3139 => x"55",
          3140 => x"19",
          3141 => x"51",
          3142 => x"91",
          3143 => x"55",
          3144 => x"ff",
          3145 => x"ff",
          3146 => x"38",
          3147 => x"0c",
          3148 => x"52",
          3149 => x"cb",
          3150 => x"88",
          3151 => x"ff",
          3152 => x"ca",
          3153 => x"7c",
          3154 => x"57",
          3155 => x"80",
          3156 => x"1a",
          3157 => x"22",
          3158 => x"75",
          3159 => x"38",
          3160 => x"58",
          3161 => x"53",
          3162 => x"1b",
          3163 => x"88",
          3164 => x"88",
          3165 => x"38",
          3166 => x"33",
          3167 => x"80",
          3168 => x"b0",
          3169 => x"31",
          3170 => x"27",
          3171 => x"80",
          3172 => x"52",
          3173 => x"77",
          3174 => x"7d",
          3175 => x"e0",
          3176 => x"2b",
          3177 => x"76",
          3178 => x"94",
          3179 => x"ff",
          3180 => x"71",
          3181 => x"7b",
          3182 => x"38",
          3183 => x"19",
          3184 => x"51",
          3185 => x"91",
          3186 => x"fe",
          3187 => x"53",
          3188 => x"83",
          3189 => x"b4",
          3190 => x"51",
          3191 => x"7b",
          3192 => x"08",
          3193 => x"76",
          3194 => x"08",
          3195 => x"0c",
          3196 => x"f3",
          3197 => x"75",
          3198 => x"0c",
          3199 => x"04",
          3200 => x"60",
          3201 => x"40",
          3202 => x"80",
          3203 => x"3d",
          3204 => x"77",
          3205 => x"3f",
          3206 => x"08",
          3207 => x"88",
          3208 => x"91",
          3209 => x"74",
          3210 => x"38",
          3211 => x"b8",
          3212 => x"33",
          3213 => x"70",
          3214 => x"56",
          3215 => x"74",
          3216 => x"a4",
          3217 => x"82",
          3218 => x"34",
          3219 => x"98",
          3220 => x"91",
          3221 => x"56",
          3222 => x"94",
          3223 => x"11",
          3224 => x"76",
          3225 => x"75",
          3226 => x"80",
          3227 => x"38",
          3228 => x"70",
          3229 => x"56",
          3230 => x"fd",
          3231 => x"11",
          3232 => x"77",
          3233 => x"5c",
          3234 => x"38",
          3235 => x"88",
          3236 => x"74",
          3237 => x"52",
          3238 => x"18",
          3239 => x"51",
          3240 => x"91",
          3241 => x"55",
          3242 => x"08",
          3243 => x"ab",
          3244 => x"2e",
          3245 => x"74",
          3246 => x"95",
          3247 => x"19",
          3248 => x"08",
          3249 => x"88",
          3250 => x"55",
          3251 => x"9c",
          3252 => x"09",
          3253 => x"38",
          3254 => x"c1",
          3255 => x"88",
          3256 => x"38",
          3257 => x"52",
          3258 => x"97",
          3259 => x"88",
          3260 => x"fe",
          3261 => x"ca",
          3262 => x"7c",
          3263 => x"57",
          3264 => x"80",
          3265 => x"1b",
          3266 => x"22",
          3267 => x"75",
          3268 => x"38",
          3269 => x"59",
          3270 => x"53",
          3271 => x"1a",
          3272 => x"be",
          3273 => x"88",
          3274 => x"38",
          3275 => x"08",
          3276 => x"56",
          3277 => x"9b",
          3278 => x"53",
          3279 => x"77",
          3280 => x"7d",
          3281 => x"16",
          3282 => x"3f",
          3283 => x"0b",
          3284 => x"78",
          3285 => x"80",
          3286 => x"18",
          3287 => x"08",
          3288 => x"7e",
          3289 => x"3f",
          3290 => x"08",
          3291 => x"7e",
          3292 => x"0c",
          3293 => x"19",
          3294 => x"08",
          3295 => x"84",
          3296 => x"57",
          3297 => x"27",
          3298 => x"56",
          3299 => x"52",
          3300 => x"f9",
          3301 => x"88",
          3302 => x"38",
          3303 => x"52",
          3304 => x"83",
          3305 => x"b4",
          3306 => x"d4",
          3307 => x"81",
          3308 => x"34",
          3309 => x"7e",
          3310 => x"0c",
          3311 => x"1a",
          3312 => x"94",
          3313 => x"1b",
          3314 => x"5e",
          3315 => x"27",
          3316 => x"55",
          3317 => x"0c",
          3318 => x"90",
          3319 => x"c0",
          3320 => x"90",
          3321 => x"56",
          3322 => x"88",
          3323 => x"0d",
          3324 => x"0d",
          3325 => x"fc",
          3326 => x"52",
          3327 => x"3f",
          3328 => x"08",
          3329 => x"88",
          3330 => x"38",
          3331 => x"70",
          3332 => x"81",
          3333 => x"55",
          3334 => x"80",
          3335 => x"16",
          3336 => x"51",
          3337 => x"91",
          3338 => x"57",
          3339 => x"08",
          3340 => x"a4",
          3341 => x"11",
          3342 => x"55",
          3343 => x"16",
          3344 => x"08",
          3345 => x"75",
          3346 => x"e8",
          3347 => x"08",
          3348 => x"51",
          3349 => x"82",
          3350 => x"52",
          3351 => x"c9",
          3352 => x"52",
          3353 => x"c9",
          3354 => x"54",
          3355 => x"15",
          3356 => x"cc",
          3357 => x"ca",
          3358 => x"17",
          3359 => x"06",
          3360 => x"90",
          3361 => x"91",
          3362 => x"8a",
          3363 => x"fc",
          3364 => x"70",
          3365 => x"d9",
          3366 => x"88",
          3367 => x"ca",
          3368 => x"38",
          3369 => x"05",
          3370 => x"f1",
          3371 => x"ca",
          3372 => x"91",
          3373 => x"87",
          3374 => x"88",
          3375 => x"72",
          3376 => x"0c",
          3377 => x"04",
          3378 => x"84",
          3379 => x"e4",
          3380 => x"80",
          3381 => x"88",
          3382 => x"38",
          3383 => x"08",
          3384 => x"34",
          3385 => x"91",
          3386 => x"83",
          3387 => x"ef",
          3388 => x"53",
          3389 => x"05",
          3390 => x"51",
          3391 => x"91",
          3392 => x"55",
          3393 => x"08",
          3394 => x"76",
          3395 => x"93",
          3396 => x"51",
          3397 => x"91",
          3398 => x"55",
          3399 => x"08",
          3400 => x"80",
          3401 => x"70",
          3402 => x"56",
          3403 => x"89",
          3404 => x"94",
          3405 => x"b2",
          3406 => x"05",
          3407 => x"2a",
          3408 => x"51",
          3409 => x"80",
          3410 => x"76",
          3411 => x"52",
          3412 => x"3f",
          3413 => x"08",
          3414 => x"8e",
          3415 => x"88",
          3416 => x"09",
          3417 => x"38",
          3418 => x"91",
          3419 => x"93",
          3420 => x"e4",
          3421 => x"6f",
          3422 => x"7a",
          3423 => x"9e",
          3424 => x"05",
          3425 => x"51",
          3426 => x"91",
          3427 => x"57",
          3428 => x"08",
          3429 => x"7b",
          3430 => x"94",
          3431 => x"55",
          3432 => x"73",
          3433 => x"ed",
          3434 => x"93",
          3435 => x"55",
          3436 => x"91",
          3437 => x"57",
          3438 => x"08",
          3439 => x"68",
          3440 => x"c9",
          3441 => x"ca",
          3442 => x"91",
          3443 => x"82",
          3444 => x"52",
          3445 => x"a3",
          3446 => x"88",
          3447 => x"52",
          3448 => x"b8",
          3449 => x"88",
          3450 => x"ca",
          3451 => x"a2",
          3452 => x"74",
          3453 => x"3f",
          3454 => x"08",
          3455 => x"88",
          3456 => x"69",
          3457 => x"d9",
          3458 => x"91",
          3459 => x"2e",
          3460 => x"52",
          3461 => x"cf",
          3462 => x"88",
          3463 => x"ca",
          3464 => x"2e",
          3465 => x"84",
          3466 => x"06",
          3467 => x"57",
          3468 => x"76",
          3469 => x"9e",
          3470 => x"05",
          3471 => x"dc",
          3472 => x"90",
          3473 => x"81",
          3474 => x"56",
          3475 => x"80",
          3476 => x"02",
          3477 => x"81",
          3478 => x"70",
          3479 => x"56",
          3480 => x"81",
          3481 => x"78",
          3482 => x"38",
          3483 => x"99",
          3484 => x"81",
          3485 => x"18",
          3486 => x"18",
          3487 => x"58",
          3488 => x"33",
          3489 => x"ee",
          3490 => x"6f",
          3491 => x"af",
          3492 => x"8d",
          3493 => x"2e",
          3494 => x"8a",
          3495 => x"6f",
          3496 => x"af",
          3497 => x"0b",
          3498 => x"33",
          3499 => x"91",
          3500 => x"70",
          3501 => x"52",
          3502 => x"56",
          3503 => x"8d",
          3504 => x"70",
          3505 => x"51",
          3506 => x"f5",
          3507 => x"54",
          3508 => x"a7",
          3509 => x"74",
          3510 => x"38",
          3511 => x"73",
          3512 => x"81",
          3513 => x"81",
          3514 => x"39",
          3515 => x"81",
          3516 => x"74",
          3517 => x"81",
          3518 => x"91",
          3519 => x"6e",
          3520 => x"59",
          3521 => x"7a",
          3522 => x"5c",
          3523 => x"26",
          3524 => x"7a",
          3525 => x"ca",
          3526 => x"3d",
          3527 => x"3d",
          3528 => x"8d",
          3529 => x"54",
          3530 => x"55",
          3531 => x"91",
          3532 => x"53",
          3533 => x"08",
          3534 => x"91",
          3535 => x"72",
          3536 => x"8c",
          3537 => x"73",
          3538 => x"38",
          3539 => x"70",
          3540 => x"81",
          3541 => x"57",
          3542 => x"73",
          3543 => x"08",
          3544 => x"94",
          3545 => x"75",
          3546 => x"97",
          3547 => x"11",
          3548 => x"2b",
          3549 => x"73",
          3550 => x"38",
          3551 => x"16",
          3552 => x"e5",
          3553 => x"88",
          3554 => x"78",
          3555 => x"55",
          3556 => x"d5",
          3557 => x"88",
          3558 => x"96",
          3559 => x"70",
          3560 => x"94",
          3561 => x"71",
          3562 => x"08",
          3563 => x"53",
          3564 => x"15",
          3565 => x"a6",
          3566 => x"74",
          3567 => x"3f",
          3568 => x"08",
          3569 => x"88",
          3570 => x"81",
          3571 => x"ca",
          3572 => x"2e",
          3573 => x"91",
          3574 => x"88",
          3575 => x"98",
          3576 => x"80",
          3577 => x"38",
          3578 => x"80",
          3579 => x"77",
          3580 => x"08",
          3581 => x"0c",
          3582 => x"70",
          3583 => x"81",
          3584 => x"5a",
          3585 => x"2e",
          3586 => x"52",
          3587 => x"f9",
          3588 => x"88",
          3589 => x"ca",
          3590 => x"38",
          3591 => x"08",
          3592 => x"73",
          3593 => x"c7",
          3594 => x"ca",
          3595 => x"73",
          3596 => x"38",
          3597 => x"af",
          3598 => x"73",
          3599 => x"27",
          3600 => x"98",
          3601 => x"a0",
          3602 => x"08",
          3603 => x"0c",
          3604 => x"06",
          3605 => x"2e",
          3606 => x"52",
          3607 => x"a3",
          3608 => x"88",
          3609 => x"82",
          3610 => x"34",
          3611 => x"c4",
          3612 => x"91",
          3613 => x"53",
          3614 => x"89",
          3615 => x"88",
          3616 => x"94",
          3617 => x"8c",
          3618 => x"27",
          3619 => x"8c",
          3620 => x"15",
          3621 => x"07",
          3622 => x"16",
          3623 => x"ff",
          3624 => x"80",
          3625 => x"77",
          3626 => x"2e",
          3627 => x"9c",
          3628 => x"53",
          3629 => x"88",
          3630 => x"0d",
          3631 => x"0d",
          3632 => x"54",
          3633 => x"81",
          3634 => x"53",
          3635 => x"05",
          3636 => x"84",
          3637 => x"e7",
          3638 => x"88",
          3639 => x"ca",
          3640 => x"ea",
          3641 => x"0c",
          3642 => x"51",
          3643 => x"91",
          3644 => x"55",
          3645 => x"08",
          3646 => x"ab",
          3647 => x"98",
          3648 => x"80",
          3649 => x"38",
          3650 => x"70",
          3651 => x"81",
          3652 => x"57",
          3653 => x"ad",
          3654 => x"08",
          3655 => x"d3",
          3656 => x"ca",
          3657 => x"17",
          3658 => x"86",
          3659 => x"17",
          3660 => x"75",
          3661 => x"3f",
          3662 => x"08",
          3663 => x"2e",
          3664 => x"85",
          3665 => x"86",
          3666 => x"2e",
          3667 => x"76",
          3668 => x"73",
          3669 => x"0c",
          3670 => x"04",
          3671 => x"76",
          3672 => x"05",
          3673 => x"53",
          3674 => x"91",
          3675 => x"87",
          3676 => x"88",
          3677 => x"86",
          3678 => x"fb",
          3679 => x"79",
          3680 => x"05",
          3681 => x"56",
          3682 => x"3f",
          3683 => x"08",
          3684 => x"88",
          3685 => x"38",
          3686 => x"91",
          3687 => x"52",
          3688 => x"f8",
          3689 => x"88",
          3690 => x"ca",
          3691 => x"88",
          3692 => x"51",
          3693 => x"91",
          3694 => x"53",
          3695 => x"08",
          3696 => x"81",
          3697 => x"80",
          3698 => x"91",
          3699 => x"a6",
          3700 => x"73",
          3701 => x"3f",
          3702 => x"51",
          3703 => x"91",
          3704 => x"84",
          3705 => x"70",
          3706 => x"2c",
          3707 => x"88",
          3708 => x"51",
          3709 => x"91",
          3710 => x"87",
          3711 => x"ee",
          3712 => x"57",
          3713 => x"3d",
          3714 => x"3d",
          3715 => x"af",
          3716 => x"88",
          3717 => x"ca",
          3718 => x"38",
          3719 => x"51",
          3720 => x"91",
          3721 => x"55",
          3722 => x"08",
          3723 => x"80",
          3724 => x"70",
          3725 => x"58",
          3726 => x"85",
          3727 => x"8d",
          3728 => x"2e",
          3729 => x"52",
          3730 => x"be",
          3731 => x"ca",
          3732 => x"3d",
          3733 => x"3d",
          3734 => x"55",
          3735 => x"92",
          3736 => x"52",
          3737 => x"de",
          3738 => x"ca",
          3739 => x"91",
          3740 => x"82",
          3741 => x"74",
          3742 => x"98",
          3743 => x"11",
          3744 => x"59",
          3745 => x"75",
          3746 => x"38",
          3747 => x"81",
          3748 => x"5b",
          3749 => x"82",
          3750 => x"39",
          3751 => x"08",
          3752 => x"59",
          3753 => x"09",
          3754 => x"38",
          3755 => x"57",
          3756 => x"3d",
          3757 => x"c1",
          3758 => x"ca",
          3759 => x"2e",
          3760 => x"ca",
          3761 => x"2e",
          3762 => x"ca",
          3763 => x"70",
          3764 => x"08",
          3765 => x"7a",
          3766 => x"7f",
          3767 => x"54",
          3768 => x"77",
          3769 => x"80",
          3770 => x"15",
          3771 => x"88",
          3772 => x"75",
          3773 => x"52",
          3774 => x"52",
          3775 => x"8d",
          3776 => x"88",
          3777 => x"ca",
          3778 => x"d6",
          3779 => x"33",
          3780 => x"1a",
          3781 => x"54",
          3782 => x"09",
          3783 => x"38",
          3784 => x"ff",
          3785 => x"91",
          3786 => x"83",
          3787 => x"70",
          3788 => x"25",
          3789 => x"59",
          3790 => x"9b",
          3791 => x"51",
          3792 => x"3f",
          3793 => x"08",
          3794 => x"70",
          3795 => x"25",
          3796 => x"59",
          3797 => x"75",
          3798 => x"7a",
          3799 => x"ff",
          3800 => x"7c",
          3801 => x"90",
          3802 => x"11",
          3803 => x"56",
          3804 => x"15",
          3805 => x"ca",
          3806 => x"3d",
          3807 => x"3d",
          3808 => x"3d",
          3809 => x"70",
          3810 => x"dd",
          3811 => x"88",
          3812 => x"ca",
          3813 => x"a8",
          3814 => x"33",
          3815 => x"a0",
          3816 => x"33",
          3817 => x"70",
          3818 => x"55",
          3819 => x"73",
          3820 => x"8e",
          3821 => x"08",
          3822 => x"18",
          3823 => x"80",
          3824 => x"38",
          3825 => x"08",
          3826 => x"08",
          3827 => x"c4",
          3828 => x"ca",
          3829 => x"88",
          3830 => x"80",
          3831 => x"17",
          3832 => x"51",
          3833 => x"3f",
          3834 => x"08",
          3835 => x"81",
          3836 => x"81",
          3837 => x"88",
          3838 => x"09",
          3839 => x"38",
          3840 => x"39",
          3841 => x"77",
          3842 => x"88",
          3843 => x"08",
          3844 => x"98",
          3845 => x"91",
          3846 => x"52",
          3847 => x"bd",
          3848 => x"88",
          3849 => x"17",
          3850 => x"0c",
          3851 => x"80",
          3852 => x"73",
          3853 => x"75",
          3854 => x"38",
          3855 => x"34",
          3856 => x"91",
          3857 => x"89",
          3858 => x"e2",
          3859 => x"53",
          3860 => x"a4",
          3861 => x"3d",
          3862 => x"3f",
          3863 => x"08",
          3864 => x"88",
          3865 => x"38",
          3866 => x"3d",
          3867 => x"3d",
          3868 => x"d1",
          3869 => x"ca",
          3870 => x"91",
          3871 => x"81",
          3872 => x"80",
          3873 => x"70",
          3874 => x"81",
          3875 => x"56",
          3876 => x"81",
          3877 => x"98",
          3878 => x"74",
          3879 => x"38",
          3880 => x"05",
          3881 => x"06",
          3882 => x"55",
          3883 => x"38",
          3884 => x"51",
          3885 => x"91",
          3886 => x"74",
          3887 => x"81",
          3888 => x"56",
          3889 => x"80",
          3890 => x"54",
          3891 => x"08",
          3892 => x"2e",
          3893 => x"73",
          3894 => x"88",
          3895 => x"52",
          3896 => x"52",
          3897 => x"3f",
          3898 => x"08",
          3899 => x"88",
          3900 => x"38",
          3901 => x"08",
          3902 => x"cc",
          3903 => x"ca",
          3904 => x"91",
          3905 => x"86",
          3906 => x"80",
          3907 => x"ca",
          3908 => x"2e",
          3909 => x"ca",
          3910 => x"c0",
          3911 => x"ce",
          3912 => x"ca",
          3913 => x"ca",
          3914 => x"70",
          3915 => x"08",
          3916 => x"51",
          3917 => x"80",
          3918 => x"73",
          3919 => x"38",
          3920 => x"52",
          3921 => x"95",
          3922 => x"88",
          3923 => x"8c",
          3924 => x"ff",
          3925 => x"91",
          3926 => x"55",
          3927 => x"88",
          3928 => x"0d",
          3929 => x"0d",
          3930 => x"3d",
          3931 => x"9a",
          3932 => x"cb",
          3933 => x"88",
          3934 => x"ca",
          3935 => x"b0",
          3936 => x"69",
          3937 => x"70",
          3938 => x"97",
          3939 => x"88",
          3940 => x"ca",
          3941 => x"38",
          3942 => x"94",
          3943 => x"88",
          3944 => x"09",
          3945 => x"88",
          3946 => x"df",
          3947 => x"85",
          3948 => x"51",
          3949 => x"74",
          3950 => x"78",
          3951 => x"8a",
          3952 => x"57",
          3953 => x"91",
          3954 => x"75",
          3955 => x"ca",
          3956 => x"38",
          3957 => x"ca",
          3958 => x"2e",
          3959 => x"83",
          3960 => x"91",
          3961 => x"ff",
          3962 => x"06",
          3963 => x"54",
          3964 => x"73",
          3965 => x"91",
          3966 => x"52",
          3967 => x"a4",
          3968 => x"88",
          3969 => x"ca",
          3970 => x"9a",
          3971 => x"a0",
          3972 => x"51",
          3973 => x"3f",
          3974 => x"0b",
          3975 => x"78",
          3976 => x"bf",
          3977 => x"88",
          3978 => x"80",
          3979 => x"ff",
          3980 => x"75",
          3981 => x"11",
          3982 => x"f8",
          3983 => x"78",
          3984 => x"80",
          3985 => x"ff",
          3986 => x"78",
          3987 => x"80",
          3988 => x"7f",
          3989 => x"d4",
          3990 => x"c9",
          3991 => x"54",
          3992 => x"15",
          3993 => x"cb",
          3994 => x"ca",
          3995 => x"91",
          3996 => x"b2",
          3997 => x"b2",
          3998 => x"96",
          3999 => x"b5",
          4000 => x"53",
          4001 => x"51",
          4002 => x"64",
          4003 => x"8b",
          4004 => x"54",
          4005 => x"15",
          4006 => x"ff",
          4007 => x"91",
          4008 => x"54",
          4009 => x"53",
          4010 => x"51",
          4011 => x"3f",
          4012 => x"88",
          4013 => x"0d",
          4014 => x"0d",
          4015 => x"05",
          4016 => x"3f",
          4017 => x"3d",
          4018 => x"52",
          4019 => x"d5",
          4020 => x"ca",
          4021 => x"91",
          4022 => x"82",
          4023 => x"4d",
          4024 => x"52",
          4025 => x"52",
          4026 => x"3f",
          4027 => x"08",
          4028 => x"88",
          4029 => x"38",
          4030 => x"05",
          4031 => x"06",
          4032 => x"73",
          4033 => x"a0",
          4034 => x"08",
          4035 => x"ff",
          4036 => x"ff",
          4037 => x"ac",
          4038 => x"92",
          4039 => x"54",
          4040 => x"3f",
          4041 => x"52",
          4042 => x"f7",
          4043 => x"88",
          4044 => x"ca",
          4045 => x"38",
          4046 => x"09",
          4047 => x"38",
          4048 => x"08",
          4049 => x"88",
          4050 => x"39",
          4051 => x"08",
          4052 => x"81",
          4053 => x"38",
          4054 => x"b1",
          4055 => x"88",
          4056 => x"ca",
          4057 => x"c8",
          4058 => x"93",
          4059 => x"ff",
          4060 => x"8d",
          4061 => x"b4",
          4062 => x"af",
          4063 => x"17",
          4064 => x"33",
          4065 => x"70",
          4066 => x"55",
          4067 => x"38",
          4068 => x"54",
          4069 => x"34",
          4070 => x"0b",
          4071 => x"8b",
          4072 => x"84",
          4073 => x"06",
          4074 => x"73",
          4075 => x"e5",
          4076 => x"2e",
          4077 => x"75",
          4078 => x"c6",
          4079 => x"ca",
          4080 => x"78",
          4081 => x"bb",
          4082 => x"91",
          4083 => x"80",
          4084 => x"38",
          4085 => x"08",
          4086 => x"ff",
          4087 => x"91",
          4088 => x"79",
          4089 => x"58",
          4090 => x"ca",
          4091 => x"c0",
          4092 => x"33",
          4093 => x"2e",
          4094 => x"99",
          4095 => x"75",
          4096 => x"c6",
          4097 => x"54",
          4098 => x"15",
          4099 => x"91",
          4100 => x"9c",
          4101 => x"c8",
          4102 => x"ca",
          4103 => x"91",
          4104 => x"8c",
          4105 => x"ff",
          4106 => x"91",
          4107 => x"55",
          4108 => x"88",
          4109 => x"0d",
          4110 => x"0d",
          4111 => x"05",
          4112 => x"05",
          4113 => x"33",
          4114 => x"53",
          4115 => x"05",
          4116 => x"51",
          4117 => x"91",
          4118 => x"55",
          4119 => x"08",
          4120 => x"78",
          4121 => x"95",
          4122 => x"51",
          4123 => x"91",
          4124 => x"55",
          4125 => x"08",
          4126 => x"80",
          4127 => x"81",
          4128 => x"86",
          4129 => x"38",
          4130 => x"61",
          4131 => x"12",
          4132 => x"7a",
          4133 => x"51",
          4134 => x"74",
          4135 => x"78",
          4136 => x"83",
          4137 => x"51",
          4138 => x"3f",
          4139 => x"08",
          4140 => x"ca",
          4141 => x"3d",
          4142 => x"3d",
          4143 => x"82",
          4144 => x"d0",
          4145 => x"3d",
          4146 => x"3f",
          4147 => x"08",
          4148 => x"88",
          4149 => x"38",
          4150 => x"52",
          4151 => x"05",
          4152 => x"3f",
          4153 => x"08",
          4154 => x"88",
          4155 => x"02",
          4156 => x"33",
          4157 => x"54",
          4158 => x"a6",
          4159 => x"22",
          4160 => x"71",
          4161 => x"53",
          4162 => x"51",
          4163 => x"3f",
          4164 => x"0b",
          4165 => x"76",
          4166 => x"b8",
          4167 => x"88",
          4168 => x"91",
          4169 => x"93",
          4170 => x"ea",
          4171 => x"6b",
          4172 => x"53",
          4173 => x"05",
          4174 => x"51",
          4175 => x"91",
          4176 => x"91",
          4177 => x"30",
          4178 => x"88",
          4179 => x"25",
          4180 => x"79",
          4181 => x"85",
          4182 => x"75",
          4183 => x"73",
          4184 => x"f9",
          4185 => x"80",
          4186 => x"8d",
          4187 => x"54",
          4188 => x"3f",
          4189 => x"08",
          4190 => x"88",
          4191 => x"38",
          4192 => x"51",
          4193 => x"91",
          4194 => x"57",
          4195 => x"08",
          4196 => x"ca",
          4197 => x"ca",
          4198 => x"5b",
          4199 => x"18",
          4200 => x"18",
          4201 => x"74",
          4202 => x"81",
          4203 => x"78",
          4204 => x"8b",
          4205 => x"54",
          4206 => x"75",
          4207 => x"38",
          4208 => x"1b",
          4209 => x"55",
          4210 => x"2e",
          4211 => x"39",
          4212 => x"09",
          4213 => x"38",
          4214 => x"80",
          4215 => x"70",
          4216 => x"25",
          4217 => x"80",
          4218 => x"38",
          4219 => x"bc",
          4220 => x"11",
          4221 => x"ff",
          4222 => x"91",
          4223 => x"57",
          4224 => x"08",
          4225 => x"70",
          4226 => x"80",
          4227 => x"83",
          4228 => x"80",
          4229 => x"84",
          4230 => x"a7",
          4231 => x"b4",
          4232 => x"ad",
          4233 => x"ca",
          4234 => x"0c",
          4235 => x"88",
          4236 => x"0d",
          4237 => x"0d",
          4238 => x"3d",
          4239 => x"52",
          4240 => x"ce",
          4241 => x"ca",
          4242 => x"ca",
          4243 => x"54",
          4244 => x"08",
          4245 => x"8b",
          4246 => x"8b",
          4247 => x"59",
          4248 => x"3f",
          4249 => x"33",
          4250 => x"06",
          4251 => x"57",
          4252 => x"81",
          4253 => x"58",
          4254 => x"06",
          4255 => x"4e",
          4256 => x"ff",
          4257 => x"91",
          4258 => x"80",
          4259 => x"6c",
          4260 => x"53",
          4261 => x"ae",
          4262 => x"ca",
          4263 => x"2e",
          4264 => x"88",
          4265 => x"6d",
          4266 => x"55",
          4267 => x"ca",
          4268 => x"ff",
          4269 => x"83",
          4270 => x"51",
          4271 => x"26",
          4272 => x"15",
          4273 => x"ff",
          4274 => x"80",
          4275 => x"87",
          4276 => x"94",
          4277 => x"74",
          4278 => x"38",
          4279 => x"ba",
          4280 => x"ae",
          4281 => x"ca",
          4282 => x"38",
          4283 => x"27",
          4284 => x"89",
          4285 => x"8b",
          4286 => x"27",
          4287 => x"55",
          4288 => x"81",
          4289 => x"8f",
          4290 => x"2a",
          4291 => x"70",
          4292 => x"34",
          4293 => x"74",
          4294 => x"05",
          4295 => x"17",
          4296 => x"70",
          4297 => x"52",
          4298 => x"73",
          4299 => x"c8",
          4300 => x"33",
          4301 => x"73",
          4302 => x"81",
          4303 => x"80",
          4304 => x"02",
          4305 => x"76",
          4306 => x"51",
          4307 => x"2e",
          4308 => x"87",
          4309 => x"57",
          4310 => x"79",
          4311 => x"80",
          4312 => x"70",
          4313 => x"ba",
          4314 => x"ca",
          4315 => x"91",
          4316 => x"80",
          4317 => x"52",
          4318 => x"bf",
          4319 => x"ca",
          4320 => x"91",
          4321 => x"8d",
          4322 => x"c4",
          4323 => x"e5",
          4324 => x"c6",
          4325 => x"88",
          4326 => x"09",
          4327 => x"cc",
          4328 => x"76",
          4329 => x"c4",
          4330 => x"74",
          4331 => x"b0",
          4332 => x"88",
          4333 => x"ca",
          4334 => x"38",
          4335 => x"ca",
          4336 => x"67",
          4337 => x"db",
          4338 => x"88",
          4339 => x"34",
          4340 => x"52",
          4341 => x"ab",
          4342 => x"54",
          4343 => x"15",
          4344 => x"ff",
          4345 => x"91",
          4346 => x"54",
          4347 => x"91",
          4348 => x"9c",
          4349 => x"f2",
          4350 => x"62",
          4351 => x"80",
          4352 => x"93",
          4353 => x"55",
          4354 => x"5e",
          4355 => x"3f",
          4356 => x"08",
          4357 => x"88",
          4358 => x"38",
          4359 => x"58",
          4360 => x"38",
          4361 => x"97",
          4362 => x"08",
          4363 => x"38",
          4364 => x"70",
          4365 => x"81",
          4366 => x"55",
          4367 => x"87",
          4368 => x"39",
          4369 => x"90",
          4370 => x"82",
          4371 => x"8a",
          4372 => x"89",
          4373 => x"7f",
          4374 => x"56",
          4375 => x"3f",
          4376 => x"06",
          4377 => x"72",
          4378 => x"91",
          4379 => x"05",
          4380 => x"7c",
          4381 => x"55",
          4382 => x"27",
          4383 => x"16",
          4384 => x"83",
          4385 => x"76",
          4386 => x"80",
          4387 => x"79",
          4388 => x"99",
          4389 => x"7f",
          4390 => x"14",
          4391 => x"83",
          4392 => x"91",
          4393 => x"81",
          4394 => x"38",
          4395 => x"08",
          4396 => x"95",
          4397 => x"88",
          4398 => x"81",
          4399 => x"7b",
          4400 => x"06",
          4401 => x"39",
          4402 => x"56",
          4403 => x"09",
          4404 => x"b9",
          4405 => x"80",
          4406 => x"80",
          4407 => x"78",
          4408 => x"7a",
          4409 => x"38",
          4410 => x"73",
          4411 => x"81",
          4412 => x"ff",
          4413 => x"74",
          4414 => x"ff",
          4415 => x"91",
          4416 => x"58",
          4417 => x"08",
          4418 => x"74",
          4419 => x"16",
          4420 => x"73",
          4421 => x"39",
          4422 => x"7e",
          4423 => x"0c",
          4424 => x"2e",
          4425 => x"88",
          4426 => x"8c",
          4427 => x"1a",
          4428 => x"07",
          4429 => x"1b",
          4430 => x"08",
          4431 => x"16",
          4432 => x"75",
          4433 => x"38",
          4434 => x"90",
          4435 => x"15",
          4436 => x"54",
          4437 => x"34",
          4438 => x"91",
          4439 => x"90",
          4440 => x"e9",
          4441 => x"6d",
          4442 => x"80",
          4443 => x"9d",
          4444 => x"5c",
          4445 => x"3f",
          4446 => x"0b",
          4447 => x"08",
          4448 => x"38",
          4449 => x"08",
          4450 => x"ca",
          4451 => x"08",
          4452 => x"80",
          4453 => x"80",
          4454 => x"ca",
          4455 => x"ff",
          4456 => x"52",
          4457 => x"a0",
          4458 => x"ca",
          4459 => x"ff",
          4460 => x"06",
          4461 => x"56",
          4462 => x"38",
          4463 => x"70",
          4464 => x"55",
          4465 => x"8b",
          4466 => x"3d",
          4467 => x"83",
          4468 => x"ff",
          4469 => x"91",
          4470 => x"99",
          4471 => x"74",
          4472 => x"38",
          4473 => x"80",
          4474 => x"ff",
          4475 => x"55",
          4476 => x"83",
          4477 => x"78",
          4478 => x"38",
          4479 => x"26",
          4480 => x"81",
          4481 => x"8b",
          4482 => x"79",
          4483 => x"80",
          4484 => x"93",
          4485 => x"39",
          4486 => x"6e",
          4487 => x"89",
          4488 => x"48",
          4489 => x"83",
          4490 => x"61",
          4491 => x"25",
          4492 => x"55",
          4493 => x"8a",
          4494 => x"3d",
          4495 => x"81",
          4496 => x"ff",
          4497 => x"81",
          4498 => x"88",
          4499 => x"38",
          4500 => x"70",
          4501 => x"ca",
          4502 => x"56",
          4503 => x"38",
          4504 => x"55",
          4505 => x"75",
          4506 => x"38",
          4507 => x"70",
          4508 => x"ff",
          4509 => x"83",
          4510 => x"78",
          4511 => x"89",
          4512 => x"81",
          4513 => x"06",
          4514 => x"80",
          4515 => x"77",
          4516 => x"74",
          4517 => x"8d",
          4518 => x"06",
          4519 => x"2e",
          4520 => x"77",
          4521 => x"93",
          4522 => x"74",
          4523 => x"cb",
          4524 => x"7d",
          4525 => x"81",
          4526 => x"38",
          4527 => x"66",
          4528 => x"81",
          4529 => x"b8",
          4530 => x"74",
          4531 => x"38",
          4532 => x"98",
          4533 => x"b8",
          4534 => x"82",
          4535 => x"57",
          4536 => x"80",
          4537 => x"76",
          4538 => x"38",
          4539 => x"51",
          4540 => x"3f",
          4541 => x"08",
          4542 => x"87",
          4543 => x"2a",
          4544 => x"5c",
          4545 => x"ca",
          4546 => x"80",
          4547 => x"44",
          4548 => x"0a",
          4549 => x"ec",
          4550 => x"39",
          4551 => x"66",
          4552 => x"81",
          4553 => x"a8",
          4554 => x"74",
          4555 => x"38",
          4556 => x"98",
          4557 => x"a8",
          4558 => x"82",
          4559 => x"57",
          4560 => x"80",
          4561 => x"76",
          4562 => x"38",
          4563 => x"51",
          4564 => x"3f",
          4565 => x"08",
          4566 => x"57",
          4567 => x"08",
          4568 => x"96",
          4569 => x"91",
          4570 => x"10",
          4571 => x"08",
          4572 => x"72",
          4573 => x"59",
          4574 => x"ff",
          4575 => x"5d",
          4576 => x"44",
          4577 => x"11",
          4578 => x"70",
          4579 => x"71",
          4580 => x"06",
          4581 => x"52",
          4582 => x"40",
          4583 => x"09",
          4584 => x"38",
          4585 => x"18",
          4586 => x"39",
          4587 => x"79",
          4588 => x"70",
          4589 => x"58",
          4590 => x"76",
          4591 => x"38",
          4592 => x"7d",
          4593 => x"70",
          4594 => x"55",
          4595 => x"3f",
          4596 => x"08",
          4597 => x"2e",
          4598 => x"9b",
          4599 => x"88",
          4600 => x"f5",
          4601 => x"38",
          4602 => x"38",
          4603 => x"59",
          4604 => x"38",
          4605 => x"7d",
          4606 => x"81",
          4607 => x"38",
          4608 => x"0b",
          4609 => x"08",
          4610 => x"78",
          4611 => x"1a",
          4612 => x"c0",
          4613 => x"74",
          4614 => x"39",
          4615 => x"55",
          4616 => x"8f",
          4617 => x"fd",
          4618 => x"ca",
          4619 => x"f5",
          4620 => x"78",
          4621 => x"79",
          4622 => x"80",
          4623 => x"f1",
          4624 => x"39",
          4625 => x"81",
          4626 => x"06",
          4627 => x"55",
          4628 => x"27",
          4629 => x"81",
          4630 => x"56",
          4631 => x"38",
          4632 => x"80",
          4633 => x"ff",
          4634 => x"8b",
          4635 => x"d0",
          4636 => x"ff",
          4637 => x"84",
          4638 => x"1b",
          4639 => x"b3",
          4640 => x"1c",
          4641 => x"ff",
          4642 => x"8e",
          4643 => x"a1",
          4644 => x"0b",
          4645 => x"7d",
          4646 => x"30",
          4647 => x"84",
          4648 => x"51",
          4649 => x"51",
          4650 => x"3f",
          4651 => x"83",
          4652 => x"90",
          4653 => x"ff",
          4654 => x"93",
          4655 => x"a0",
          4656 => x"39",
          4657 => x"1b",
          4658 => x"85",
          4659 => x"95",
          4660 => x"52",
          4661 => x"ff",
          4662 => x"81",
          4663 => x"1b",
          4664 => x"cf",
          4665 => x"9c",
          4666 => x"a0",
          4667 => x"83",
          4668 => x"06",
          4669 => x"82",
          4670 => x"52",
          4671 => x"51",
          4672 => x"3f",
          4673 => x"1b",
          4674 => x"c5",
          4675 => x"ac",
          4676 => x"a0",
          4677 => x"52",
          4678 => x"ff",
          4679 => x"86",
          4680 => x"51",
          4681 => x"3f",
          4682 => x"80",
          4683 => x"a9",
          4684 => x"1c",
          4685 => x"91",
          4686 => x"80",
          4687 => x"ae",
          4688 => x"b2",
          4689 => x"1b",
          4690 => x"85",
          4691 => x"ff",
          4692 => x"96",
          4693 => x"9f",
          4694 => x"80",
          4695 => x"34",
          4696 => x"1c",
          4697 => x"91",
          4698 => x"ab",
          4699 => x"a0",
          4700 => x"d4",
          4701 => x"fe",
          4702 => x"59",
          4703 => x"3f",
          4704 => x"53",
          4705 => x"51",
          4706 => x"3f",
          4707 => x"ca",
          4708 => x"e7",
          4709 => x"2e",
          4710 => x"80",
          4711 => x"54",
          4712 => x"53",
          4713 => x"51",
          4714 => x"3f",
          4715 => x"80",
          4716 => x"ff",
          4717 => x"84",
          4718 => x"d2",
          4719 => x"ff",
          4720 => x"86",
          4721 => x"f2",
          4722 => x"1b",
          4723 => x"81",
          4724 => x"52",
          4725 => x"51",
          4726 => x"3f",
          4727 => x"ec",
          4728 => x"9e",
          4729 => x"d4",
          4730 => x"51",
          4731 => x"3f",
          4732 => x"87",
          4733 => x"52",
          4734 => x"9a",
          4735 => x"54",
          4736 => x"7a",
          4737 => x"ff",
          4738 => x"65",
          4739 => x"7a",
          4740 => x"8f",
          4741 => x"80",
          4742 => x"2e",
          4743 => x"9a",
          4744 => x"7a",
          4745 => x"a9",
          4746 => x"84",
          4747 => x"9e",
          4748 => x"0a",
          4749 => x"51",
          4750 => x"ff",
          4751 => x"7d",
          4752 => x"38",
          4753 => x"52",
          4754 => x"9e",
          4755 => x"55",
          4756 => x"62",
          4757 => x"74",
          4758 => x"75",
          4759 => x"7e",
          4760 => x"fe",
          4761 => x"88",
          4762 => x"38",
          4763 => x"91",
          4764 => x"52",
          4765 => x"9e",
          4766 => x"16",
          4767 => x"56",
          4768 => x"38",
          4769 => x"77",
          4770 => x"8d",
          4771 => x"7d",
          4772 => x"38",
          4773 => x"57",
          4774 => x"83",
          4775 => x"76",
          4776 => x"7a",
          4777 => x"ff",
          4778 => x"91",
          4779 => x"81",
          4780 => x"16",
          4781 => x"56",
          4782 => x"38",
          4783 => x"83",
          4784 => x"86",
          4785 => x"ff",
          4786 => x"38",
          4787 => x"82",
          4788 => x"81",
          4789 => x"06",
          4790 => x"fe",
          4791 => x"53",
          4792 => x"51",
          4793 => x"3f",
          4794 => x"52",
          4795 => x"9c",
          4796 => x"be",
          4797 => x"75",
          4798 => x"81",
          4799 => x"0b",
          4800 => x"77",
          4801 => x"75",
          4802 => x"60",
          4803 => x"80",
          4804 => x"75",
          4805 => x"d1",
          4806 => x"85",
          4807 => x"ca",
          4808 => x"2a",
          4809 => x"75",
          4810 => x"91",
          4811 => x"87",
          4812 => x"52",
          4813 => x"51",
          4814 => x"3f",
          4815 => x"ca",
          4816 => x"9c",
          4817 => x"54",
          4818 => x"52",
          4819 => x"98",
          4820 => x"56",
          4821 => x"08",
          4822 => x"53",
          4823 => x"51",
          4824 => x"3f",
          4825 => x"ca",
          4826 => x"38",
          4827 => x"56",
          4828 => x"56",
          4829 => x"ca",
          4830 => x"75",
          4831 => x"0c",
          4832 => x"04",
          4833 => x"73",
          4834 => x"26",
          4835 => x"71",
          4836 => x"b3",
          4837 => x"71",
          4838 => x"bb",
          4839 => x"80",
          4840 => x"e4",
          4841 => x"39",
          4842 => x"51",
          4843 => x"91",
          4844 => x"80",
          4845 => x"bc",
          4846 => x"e4",
          4847 => x"ac",
          4848 => x"39",
          4849 => x"51",
          4850 => x"91",
          4851 => x"80",
          4852 => x"bc",
          4853 => x"c8",
          4854 => x"80",
          4855 => x"39",
          4856 => x"51",
          4857 => x"bd",
          4858 => x"39",
          4859 => x"51",
          4860 => x"bd",
          4861 => x"39",
          4862 => x"51",
          4863 => x"be",
          4864 => x"39",
          4865 => x"51",
          4866 => x"be",
          4867 => x"39",
          4868 => x"51",
          4869 => x"bf",
          4870 => x"39",
          4871 => x"51",
          4872 => x"3f",
          4873 => x"04",
          4874 => x"77",
          4875 => x"74",
          4876 => x"8a",
          4877 => x"75",
          4878 => x"51",
          4879 => x"e8",
          4880 => x"fe",
          4881 => x"91",
          4882 => x"52",
          4883 => x"f2",
          4884 => x"ca",
          4885 => x"79",
          4886 => x"91",
          4887 => x"ff",
          4888 => x"87",
          4889 => x"f5",
          4890 => x"7f",
          4891 => x"05",
          4892 => x"33",
          4893 => x"66",
          4894 => x"5a",
          4895 => x"78",
          4896 => x"c4",
          4897 => x"fa",
          4898 => x"cc",
          4899 => x"8e",
          4900 => x"74",
          4901 => x"fc",
          4902 => x"2e",
          4903 => x"a0",
          4904 => x"80",
          4905 => x"16",
          4906 => x"27",
          4907 => x"22",
          4908 => x"d0",
          4909 => x"ca",
          4910 => x"91",
          4911 => x"ff",
          4912 => x"82",
          4913 => x"c3",
          4914 => x"53",
          4915 => x"8e",
          4916 => x"52",
          4917 => x"51",
          4918 => x"3f",
          4919 => x"bf",
          4920 => x"86",
          4921 => x"15",
          4922 => x"74",
          4923 => x"78",
          4924 => x"72",
          4925 => x"bf",
          4926 => x"8c",
          4927 => x"39",
          4928 => x"51",
          4929 => x"3f",
          4930 => x"a0",
          4931 => x"8d",
          4932 => x"39",
          4933 => x"51",
          4934 => x"3f",
          4935 => x"77",
          4936 => x"74",
          4937 => x"79",
          4938 => x"55",
          4939 => x"27",
          4940 => x"80",
          4941 => x"73",
          4942 => x"85",
          4943 => x"83",
          4944 => x"fe",
          4945 => x"81",
          4946 => x"39",
          4947 => x"51",
          4948 => x"3f",
          4949 => x"1a",
          4950 => x"fd",
          4951 => x"ca",
          4952 => x"2b",
          4953 => x"51",
          4954 => x"2e",
          4955 => x"a5",
          4956 => x"fb",
          4957 => x"88",
          4958 => x"70",
          4959 => x"a0",
          4960 => x"70",
          4961 => x"2a",
          4962 => x"51",
          4963 => x"2e",
          4964 => x"dd",
          4965 => x"2e",
          4966 => x"85",
          4967 => x"8c",
          4968 => x"53",
          4969 => x"fd",
          4970 => x"53",
          4971 => x"88",
          4972 => x"0d",
          4973 => x"0d",
          4974 => x"05",
          4975 => x"33",
          4976 => x"70",
          4977 => x"25",
          4978 => x"74",
          4979 => x"51",
          4980 => x"56",
          4981 => x"80",
          4982 => x"53",
          4983 => x"3d",
          4984 => x"c0",
          4985 => x"ca",
          4986 => x"91",
          4987 => x"b8",
          4988 => x"88",
          4989 => x"98",
          4990 => x"ca",
          4991 => x"96",
          4992 => x"54",
          4993 => x"77",
          4994 => x"c4",
          4995 => x"ca",
          4996 => x"91",
          4997 => x"90",
          4998 => x"74",
          4999 => x"38",
          5000 => x"19",
          5001 => x"39",
          5002 => x"05",
          5003 => x"3f",
          5004 => x"77",
          5005 => x"51",
          5006 => x"2e",
          5007 => x"80",
          5008 => x"91",
          5009 => x"87",
          5010 => x"08",
          5011 => x"fb",
          5012 => x"57",
          5013 => x"88",
          5014 => x"0d",
          5015 => x"0d",
          5016 => x"05",
          5017 => x"57",
          5018 => x"80",
          5019 => x"79",
          5020 => x"3f",
          5021 => x"08",
          5022 => x"80",
          5023 => x"75",
          5024 => x"38",
          5025 => x"55",
          5026 => x"ca",
          5027 => x"52",
          5028 => x"2d",
          5029 => x"08",
          5030 => x"77",
          5031 => x"ca",
          5032 => x"3d",
          5033 => x"3d",
          5034 => x"05",
          5035 => x"80",
          5036 => x"88",
          5037 => x"88",
          5038 => x"c7",
          5039 => x"ff",
          5040 => x"91",
          5041 => x"91",
          5042 => x"91",
          5043 => x"52",
          5044 => x"51",
          5045 => x"3f",
          5046 => x"85",
          5047 => x"92",
          5048 => x"0d",
          5049 => x"0d",
          5050 => x"80",
          5051 => x"80",
          5052 => x"51",
          5053 => x"3f",
          5054 => x"51",
          5055 => x"3f",
          5056 => x"f5",
          5057 => x"81",
          5058 => x"06",
          5059 => x"80",
          5060 => x"81",
          5061 => x"eb",
          5062 => x"e0",
          5063 => x"e3",
          5064 => x"fe",
          5065 => x"72",
          5066 => x"81",
          5067 => x"71",
          5068 => x"38",
          5069 => x"f5",
          5070 => x"c0",
          5071 => x"f7",
          5072 => x"51",
          5073 => x"3f",
          5074 => x"70",
          5075 => x"52",
          5076 => x"95",
          5077 => x"fe",
          5078 => x"91",
          5079 => x"fe",
          5080 => x"80",
          5081 => x"9b",
          5082 => x"2a",
          5083 => x"51",
          5084 => x"2e",
          5085 => x"51",
          5086 => x"3f",
          5087 => x"51",
          5088 => x"3f",
          5089 => x"f4",
          5090 => x"85",
          5091 => x"06",
          5092 => x"80",
          5093 => x"81",
          5094 => x"e7",
          5095 => x"ac",
          5096 => x"df",
          5097 => x"fe",
          5098 => x"72",
          5099 => x"81",
          5100 => x"71",
          5101 => x"38",
          5102 => x"f4",
          5103 => x"c1",
          5104 => x"f6",
          5105 => x"51",
          5106 => x"3f",
          5107 => x"70",
          5108 => x"52",
          5109 => x"95",
          5110 => x"fe",
          5111 => x"91",
          5112 => x"fe",
          5113 => x"80",
          5114 => x"97",
          5115 => x"2a",
          5116 => x"51",
          5117 => x"2e",
          5118 => x"51",
          5119 => x"3f",
          5120 => x"51",
          5121 => x"3f",
          5122 => x"f3",
          5123 => x"ff",
          5124 => x"3d",
          5125 => x"3d",
          5126 => x"08",
          5127 => x"57",
          5128 => x"80",
          5129 => x"39",
          5130 => x"85",
          5131 => x"80",
          5132 => x"14",
          5133 => x"33",
          5134 => x"06",
          5135 => x"74",
          5136 => x"38",
          5137 => x"80",
          5138 => x"72",
          5139 => x"81",
          5140 => x"72",
          5141 => x"81",
          5142 => x"80",
          5143 => x"05",
          5144 => x"56",
          5145 => x"91",
          5146 => x"77",
          5147 => x"08",
          5148 => x"ed",
          5149 => x"ca",
          5150 => x"38",
          5151 => x"53",
          5152 => x"ff",
          5153 => x"16",
          5154 => x"06",
          5155 => x"76",
          5156 => x"ff",
          5157 => x"ca",
          5158 => x"3d",
          5159 => x"3d",
          5160 => x"71",
          5161 => x"0c",
          5162 => x"52",
          5163 => x"8a",
          5164 => x"ca",
          5165 => x"ff",
          5166 => x"7c",
          5167 => x"06",
          5168 => x"c2",
          5169 => x"3d",
          5170 => x"ff",
          5171 => x"7b",
          5172 => x"91",
          5173 => x"ff",
          5174 => x"91",
          5175 => x"7c",
          5176 => x"91",
          5177 => x"90",
          5178 => x"70",
          5179 => x"c2",
          5180 => x"fe",
          5181 => x"3d",
          5182 => x"80",
          5183 => x"52",
          5184 => x"eb",
          5185 => x"f8",
          5186 => x"ff",
          5187 => x"b7",
          5188 => x"05",
          5189 => x"3f",
          5190 => x"08",
          5191 => x"90",
          5192 => x"78",
          5193 => x"8a",
          5194 => x"80",
          5195 => x"e0",
          5196 => x"2e",
          5197 => x"78",
          5198 => x"38",
          5199 => x"82",
          5200 => x"84",
          5201 => x"78",
          5202 => x"a2",
          5203 => x"2e",
          5204 => x"8e",
          5205 => x"94",
          5206 => x"38",
          5207 => x"83",
          5208 => x"e2",
          5209 => x"2e",
          5210 => x"78",
          5211 => x"38",
          5212 => x"84",
          5213 => x"bd",
          5214 => x"38",
          5215 => x"78",
          5216 => x"86",
          5217 => x"80",
          5218 => x"cf",
          5219 => x"39",
          5220 => x"2e",
          5221 => x"78",
          5222 => x"b0",
          5223 => x"d1",
          5224 => x"38",
          5225 => x"24",
          5226 => x"80",
          5227 => x"83",
          5228 => x"d0",
          5229 => x"38",
          5230 => x"78",
          5231 => x"8c",
          5232 => x"80",
          5233 => x"d6",
          5234 => x"39",
          5235 => x"2e",
          5236 => x"78",
          5237 => x"92",
          5238 => x"f9",
          5239 => x"38",
          5240 => x"2e",
          5241 => x"8d",
          5242 => x"81",
          5243 => x"cf",
          5244 => x"87",
          5245 => x"38",
          5246 => x"b7",
          5247 => x"11",
          5248 => x"05",
          5249 => x"ef",
          5250 => x"88",
          5251 => x"91",
          5252 => x"8e",
          5253 => x"3d",
          5254 => x"53",
          5255 => x"51",
          5256 => x"3f",
          5257 => x"08",
          5258 => x"38",
          5259 => x"83",
          5260 => x"02",
          5261 => x"33",
          5262 => x"cf",
          5263 => x"ff",
          5264 => x"91",
          5265 => x"81",
          5266 => x"78",
          5267 => x"c2",
          5268 => x"fb",
          5269 => x"5d",
          5270 => x"91",
          5271 => x"8b",
          5272 => x"3d",
          5273 => x"53",
          5274 => x"51",
          5275 => x"3f",
          5276 => x"08",
          5277 => x"f6",
          5278 => x"80",
          5279 => x"cf",
          5280 => x"ff",
          5281 => x"91",
          5282 => x"52",
          5283 => x"51",
          5284 => x"b7",
          5285 => x"11",
          5286 => x"05",
          5287 => x"d7",
          5288 => x"88",
          5289 => x"87",
          5290 => x"26",
          5291 => x"b7",
          5292 => x"11",
          5293 => x"05",
          5294 => x"bb",
          5295 => x"88",
          5296 => x"91",
          5297 => x"43",
          5298 => x"c3",
          5299 => x"51",
          5300 => x"3f",
          5301 => x"05",
          5302 => x"52",
          5303 => x"29",
          5304 => x"05",
          5305 => x"d5",
          5306 => x"88",
          5307 => x"38",
          5308 => x"51",
          5309 => x"3f",
          5310 => x"f2",
          5311 => x"fe",
          5312 => x"fe",
          5313 => x"91",
          5314 => x"b8",
          5315 => x"05",
          5316 => x"eb",
          5317 => x"53",
          5318 => x"08",
          5319 => x"f5",
          5320 => x"d5",
          5321 => x"fe",
          5322 => x"fe",
          5323 => x"91",
          5324 => x"b8",
          5325 => x"05",
          5326 => x"ea",
          5327 => x"ca",
          5328 => x"3d",
          5329 => x"52",
          5330 => x"ca",
          5331 => x"88",
          5332 => x"fe",
          5333 => x"59",
          5334 => x"3f",
          5335 => x"58",
          5336 => x"57",
          5337 => x"55",
          5338 => x"08",
          5339 => x"54",
          5340 => x"52",
          5341 => x"e5",
          5342 => x"88",
          5343 => x"fa",
          5344 => x"ca",
          5345 => x"ef",
          5346 => x"e2",
          5347 => x"fe",
          5348 => x"fe",
          5349 => x"ff",
          5350 => x"91",
          5351 => x"80",
          5352 => x"38",
          5353 => x"f0",
          5354 => x"f8",
          5355 => x"80",
          5356 => x"ca",
          5357 => x"2e",
          5358 => x"b7",
          5359 => x"11",
          5360 => x"05",
          5361 => x"af",
          5362 => x"88",
          5363 => x"91",
          5364 => x"42",
          5365 => x"51",
          5366 => x"3f",
          5367 => x"5a",
          5368 => x"81",
          5369 => x"59",
          5370 => x"84",
          5371 => x"7a",
          5372 => x"38",
          5373 => x"b7",
          5374 => x"11",
          5375 => x"05",
          5376 => x"f3",
          5377 => x"88",
          5378 => x"f9",
          5379 => x"3d",
          5380 => x"53",
          5381 => x"51",
          5382 => x"3f",
          5383 => x"08",
          5384 => x"ca",
          5385 => x"fe",
          5386 => x"fe",
          5387 => x"fe",
          5388 => x"91",
          5389 => x"80",
          5390 => x"38",
          5391 => x"51",
          5392 => x"3f",
          5393 => x"63",
          5394 => x"38",
          5395 => x"70",
          5396 => x"33",
          5397 => x"81",
          5398 => x"39",
          5399 => x"f4",
          5400 => x"f8",
          5401 => x"ff",
          5402 => x"ca",
          5403 => x"2e",
          5404 => x"b7",
          5405 => x"11",
          5406 => x"05",
          5407 => x"f7",
          5408 => x"88",
          5409 => x"f8",
          5410 => x"3d",
          5411 => x"53",
          5412 => x"51",
          5413 => x"3f",
          5414 => x"08",
          5415 => x"ce",
          5416 => x"c4",
          5417 => x"f6",
          5418 => x"79",
          5419 => x"38",
          5420 => x"7b",
          5421 => x"5b",
          5422 => x"92",
          5423 => x"7a",
          5424 => x"53",
          5425 => x"c3",
          5426 => x"fc",
          5427 => x"1a",
          5428 => x"43",
          5429 => x"91",
          5430 => x"86",
          5431 => x"3d",
          5432 => x"53",
          5433 => x"51",
          5434 => x"3f",
          5435 => x"08",
          5436 => x"91",
          5437 => x"59",
          5438 => x"88",
          5439 => x"e4",
          5440 => x"39",
          5441 => x"33",
          5442 => x"2e",
          5443 => x"c6",
          5444 => x"a2",
          5445 => x"93",
          5446 => x"8b",
          5447 => x"94",
          5448 => x"80",
          5449 => x"91",
          5450 => x"44",
          5451 => x"c7",
          5452 => x"80",
          5453 => x"3d",
          5454 => x"53",
          5455 => x"51",
          5456 => x"3f",
          5457 => x"08",
          5458 => x"91",
          5459 => x"59",
          5460 => x"88",
          5461 => x"e8",
          5462 => x"39",
          5463 => x"33",
          5464 => x"2e",
          5465 => x"c6",
          5466 => x"a1",
          5467 => x"93",
          5468 => x"8b",
          5469 => x"94",
          5470 => x"80",
          5471 => x"91",
          5472 => x"43",
          5473 => x"c7",
          5474 => x"05",
          5475 => x"fe",
          5476 => x"fe",
          5477 => x"fe",
          5478 => x"91",
          5479 => x"80",
          5480 => x"80",
          5481 => x"79",
          5482 => x"38",
          5483 => x"90",
          5484 => x"78",
          5485 => x"38",
          5486 => x"83",
          5487 => x"91",
          5488 => x"fe",
          5489 => x"a0",
          5490 => x"61",
          5491 => x"63",
          5492 => x"3f",
          5493 => x"51",
          5494 => x"b7",
          5495 => x"11",
          5496 => x"05",
          5497 => x"8f",
          5498 => x"88",
          5499 => x"f5",
          5500 => x"3d",
          5501 => x"53",
          5502 => x"51",
          5503 => x"3f",
          5504 => x"08",
          5505 => x"38",
          5506 => x"80",
          5507 => x"79",
          5508 => x"05",
          5509 => x"fe",
          5510 => x"fe",
          5511 => x"fe",
          5512 => x"91",
          5513 => x"e0",
          5514 => x"39",
          5515 => x"54",
          5516 => x"8c",
          5517 => x"ca",
          5518 => x"52",
          5519 => x"fa",
          5520 => x"45",
          5521 => x"78",
          5522 => x"a2",
          5523 => x"27",
          5524 => x"3d",
          5525 => x"53",
          5526 => x"51",
          5527 => x"3f",
          5528 => x"08",
          5529 => x"38",
          5530 => x"80",
          5531 => x"79",
          5532 => x"05",
          5533 => x"39",
          5534 => x"51",
          5535 => x"3f",
          5536 => x"b7",
          5537 => x"11",
          5538 => x"05",
          5539 => x"d9",
          5540 => x"88",
          5541 => x"f4",
          5542 => x"3d",
          5543 => x"53",
          5544 => x"51",
          5545 => x"3f",
          5546 => x"08",
          5547 => x"38",
          5548 => x"be",
          5549 => x"70",
          5550 => x"23",
          5551 => x"3d",
          5552 => x"53",
          5553 => x"51",
          5554 => x"3f",
          5555 => x"08",
          5556 => x"9a",
          5557 => x"22",
          5558 => x"c4",
          5559 => x"f8",
          5560 => x"f8",
          5561 => x"fe",
          5562 => x"79",
          5563 => x"59",
          5564 => x"f3",
          5565 => x"9f",
          5566 => x"60",
          5567 => x"d5",
          5568 => x"fe",
          5569 => x"fe",
          5570 => x"fe",
          5571 => x"91",
          5572 => x"80",
          5573 => x"60",
          5574 => x"05",
          5575 => x"82",
          5576 => x"78",
          5577 => x"39",
          5578 => x"51",
          5579 => x"3f",
          5580 => x"b7",
          5581 => x"11",
          5582 => x"05",
          5583 => x"a9",
          5584 => x"88",
          5585 => x"f3",
          5586 => x"3d",
          5587 => x"53",
          5588 => x"51",
          5589 => x"3f",
          5590 => x"08",
          5591 => x"38",
          5592 => x"0c",
          5593 => x"05",
          5594 => x"fe",
          5595 => x"fe",
          5596 => x"fe",
          5597 => x"91",
          5598 => x"e4",
          5599 => x"39",
          5600 => x"54",
          5601 => x"ac",
          5602 => x"f6",
          5603 => x"52",
          5604 => x"f7",
          5605 => x"45",
          5606 => x"78",
          5607 => x"ce",
          5608 => x"27",
          5609 => x"3d",
          5610 => x"53",
          5611 => x"51",
          5612 => x"3f",
          5613 => x"08",
          5614 => x"38",
          5615 => x"52",
          5616 => x"51",
          5617 => x"3f",
          5618 => x"0c",
          5619 => x"05",
          5620 => x"39",
          5621 => x"51",
          5622 => x"3f",
          5623 => x"91",
          5624 => x"fe",
          5625 => x"82",
          5626 => x"a6",
          5627 => x"39",
          5628 => x"51",
          5629 => x"3f",
          5630 => x"ee",
          5631 => x"ee",
          5632 => x"81",
          5633 => x"94",
          5634 => x"80",
          5635 => x"c0",
          5636 => x"91",
          5637 => x"fe",
          5638 => x"f1",
          5639 => x"c4",
          5640 => x"ef",
          5641 => x"80",
          5642 => x"c0",
          5643 => x"8c",
          5644 => x"87",
          5645 => x"0c",
          5646 => x"b7",
          5647 => x"11",
          5648 => x"05",
          5649 => x"af",
          5650 => x"88",
          5651 => x"f1",
          5652 => x"52",
          5653 => x"51",
          5654 => x"3f",
          5655 => x"04",
          5656 => x"f4",
          5657 => x"f8",
          5658 => x"f7",
          5659 => x"ca",
          5660 => x"2e",
          5661 => x"63",
          5662 => x"ac",
          5663 => x"82",
          5664 => x"78",
          5665 => x"88",
          5666 => x"ca",
          5667 => x"2e",
          5668 => x"91",
          5669 => x"52",
          5670 => x"51",
          5671 => x"3f",
          5672 => x"91",
          5673 => x"fe",
          5674 => x"fe",
          5675 => x"f0",
          5676 => x"c6",
          5677 => x"ee",
          5678 => x"59",
          5679 => x"fe",
          5680 => x"f0",
          5681 => x"70",
          5682 => x"78",
          5683 => x"9e",
          5684 => x"2e",
          5685 => x"7c",
          5686 => x"cc",
          5687 => x"fe",
          5688 => x"fe",
          5689 => x"91",
          5690 => x"91",
          5691 => x"55",
          5692 => x"54",
          5693 => x"c6",
          5694 => x"3d",
          5695 => x"fe",
          5696 => x"91",
          5697 => x"91",
          5698 => x"80",
          5699 => x"11",
          5700 => x"55",
          5701 => x"80",
          5702 => x"80",
          5703 => x"51",
          5704 => x"91",
          5705 => x"5e",
          5706 => x"7c",
          5707 => x"59",
          5708 => x"7d",
          5709 => x"81",
          5710 => x"38",
          5711 => x"51",
          5712 => x"3f",
          5713 => x"80",
          5714 => x"0b",
          5715 => x"34",
          5716 => x"0b",
          5717 => x"0c",
          5718 => x"0b",
          5719 => x"0c",
          5720 => x"3f",
          5721 => x"3f",
          5722 => x"51",
          5723 => x"3f",
          5724 => x"51",
          5725 => x"3f",
          5726 => x"51",
          5727 => x"3f",
          5728 => x"a2",
          5729 => x"3f",
          5730 => x"04",
          5731 => x"04",
          5732 => x"04",
          5733 => x"04",
          5734 => x"04",
          5735 => x"04",
          5736 => x"04",
          5737 => x"04",
          5738 => x"04",
          5739 => x"04",
          5740 => x"04",
          5741 => x"04",
          5742 => x"04",
          5743 => x"04",
          5744 => x"04",
          5745 => x"04",
          5746 => x"04",
          5747 => x"04",
          5748 => x"04",
          5749 => x"04",
          5750 => x"04",
          5751 => x"04",
          5752 => x"04",
          5753 => x"04",
          5754 => x"04",
          5755 => x"64",
          5756 => x"2f",
          5757 => x"25",
          5758 => x"64",
          5759 => x"2e",
          5760 => x"64",
          5761 => x"6f",
          5762 => x"6f",
          5763 => x"67",
          5764 => x"74",
          5765 => x"00",
          5766 => x"28",
          5767 => x"6d",
          5768 => x"43",
          5769 => x"6e",
          5770 => x"29",
          5771 => x"0a",
          5772 => x"69",
          5773 => x"20",
          5774 => x"6c",
          5775 => x"6e",
          5776 => x"3a",
          5777 => x"20",
          5778 => x"4e",
          5779 => x"42",
          5780 => x"20",
          5781 => x"61",
          5782 => x"25",
          5783 => x"2c",
          5784 => x"7a",
          5785 => x"30",
          5786 => x"2e",
          5787 => x"20",
          5788 => x"52",
          5789 => x"28",
          5790 => x"72",
          5791 => x"30",
          5792 => x"20",
          5793 => x"65",
          5794 => x"38",
          5795 => x"0a",
          5796 => x"20",
          5797 => x"41",
          5798 => x"53",
          5799 => x"74",
          5800 => x"38",
          5801 => x"53",
          5802 => x"3d",
          5803 => x"58",
          5804 => x"00",
          5805 => x"20",
          5806 => x"4f",
          5807 => x"0a",
          5808 => x"20",
          5809 => x"53",
          5810 => x"00",
          5811 => x"20",
          5812 => x"50",
          5813 => x"00",
          5814 => x"20",
          5815 => x"44",
          5816 => x"72",
          5817 => x"44",
          5818 => x"63",
          5819 => x"25",
          5820 => x"29",
          5821 => x"00",
          5822 => x"20",
          5823 => x"4e",
          5824 => x"52",
          5825 => x"20",
          5826 => x"54",
          5827 => x"4c",
          5828 => x"00",
          5829 => x"20",
          5830 => x"49",
          5831 => x"31",
          5832 => x"69",
          5833 => x"73",
          5834 => x"31",
          5835 => x"0a",
          5836 => x"64",
          5837 => x"73",
          5838 => x"3a",
          5839 => x"20",
          5840 => x"50",
          5841 => x"65",
          5842 => x"20",
          5843 => x"74",
          5844 => x"41",
          5845 => x"65",
          5846 => x"3d",
          5847 => x"38",
          5848 => x"00",
          5849 => x"20",
          5850 => x"50",
          5851 => x"65",
          5852 => x"79",
          5853 => x"61",
          5854 => x"41",
          5855 => x"65",
          5856 => x"3d",
          5857 => x"38",
          5858 => x"00",
          5859 => x"20",
          5860 => x"74",
          5861 => x"20",
          5862 => x"72",
          5863 => x"64",
          5864 => x"73",
          5865 => x"20",
          5866 => x"3d",
          5867 => x"38",
          5868 => x"00",
          5869 => x"20",
          5870 => x"50",
          5871 => x"64",
          5872 => x"20",
          5873 => x"20",
          5874 => x"20",
          5875 => x"20",
          5876 => x"3d",
          5877 => x"38",
          5878 => x"00",
          5879 => x"20",
          5880 => x"79",
          5881 => x"6d",
          5882 => x"6f",
          5883 => x"46",
          5884 => x"20",
          5885 => x"20",
          5886 => x"3d",
          5887 => x"38",
          5888 => x"00",
          5889 => x"6d",
          5890 => x"00",
          5891 => x"65",
          5892 => x"6d",
          5893 => x"6c",
          5894 => x"00",
          5895 => x"56",
          5896 => x"56",
          5897 => x"6e",
          5898 => x"6e",
          5899 => x"77",
          5900 => x"44",
          5901 => x"2a",
          5902 => x"3b",
          5903 => x"3f",
          5904 => x"7f",
          5905 => x"41",
          5906 => x"41",
          5907 => x"00",
          5908 => x"fe",
          5909 => x"44",
          5910 => x"2e",
          5911 => x"4f",
          5912 => x"4d",
          5913 => x"20",
          5914 => x"54",
          5915 => x"20",
          5916 => x"4f",
          5917 => x"4d",
          5918 => x"20",
          5919 => x"54",
          5920 => x"20",
          5921 => x"04",
          5922 => x"00",
          5923 => x"00",
          5924 => x"00",
          5925 => x"9a",
          5926 => x"41",
          5927 => x"45",
          5928 => x"49",
          5929 => x"92",
          5930 => x"4f",
          5931 => x"99",
          5932 => x"9d",
          5933 => x"49",
          5934 => x"a5",
          5935 => x"a9",
          5936 => x"ad",
          5937 => x"b1",
          5938 => x"b5",
          5939 => x"b9",
          5940 => x"bd",
          5941 => x"c1",
          5942 => x"c5",
          5943 => x"c9",
          5944 => x"cd",
          5945 => x"d1",
          5946 => x"d5",
          5947 => x"d9",
          5948 => x"dd",
          5949 => x"e1",
          5950 => x"e5",
          5951 => x"e9",
          5952 => x"ed",
          5953 => x"f1",
          5954 => x"f5",
          5955 => x"f9",
          5956 => x"fd",
          5957 => x"2e",
          5958 => x"5b",
          5959 => x"22",
          5960 => x"3e",
          5961 => x"00",
          5962 => x"01",
          5963 => x"10",
          5964 => x"00",
          5965 => x"00",
          5966 => x"01",
          5967 => x"04",
          5968 => x"10",
          5969 => x"00",
          5970 => x"69",
          5971 => x"00",
          5972 => x"69",
          5973 => x"6c",
          5974 => x"69",
          5975 => x"00",
          5976 => x"6c",
          5977 => x"00",
          5978 => x"65",
          5979 => x"00",
          5980 => x"63",
          5981 => x"72",
          5982 => x"63",
          5983 => x"00",
          5984 => x"64",
          5985 => x"00",
          5986 => x"64",
          5987 => x"00",
          5988 => x"65",
          5989 => x"65",
          5990 => x"65",
          5991 => x"69",
          5992 => x"69",
          5993 => x"66",
          5994 => x"66",
          5995 => x"61",
          5996 => x"00",
          5997 => x"6d",
          5998 => x"65",
          5999 => x"72",
          6000 => x"65",
          6001 => x"00",
          6002 => x"6e",
          6003 => x"00",
          6004 => x"65",
          6005 => x"00",
          6006 => x"69",
          6007 => x"45",
          6008 => x"72",
          6009 => x"6e",
          6010 => x"6e",
          6011 => x"65",
          6012 => x"72",
          6013 => x"00",
          6014 => x"69",
          6015 => x"6e",
          6016 => x"72",
          6017 => x"79",
          6018 => x"00",
          6019 => x"6f",
          6020 => x"6c",
          6021 => x"6f",
          6022 => x"2e",
          6023 => x"6f",
          6024 => x"74",
          6025 => x"6f",
          6026 => x"2e",
          6027 => x"6e",
          6028 => x"69",
          6029 => x"69",
          6030 => x"61",
          6031 => x"0a",
          6032 => x"63",
          6033 => x"73",
          6034 => x"6e",
          6035 => x"2e",
          6036 => x"69",
          6037 => x"61",
          6038 => x"61",
          6039 => x"65",
          6040 => x"74",
          6041 => x"00",
          6042 => x"69",
          6043 => x"68",
          6044 => x"6c",
          6045 => x"6e",
          6046 => x"69",
          6047 => x"00",
          6048 => x"44",
          6049 => x"20",
          6050 => x"74",
          6051 => x"72",
          6052 => x"63",
          6053 => x"2e",
          6054 => x"72",
          6055 => x"20",
          6056 => x"62",
          6057 => x"69",
          6058 => x"6e",
          6059 => x"69",
          6060 => x"00",
          6061 => x"69",
          6062 => x"6e",
          6063 => x"65",
          6064 => x"6c",
          6065 => x"0a",
          6066 => x"6f",
          6067 => x"6d",
          6068 => x"69",
          6069 => x"20",
          6070 => x"65",
          6071 => x"74",
          6072 => x"66",
          6073 => x"64",
          6074 => x"20",
          6075 => x"6b",
          6076 => x"00",
          6077 => x"6f",
          6078 => x"74",
          6079 => x"6f",
          6080 => x"64",
          6081 => x"00",
          6082 => x"69",
          6083 => x"75",
          6084 => x"6f",
          6085 => x"61",
          6086 => x"6e",
          6087 => x"6e",
          6088 => x"6c",
          6089 => x"0a",
          6090 => x"69",
          6091 => x"69",
          6092 => x"6f",
          6093 => x"64",
          6094 => x"00",
          6095 => x"6e",
          6096 => x"66",
          6097 => x"65",
          6098 => x"6d",
          6099 => x"72",
          6100 => x"00",
          6101 => x"6f",
          6102 => x"61",
          6103 => x"6f",
          6104 => x"20",
          6105 => x"65",
          6106 => x"00",
          6107 => x"61",
          6108 => x"65",
          6109 => x"73",
          6110 => x"63",
          6111 => x"65",
          6112 => x"0a",
          6113 => x"75",
          6114 => x"73",
          6115 => x"00",
          6116 => x"6e",
          6117 => x"77",
          6118 => x"72",
          6119 => x"2e",
          6120 => x"25",
          6121 => x"62",
          6122 => x"73",
          6123 => x"20",
          6124 => x"25",
          6125 => x"62",
          6126 => x"73",
          6127 => x"63",
          6128 => x"00",
          6129 => x"30",
          6130 => x"00",
          6131 => x"20",
          6132 => x"30",
          6133 => x"00",
          6134 => x"20",
          6135 => x"20",
          6136 => x"00",
          6137 => x"30",
          6138 => x"00",
          6139 => x"20",
          6140 => x"7c",
          6141 => x"0d",
          6142 => x"65",
          6143 => x"00",
          6144 => x"50",
          6145 => x"00",
          6146 => x"2a",
          6147 => x"73",
          6148 => x"00",
          6149 => x"38",
          6150 => x"2f",
          6151 => x"39",
          6152 => x"31",
          6153 => x"00",
          6154 => x"5a",
          6155 => x"20",
          6156 => x"20",
          6157 => x"78",
          6158 => x"73",
          6159 => x"20",
          6160 => x"0a",
          6161 => x"50",
          6162 => x"20",
          6163 => x"65",
          6164 => x"70",
          6165 => x"61",
          6166 => x"65",
          6167 => x"00",
          6168 => x"69",
          6169 => x"20",
          6170 => x"65",
          6171 => x"70",
          6172 => x"00",
          6173 => x"53",
          6174 => x"6e",
          6175 => x"72",
          6176 => x"0a",
          6177 => x"4f",
          6178 => x"20",
          6179 => x"69",
          6180 => x"72",
          6181 => x"74",
          6182 => x"4f",
          6183 => x"20",
          6184 => x"69",
          6185 => x"72",
          6186 => x"74",
          6187 => x"41",
          6188 => x"20",
          6189 => x"69",
          6190 => x"72",
          6191 => x"74",
          6192 => x"41",
          6193 => x"20",
          6194 => x"69",
          6195 => x"72",
          6196 => x"74",
          6197 => x"41",
          6198 => x"20",
          6199 => x"69",
          6200 => x"72",
          6201 => x"74",
          6202 => x"41",
          6203 => x"20",
          6204 => x"69",
          6205 => x"72",
          6206 => x"74",
          6207 => x"65",
          6208 => x"6e",
          6209 => x"70",
          6210 => x"6d",
          6211 => x"2e",
          6212 => x"00",
          6213 => x"6e",
          6214 => x"69",
          6215 => x"74",
          6216 => x"72",
          6217 => x"0a",
          6218 => x"3a",
          6219 => x"61",
          6220 => x"64",
          6221 => x"20",
          6222 => x"74",
          6223 => x"69",
          6224 => x"73",
          6225 => x"61",
          6226 => x"30",
          6227 => x"6c",
          6228 => x"65",
          6229 => x"69",
          6230 => x"61",
          6231 => x"6c",
          6232 => x"0a",
          6233 => x"20",
          6234 => x"61",
          6235 => x"69",
          6236 => x"69",
          6237 => x"00",
          6238 => x"6e",
          6239 => x"61",
          6240 => x"65",
          6241 => x"00",
          6242 => x"61",
          6243 => x"64",
          6244 => x"20",
          6245 => x"74",
          6246 => x"69",
          6247 => x"0a",
          6248 => x"63",
          6249 => x"0a",
          6250 => x"75",
          6251 => x"6c",
          6252 => x"69",
          6253 => x"2e",
          6254 => x"6f",
          6255 => x"6e",
          6256 => x"2e",
          6257 => x"6f",
          6258 => x"72",
          6259 => x"2e",
          6260 => x"00",
          6261 => x"30",
          6262 => x"28",
          6263 => x"78",
          6264 => x"25",
          6265 => x"78",
          6266 => x"38",
          6267 => x"00",
          6268 => x"75",
          6269 => x"4d",
          6270 => x"72",
          6271 => x"00",
          6272 => x"43",
          6273 => x"6c",
          6274 => x"2e",
          6275 => x"30",
          6276 => x"25",
          6277 => x"2d",
          6278 => x"3f",
          6279 => x"00",
          6280 => x"30",
          6281 => x"25",
          6282 => x"2d",
          6283 => x"30",
          6284 => x"25",
          6285 => x"2d",
          6286 => x"69",
          6287 => x"6c",
          6288 => x"20",
          6289 => x"65",
          6290 => x"70",
          6291 => x"00",
          6292 => x"6e",
          6293 => x"69",
          6294 => x"69",
          6295 => x"72",
          6296 => x"74",
          6297 => x"00",
          6298 => x"69",
          6299 => x"6c",
          6300 => x"75",
          6301 => x"20",
          6302 => x"6f",
          6303 => x"6e",
          6304 => x"69",
          6305 => x"75",
          6306 => x"20",
          6307 => x"6f",
          6308 => x"78",
          6309 => x"74",
          6310 => x"20",
          6311 => x"65",
          6312 => x"25",
          6313 => x"20",
          6314 => x"0a",
          6315 => x"61",
          6316 => x"6e",
          6317 => x"6f",
          6318 => x"40",
          6319 => x"38",
          6320 => x"2e",
          6321 => x"00",
          6322 => x"61",
          6323 => x"72",
          6324 => x"72",
          6325 => x"20",
          6326 => x"65",
          6327 => x"64",
          6328 => x"00",
          6329 => x"65",
          6330 => x"72",
          6331 => x"67",
          6332 => x"70",
          6333 => x"61",
          6334 => x"6e",
          6335 => x"0a",
          6336 => x"6f",
          6337 => x"72",
          6338 => x"6f",
          6339 => x"67",
          6340 => x"0a",
          6341 => x"50",
          6342 => x"69",
          6343 => x"64",
          6344 => x"73",
          6345 => x"2e",
          6346 => x"00",
          6347 => x"61",
          6348 => x"6f",
          6349 => x"6e",
          6350 => x"00",
          6351 => x"75",
          6352 => x"6e",
          6353 => x"2e",
          6354 => x"6e",
          6355 => x"69",
          6356 => x"69",
          6357 => x"72",
          6358 => x"74",
          6359 => x"2e",
          6360 => x"00",
          6361 => x"00",
          6362 => x"00",
          6363 => x"00",
          6364 => x"00",
          6365 => x"01",
          6366 => x"00",
          6367 => x"00",
          6368 => x"00",
          6369 => x"00",
          6370 => x"00",
          6371 => x"f5",
          6372 => x"01",
          6373 => x"01",
          6374 => x"01",
          6375 => x"00",
          6376 => x"00",
          6377 => x"00",
          6378 => x"04",
          6379 => x"02",
          6380 => x"00",
          6381 => x"00",
          6382 => x"04",
          6383 => x"04",
          6384 => x"00",
          6385 => x"00",
          6386 => x"04",
          6387 => x"14",
          6388 => x"00",
          6389 => x"00",
          6390 => x"04",
          6391 => x"2b",
          6392 => x"00",
          6393 => x"00",
          6394 => x"04",
          6395 => x"30",
          6396 => x"00",
          6397 => x"00",
          6398 => x"04",
          6399 => x"3c",
          6400 => x"00",
          6401 => x"00",
          6402 => x"04",
          6403 => x"3d",
          6404 => x"00",
          6405 => x"00",
          6406 => x"04",
          6407 => x"3f",
          6408 => x"00",
          6409 => x"00",
          6410 => x"04",
          6411 => x"40",
          6412 => x"00",
          6413 => x"00",
          6414 => x"04",
          6415 => x"41",
          6416 => x"00",
          6417 => x"00",
          6418 => x"04",
          6419 => x"42",
          6420 => x"00",
          6421 => x"00",
          6422 => x"04",
          6423 => x"43",
          6424 => x"00",
          6425 => x"00",
          6426 => x"04",
          6427 => x"50",
          6428 => x"00",
          6429 => x"00",
          6430 => x"04",
          6431 => x"51",
          6432 => x"00",
          6433 => x"00",
          6434 => x"04",
          6435 => x"54",
          6436 => x"00",
          6437 => x"00",
          6438 => x"04",
          6439 => x"55",
          6440 => x"00",
          6441 => x"00",
          6442 => x"04",
          6443 => x"79",
          6444 => x"00",
          6445 => x"00",
          6446 => x"04",
          6447 => x"78",
          6448 => x"00",
          6449 => x"00",
          6450 => x"04",
          6451 => x"82",
          6452 => x"00",
          6453 => x"00",
          6454 => x"04",
          6455 => x"83",
          6456 => x"00",
          6457 => x"00",
          6458 => x"04",
          6459 => x"85",
          6460 => x"00",
          6461 => x"00",
          6462 => x"04",
          6463 => x"87",
          6464 => x"00",
          6465 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"90",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"90",
            11 => x"0b",
            12 => x"96",
            13 => x"90",
            14 => x"0b",
            15 => x"b8",
            16 => x"90",
            17 => x"0b",
            18 => x"da",
            19 => x"90",
            20 => x"0b",
            21 => x"fc",
            22 => x"90",
            23 => x"0b",
            24 => x"9e",
            25 => x"90",
            26 => x"0b",
            27 => x"c0",
            28 => x"90",
            29 => x"0b",
            30 => x"e2",
            31 => x"90",
            32 => x"0b",
            33 => x"84",
            34 => x"90",
            35 => x"0b",
            36 => x"a6",
            37 => x"90",
            38 => x"0b",
            39 => x"c8",
            40 => x"90",
            41 => x"0b",
            42 => x"ea",
            43 => x"90",
            44 => x"0b",
            45 => x"8c",
            46 => x"90",
            47 => x"0b",
            48 => x"ae",
            49 => x"90",
            50 => x"0b",
            51 => x"d0",
            52 => x"90",
            53 => x"0b",
            54 => x"f2",
            55 => x"90",
            56 => x"0b",
            57 => x"94",
            58 => x"90",
            59 => x"0b",
            60 => x"b6",
            61 => x"90",
            62 => x"0b",
            63 => x"d8",
            64 => x"90",
            65 => x"0b",
            66 => x"fa",
            67 => x"90",
            68 => x"0b",
            69 => x"9c",
            70 => x"90",
            71 => x"0b",
            72 => x"be",
            73 => x"90",
            74 => x"0b",
            75 => x"e0",
            76 => x"90",
            77 => x"0b",
            78 => x"82",
            79 => x"90",
            80 => x"0b",
            81 => x"a4",
            82 => x"90",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"04",
           130 => x"0c",
           131 => x"2d",
           132 => x"08",
           133 => x"90",
           134 => x"94",
           135 => x"bf",
           136 => x"94",
           137 => x"80",
           138 => x"ca",
           139 => x"9f",
           140 => x"ca",
           141 => x"c0",
           142 => x"91",
           143 => x"90",
           144 => x"91",
           145 => x"88",
           146 => x"04",
           147 => x"0c",
           148 => x"2d",
           149 => x"08",
           150 => x"90",
           151 => x"94",
           152 => x"d8",
           153 => x"94",
           154 => x"80",
           155 => x"ca",
           156 => x"a0",
           157 => x"ca",
           158 => x"c0",
           159 => x"91",
           160 => x"90",
           161 => x"91",
           162 => x"88",
           163 => x"04",
           164 => x"0c",
           165 => x"2d",
           166 => x"08",
           167 => x"90",
           168 => x"94",
           169 => x"80",
           170 => x"94",
           171 => x"80",
           172 => x"ca",
           173 => x"a6",
           174 => x"ca",
           175 => x"c0",
           176 => x"91",
           177 => x"90",
           178 => x"91",
           179 => x"88",
           180 => x"04",
           181 => x"0c",
           182 => x"2d",
           183 => x"08",
           184 => x"90",
           185 => x"94",
           186 => x"ed",
           187 => x"94",
           188 => x"80",
           189 => x"ca",
           190 => x"90",
           191 => x"ca",
           192 => x"c0",
           193 => x"91",
           194 => x"90",
           195 => x"91",
           196 => x"88",
           197 => x"04",
           198 => x"0c",
           199 => x"2d",
           200 => x"08",
           201 => x"90",
           202 => x"94",
           203 => x"9c",
           204 => x"94",
           205 => x"80",
           206 => x"ca",
           207 => x"e9",
           208 => x"ca",
           209 => x"c0",
           210 => x"91",
           211 => x"90",
           212 => x"91",
           213 => x"88",
           214 => x"04",
           215 => x"0c",
           216 => x"2d",
           217 => x"08",
           218 => x"90",
           219 => x"94",
           220 => x"9c",
           221 => x"94",
           222 => x"80",
           223 => x"ca",
           224 => x"f6",
           225 => x"ca",
           226 => x"c0",
           227 => x"91",
           228 => x"90",
           229 => x"91",
           230 => x"88",
           231 => x"04",
           232 => x"0c",
           233 => x"2d",
           234 => x"08",
           235 => x"90",
           236 => x"94",
           237 => x"da",
           238 => x"94",
           239 => x"80",
           240 => x"ca",
           241 => x"f2",
           242 => x"ca",
           243 => x"c0",
           244 => x"91",
           245 => x"90",
           246 => x"91",
           247 => x"88",
           248 => x"04",
           249 => x"0c",
           250 => x"2d",
           251 => x"08",
           252 => x"90",
           253 => x"94",
           254 => x"b7",
           255 => x"94",
           256 => x"80",
           257 => x"ca",
           258 => x"f3",
           259 => x"ca",
           260 => x"c0",
           261 => x"91",
           262 => x"91",
           263 => x"91",
           264 => x"88",
           265 => x"04",
           266 => x"0c",
           267 => x"2d",
           268 => x"08",
           269 => x"90",
           270 => x"94",
           271 => x"ed",
           272 => x"94",
           273 => x"80",
           274 => x"ca",
           275 => x"e9",
           276 => x"ca",
           277 => x"c0",
           278 => x"91",
           279 => x"90",
           280 => x"91",
           281 => x"88",
           282 => x"04",
           283 => x"0c",
           284 => x"2d",
           285 => x"08",
           286 => x"90",
           287 => x"94",
           288 => x"a9",
           289 => x"94",
           290 => x"80",
           291 => x"ca",
           292 => x"84",
           293 => x"ca",
           294 => x"c0",
           295 => x"91",
           296 => x"91",
           297 => x"91",
           298 => x"88",
           299 => x"04",
           300 => x"0c",
           301 => x"2d",
           302 => x"08",
           303 => x"90",
           304 => x"94",
           305 => x"e1",
           306 => x"94",
           307 => x"80",
           308 => x"ca",
           309 => x"ac",
           310 => x"ca",
           311 => x"c0",
           312 => x"91",
           313 => x"90",
           314 => x"91",
           315 => x"88",
           316 => x"04",
           317 => x"0c",
           318 => x"2d",
           319 => x"08",
           320 => x"90",
           321 => x"94",
           322 => x"b2",
           323 => x"94",
           324 => x"80",
           325 => x"ca",
           326 => x"91",
           327 => x"ca",
           328 => x"c0",
           329 => x"91",
           330 => x"90",
           331 => x"91",
           332 => x"88",
           333 => x"04",
           334 => x"0c",
           335 => x"2d",
           336 => x"08",
           337 => x"90",
           338 => x"88",
           339 => x"8c",
           340 => x"80",
           341 => x"05",
           342 => x"0b",
           343 => x"04",
           344 => x"51",
           345 => x"04",
           346 => x"ca",
           347 => x"91",
           348 => x"fd",
           349 => x"53",
           350 => x"08",
           351 => x"52",
           352 => x"08",
           353 => x"51",
           354 => x"91",
           355 => x"70",
           356 => x"0c",
           357 => x"0d",
           358 => x"0c",
           359 => x"94",
           360 => x"ca",
           361 => x"3d",
           362 => x"91",
           363 => x"8c",
           364 => x"91",
           365 => x"88",
           366 => x"93",
           367 => x"88",
           368 => x"ca",
           369 => x"85",
           370 => x"ca",
           371 => x"91",
           372 => x"02",
           373 => x"0c",
           374 => x"81",
           375 => x"94",
           376 => x"0c",
           377 => x"ca",
           378 => x"05",
           379 => x"94",
           380 => x"08",
           381 => x"08",
           382 => x"27",
           383 => x"ca",
           384 => x"05",
           385 => x"ae",
           386 => x"91",
           387 => x"8c",
           388 => x"a2",
           389 => x"94",
           390 => x"08",
           391 => x"94",
           392 => x"0c",
           393 => x"08",
           394 => x"10",
           395 => x"08",
           396 => x"ff",
           397 => x"ca",
           398 => x"05",
           399 => x"80",
           400 => x"ca",
           401 => x"05",
           402 => x"94",
           403 => x"08",
           404 => x"91",
           405 => x"88",
           406 => x"ca",
           407 => x"05",
           408 => x"ca",
           409 => x"05",
           410 => x"94",
           411 => x"08",
           412 => x"08",
           413 => x"07",
           414 => x"08",
           415 => x"91",
           416 => x"fc",
           417 => x"2a",
           418 => x"08",
           419 => x"91",
           420 => x"8c",
           421 => x"2a",
           422 => x"08",
           423 => x"ff",
           424 => x"ca",
           425 => x"05",
           426 => x"93",
           427 => x"94",
           428 => x"08",
           429 => x"94",
           430 => x"0c",
           431 => x"91",
           432 => x"f8",
           433 => x"91",
           434 => x"f4",
           435 => x"91",
           436 => x"f4",
           437 => x"ca",
           438 => x"3d",
           439 => x"94",
           440 => x"3d",
           441 => x"71",
           442 => x"9f",
           443 => x"55",
           444 => x"72",
           445 => x"74",
           446 => x"70",
           447 => x"38",
           448 => x"71",
           449 => x"38",
           450 => x"81",
           451 => x"ff",
           452 => x"ff",
           453 => x"06",
           454 => x"91",
           455 => x"86",
           456 => x"74",
           457 => x"75",
           458 => x"90",
           459 => x"54",
           460 => x"27",
           461 => x"71",
           462 => x"53",
           463 => x"70",
           464 => x"0c",
           465 => x"84",
           466 => x"72",
           467 => x"05",
           468 => x"12",
           469 => x"26",
           470 => x"72",
           471 => x"72",
           472 => x"05",
           473 => x"12",
           474 => x"26",
           475 => x"53",
           476 => x"fb",
           477 => x"79",
           478 => x"83",
           479 => x"52",
           480 => x"71",
           481 => x"54",
           482 => x"73",
           483 => x"c6",
           484 => x"54",
           485 => x"70",
           486 => x"52",
           487 => x"2e",
           488 => x"33",
           489 => x"2e",
           490 => x"95",
           491 => x"81",
           492 => x"70",
           493 => x"54",
           494 => x"70",
           495 => x"33",
           496 => x"ff",
           497 => x"ff",
           498 => x"31",
           499 => x"0c",
           500 => x"3d",
           501 => x"09",
           502 => x"fd",
           503 => x"70",
           504 => x"81",
           505 => x"51",
           506 => x"38",
           507 => x"16",
           508 => x"56",
           509 => x"08",
           510 => x"73",
           511 => x"ff",
           512 => x"0b",
           513 => x"0c",
           514 => x"04",
           515 => x"80",
           516 => x"71",
           517 => x"87",
           518 => x"ca",
           519 => x"ff",
           520 => x"ff",
           521 => x"72",
           522 => x"38",
           523 => x"88",
           524 => x"0d",
           525 => x"0d",
           526 => x"70",
           527 => x"71",
           528 => x"ca",
           529 => x"51",
           530 => x"09",
           531 => x"38",
           532 => x"f1",
           533 => x"84",
           534 => x"53",
           535 => x"70",
           536 => x"53",
           537 => x"a0",
           538 => x"81",
           539 => x"2e",
           540 => x"e5",
           541 => x"ff",
           542 => x"a0",
           543 => x"06",
           544 => x"73",
           545 => x"55",
           546 => x"0c",
           547 => x"91",
           548 => x"87",
           549 => x"fc",
           550 => x"53",
           551 => x"2e",
           552 => x"3d",
           553 => x"72",
           554 => x"3f",
           555 => x"08",
           556 => x"53",
           557 => x"53",
           558 => x"88",
           559 => x"0d",
           560 => x"0d",
           561 => x"33",
           562 => x"53",
           563 => x"8b",
           564 => x"38",
           565 => x"ff",
           566 => x"52",
           567 => x"81",
           568 => x"13",
           569 => x"52",
           570 => x"80",
           571 => x"13",
           572 => x"52",
           573 => x"80",
           574 => x"13",
           575 => x"52",
           576 => x"80",
           577 => x"13",
           578 => x"52",
           579 => x"26",
           580 => x"8a",
           581 => x"87",
           582 => x"e7",
           583 => x"38",
           584 => x"c0",
           585 => x"72",
           586 => x"98",
           587 => x"13",
           588 => x"98",
           589 => x"13",
           590 => x"98",
           591 => x"13",
           592 => x"98",
           593 => x"13",
           594 => x"98",
           595 => x"13",
           596 => x"98",
           597 => x"87",
           598 => x"0c",
           599 => x"98",
           600 => x"0b",
           601 => x"9c",
           602 => x"71",
           603 => x"0c",
           604 => x"04",
           605 => x"7f",
           606 => x"98",
           607 => x"7d",
           608 => x"98",
           609 => x"7d",
           610 => x"c0",
           611 => x"5a",
           612 => x"34",
           613 => x"b4",
           614 => x"83",
           615 => x"c0",
           616 => x"5a",
           617 => x"34",
           618 => x"ac",
           619 => x"85",
           620 => x"c0",
           621 => x"5a",
           622 => x"34",
           623 => x"a4",
           624 => x"88",
           625 => x"c0",
           626 => x"5a",
           627 => x"23",
           628 => x"79",
           629 => x"06",
           630 => x"ff",
           631 => x"86",
           632 => x"85",
           633 => x"84",
           634 => x"83",
           635 => x"82",
           636 => x"7d",
           637 => x"06",
           638 => x"ec",
           639 => x"3f",
           640 => x"04",
           641 => x"02",
           642 => x"70",
           643 => x"2a",
           644 => x"70",
           645 => x"c6",
           646 => x"3d",
           647 => x"3d",
           648 => x"0b",
           649 => x"33",
           650 => x"06",
           651 => x"87",
           652 => x"51",
           653 => x"86",
           654 => x"94",
           655 => x"08",
           656 => x"70",
           657 => x"54",
           658 => x"2e",
           659 => x"91",
           660 => x"06",
           661 => x"d7",
           662 => x"32",
           663 => x"51",
           664 => x"2e",
           665 => x"93",
           666 => x"06",
           667 => x"ff",
           668 => x"81",
           669 => x"87",
           670 => x"52",
           671 => x"86",
           672 => x"94",
           673 => x"72",
           674 => x"ca",
           675 => x"3d",
           676 => x"3d",
           677 => x"05",
           678 => x"91",
           679 => x"70",
           680 => x"57",
           681 => x"c0",
           682 => x"74",
           683 => x"38",
           684 => x"94",
           685 => x"70",
           686 => x"81",
           687 => x"52",
           688 => x"8c",
           689 => x"2a",
           690 => x"51",
           691 => x"38",
           692 => x"70",
           693 => x"51",
           694 => x"8d",
           695 => x"2a",
           696 => x"51",
           697 => x"be",
           698 => x"ff",
           699 => x"c0",
           700 => x"70",
           701 => x"38",
           702 => x"90",
           703 => x"0c",
           704 => x"04",
           705 => x"79",
           706 => x"33",
           707 => x"06",
           708 => x"70",
           709 => x"fe",
           710 => x"ff",
           711 => x"0b",
           712 => x"e0",
           713 => x"ff",
           714 => x"55",
           715 => x"94",
           716 => x"80",
           717 => x"87",
           718 => x"51",
           719 => x"96",
           720 => x"06",
           721 => x"70",
           722 => x"38",
           723 => x"70",
           724 => x"51",
           725 => x"72",
           726 => x"81",
           727 => x"70",
           728 => x"38",
           729 => x"70",
           730 => x"51",
           731 => x"38",
           732 => x"06",
           733 => x"94",
           734 => x"80",
           735 => x"87",
           736 => x"52",
           737 => x"81",
           738 => x"70",
           739 => x"53",
           740 => x"ff",
           741 => x"91",
           742 => x"89",
           743 => x"fe",
           744 => x"0b",
           745 => x"33",
           746 => x"06",
           747 => x"c0",
           748 => x"72",
           749 => x"38",
           750 => x"94",
           751 => x"70",
           752 => x"81",
           753 => x"51",
           754 => x"e2",
           755 => x"ff",
           756 => x"c0",
           757 => x"70",
           758 => x"38",
           759 => x"90",
           760 => x"70",
           761 => x"91",
           762 => x"51",
           763 => x"04",
           764 => x"0b",
           765 => x"e0",
           766 => x"ff",
           767 => x"87",
           768 => x"52",
           769 => x"86",
           770 => x"94",
           771 => x"08",
           772 => x"70",
           773 => x"51",
           774 => x"70",
           775 => x"38",
           776 => x"06",
           777 => x"94",
           778 => x"80",
           779 => x"87",
           780 => x"52",
           781 => x"98",
           782 => x"2c",
           783 => x"71",
           784 => x"0c",
           785 => x"04",
           786 => x"87",
           787 => x"08",
           788 => x"8a",
           789 => x"70",
           790 => x"93",
           791 => x"9e",
           792 => x"c6",
           793 => x"c0",
           794 => x"91",
           795 => x"87",
           796 => x"08",
           797 => x"0c",
           798 => x"90",
           799 => x"f0",
           800 => x"9e",
           801 => x"c6",
           802 => x"c0",
           803 => x"91",
           804 => x"87",
           805 => x"08",
           806 => x"0c",
           807 => x"a8",
           808 => x"80",
           809 => x"9e",
           810 => x"c7",
           811 => x"c0",
           812 => x"51",
           813 => x"88",
           814 => x"9e",
           815 => x"c7",
           816 => x"0b",
           817 => x"34",
           818 => x"c0",
           819 => x"70",
           820 => x"51",
           821 => x"80",
           822 => x"81",
           823 => x"c7",
           824 => x"0b",
           825 => x"88",
           826 => x"80",
           827 => x"52",
           828 => x"2e",
           829 => x"52",
           830 => x"92",
           831 => x"87",
           832 => x"08",
           833 => x"80",
           834 => x"52",
           835 => x"83",
           836 => x"71",
           837 => x"34",
           838 => x"c0",
           839 => x"70",
           840 => x"51",
           841 => x"80",
           842 => x"81",
           843 => x"c7",
           844 => x"0b",
           845 => x"88",
           846 => x"80",
           847 => x"52",
           848 => x"83",
           849 => x"71",
           850 => x"34",
           851 => x"c0",
           852 => x"70",
           853 => x"51",
           854 => x"80",
           855 => x"81",
           856 => x"c7",
           857 => x"0b",
           858 => x"88",
           859 => x"80",
           860 => x"52",
           861 => x"83",
           862 => x"71",
           863 => x"34",
           864 => x"c0",
           865 => x"70",
           866 => x"51",
           867 => x"80",
           868 => x"81",
           869 => x"c7",
           870 => x"c0",
           871 => x"70",
           872 => x"70",
           873 => x"51",
           874 => x"c7",
           875 => x"0b",
           876 => x"88",
           877 => x"06",
           878 => x"70",
           879 => x"38",
           880 => x"91",
           881 => x"80",
           882 => x"9e",
           883 => x"88",
           884 => x"52",
           885 => x"83",
           886 => x"71",
           887 => x"34",
           888 => x"88",
           889 => x"06",
           890 => x"91",
           891 => x"83",
           892 => x"fd",
           893 => x"b4",
           894 => x"a3",
           895 => x"90",
           896 => x"80",
           897 => x"91",
           898 => x"84",
           899 => x"b4",
           900 => x"8b",
           901 => x"91",
           902 => x"80",
           903 => x"91",
           904 => x"53",
           905 => x"08",
           906 => x"c4",
           907 => x"3f",
           908 => x"33",
           909 => x"2e",
           910 => x"c6",
           911 => x"91",
           912 => x"52",
           913 => x"51",
           914 => x"91",
           915 => x"54",
           916 => x"91",
           917 => x"54",
           918 => x"92",
           919 => x"f8",
           920 => x"c6",
           921 => x"91",
           922 => x"89",
           923 => x"c7",
           924 => x"73",
           925 => x"38",
           926 => x"51",
           927 => x"91",
           928 => x"54",
           929 => x"88",
           930 => x"c0",
           931 => x"3f",
           932 => x"33",
           933 => x"2e",
           934 => x"b5",
           935 => x"ff",
           936 => x"98",
           937 => x"80",
           938 => x"91",
           939 => x"52",
           940 => x"51",
           941 => x"91",
           942 => x"54",
           943 => x"88",
           944 => x"f8",
           945 => x"3f",
           946 => x"33",
           947 => x"2e",
           948 => x"c7",
           949 => x"91",
           950 => x"88",
           951 => x"b6",
           952 => x"bb",
           953 => x"fc",
           954 => x"b6",
           955 => x"93",
           956 => x"80",
           957 => x"b6",
           958 => x"87",
           959 => x"84",
           960 => x"b7",
           961 => x"fb",
           962 => x"88",
           963 => x"b7",
           964 => x"ef",
           965 => x"8c",
           966 => x"b7",
           967 => x"e3",
           968 => x"0d",
           969 => x"0d",
           970 => x"33",
           971 => x"71",
           972 => x"38",
           973 => x"0b",
           974 => x"88",
           975 => x"08",
           976 => x"84",
           977 => x"91",
           978 => x"97",
           979 => x"94",
           980 => x"91",
           981 => x"8b",
           982 => x"a0",
           983 => x"91",
           984 => x"f7",
           985 => x"3d",
           986 => x"88",
           987 => x"80",
           988 => x"96",
           989 => x"ff",
           990 => x"c0",
           991 => x"08",
           992 => x"72",
           993 => x"07",
           994 => x"a0",
           995 => x"83",
           996 => x"ff",
           997 => x"c0",
           998 => x"08",
           999 => x"0c",
          1000 => x"0c",
          1001 => x"91",
          1002 => x"06",
          1003 => x"a0",
          1004 => x"51",
          1005 => x"04",
          1006 => x"08",
          1007 => x"84",
          1008 => x"3d",
          1009 => x"05",
          1010 => x"8a",
          1011 => x"06",
          1012 => x"51",
          1013 => x"ca",
          1014 => x"71",
          1015 => x"38",
          1016 => x"91",
          1017 => x"81",
          1018 => x"a0",
          1019 => x"91",
          1020 => x"52",
          1021 => x"85",
          1022 => x"71",
          1023 => x"0d",
          1024 => x"0d",
          1025 => x"33",
          1026 => x"08",
          1027 => x"98",
          1028 => x"ff",
          1029 => x"91",
          1030 => x"84",
          1031 => x"fd",
          1032 => x"54",
          1033 => x"81",
          1034 => x"53",
          1035 => x"8e",
          1036 => x"ff",
          1037 => x"14",
          1038 => x"3f",
          1039 => x"3d",
          1040 => x"3d",
          1041 => x"ca",
          1042 => x"91",
          1043 => x"56",
          1044 => x"70",
          1045 => x"53",
          1046 => x"2e",
          1047 => x"81",
          1048 => x"81",
          1049 => x"da",
          1050 => x"74",
          1051 => x"0c",
          1052 => x"04",
          1053 => x"66",
          1054 => x"78",
          1055 => x"5a",
          1056 => x"80",
          1057 => x"38",
          1058 => x"09",
          1059 => x"de",
          1060 => x"7a",
          1061 => x"5c",
          1062 => x"5b",
          1063 => x"09",
          1064 => x"38",
          1065 => x"39",
          1066 => x"09",
          1067 => x"38",
          1068 => x"70",
          1069 => x"33",
          1070 => x"2e",
          1071 => x"92",
          1072 => x"19",
          1073 => x"70",
          1074 => x"33",
          1075 => x"53",
          1076 => x"16",
          1077 => x"26",
          1078 => x"88",
          1079 => x"05",
          1080 => x"05",
          1081 => x"05",
          1082 => x"5b",
          1083 => x"80",
          1084 => x"30",
          1085 => x"80",
          1086 => x"cc",
          1087 => x"70",
          1088 => x"25",
          1089 => x"54",
          1090 => x"53",
          1091 => x"8c",
          1092 => x"07",
          1093 => x"05",
          1094 => x"5a",
          1095 => x"83",
          1096 => x"54",
          1097 => x"27",
          1098 => x"16",
          1099 => x"06",
          1100 => x"80",
          1101 => x"aa",
          1102 => x"cf",
          1103 => x"73",
          1104 => x"81",
          1105 => x"80",
          1106 => x"38",
          1107 => x"2e",
          1108 => x"81",
          1109 => x"80",
          1110 => x"8a",
          1111 => x"39",
          1112 => x"2e",
          1113 => x"73",
          1114 => x"8a",
          1115 => x"d3",
          1116 => x"80",
          1117 => x"80",
          1118 => x"ee",
          1119 => x"39",
          1120 => x"71",
          1121 => x"53",
          1122 => x"54",
          1123 => x"2e",
          1124 => x"15",
          1125 => x"33",
          1126 => x"72",
          1127 => x"81",
          1128 => x"39",
          1129 => x"56",
          1130 => x"27",
          1131 => x"51",
          1132 => x"75",
          1133 => x"72",
          1134 => x"38",
          1135 => x"df",
          1136 => x"16",
          1137 => x"7b",
          1138 => x"38",
          1139 => x"f2",
          1140 => x"77",
          1141 => x"12",
          1142 => x"53",
          1143 => x"5c",
          1144 => x"5c",
          1145 => x"5c",
          1146 => x"5c",
          1147 => x"51",
          1148 => x"fd",
          1149 => x"82",
          1150 => x"06",
          1151 => x"80",
          1152 => x"77",
          1153 => x"53",
          1154 => x"18",
          1155 => x"72",
          1156 => x"c4",
          1157 => x"70",
          1158 => x"25",
          1159 => x"55",
          1160 => x"8d",
          1161 => x"2e",
          1162 => x"30",
          1163 => x"5b",
          1164 => x"8f",
          1165 => x"7b",
          1166 => x"e6",
          1167 => x"ca",
          1168 => x"ff",
          1169 => x"75",
          1170 => x"9e",
          1171 => x"88",
          1172 => x"74",
          1173 => x"a7",
          1174 => x"80",
          1175 => x"38",
          1176 => x"72",
          1177 => x"54",
          1178 => x"72",
          1179 => x"05",
          1180 => x"17",
          1181 => x"77",
          1182 => x"51",
          1183 => x"9f",
          1184 => x"72",
          1185 => x"79",
          1186 => x"81",
          1187 => x"72",
          1188 => x"38",
          1189 => x"05",
          1190 => x"ad",
          1191 => x"17",
          1192 => x"81",
          1193 => x"b0",
          1194 => x"38",
          1195 => x"81",
          1196 => x"06",
          1197 => x"9f",
          1198 => x"55",
          1199 => x"97",
          1200 => x"f9",
          1201 => x"81",
          1202 => x"8b",
          1203 => x"16",
          1204 => x"73",
          1205 => x"96",
          1206 => x"e0",
          1207 => x"17",
          1208 => x"33",
          1209 => x"f9",
          1210 => x"f2",
          1211 => x"16",
          1212 => x"7b",
          1213 => x"38",
          1214 => x"c6",
          1215 => x"96",
          1216 => x"fd",
          1217 => x"3d",
          1218 => x"05",
          1219 => x"52",
          1220 => x"e0",
          1221 => x"0d",
          1222 => x"0d",
          1223 => x"a0",
          1224 => x"88",
          1225 => x"51",
          1226 => x"91",
          1227 => x"53",
          1228 => x"80",
          1229 => x"a0",
          1230 => x"0d",
          1231 => x"0d",
          1232 => x"08",
          1233 => x"98",
          1234 => x"88",
          1235 => x"52",
          1236 => x"3f",
          1237 => x"98",
          1238 => x"0d",
          1239 => x"0d",
          1240 => x"ca",
          1241 => x"56",
          1242 => x"80",
          1243 => x"2e",
          1244 => x"91",
          1245 => x"52",
          1246 => x"ca",
          1247 => x"ff",
          1248 => x"80",
          1249 => x"38",
          1250 => x"b9",
          1251 => x"32",
          1252 => x"80",
          1253 => x"52",
          1254 => x"8b",
          1255 => x"2e",
          1256 => x"14",
          1257 => x"9f",
          1258 => x"38",
          1259 => x"73",
          1260 => x"38",
          1261 => x"72",
          1262 => x"14",
          1263 => x"f8",
          1264 => x"af",
          1265 => x"52",
          1266 => x"8a",
          1267 => x"3f",
          1268 => x"91",
          1269 => x"87",
          1270 => x"fe",
          1271 => x"ca",
          1272 => x"91",
          1273 => x"77",
          1274 => x"53",
          1275 => x"72",
          1276 => x"0c",
          1277 => x"04",
          1278 => x"7a",
          1279 => x"80",
          1280 => x"58",
          1281 => x"33",
          1282 => x"a0",
          1283 => x"06",
          1284 => x"13",
          1285 => x"39",
          1286 => x"09",
          1287 => x"38",
          1288 => x"11",
          1289 => x"08",
          1290 => x"54",
          1291 => x"2e",
          1292 => x"80",
          1293 => x"08",
          1294 => x"0c",
          1295 => x"33",
          1296 => x"80",
          1297 => x"38",
          1298 => x"80",
          1299 => x"38",
          1300 => x"57",
          1301 => x"0c",
          1302 => x"33",
          1303 => x"39",
          1304 => x"74",
          1305 => x"38",
          1306 => x"80",
          1307 => x"89",
          1308 => x"38",
          1309 => x"d0",
          1310 => x"55",
          1311 => x"80",
          1312 => x"39",
          1313 => x"d9",
          1314 => x"80",
          1315 => x"27",
          1316 => x"80",
          1317 => x"89",
          1318 => x"70",
          1319 => x"55",
          1320 => x"70",
          1321 => x"55",
          1322 => x"27",
          1323 => x"14",
          1324 => x"06",
          1325 => x"74",
          1326 => x"73",
          1327 => x"38",
          1328 => x"14",
          1329 => x"05",
          1330 => x"08",
          1331 => x"54",
          1332 => x"39",
          1333 => x"84",
          1334 => x"55",
          1335 => x"81",
          1336 => x"ca",
          1337 => x"3d",
          1338 => x"3d",
          1339 => x"5a",
          1340 => x"7a",
          1341 => x"08",
          1342 => x"53",
          1343 => x"09",
          1344 => x"38",
          1345 => x"0c",
          1346 => x"ad",
          1347 => x"06",
          1348 => x"76",
          1349 => x"0c",
          1350 => x"33",
          1351 => x"73",
          1352 => x"81",
          1353 => x"38",
          1354 => x"05",
          1355 => x"08",
          1356 => x"53",
          1357 => x"2e",
          1358 => x"57",
          1359 => x"2e",
          1360 => x"39",
          1361 => x"13",
          1362 => x"08",
          1363 => x"53",
          1364 => x"55",
          1365 => x"80",
          1366 => x"14",
          1367 => x"88",
          1368 => x"27",
          1369 => x"eb",
          1370 => x"53",
          1371 => x"89",
          1372 => x"38",
          1373 => x"55",
          1374 => x"8a",
          1375 => x"a0",
          1376 => x"c2",
          1377 => x"74",
          1378 => x"e0",
          1379 => x"ff",
          1380 => x"d0",
          1381 => x"ff",
          1382 => x"90",
          1383 => x"38",
          1384 => x"81",
          1385 => x"53",
          1386 => x"ca",
          1387 => x"27",
          1388 => x"77",
          1389 => x"08",
          1390 => x"0c",
          1391 => x"33",
          1392 => x"ff",
          1393 => x"80",
          1394 => x"74",
          1395 => x"79",
          1396 => x"74",
          1397 => x"0c",
          1398 => x"04",
          1399 => x"02",
          1400 => x"51",
          1401 => x"72",
          1402 => x"91",
          1403 => x"33",
          1404 => x"ca",
          1405 => x"3d",
          1406 => x"3d",
          1407 => x"05",
          1408 => x"05",
          1409 => x"56",
          1410 => x"72",
          1411 => x"e0",
          1412 => x"2b",
          1413 => x"8c",
          1414 => x"88",
          1415 => x"2e",
          1416 => x"88",
          1417 => x"0c",
          1418 => x"8c",
          1419 => x"71",
          1420 => x"87",
          1421 => x"0c",
          1422 => x"08",
          1423 => x"51",
          1424 => x"2e",
          1425 => x"c0",
          1426 => x"51",
          1427 => x"71",
          1428 => x"80",
          1429 => x"92",
          1430 => x"98",
          1431 => x"70",
          1432 => x"38",
          1433 => x"a4",
          1434 => x"c7",
          1435 => x"51",
          1436 => x"88",
          1437 => x"0d",
          1438 => x"0d",
          1439 => x"02",
          1440 => x"05",
          1441 => x"58",
          1442 => x"52",
          1443 => x"3f",
          1444 => x"08",
          1445 => x"54",
          1446 => x"be",
          1447 => x"75",
          1448 => x"c0",
          1449 => x"87",
          1450 => x"12",
          1451 => x"84",
          1452 => x"40",
          1453 => x"85",
          1454 => x"98",
          1455 => x"7d",
          1456 => x"0c",
          1457 => x"85",
          1458 => x"06",
          1459 => x"71",
          1460 => x"38",
          1461 => x"71",
          1462 => x"05",
          1463 => x"19",
          1464 => x"a2",
          1465 => x"71",
          1466 => x"38",
          1467 => x"83",
          1468 => x"38",
          1469 => x"8a",
          1470 => x"98",
          1471 => x"71",
          1472 => x"c0",
          1473 => x"52",
          1474 => x"87",
          1475 => x"80",
          1476 => x"81",
          1477 => x"c0",
          1478 => x"53",
          1479 => x"82",
          1480 => x"71",
          1481 => x"1a",
          1482 => x"84",
          1483 => x"19",
          1484 => x"06",
          1485 => x"79",
          1486 => x"38",
          1487 => x"80",
          1488 => x"87",
          1489 => x"26",
          1490 => x"73",
          1491 => x"06",
          1492 => x"2e",
          1493 => x"52",
          1494 => x"91",
          1495 => x"8f",
          1496 => x"f3",
          1497 => x"62",
          1498 => x"05",
          1499 => x"57",
          1500 => x"83",
          1501 => x"52",
          1502 => x"3f",
          1503 => x"08",
          1504 => x"54",
          1505 => x"2e",
          1506 => x"81",
          1507 => x"74",
          1508 => x"c0",
          1509 => x"87",
          1510 => x"12",
          1511 => x"84",
          1512 => x"5f",
          1513 => x"0b",
          1514 => x"8c",
          1515 => x"0c",
          1516 => x"80",
          1517 => x"70",
          1518 => x"81",
          1519 => x"54",
          1520 => x"8c",
          1521 => x"81",
          1522 => x"7c",
          1523 => x"58",
          1524 => x"70",
          1525 => x"52",
          1526 => x"8a",
          1527 => x"98",
          1528 => x"71",
          1529 => x"c0",
          1530 => x"52",
          1531 => x"87",
          1532 => x"80",
          1533 => x"81",
          1534 => x"c0",
          1535 => x"53",
          1536 => x"82",
          1537 => x"71",
          1538 => x"19",
          1539 => x"81",
          1540 => x"ff",
          1541 => x"19",
          1542 => x"78",
          1543 => x"38",
          1544 => x"80",
          1545 => x"87",
          1546 => x"26",
          1547 => x"73",
          1548 => x"06",
          1549 => x"2e",
          1550 => x"52",
          1551 => x"91",
          1552 => x"8f",
          1553 => x"f6",
          1554 => x"02",
          1555 => x"05",
          1556 => x"05",
          1557 => x"71",
          1558 => x"57",
          1559 => x"91",
          1560 => x"81",
          1561 => x"54",
          1562 => x"38",
          1563 => x"c0",
          1564 => x"81",
          1565 => x"2e",
          1566 => x"71",
          1567 => x"38",
          1568 => x"87",
          1569 => x"11",
          1570 => x"80",
          1571 => x"80",
          1572 => x"83",
          1573 => x"38",
          1574 => x"72",
          1575 => x"2a",
          1576 => x"51",
          1577 => x"80",
          1578 => x"87",
          1579 => x"08",
          1580 => x"38",
          1581 => x"8c",
          1582 => x"96",
          1583 => x"0c",
          1584 => x"8c",
          1585 => x"08",
          1586 => x"51",
          1587 => x"38",
          1588 => x"56",
          1589 => x"80",
          1590 => x"85",
          1591 => x"77",
          1592 => x"83",
          1593 => x"75",
          1594 => x"ca",
          1595 => x"3d",
          1596 => x"3d",
          1597 => x"11",
          1598 => x"71",
          1599 => x"91",
          1600 => x"53",
          1601 => x"0d",
          1602 => x"0d",
          1603 => x"33",
          1604 => x"71",
          1605 => x"88",
          1606 => x"14",
          1607 => x"07",
          1608 => x"33",
          1609 => x"ca",
          1610 => x"53",
          1611 => x"52",
          1612 => x"04",
          1613 => x"73",
          1614 => x"92",
          1615 => x"52",
          1616 => x"81",
          1617 => x"70",
          1618 => x"70",
          1619 => x"3d",
          1620 => x"3d",
          1621 => x"52",
          1622 => x"70",
          1623 => x"34",
          1624 => x"51",
          1625 => x"81",
          1626 => x"70",
          1627 => x"70",
          1628 => x"05",
          1629 => x"88",
          1630 => x"72",
          1631 => x"0d",
          1632 => x"0d",
          1633 => x"54",
          1634 => x"80",
          1635 => x"71",
          1636 => x"53",
          1637 => x"81",
          1638 => x"ff",
          1639 => x"39",
          1640 => x"04",
          1641 => x"75",
          1642 => x"52",
          1643 => x"70",
          1644 => x"34",
          1645 => x"70",
          1646 => x"3d",
          1647 => x"3d",
          1648 => x"79",
          1649 => x"74",
          1650 => x"56",
          1651 => x"81",
          1652 => x"71",
          1653 => x"16",
          1654 => x"52",
          1655 => x"86",
          1656 => x"2e",
          1657 => x"91",
          1658 => x"86",
          1659 => x"fe",
          1660 => x"76",
          1661 => x"39",
          1662 => x"8a",
          1663 => x"51",
          1664 => x"71",
          1665 => x"33",
          1666 => x"0c",
          1667 => x"04",
          1668 => x"ca",
          1669 => x"80",
          1670 => x"88",
          1671 => x"3d",
          1672 => x"80",
          1673 => x"33",
          1674 => x"7a",
          1675 => x"38",
          1676 => x"16",
          1677 => x"16",
          1678 => x"17",
          1679 => x"fa",
          1680 => x"ca",
          1681 => x"2e",
          1682 => x"b7",
          1683 => x"88",
          1684 => x"34",
          1685 => x"70",
          1686 => x"31",
          1687 => x"59",
          1688 => x"77",
          1689 => x"82",
          1690 => x"74",
          1691 => x"81",
          1692 => x"81",
          1693 => x"53",
          1694 => x"16",
          1695 => x"e3",
          1696 => x"81",
          1697 => x"ca",
          1698 => x"3d",
          1699 => x"3d",
          1700 => x"56",
          1701 => x"74",
          1702 => x"2e",
          1703 => x"51",
          1704 => x"91",
          1705 => x"57",
          1706 => x"08",
          1707 => x"54",
          1708 => x"16",
          1709 => x"33",
          1710 => x"3f",
          1711 => x"08",
          1712 => x"38",
          1713 => x"57",
          1714 => x"0c",
          1715 => x"88",
          1716 => x"0d",
          1717 => x"0d",
          1718 => x"57",
          1719 => x"91",
          1720 => x"58",
          1721 => x"08",
          1722 => x"76",
          1723 => x"83",
          1724 => x"06",
          1725 => x"84",
          1726 => x"78",
          1727 => x"81",
          1728 => x"38",
          1729 => x"91",
          1730 => x"52",
          1731 => x"52",
          1732 => x"3f",
          1733 => x"52",
          1734 => x"51",
          1735 => x"84",
          1736 => x"d2",
          1737 => x"fc",
          1738 => x"8a",
          1739 => x"52",
          1740 => x"51",
          1741 => x"90",
          1742 => x"84",
          1743 => x"fc",
          1744 => x"17",
          1745 => x"a0",
          1746 => x"86",
          1747 => x"08",
          1748 => x"b0",
          1749 => x"55",
          1750 => x"81",
          1751 => x"f8",
          1752 => x"84",
          1753 => x"53",
          1754 => x"17",
          1755 => x"d7",
          1756 => x"88",
          1757 => x"83",
          1758 => x"77",
          1759 => x"0c",
          1760 => x"04",
          1761 => x"77",
          1762 => x"12",
          1763 => x"55",
          1764 => x"56",
          1765 => x"8d",
          1766 => x"22",
          1767 => x"ac",
          1768 => x"57",
          1769 => x"ca",
          1770 => x"3d",
          1771 => x"3d",
          1772 => x"70",
          1773 => x"57",
          1774 => x"81",
          1775 => x"98",
          1776 => x"81",
          1777 => x"74",
          1778 => x"72",
          1779 => x"f5",
          1780 => x"24",
          1781 => x"81",
          1782 => x"81",
          1783 => x"83",
          1784 => x"38",
          1785 => x"76",
          1786 => x"70",
          1787 => x"16",
          1788 => x"74",
          1789 => x"96",
          1790 => x"88",
          1791 => x"38",
          1792 => x"06",
          1793 => x"33",
          1794 => x"89",
          1795 => x"08",
          1796 => x"54",
          1797 => x"fc",
          1798 => x"ca",
          1799 => x"fe",
          1800 => x"ff",
          1801 => x"11",
          1802 => x"2b",
          1803 => x"81",
          1804 => x"2a",
          1805 => x"51",
          1806 => x"e2",
          1807 => x"ff",
          1808 => x"da",
          1809 => x"2a",
          1810 => x"05",
          1811 => x"fc",
          1812 => x"ca",
          1813 => x"c6",
          1814 => x"83",
          1815 => x"05",
          1816 => x"f9",
          1817 => x"ca",
          1818 => x"ff",
          1819 => x"ae",
          1820 => x"2a",
          1821 => x"05",
          1822 => x"fc",
          1823 => x"ca",
          1824 => x"38",
          1825 => x"83",
          1826 => x"05",
          1827 => x"f8",
          1828 => x"ca",
          1829 => x"0a",
          1830 => x"39",
          1831 => x"91",
          1832 => x"89",
          1833 => x"f8",
          1834 => x"7c",
          1835 => x"56",
          1836 => x"77",
          1837 => x"38",
          1838 => x"08",
          1839 => x"38",
          1840 => x"72",
          1841 => x"9d",
          1842 => x"24",
          1843 => x"81",
          1844 => x"82",
          1845 => x"83",
          1846 => x"38",
          1847 => x"76",
          1848 => x"70",
          1849 => x"18",
          1850 => x"76",
          1851 => x"9e",
          1852 => x"88",
          1853 => x"ca",
          1854 => x"d9",
          1855 => x"ff",
          1856 => x"05",
          1857 => x"81",
          1858 => x"54",
          1859 => x"80",
          1860 => x"77",
          1861 => x"f0",
          1862 => x"8f",
          1863 => x"51",
          1864 => x"34",
          1865 => x"17",
          1866 => x"2a",
          1867 => x"05",
          1868 => x"fa",
          1869 => x"ca",
          1870 => x"91",
          1871 => x"81",
          1872 => x"83",
          1873 => x"b4",
          1874 => x"2a",
          1875 => x"8f",
          1876 => x"2a",
          1877 => x"f0",
          1878 => x"06",
          1879 => x"72",
          1880 => x"ec",
          1881 => x"2a",
          1882 => x"05",
          1883 => x"fa",
          1884 => x"ca",
          1885 => x"91",
          1886 => x"80",
          1887 => x"83",
          1888 => x"52",
          1889 => x"fe",
          1890 => x"b4",
          1891 => x"a4",
          1892 => x"76",
          1893 => x"17",
          1894 => x"75",
          1895 => x"3f",
          1896 => x"08",
          1897 => x"88",
          1898 => x"77",
          1899 => x"77",
          1900 => x"fc",
          1901 => x"b4",
          1902 => x"51",
          1903 => x"c9",
          1904 => x"88",
          1905 => x"06",
          1906 => x"72",
          1907 => x"3f",
          1908 => x"17",
          1909 => x"ca",
          1910 => x"3d",
          1911 => x"3d",
          1912 => x"7e",
          1913 => x"56",
          1914 => x"75",
          1915 => x"74",
          1916 => x"27",
          1917 => x"80",
          1918 => x"ff",
          1919 => x"75",
          1920 => x"3f",
          1921 => x"08",
          1922 => x"88",
          1923 => x"38",
          1924 => x"54",
          1925 => x"81",
          1926 => x"39",
          1927 => x"08",
          1928 => x"39",
          1929 => x"51",
          1930 => x"91",
          1931 => x"58",
          1932 => x"08",
          1933 => x"c7",
          1934 => x"88",
          1935 => x"d2",
          1936 => x"88",
          1937 => x"cf",
          1938 => x"74",
          1939 => x"fc",
          1940 => x"ca",
          1941 => x"38",
          1942 => x"fe",
          1943 => x"08",
          1944 => x"74",
          1945 => x"38",
          1946 => x"17",
          1947 => x"33",
          1948 => x"73",
          1949 => x"77",
          1950 => x"26",
          1951 => x"80",
          1952 => x"ca",
          1953 => x"3d",
          1954 => x"3d",
          1955 => x"71",
          1956 => x"5b",
          1957 => x"8c",
          1958 => x"77",
          1959 => x"38",
          1960 => x"78",
          1961 => x"81",
          1962 => x"79",
          1963 => x"f9",
          1964 => x"55",
          1965 => x"88",
          1966 => x"e0",
          1967 => x"88",
          1968 => x"ca",
          1969 => x"2e",
          1970 => x"98",
          1971 => x"ca",
          1972 => x"82",
          1973 => x"58",
          1974 => x"70",
          1975 => x"80",
          1976 => x"38",
          1977 => x"09",
          1978 => x"e2",
          1979 => x"56",
          1980 => x"76",
          1981 => x"82",
          1982 => x"7a",
          1983 => x"3f",
          1984 => x"ca",
          1985 => x"2e",
          1986 => x"86",
          1987 => x"88",
          1988 => x"ca",
          1989 => x"70",
          1990 => x"07",
          1991 => x"7c",
          1992 => x"88",
          1993 => x"51",
          1994 => x"81",
          1995 => x"ca",
          1996 => x"2e",
          1997 => x"17",
          1998 => x"74",
          1999 => x"73",
          2000 => x"27",
          2001 => x"58",
          2002 => x"80",
          2003 => x"56",
          2004 => x"98",
          2005 => x"26",
          2006 => x"56",
          2007 => x"81",
          2008 => x"52",
          2009 => x"c6",
          2010 => x"88",
          2011 => x"b8",
          2012 => x"91",
          2013 => x"81",
          2014 => x"06",
          2015 => x"ca",
          2016 => x"91",
          2017 => x"09",
          2018 => x"72",
          2019 => x"70",
          2020 => x"51",
          2021 => x"80",
          2022 => x"78",
          2023 => x"06",
          2024 => x"73",
          2025 => x"39",
          2026 => x"52",
          2027 => x"f7",
          2028 => x"88",
          2029 => x"88",
          2030 => x"91",
          2031 => x"07",
          2032 => x"55",
          2033 => x"2e",
          2034 => x"80",
          2035 => x"75",
          2036 => x"76",
          2037 => x"3f",
          2038 => x"08",
          2039 => x"38",
          2040 => x"0c",
          2041 => x"fe",
          2042 => x"08",
          2043 => x"74",
          2044 => x"ff",
          2045 => x"0c",
          2046 => x"81",
          2047 => x"84",
          2048 => x"39",
          2049 => x"81",
          2050 => x"8c",
          2051 => x"8c",
          2052 => x"88",
          2053 => x"39",
          2054 => x"55",
          2055 => x"88",
          2056 => x"0d",
          2057 => x"0d",
          2058 => x"55",
          2059 => x"91",
          2060 => x"58",
          2061 => x"ca",
          2062 => x"d8",
          2063 => x"74",
          2064 => x"3f",
          2065 => x"08",
          2066 => x"08",
          2067 => x"59",
          2068 => x"77",
          2069 => x"70",
          2070 => x"c8",
          2071 => x"84",
          2072 => x"56",
          2073 => x"58",
          2074 => x"97",
          2075 => x"75",
          2076 => x"52",
          2077 => x"51",
          2078 => x"91",
          2079 => x"80",
          2080 => x"8a",
          2081 => x"32",
          2082 => x"72",
          2083 => x"2a",
          2084 => x"56",
          2085 => x"88",
          2086 => x"0d",
          2087 => x"0d",
          2088 => x"08",
          2089 => x"74",
          2090 => x"26",
          2091 => x"74",
          2092 => x"72",
          2093 => x"74",
          2094 => x"88",
          2095 => x"73",
          2096 => x"33",
          2097 => x"27",
          2098 => x"16",
          2099 => x"9b",
          2100 => x"2a",
          2101 => x"88",
          2102 => x"58",
          2103 => x"80",
          2104 => x"16",
          2105 => x"0c",
          2106 => x"8a",
          2107 => x"89",
          2108 => x"72",
          2109 => x"38",
          2110 => x"51",
          2111 => x"91",
          2112 => x"54",
          2113 => x"08",
          2114 => x"38",
          2115 => x"ca",
          2116 => x"8b",
          2117 => x"08",
          2118 => x"08",
          2119 => x"82",
          2120 => x"74",
          2121 => x"cb",
          2122 => x"75",
          2123 => x"3f",
          2124 => x"08",
          2125 => x"73",
          2126 => x"98",
          2127 => x"82",
          2128 => x"2e",
          2129 => x"39",
          2130 => x"39",
          2131 => x"13",
          2132 => x"74",
          2133 => x"16",
          2134 => x"18",
          2135 => x"77",
          2136 => x"0c",
          2137 => x"04",
          2138 => x"7a",
          2139 => x"12",
          2140 => x"59",
          2141 => x"80",
          2142 => x"86",
          2143 => x"98",
          2144 => x"14",
          2145 => x"55",
          2146 => x"81",
          2147 => x"83",
          2148 => x"77",
          2149 => x"81",
          2150 => x"0c",
          2151 => x"55",
          2152 => x"76",
          2153 => x"17",
          2154 => x"74",
          2155 => x"9b",
          2156 => x"39",
          2157 => x"ff",
          2158 => x"2a",
          2159 => x"81",
          2160 => x"52",
          2161 => x"e6",
          2162 => x"88",
          2163 => x"55",
          2164 => x"ca",
          2165 => x"80",
          2166 => x"55",
          2167 => x"08",
          2168 => x"f4",
          2169 => x"08",
          2170 => x"08",
          2171 => x"38",
          2172 => x"77",
          2173 => x"84",
          2174 => x"39",
          2175 => x"52",
          2176 => x"86",
          2177 => x"88",
          2178 => x"55",
          2179 => x"08",
          2180 => x"c4",
          2181 => x"91",
          2182 => x"81",
          2183 => x"81",
          2184 => x"88",
          2185 => x"b0",
          2186 => x"88",
          2187 => x"51",
          2188 => x"91",
          2189 => x"a0",
          2190 => x"15",
          2191 => x"75",
          2192 => x"3f",
          2193 => x"08",
          2194 => x"76",
          2195 => x"77",
          2196 => x"9c",
          2197 => x"55",
          2198 => x"88",
          2199 => x"0d",
          2200 => x"0d",
          2201 => x"08",
          2202 => x"80",
          2203 => x"fc",
          2204 => x"ca",
          2205 => x"91",
          2206 => x"80",
          2207 => x"ca",
          2208 => x"98",
          2209 => x"78",
          2210 => x"3f",
          2211 => x"08",
          2212 => x"88",
          2213 => x"38",
          2214 => x"08",
          2215 => x"70",
          2216 => x"58",
          2217 => x"2e",
          2218 => x"83",
          2219 => x"91",
          2220 => x"55",
          2221 => x"81",
          2222 => x"07",
          2223 => x"2e",
          2224 => x"16",
          2225 => x"2e",
          2226 => x"88",
          2227 => x"91",
          2228 => x"56",
          2229 => x"51",
          2230 => x"91",
          2231 => x"54",
          2232 => x"08",
          2233 => x"9b",
          2234 => x"2e",
          2235 => x"83",
          2236 => x"73",
          2237 => x"0c",
          2238 => x"04",
          2239 => x"76",
          2240 => x"54",
          2241 => x"91",
          2242 => x"83",
          2243 => x"76",
          2244 => x"53",
          2245 => x"2e",
          2246 => x"90",
          2247 => x"51",
          2248 => x"91",
          2249 => x"90",
          2250 => x"53",
          2251 => x"88",
          2252 => x"0d",
          2253 => x"0d",
          2254 => x"83",
          2255 => x"54",
          2256 => x"55",
          2257 => x"3f",
          2258 => x"51",
          2259 => x"2e",
          2260 => x"8b",
          2261 => x"2a",
          2262 => x"51",
          2263 => x"86",
          2264 => x"f7",
          2265 => x"7d",
          2266 => x"75",
          2267 => x"98",
          2268 => x"2e",
          2269 => x"98",
          2270 => x"78",
          2271 => x"3f",
          2272 => x"08",
          2273 => x"88",
          2274 => x"38",
          2275 => x"70",
          2276 => x"73",
          2277 => x"58",
          2278 => x"8b",
          2279 => x"bf",
          2280 => x"ff",
          2281 => x"53",
          2282 => x"34",
          2283 => x"08",
          2284 => x"e5",
          2285 => x"81",
          2286 => x"2e",
          2287 => x"70",
          2288 => x"57",
          2289 => x"9e",
          2290 => x"2e",
          2291 => x"ca",
          2292 => x"df",
          2293 => x"72",
          2294 => x"81",
          2295 => x"76",
          2296 => x"2e",
          2297 => x"52",
          2298 => x"fc",
          2299 => x"88",
          2300 => x"ca",
          2301 => x"38",
          2302 => x"fe",
          2303 => x"39",
          2304 => x"16",
          2305 => x"ca",
          2306 => x"3d",
          2307 => x"3d",
          2308 => x"08",
          2309 => x"52",
          2310 => x"c5",
          2311 => x"88",
          2312 => x"ca",
          2313 => x"38",
          2314 => x"52",
          2315 => x"de",
          2316 => x"88",
          2317 => x"ca",
          2318 => x"38",
          2319 => x"ca",
          2320 => x"9c",
          2321 => x"ea",
          2322 => x"53",
          2323 => x"9c",
          2324 => x"ea",
          2325 => x"0b",
          2326 => x"74",
          2327 => x"0c",
          2328 => x"04",
          2329 => x"75",
          2330 => x"12",
          2331 => x"53",
          2332 => x"9a",
          2333 => x"88",
          2334 => x"9c",
          2335 => x"e5",
          2336 => x"0b",
          2337 => x"85",
          2338 => x"fa",
          2339 => x"7a",
          2340 => x"0b",
          2341 => x"98",
          2342 => x"2e",
          2343 => x"80",
          2344 => x"55",
          2345 => x"17",
          2346 => x"33",
          2347 => x"51",
          2348 => x"2e",
          2349 => x"85",
          2350 => x"06",
          2351 => x"e5",
          2352 => x"2e",
          2353 => x"8b",
          2354 => x"70",
          2355 => x"34",
          2356 => x"71",
          2357 => x"05",
          2358 => x"15",
          2359 => x"27",
          2360 => x"15",
          2361 => x"80",
          2362 => x"34",
          2363 => x"52",
          2364 => x"88",
          2365 => x"17",
          2366 => x"52",
          2367 => x"3f",
          2368 => x"08",
          2369 => x"12",
          2370 => x"3f",
          2371 => x"08",
          2372 => x"98",
          2373 => x"da",
          2374 => x"88",
          2375 => x"23",
          2376 => x"04",
          2377 => x"7f",
          2378 => x"5b",
          2379 => x"33",
          2380 => x"73",
          2381 => x"38",
          2382 => x"80",
          2383 => x"38",
          2384 => x"8c",
          2385 => x"08",
          2386 => x"aa",
          2387 => x"41",
          2388 => x"33",
          2389 => x"73",
          2390 => x"81",
          2391 => x"81",
          2392 => x"dc",
          2393 => x"70",
          2394 => x"07",
          2395 => x"73",
          2396 => x"88",
          2397 => x"70",
          2398 => x"73",
          2399 => x"38",
          2400 => x"ab",
          2401 => x"52",
          2402 => x"91",
          2403 => x"88",
          2404 => x"98",
          2405 => x"61",
          2406 => x"5a",
          2407 => x"a0",
          2408 => x"e7",
          2409 => x"70",
          2410 => x"79",
          2411 => x"73",
          2412 => x"81",
          2413 => x"38",
          2414 => x"33",
          2415 => x"ae",
          2416 => x"70",
          2417 => x"82",
          2418 => x"51",
          2419 => x"54",
          2420 => x"79",
          2421 => x"74",
          2422 => x"57",
          2423 => x"af",
          2424 => x"70",
          2425 => x"51",
          2426 => x"dc",
          2427 => x"73",
          2428 => x"38",
          2429 => x"82",
          2430 => x"19",
          2431 => x"54",
          2432 => x"82",
          2433 => x"54",
          2434 => x"78",
          2435 => x"81",
          2436 => x"54",
          2437 => x"81",
          2438 => x"af",
          2439 => x"77",
          2440 => x"70",
          2441 => x"25",
          2442 => x"07",
          2443 => x"51",
          2444 => x"2e",
          2445 => x"39",
          2446 => x"80",
          2447 => x"33",
          2448 => x"73",
          2449 => x"81",
          2450 => x"81",
          2451 => x"dc",
          2452 => x"70",
          2453 => x"07",
          2454 => x"73",
          2455 => x"b5",
          2456 => x"2e",
          2457 => x"83",
          2458 => x"76",
          2459 => x"07",
          2460 => x"2e",
          2461 => x"8b",
          2462 => x"77",
          2463 => x"30",
          2464 => x"71",
          2465 => x"53",
          2466 => x"55",
          2467 => x"38",
          2468 => x"5c",
          2469 => x"75",
          2470 => x"73",
          2471 => x"38",
          2472 => x"06",
          2473 => x"11",
          2474 => x"75",
          2475 => x"3f",
          2476 => x"08",
          2477 => x"38",
          2478 => x"33",
          2479 => x"54",
          2480 => x"e6",
          2481 => x"ca",
          2482 => x"2e",
          2483 => x"ff",
          2484 => x"74",
          2485 => x"38",
          2486 => x"75",
          2487 => x"17",
          2488 => x"57",
          2489 => x"a7",
          2490 => x"91",
          2491 => x"e5",
          2492 => x"ca",
          2493 => x"38",
          2494 => x"54",
          2495 => x"89",
          2496 => x"70",
          2497 => x"57",
          2498 => x"54",
          2499 => x"81",
          2500 => x"f7",
          2501 => x"7e",
          2502 => x"2e",
          2503 => x"33",
          2504 => x"e5",
          2505 => x"06",
          2506 => x"7a",
          2507 => x"a0",
          2508 => x"38",
          2509 => x"55",
          2510 => x"84",
          2511 => x"39",
          2512 => x"8b",
          2513 => x"7b",
          2514 => x"7a",
          2515 => x"3f",
          2516 => x"08",
          2517 => x"88",
          2518 => x"38",
          2519 => x"52",
          2520 => x"aa",
          2521 => x"88",
          2522 => x"ca",
          2523 => x"c2",
          2524 => x"08",
          2525 => x"55",
          2526 => x"ff",
          2527 => x"15",
          2528 => x"54",
          2529 => x"34",
          2530 => x"70",
          2531 => x"81",
          2532 => x"58",
          2533 => x"8b",
          2534 => x"74",
          2535 => x"3f",
          2536 => x"08",
          2537 => x"38",
          2538 => x"51",
          2539 => x"ff",
          2540 => x"ab",
          2541 => x"55",
          2542 => x"bb",
          2543 => x"2e",
          2544 => x"80",
          2545 => x"85",
          2546 => x"06",
          2547 => x"58",
          2548 => x"80",
          2549 => x"75",
          2550 => x"73",
          2551 => x"b5",
          2552 => x"0b",
          2553 => x"80",
          2554 => x"39",
          2555 => x"54",
          2556 => x"85",
          2557 => x"75",
          2558 => x"81",
          2559 => x"73",
          2560 => x"1b",
          2561 => x"2a",
          2562 => x"51",
          2563 => x"80",
          2564 => x"90",
          2565 => x"ff",
          2566 => x"05",
          2567 => x"f5",
          2568 => x"ca",
          2569 => x"1c",
          2570 => x"39",
          2571 => x"88",
          2572 => x"0d",
          2573 => x"0d",
          2574 => x"7b",
          2575 => x"73",
          2576 => x"55",
          2577 => x"2e",
          2578 => x"75",
          2579 => x"57",
          2580 => x"26",
          2581 => x"ba",
          2582 => x"70",
          2583 => x"ba",
          2584 => x"06",
          2585 => x"73",
          2586 => x"70",
          2587 => x"51",
          2588 => x"89",
          2589 => x"82",
          2590 => x"ff",
          2591 => x"56",
          2592 => x"2e",
          2593 => x"80",
          2594 => x"84",
          2595 => x"08",
          2596 => x"76",
          2597 => x"58",
          2598 => x"81",
          2599 => x"ff",
          2600 => x"53",
          2601 => x"26",
          2602 => x"13",
          2603 => x"06",
          2604 => x"9f",
          2605 => x"99",
          2606 => x"e0",
          2607 => x"ff",
          2608 => x"72",
          2609 => x"2a",
          2610 => x"72",
          2611 => x"06",
          2612 => x"ff",
          2613 => x"30",
          2614 => x"70",
          2615 => x"07",
          2616 => x"9f",
          2617 => x"54",
          2618 => x"80",
          2619 => x"81",
          2620 => x"59",
          2621 => x"25",
          2622 => x"8b",
          2623 => x"24",
          2624 => x"76",
          2625 => x"78",
          2626 => x"91",
          2627 => x"51",
          2628 => x"88",
          2629 => x"0d",
          2630 => x"0d",
          2631 => x"0b",
          2632 => x"ff",
          2633 => x"0c",
          2634 => x"51",
          2635 => x"84",
          2636 => x"88",
          2637 => x"38",
          2638 => x"51",
          2639 => x"91",
          2640 => x"83",
          2641 => x"54",
          2642 => x"82",
          2643 => x"09",
          2644 => x"e3",
          2645 => x"b4",
          2646 => x"57",
          2647 => x"2e",
          2648 => x"83",
          2649 => x"74",
          2650 => x"70",
          2651 => x"25",
          2652 => x"51",
          2653 => x"38",
          2654 => x"2e",
          2655 => x"b5",
          2656 => x"91",
          2657 => x"80",
          2658 => x"e0",
          2659 => x"ca",
          2660 => x"91",
          2661 => x"80",
          2662 => x"85",
          2663 => x"c8",
          2664 => x"16",
          2665 => x"3f",
          2666 => x"08",
          2667 => x"88",
          2668 => x"83",
          2669 => x"74",
          2670 => x"0c",
          2671 => x"04",
          2672 => x"61",
          2673 => x"80",
          2674 => x"58",
          2675 => x"0c",
          2676 => x"e1",
          2677 => x"88",
          2678 => x"56",
          2679 => x"ca",
          2680 => x"86",
          2681 => x"ca",
          2682 => x"29",
          2683 => x"05",
          2684 => x"53",
          2685 => x"80",
          2686 => x"38",
          2687 => x"76",
          2688 => x"74",
          2689 => x"72",
          2690 => x"38",
          2691 => x"51",
          2692 => x"91",
          2693 => x"81",
          2694 => x"81",
          2695 => x"72",
          2696 => x"80",
          2697 => x"38",
          2698 => x"70",
          2699 => x"53",
          2700 => x"86",
          2701 => x"a7",
          2702 => x"34",
          2703 => x"34",
          2704 => x"14",
          2705 => x"b2",
          2706 => x"88",
          2707 => x"06",
          2708 => x"54",
          2709 => x"72",
          2710 => x"76",
          2711 => x"38",
          2712 => x"70",
          2713 => x"53",
          2714 => x"85",
          2715 => x"70",
          2716 => x"5b",
          2717 => x"91",
          2718 => x"81",
          2719 => x"76",
          2720 => x"81",
          2721 => x"38",
          2722 => x"56",
          2723 => x"83",
          2724 => x"70",
          2725 => x"80",
          2726 => x"83",
          2727 => x"dc",
          2728 => x"ca",
          2729 => x"76",
          2730 => x"05",
          2731 => x"16",
          2732 => x"56",
          2733 => x"d7",
          2734 => x"8d",
          2735 => x"72",
          2736 => x"54",
          2737 => x"57",
          2738 => x"95",
          2739 => x"73",
          2740 => x"3f",
          2741 => x"08",
          2742 => x"57",
          2743 => x"89",
          2744 => x"56",
          2745 => x"d7",
          2746 => x"76",
          2747 => x"f1",
          2748 => x"76",
          2749 => x"e9",
          2750 => x"51",
          2751 => x"91",
          2752 => x"83",
          2753 => x"53",
          2754 => x"2e",
          2755 => x"84",
          2756 => x"ca",
          2757 => x"da",
          2758 => x"88",
          2759 => x"ff",
          2760 => x"8d",
          2761 => x"14",
          2762 => x"3f",
          2763 => x"08",
          2764 => x"15",
          2765 => x"14",
          2766 => x"34",
          2767 => x"33",
          2768 => x"81",
          2769 => x"54",
          2770 => x"72",
          2771 => x"91",
          2772 => x"ff",
          2773 => x"29",
          2774 => x"33",
          2775 => x"72",
          2776 => x"72",
          2777 => x"38",
          2778 => x"06",
          2779 => x"2e",
          2780 => x"56",
          2781 => x"80",
          2782 => x"da",
          2783 => x"ca",
          2784 => x"91",
          2785 => x"88",
          2786 => x"8f",
          2787 => x"56",
          2788 => x"38",
          2789 => x"51",
          2790 => x"91",
          2791 => x"83",
          2792 => x"55",
          2793 => x"80",
          2794 => x"da",
          2795 => x"ca",
          2796 => x"80",
          2797 => x"da",
          2798 => x"ca",
          2799 => x"ff",
          2800 => x"8d",
          2801 => x"2e",
          2802 => x"88",
          2803 => x"14",
          2804 => x"05",
          2805 => x"75",
          2806 => x"38",
          2807 => x"52",
          2808 => x"51",
          2809 => x"3f",
          2810 => x"08",
          2811 => x"88",
          2812 => x"82",
          2813 => x"ca",
          2814 => x"ff",
          2815 => x"26",
          2816 => x"57",
          2817 => x"f5",
          2818 => x"82",
          2819 => x"f5",
          2820 => x"81",
          2821 => x"8d",
          2822 => x"2e",
          2823 => x"82",
          2824 => x"16",
          2825 => x"16",
          2826 => x"70",
          2827 => x"7a",
          2828 => x"0c",
          2829 => x"83",
          2830 => x"06",
          2831 => x"de",
          2832 => x"ae",
          2833 => x"88",
          2834 => x"ff",
          2835 => x"56",
          2836 => x"38",
          2837 => x"38",
          2838 => x"51",
          2839 => x"91",
          2840 => x"a8",
          2841 => x"82",
          2842 => x"39",
          2843 => x"80",
          2844 => x"38",
          2845 => x"15",
          2846 => x"53",
          2847 => x"8d",
          2848 => x"15",
          2849 => x"76",
          2850 => x"51",
          2851 => x"13",
          2852 => x"8d",
          2853 => x"15",
          2854 => x"c5",
          2855 => x"90",
          2856 => x"0b",
          2857 => x"ff",
          2858 => x"15",
          2859 => x"2e",
          2860 => x"81",
          2861 => x"e4",
          2862 => x"b6",
          2863 => x"88",
          2864 => x"ff",
          2865 => x"81",
          2866 => x"06",
          2867 => x"81",
          2868 => x"51",
          2869 => x"91",
          2870 => x"80",
          2871 => x"ca",
          2872 => x"15",
          2873 => x"14",
          2874 => x"3f",
          2875 => x"08",
          2876 => x"06",
          2877 => x"d4",
          2878 => x"81",
          2879 => x"38",
          2880 => x"d8",
          2881 => x"ca",
          2882 => x"8b",
          2883 => x"2e",
          2884 => x"b3",
          2885 => x"14",
          2886 => x"3f",
          2887 => x"08",
          2888 => x"e4",
          2889 => x"81",
          2890 => x"84",
          2891 => x"d7",
          2892 => x"ca",
          2893 => x"15",
          2894 => x"14",
          2895 => x"3f",
          2896 => x"08",
          2897 => x"76",
          2898 => x"ca",
          2899 => x"05",
          2900 => x"ca",
          2901 => x"86",
          2902 => x"0b",
          2903 => x"80",
          2904 => x"ca",
          2905 => x"3d",
          2906 => x"3d",
          2907 => x"89",
          2908 => x"2e",
          2909 => x"08",
          2910 => x"2e",
          2911 => x"33",
          2912 => x"2e",
          2913 => x"13",
          2914 => x"22",
          2915 => x"76",
          2916 => x"06",
          2917 => x"13",
          2918 => x"c0",
          2919 => x"88",
          2920 => x"52",
          2921 => x"71",
          2922 => x"55",
          2923 => x"53",
          2924 => x"0c",
          2925 => x"ca",
          2926 => x"3d",
          2927 => x"3d",
          2928 => x"05",
          2929 => x"89",
          2930 => x"52",
          2931 => x"3f",
          2932 => x"0b",
          2933 => x"08",
          2934 => x"91",
          2935 => x"84",
          2936 => x"a4",
          2937 => x"55",
          2938 => x"2e",
          2939 => x"74",
          2940 => x"73",
          2941 => x"38",
          2942 => x"78",
          2943 => x"54",
          2944 => x"92",
          2945 => x"89",
          2946 => x"84",
          2947 => x"b0",
          2948 => x"88",
          2949 => x"91",
          2950 => x"88",
          2951 => x"eb",
          2952 => x"02",
          2953 => x"e7",
          2954 => x"59",
          2955 => x"80",
          2956 => x"38",
          2957 => x"70",
          2958 => x"d0",
          2959 => x"3d",
          2960 => x"58",
          2961 => x"91",
          2962 => x"55",
          2963 => x"08",
          2964 => x"7a",
          2965 => x"8c",
          2966 => x"56",
          2967 => x"91",
          2968 => x"55",
          2969 => x"08",
          2970 => x"80",
          2971 => x"70",
          2972 => x"57",
          2973 => x"83",
          2974 => x"77",
          2975 => x"73",
          2976 => x"ab",
          2977 => x"2e",
          2978 => x"84",
          2979 => x"06",
          2980 => x"51",
          2981 => x"91",
          2982 => x"55",
          2983 => x"b2",
          2984 => x"06",
          2985 => x"b8",
          2986 => x"2a",
          2987 => x"51",
          2988 => x"2e",
          2989 => x"55",
          2990 => x"77",
          2991 => x"74",
          2992 => x"77",
          2993 => x"81",
          2994 => x"73",
          2995 => x"af",
          2996 => x"7a",
          2997 => x"3f",
          2998 => x"08",
          2999 => x"b2",
          3000 => x"8e",
          3001 => x"ea",
          3002 => x"a0",
          3003 => x"34",
          3004 => x"52",
          3005 => x"bd",
          3006 => x"62",
          3007 => x"d4",
          3008 => x"54",
          3009 => x"15",
          3010 => x"2e",
          3011 => x"7a",
          3012 => x"51",
          3013 => x"75",
          3014 => x"d4",
          3015 => x"be",
          3016 => x"88",
          3017 => x"ca",
          3018 => x"ca",
          3019 => x"74",
          3020 => x"02",
          3021 => x"70",
          3022 => x"81",
          3023 => x"56",
          3024 => x"86",
          3025 => x"82",
          3026 => x"81",
          3027 => x"06",
          3028 => x"80",
          3029 => x"75",
          3030 => x"73",
          3031 => x"38",
          3032 => x"92",
          3033 => x"7a",
          3034 => x"3f",
          3035 => x"08",
          3036 => x"8c",
          3037 => x"55",
          3038 => x"08",
          3039 => x"77",
          3040 => x"81",
          3041 => x"73",
          3042 => x"38",
          3043 => x"07",
          3044 => x"11",
          3045 => x"0c",
          3046 => x"0c",
          3047 => x"52",
          3048 => x"3f",
          3049 => x"08",
          3050 => x"08",
          3051 => x"63",
          3052 => x"5a",
          3053 => x"91",
          3054 => x"91",
          3055 => x"8c",
          3056 => x"7a",
          3057 => x"17",
          3058 => x"23",
          3059 => x"34",
          3060 => x"1a",
          3061 => x"9c",
          3062 => x"0b",
          3063 => x"77",
          3064 => x"81",
          3065 => x"73",
          3066 => x"8d",
          3067 => x"88",
          3068 => x"81",
          3069 => x"ca",
          3070 => x"1a",
          3071 => x"22",
          3072 => x"7b",
          3073 => x"a8",
          3074 => x"78",
          3075 => x"3f",
          3076 => x"08",
          3077 => x"88",
          3078 => x"83",
          3079 => x"91",
          3080 => x"ff",
          3081 => x"06",
          3082 => x"55",
          3083 => x"56",
          3084 => x"76",
          3085 => x"51",
          3086 => x"27",
          3087 => x"70",
          3088 => x"5a",
          3089 => x"76",
          3090 => x"74",
          3091 => x"83",
          3092 => x"73",
          3093 => x"38",
          3094 => x"51",
          3095 => x"91",
          3096 => x"85",
          3097 => x"8e",
          3098 => x"2a",
          3099 => x"08",
          3100 => x"0c",
          3101 => x"79",
          3102 => x"73",
          3103 => x"0c",
          3104 => x"04",
          3105 => x"60",
          3106 => x"40",
          3107 => x"80",
          3108 => x"3d",
          3109 => x"78",
          3110 => x"3f",
          3111 => x"08",
          3112 => x"88",
          3113 => x"91",
          3114 => x"74",
          3115 => x"38",
          3116 => x"c4",
          3117 => x"33",
          3118 => x"87",
          3119 => x"2e",
          3120 => x"95",
          3121 => x"91",
          3122 => x"56",
          3123 => x"81",
          3124 => x"34",
          3125 => x"a0",
          3126 => x"08",
          3127 => x"31",
          3128 => x"27",
          3129 => x"5c",
          3130 => x"82",
          3131 => x"19",
          3132 => x"ff",
          3133 => x"74",
          3134 => x"7e",
          3135 => x"ff",
          3136 => x"2a",
          3137 => x"79",
          3138 => x"87",
          3139 => x"08",
          3140 => x"98",
          3141 => x"78",
          3142 => x"3f",
          3143 => x"08",
          3144 => x"27",
          3145 => x"74",
          3146 => x"a3",
          3147 => x"1a",
          3148 => x"08",
          3149 => x"d4",
          3150 => x"ca",
          3151 => x"2e",
          3152 => x"91",
          3153 => x"1a",
          3154 => x"59",
          3155 => x"2e",
          3156 => x"77",
          3157 => x"11",
          3158 => x"55",
          3159 => x"85",
          3160 => x"31",
          3161 => x"76",
          3162 => x"81",
          3163 => x"ca",
          3164 => x"ca",
          3165 => x"d7",
          3166 => x"11",
          3167 => x"74",
          3168 => x"38",
          3169 => x"77",
          3170 => x"78",
          3171 => x"84",
          3172 => x"16",
          3173 => x"08",
          3174 => x"2b",
          3175 => x"cf",
          3176 => x"89",
          3177 => x"39",
          3178 => x"0c",
          3179 => x"83",
          3180 => x"80",
          3181 => x"55",
          3182 => x"83",
          3183 => x"9c",
          3184 => x"7e",
          3185 => x"3f",
          3186 => x"08",
          3187 => x"75",
          3188 => x"08",
          3189 => x"1f",
          3190 => x"7c",
          3191 => x"3f",
          3192 => x"7e",
          3193 => x"0c",
          3194 => x"1b",
          3195 => x"1c",
          3196 => x"fd",
          3197 => x"56",
          3198 => x"88",
          3199 => x"0d",
          3200 => x"0d",
          3201 => x"64",
          3202 => x"58",
          3203 => x"90",
          3204 => x"52",
          3205 => x"d2",
          3206 => x"88",
          3207 => x"ca",
          3208 => x"38",
          3209 => x"55",
          3210 => x"86",
          3211 => x"83",
          3212 => x"18",
          3213 => x"2a",
          3214 => x"51",
          3215 => x"56",
          3216 => x"83",
          3217 => x"39",
          3218 => x"19",
          3219 => x"83",
          3220 => x"0b",
          3221 => x"81",
          3222 => x"39",
          3223 => x"7c",
          3224 => x"74",
          3225 => x"38",
          3226 => x"7b",
          3227 => x"ec",
          3228 => x"08",
          3229 => x"06",
          3230 => x"81",
          3231 => x"8a",
          3232 => x"05",
          3233 => x"06",
          3234 => x"bf",
          3235 => x"38",
          3236 => x"55",
          3237 => x"7a",
          3238 => x"98",
          3239 => x"77",
          3240 => x"3f",
          3241 => x"08",
          3242 => x"88",
          3243 => x"82",
          3244 => x"81",
          3245 => x"38",
          3246 => x"ff",
          3247 => x"98",
          3248 => x"18",
          3249 => x"74",
          3250 => x"7e",
          3251 => x"08",
          3252 => x"2e",
          3253 => x"8d",
          3254 => x"ce",
          3255 => x"ca",
          3256 => x"ee",
          3257 => x"08",
          3258 => x"d1",
          3259 => x"ca",
          3260 => x"2e",
          3261 => x"91",
          3262 => x"1b",
          3263 => x"5a",
          3264 => x"2e",
          3265 => x"78",
          3266 => x"11",
          3267 => x"55",
          3268 => x"85",
          3269 => x"31",
          3270 => x"76",
          3271 => x"81",
          3272 => x"c8",
          3273 => x"ca",
          3274 => x"a6",
          3275 => x"11",
          3276 => x"56",
          3277 => x"27",
          3278 => x"80",
          3279 => x"08",
          3280 => x"2b",
          3281 => x"b4",
          3282 => x"b5",
          3283 => x"80",
          3284 => x"34",
          3285 => x"56",
          3286 => x"8c",
          3287 => x"19",
          3288 => x"38",
          3289 => x"b6",
          3290 => x"88",
          3291 => x"38",
          3292 => x"12",
          3293 => x"9c",
          3294 => x"18",
          3295 => x"06",
          3296 => x"31",
          3297 => x"76",
          3298 => x"7b",
          3299 => x"08",
          3300 => x"cd",
          3301 => x"ca",
          3302 => x"b6",
          3303 => x"7c",
          3304 => x"08",
          3305 => x"1f",
          3306 => x"cb",
          3307 => x"55",
          3308 => x"16",
          3309 => x"31",
          3310 => x"7f",
          3311 => x"94",
          3312 => x"70",
          3313 => x"8c",
          3314 => x"58",
          3315 => x"76",
          3316 => x"75",
          3317 => x"19",
          3318 => x"39",
          3319 => x"80",
          3320 => x"74",
          3321 => x"80",
          3322 => x"ca",
          3323 => x"3d",
          3324 => x"3d",
          3325 => x"3d",
          3326 => x"70",
          3327 => x"ea",
          3328 => x"88",
          3329 => x"ca",
          3330 => x"fb",
          3331 => x"33",
          3332 => x"70",
          3333 => x"55",
          3334 => x"2e",
          3335 => x"a0",
          3336 => x"78",
          3337 => x"3f",
          3338 => x"08",
          3339 => x"88",
          3340 => x"38",
          3341 => x"8b",
          3342 => x"07",
          3343 => x"8b",
          3344 => x"16",
          3345 => x"52",
          3346 => x"dd",
          3347 => x"16",
          3348 => x"15",
          3349 => x"3f",
          3350 => x"0a",
          3351 => x"51",
          3352 => x"76",
          3353 => x"51",
          3354 => x"78",
          3355 => x"83",
          3356 => x"51",
          3357 => x"91",
          3358 => x"90",
          3359 => x"bf",
          3360 => x"73",
          3361 => x"76",
          3362 => x"0c",
          3363 => x"04",
          3364 => x"76",
          3365 => x"fe",
          3366 => x"ca",
          3367 => x"91",
          3368 => x"9c",
          3369 => x"fc",
          3370 => x"51",
          3371 => x"91",
          3372 => x"53",
          3373 => x"08",
          3374 => x"ca",
          3375 => x"0c",
          3376 => x"88",
          3377 => x"0d",
          3378 => x"0d",
          3379 => x"e6",
          3380 => x"52",
          3381 => x"ca",
          3382 => x"8b",
          3383 => x"88",
          3384 => x"b8",
          3385 => x"71",
          3386 => x"0c",
          3387 => x"04",
          3388 => x"80",
          3389 => x"d0",
          3390 => x"3d",
          3391 => x"3f",
          3392 => x"08",
          3393 => x"88",
          3394 => x"38",
          3395 => x"52",
          3396 => x"05",
          3397 => x"3f",
          3398 => x"08",
          3399 => x"88",
          3400 => x"02",
          3401 => x"33",
          3402 => x"55",
          3403 => x"25",
          3404 => x"7a",
          3405 => x"54",
          3406 => x"a2",
          3407 => x"84",
          3408 => x"06",
          3409 => x"73",
          3410 => x"38",
          3411 => x"70",
          3412 => x"a8",
          3413 => x"88",
          3414 => x"0c",
          3415 => x"ca",
          3416 => x"2e",
          3417 => x"83",
          3418 => x"74",
          3419 => x"0c",
          3420 => x"04",
          3421 => x"6f",
          3422 => x"80",
          3423 => x"53",
          3424 => x"b8",
          3425 => x"3d",
          3426 => x"3f",
          3427 => x"08",
          3428 => x"88",
          3429 => x"38",
          3430 => x"7c",
          3431 => x"47",
          3432 => x"54",
          3433 => x"81",
          3434 => x"52",
          3435 => x"52",
          3436 => x"3f",
          3437 => x"08",
          3438 => x"88",
          3439 => x"38",
          3440 => x"51",
          3441 => x"91",
          3442 => x"57",
          3443 => x"08",
          3444 => x"69",
          3445 => x"da",
          3446 => x"ca",
          3447 => x"76",
          3448 => x"d5",
          3449 => x"ca",
          3450 => x"91",
          3451 => x"82",
          3452 => x"52",
          3453 => x"eb",
          3454 => x"88",
          3455 => x"ca",
          3456 => x"38",
          3457 => x"51",
          3458 => x"73",
          3459 => x"08",
          3460 => x"76",
          3461 => x"d6",
          3462 => x"ca",
          3463 => x"91",
          3464 => x"80",
          3465 => x"76",
          3466 => x"81",
          3467 => x"82",
          3468 => x"39",
          3469 => x"38",
          3470 => x"bc",
          3471 => x"51",
          3472 => x"76",
          3473 => x"11",
          3474 => x"51",
          3475 => x"73",
          3476 => x"38",
          3477 => x"55",
          3478 => x"16",
          3479 => x"56",
          3480 => x"38",
          3481 => x"73",
          3482 => x"90",
          3483 => x"2e",
          3484 => x"16",
          3485 => x"ff",
          3486 => x"ff",
          3487 => x"58",
          3488 => x"74",
          3489 => x"75",
          3490 => x"18",
          3491 => x"58",
          3492 => x"fe",
          3493 => x"7b",
          3494 => x"06",
          3495 => x"18",
          3496 => x"58",
          3497 => x"80",
          3498 => x"b8",
          3499 => x"29",
          3500 => x"05",
          3501 => x"33",
          3502 => x"56",
          3503 => x"2e",
          3504 => x"16",
          3505 => x"33",
          3506 => x"73",
          3507 => x"16",
          3508 => x"26",
          3509 => x"55",
          3510 => x"91",
          3511 => x"54",
          3512 => x"70",
          3513 => x"34",
          3514 => x"ec",
          3515 => x"70",
          3516 => x"34",
          3517 => x"09",
          3518 => x"38",
          3519 => x"39",
          3520 => x"19",
          3521 => x"33",
          3522 => x"05",
          3523 => x"78",
          3524 => x"80",
          3525 => x"91",
          3526 => x"9e",
          3527 => x"f7",
          3528 => x"7d",
          3529 => x"05",
          3530 => x"57",
          3531 => x"3f",
          3532 => x"08",
          3533 => x"88",
          3534 => x"38",
          3535 => x"53",
          3536 => x"38",
          3537 => x"54",
          3538 => x"92",
          3539 => x"33",
          3540 => x"70",
          3541 => x"54",
          3542 => x"38",
          3543 => x"15",
          3544 => x"70",
          3545 => x"58",
          3546 => x"82",
          3547 => x"8a",
          3548 => x"89",
          3549 => x"53",
          3550 => x"b7",
          3551 => x"ff",
          3552 => x"9b",
          3553 => x"ca",
          3554 => x"15",
          3555 => x"53",
          3556 => x"9b",
          3557 => x"ca",
          3558 => x"26",
          3559 => x"30",
          3560 => x"70",
          3561 => x"77",
          3562 => x"18",
          3563 => x"51",
          3564 => x"88",
          3565 => x"73",
          3566 => x"52",
          3567 => x"ca",
          3568 => x"88",
          3569 => x"ca",
          3570 => x"2e",
          3571 => x"91",
          3572 => x"ff",
          3573 => x"38",
          3574 => x"08",
          3575 => x"73",
          3576 => x"73",
          3577 => x"9c",
          3578 => x"27",
          3579 => x"75",
          3580 => x"16",
          3581 => x"17",
          3582 => x"33",
          3583 => x"70",
          3584 => x"55",
          3585 => x"80",
          3586 => x"73",
          3587 => x"cc",
          3588 => x"ca",
          3589 => x"91",
          3590 => x"94",
          3591 => x"88",
          3592 => x"39",
          3593 => x"51",
          3594 => x"91",
          3595 => x"54",
          3596 => x"be",
          3597 => x"27",
          3598 => x"53",
          3599 => x"08",
          3600 => x"73",
          3601 => x"ff",
          3602 => x"15",
          3603 => x"16",
          3604 => x"ff",
          3605 => x"80",
          3606 => x"73",
          3607 => x"c6",
          3608 => x"ca",
          3609 => x"38",
          3610 => x"16",
          3611 => x"80",
          3612 => x"0b",
          3613 => x"81",
          3614 => x"75",
          3615 => x"ca",
          3616 => x"58",
          3617 => x"54",
          3618 => x"74",
          3619 => x"73",
          3620 => x"90",
          3621 => x"c0",
          3622 => x"90",
          3623 => x"83",
          3624 => x"72",
          3625 => x"38",
          3626 => x"08",
          3627 => x"77",
          3628 => x"80",
          3629 => x"ca",
          3630 => x"3d",
          3631 => x"3d",
          3632 => x"89",
          3633 => x"2e",
          3634 => x"80",
          3635 => x"fc",
          3636 => x"3d",
          3637 => x"e1",
          3638 => x"ca",
          3639 => x"91",
          3640 => x"80",
          3641 => x"76",
          3642 => x"75",
          3643 => x"3f",
          3644 => x"08",
          3645 => x"88",
          3646 => x"38",
          3647 => x"70",
          3648 => x"57",
          3649 => x"a2",
          3650 => x"33",
          3651 => x"70",
          3652 => x"55",
          3653 => x"2e",
          3654 => x"16",
          3655 => x"51",
          3656 => x"91",
          3657 => x"88",
          3658 => x"54",
          3659 => x"84",
          3660 => x"52",
          3661 => x"e5",
          3662 => x"88",
          3663 => x"84",
          3664 => x"06",
          3665 => x"55",
          3666 => x"80",
          3667 => x"80",
          3668 => x"54",
          3669 => x"88",
          3670 => x"0d",
          3671 => x"0d",
          3672 => x"fc",
          3673 => x"52",
          3674 => x"3f",
          3675 => x"08",
          3676 => x"ca",
          3677 => x"0c",
          3678 => x"04",
          3679 => x"77",
          3680 => x"fc",
          3681 => x"53",
          3682 => x"de",
          3683 => x"88",
          3684 => x"ca",
          3685 => x"df",
          3686 => x"38",
          3687 => x"08",
          3688 => x"cd",
          3689 => x"ca",
          3690 => x"80",
          3691 => x"ca",
          3692 => x"73",
          3693 => x"3f",
          3694 => x"08",
          3695 => x"88",
          3696 => x"09",
          3697 => x"38",
          3698 => x"39",
          3699 => x"08",
          3700 => x"52",
          3701 => x"b3",
          3702 => x"73",
          3703 => x"3f",
          3704 => x"08",
          3705 => x"30",
          3706 => x"9f",
          3707 => x"ca",
          3708 => x"51",
          3709 => x"72",
          3710 => x"0c",
          3711 => x"04",
          3712 => x"65",
          3713 => x"89",
          3714 => x"96",
          3715 => x"df",
          3716 => x"ca",
          3717 => x"91",
          3718 => x"b2",
          3719 => x"75",
          3720 => x"3f",
          3721 => x"08",
          3722 => x"88",
          3723 => x"02",
          3724 => x"33",
          3725 => x"55",
          3726 => x"25",
          3727 => x"55",
          3728 => x"80",
          3729 => x"76",
          3730 => x"d4",
          3731 => x"91",
          3732 => x"94",
          3733 => x"f0",
          3734 => x"65",
          3735 => x"53",
          3736 => x"05",
          3737 => x"51",
          3738 => x"91",
          3739 => x"5b",
          3740 => x"08",
          3741 => x"7c",
          3742 => x"08",
          3743 => x"fe",
          3744 => x"08",
          3745 => x"55",
          3746 => x"91",
          3747 => x"0c",
          3748 => x"81",
          3749 => x"39",
          3750 => x"c7",
          3751 => x"88",
          3752 => x"55",
          3753 => x"2e",
          3754 => x"bf",
          3755 => x"5f",
          3756 => x"92",
          3757 => x"51",
          3758 => x"91",
          3759 => x"ff",
          3760 => x"91",
          3761 => x"81",
          3762 => x"91",
          3763 => x"30",
          3764 => x"88",
          3765 => x"25",
          3766 => x"19",
          3767 => x"5a",
          3768 => x"08",
          3769 => x"38",
          3770 => x"a4",
          3771 => x"ca",
          3772 => x"58",
          3773 => x"77",
          3774 => x"7d",
          3775 => x"bf",
          3776 => x"ca",
          3777 => x"91",
          3778 => x"80",
          3779 => x"70",
          3780 => x"ff",
          3781 => x"56",
          3782 => x"2e",
          3783 => x"9e",
          3784 => x"51",
          3785 => x"3f",
          3786 => x"08",
          3787 => x"06",
          3788 => x"80",
          3789 => x"19",
          3790 => x"54",
          3791 => x"14",
          3792 => x"c5",
          3793 => x"88",
          3794 => x"06",
          3795 => x"80",
          3796 => x"19",
          3797 => x"54",
          3798 => x"06",
          3799 => x"79",
          3800 => x"78",
          3801 => x"79",
          3802 => x"84",
          3803 => x"07",
          3804 => x"84",
          3805 => x"91",
          3806 => x"92",
          3807 => x"f9",
          3808 => x"8a",
          3809 => x"53",
          3810 => x"e3",
          3811 => x"ca",
          3812 => x"91",
          3813 => x"81",
          3814 => x"17",
          3815 => x"81",
          3816 => x"17",
          3817 => x"2a",
          3818 => x"51",
          3819 => x"55",
          3820 => x"81",
          3821 => x"17",
          3822 => x"8c",
          3823 => x"81",
          3824 => x"9b",
          3825 => x"88",
          3826 => x"17",
          3827 => x"51",
          3828 => x"91",
          3829 => x"74",
          3830 => x"56",
          3831 => x"98",
          3832 => x"76",
          3833 => x"c6",
          3834 => x"88",
          3835 => x"09",
          3836 => x"38",
          3837 => x"ca",
          3838 => x"2e",
          3839 => x"85",
          3840 => x"a3",
          3841 => x"38",
          3842 => x"ca",
          3843 => x"15",
          3844 => x"38",
          3845 => x"53",
          3846 => x"08",
          3847 => x"c3",
          3848 => x"ca",
          3849 => x"94",
          3850 => x"18",
          3851 => x"33",
          3852 => x"54",
          3853 => x"34",
          3854 => x"85",
          3855 => x"18",
          3856 => x"74",
          3857 => x"0c",
          3858 => x"04",
          3859 => x"82",
          3860 => x"ff",
          3861 => x"a1",
          3862 => x"e4",
          3863 => x"88",
          3864 => x"ca",
          3865 => x"f5",
          3866 => x"a1",
          3867 => x"95",
          3868 => x"58",
          3869 => x"91",
          3870 => x"55",
          3871 => x"08",
          3872 => x"02",
          3873 => x"33",
          3874 => x"70",
          3875 => x"55",
          3876 => x"73",
          3877 => x"75",
          3878 => x"80",
          3879 => x"bd",
          3880 => x"d6",
          3881 => x"81",
          3882 => x"87",
          3883 => x"ad",
          3884 => x"78",
          3885 => x"3f",
          3886 => x"08",
          3887 => x"70",
          3888 => x"55",
          3889 => x"2e",
          3890 => x"78",
          3891 => x"88",
          3892 => x"08",
          3893 => x"38",
          3894 => x"ca",
          3895 => x"76",
          3896 => x"70",
          3897 => x"b5",
          3898 => x"88",
          3899 => x"ca",
          3900 => x"e9",
          3901 => x"88",
          3902 => x"51",
          3903 => x"91",
          3904 => x"55",
          3905 => x"08",
          3906 => x"55",
          3907 => x"91",
          3908 => x"84",
          3909 => x"91",
          3910 => x"80",
          3911 => x"51",
          3912 => x"91",
          3913 => x"91",
          3914 => x"30",
          3915 => x"88",
          3916 => x"25",
          3917 => x"75",
          3918 => x"38",
          3919 => x"8f",
          3920 => x"75",
          3921 => x"c1",
          3922 => x"ca",
          3923 => x"74",
          3924 => x"51",
          3925 => x"3f",
          3926 => x"08",
          3927 => x"ca",
          3928 => x"3d",
          3929 => x"3d",
          3930 => x"99",
          3931 => x"52",
          3932 => x"d8",
          3933 => x"ca",
          3934 => x"91",
          3935 => x"82",
          3936 => x"5e",
          3937 => x"3d",
          3938 => x"cf",
          3939 => x"ca",
          3940 => x"91",
          3941 => x"86",
          3942 => x"82",
          3943 => x"ca",
          3944 => x"2e",
          3945 => x"82",
          3946 => x"80",
          3947 => x"70",
          3948 => x"06",
          3949 => x"54",
          3950 => x"38",
          3951 => x"52",
          3952 => x"52",
          3953 => x"3f",
          3954 => x"08",
          3955 => x"91",
          3956 => x"83",
          3957 => x"91",
          3958 => x"81",
          3959 => x"06",
          3960 => x"54",
          3961 => x"08",
          3962 => x"81",
          3963 => x"81",
          3964 => x"39",
          3965 => x"38",
          3966 => x"08",
          3967 => x"c4",
          3968 => x"ca",
          3969 => x"91",
          3970 => x"81",
          3971 => x"53",
          3972 => x"19",
          3973 => x"8c",
          3974 => x"ae",
          3975 => x"34",
          3976 => x"0b",
          3977 => x"82",
          3978 => x"52",
          3979 => x"51",
          3980 => x"3f",
          3981 => x"b4",
          3982 => x"c9",
          3983 => x"53",
          3984 => x"53",
          3985 => x"51",
          3986 => x"3f",
          3987 => x"0b",
          3988 => x"34",
          3989 => x"80",
          3990 => x"51",
          3991 => x"78",
          3992 => x"83",
          3993 => x"51",
          3994 => x"91",
          3995 => x"54",
          3996 => x"08",
          3997 => x"88",
          3998 => x"64",
          3999 => x"ff",
          4000 => x"75",
          4001 => x"78",
          4002 => x"3f",
          4003 => x"0b",
          4004 => x"78",
          4005 => x"83",
          4006 => x"51",
          4007 => x"3f",
          4008 => x"08",
          4009 => x"80",
          4010 => x"76",
          4011 => x"ae",
          4012 => x"ca",
          4013 => x"3d",
          4014 => x"3d",
          4015 => x"84",
          4016 => x"f1",
          4017 => x"a8",
          4018 => x"05",
          4019 => x"51",
          4020 => x"91",
          4021 => x"55",
          4022 => x"08",
          4023 => x"78",
          4024 => x"08",
          4025 => x"70",
          4026 => x"b8",
          4027 => x"88",
          4028 => x"ca",
          4029 => x"b9",
          4030 => x"9b",
          4031 => x"a0",
          4032 => x"55",
          4033 => x"38",
          4034 => x"3d",
          4035 => x"3d",
          4036 => x"51",
          4037 => x"3f",
          4038 => x"52",
          4039 => x"52",
          4040 => x"dd",
          4041 => x"08",
          4042 => x"cb",
          4043 => x"ca",
          4044 => x"91",
          4045 => x"95",
          4046 => x"2e",
          4047 => x"88",
          4048 => x"3d",
          4049 => x"38",
          4050 => x"e5",
          4051 => x"88",
          4052 => x"09",
          4053 => x"b8",
          4054 => x"c9",
          4055 => x"ca",
          4056 => x"91",
          4057 => x"81",
          4058 => x"56",
          4059 => x"3d",
          4060 => x"52",
          4061 => x"ff",
          4062 => x"02",
          4063 => x"8b",
          4064 => x"16",
          4065 => x"2a",
          4066 => x"51",
          4067 => x"89",
          4068 => x"07",
          4069 => x"17",
          4070 => x"81",
          4071 => x"34",
          4072 => x"70",
          4073 => x"81",
          4074 => x"55",
          4075 => x"80",
          4076 => x"64",
          4077 => x"38",
          4078 => x"51",
          4079 => x"91",
          4080 => x"52",
          4081 => x"b7",
          4082 => x"55",
          4083 => x"08",
          4084 => x"dd",
          4085 => x"88",
          4086 => x"51",
          4087 => x"3f",
          4088 => x"08",
          4089 => x"11",
          4090 => x"91",
          4091 => x"80",
          4092 => x"16",
          4093 => x"ae",
          4094 => x"06",
          4095 => x"53",
          4096 => x"51",
          4097 => x"78",
          4098 => x"83",
          4099 => x"39",
          4100 => x"08",
          4101 => x"51",
          4102 => x"91",
          4103 => x"55",
          4104 => x"08",
          4105 => x"51",
          4106 => x"3f",
          4107 => x"08",
          4108 => x"ca",
          4109 => x"3d",
          4110 => x"3d",
          4111 => x"db",
          4112 => x"84",
          4113 => x"05",
          4114 => x"82",
          4115 => x"d0",
          4116 => x"3d",
          4117 => x"3f",
          4118 => x"08",
          4119 => x"88",
          4120 => x"38",
          4121 => x"52",
          4122 => x"05",
          4123 => x"3f",
          4124 => x"08",
          4125 => x"88",
          4126 => x"02",
          4127 => x"33",
          4128 => x"54",
          4129 => x"aa",
          4130 => x"06",
          4131 => x"8b",
          4132 => x"06",
          4133 => x"07",
          4134 => x"56",
          4135 => x"34",
          4136 => x"0b",
          4137 => x"78",
          4138 => x"a9",
          4139 => x"88",
          4140 => x"91",
          4141 => x"95",
          4142 => x"ef",
          4143 => x"56",
          4144 => x"3d",
          4145 => x"94",
          4146 => x"f4",
          4147 => x"88",
          4148 => x"ca",
          4149 => x"cb",
          4150 => x"63",
          4151 => x"d4",
          4152 => x"c0",
          4153 => x"88",
          4154 => x"ca",
          4155 => x"38",
          4156 => x"05",
          4157 => x"06",
          4158 => x"73",
          4159 => x"16",
          4160 => x"22",
          4161 => x"07",
          4162 => x"1f",
          4163 => x"c2",
          4164 => x"81",
          4165 => x"34",
          4166 => x"b3",
          4167 => x"ca",
          4168 => x"74",
          4169 => x"0c",
          4170 => x"04",
          4171 => x"69",
          4172 => x"80",
          4173 => x"d0",
          4174 => x"3d",
          4175 => x"3f",
          4176 => x"08",
          4177 => x"08",
          4178 => x"ca",
          4179 => x"80",
          4180 => x"57",
          4181 => x"81",
          4182 => x"70",
          4183 => x"55",
          4184 => x"80",
          4185 => x"5d",
          4186 => x"52",
          4187 => x"52",
          4188 => x"a9",
          4189 => x"88",
          4190 => x"ca",
          4191 => x"d1",
          4192 => x"73",
          4193 => x"3f",
          4194 => x"08",
          4195 => x"88",
          4196 => x"91",
          4197 => x"91",
          4198 => x"65",
          4199 => x"78",
          4200 => x"7b",
          4201 => x"55",
          4202 => x"34",
          4203 => x"8a",
          4204 => x"38",
          4205 => x"1a",
          4206 => x"34",
          4207 => x"9e",
          4208 => x"70",
          4209 => x"51",
          4210 => x"a0",
          4211 => x"8e",
          4212 => x"2e",
          4213 => x"86",
          4214 => x"34",
          4215 => x"30",
          4216 => x"80",
          4217 => x"7a",
          4218 => x"c1",
          4219 => x"2e",
          4220 => x"a0",
          4221 => x"51",
          4222 => x"3f",
          4223 => x"08",
          4224 => x"88",
          4225 => x"7b",
          4226 => x"55",
          4227 => x"73",
          4228 => x"38",
          4229 => x"73",
          4230 => x"38",
          4231 => x"15",
          4232 => x"ff",
          4233 => x"91",
          4234 => x"7b",
          4235 => x"ca",
          4236 => x"3d",
          4237 => x"3d",
          4238 => x"9c",
          4239 => x"05",
          4240 => x"51",
          4241 => x"91",
          4242 => x"91",
          4243 => x"56",
          4244 => x"88",
          4245 => x"38",
          4246 => x"52",
          4247 => x"52",
          4248 => x"c0",
          4249 => x"70",
          4250 => x"ff",
          4251 => x"55",
          4252 => x"27",
          4253 => x"78",
          4254 => x"ff",
          4255 => x"05",
          4256 => x"55",
          4257 => x"3f",
          4258 => x"08",
          4259 => x"38",
          4260 => x"70",
          4261 => x"ff",
          4262 => x"91",
          4263 => x"80",
          4264 => x"74",
          4265 => x"07",
          4266 => x"4e",
          4267 => x"91",
          4268 => x"55",
          4269 => x"70",
          4270 => x"06",
          4271 => x"99",
          4272 => x"e0",
          4273 => x"ff",
          4274 => x"54",
          4275 => x"27",
          4276 => x"b8",
          4277 => x"55",
          4278 => x"a3",
          4279 => x"91",
          4280 => x"ff",
          4281 => x"91",
          4282 => x"93",
          4283 => x"75",
          4284 => x"76",
          4285 => x"38",
          4286 => x"77",
          4287 => x"86",
          4288 => x"39",
          4289 => x"27",
          4290 => x"88",
          4291 => x"78",
          4292 => x"5a",
          4293 => x"57",
          4294 => x"81",
          4295 => x"81",
          4296 => x"33",
          4297 => x"06",
          4298 => x"57",
          4299 => x"fe",
          4300 => x"3d",
          4301 => x"55",
          4302 => x"2e",
          4303 => x"76",
          4304 => x"38",
          4305 => x"55",
          4306 => x"33",
          4307 => x"a0",
          4308 => x"06",
          4309 => x"17",
          4310 => x"38",
          4311 => x"43",
          4312 => x"3d",
          4313 => x"ff",
          4314 => x"91",
          4315 => x"54",
          4316 => x"08",
          4317 => x"81",
          4318 => x"ff",
          4319 => x"91",
          4320 => x"54",
          4321 => x"08",
          4322 => x"80",
          4323 => x"54",
          4324 => x"80",
          4325 => x"ca",
          4326 => x"2e",
          4327 => x"80",
          4328 => x"54",
          4329 => x"80",
          4330 => x"52",
          4331 => x"bd",
          4332 => x"ca",
          4333 => x"91",
          4334 => x"b1",
          4335 => x"91",
          4336 => x"52",
          4337 => x"ab",
          4338 => x"54",
          4339 => x"15",
          4340 => x"78",
          4341 => x"ff",
          4342 => x"79",
          4343 => x"83",
          4344 => x"51",
          4345 => x"3f",
          4346 => x"08",
          4347 => x"74",
          4348 => x"0c",
          4349 => x"04",
          4350 => x"60",
          4351 => x"05",
          4352 => x"33",
          4353 => x"05",
          4354 => x"40",
          4355 => x"da",
          4356 => x"88",
          4357 => x"ca",
          4358 => x"bd",
          4359 => x"33",
          4360 => x"b5",
          4361 => x"2e",
          4362 => x"1a",
          4363 => x"90",
          4364 => x"33",
          4365 => x"70",
          4366 => x"55",
          4367 => x"38",
          4368 => x"97",
          4369 => x"82",
          4370 => x"58",
          4371 => x"7e",
          4372 => x"70",
          4373 => x"55",
          4374 => x"56",
          4375 => x"8a",
          4376 => x"7d",
          4377 => x"70",
          4378 => x"2a",
          4379 => x"08",
          4380 => x"08",
          4381 => x"5d",
          4382 => x"77",
          4383 => x"98",
          4384 => x"26",
          4385 => x"57",
          4386 => x"59",
          4387 => x"52",
          4388 => x"ae",
          4389 => x"15",
          4390 => x"98",
          4391 => x"26",
          4392 => x"55",
          4393 => x"08",
          4394 => x"99",
          4395 => x"88",
          4396 => x"ff",
          4397 => x"ca",
          4398 => x"38",
          4399 => x"75",
          4400 => x"81",
          4401 => x"93",
          4402 => x"80",
          4403 => x"2e",
          4404 => x"ff",
          4405 => x"58",
          4406 => x"7d",
          4407 => x"38",
          4408 => x"55",
          4409 => x"b4",
          4410 => x"56",
          4411 => x"09",
          4412 => x"38",
          4413 => x"53",
          4414 => x"51",
          4415 => x"3f",
          4416 => x"08",
          4417 => x"88",
          4418 => x"38",
          4419 => x"ff",
          4420 => x"5c",
          4421 => x"84",
          4422 => x"5c",
          4423 => x"12",
          4424 => x"80",
          4425 => x"78",
          4426 => x"7c",
          4427 => x"90",
          4428 => x"c0",
          4429 => x"90",
          4430 => x"15",
          4431 => x"90",
          4432 => x"54",
          4433 => x"91",
          4434 => x"31",
          4435 => x"84",
          4436 => x"07",
          4437 => x"16",
          4438 => x"73",
          4439 => x"0c",
          4440 => x"04",
          4441 => x"6b",
          4442 => x"05",
          4443 => x"33",
          4444 => x"5a",
          4445 => x"bd",
          4446 => x"80",
          4447 => x"88",
          4448 => x"f8",
          4449 => x"88",
          4450 => x"91",
          4451 => x"70",
          4452 => x"74",
          4453 => x"38",
          4454 => x"91",
          4455 => x"81",
          4456 => x"81",
          4457 => x"ff",
          4458 => x"91",
          4459 => x"81",
          4460 => x"81",
          4461 => x"83",
          4462 => x"c0",
          4463 => x"2a",
          4464 => x"51",
          4465 => x"74",
          4466 => x"99",
          4467 => x"53",
          4468 => x"51",
          4469 => x"3f",
          4470 => x"08",
          4471 => x"55",
          4472 => x"92",
          4473 => x"80",
          4474 => x"38",
          4475 => x"06",
          4476 => x"2e",
          4477 => x"48",
          4478 => x"87",
          4479 => x"79",
          4480 => x"78",
          4481 => x"26",
          4482 => x"19",
          4483 => x"74",
          4484 => x"38",
          4485 => x"e4",
          4486 => x"2a",
          4487 => x"70",
          4488 => x"59",
          4489 => x"7a",
          4490 => x"56",
          4491 => x"80",
          4492 => x"51",
          4493 => x"74",
          4494 => x"99",
          4495 => x"53",
          4496 => x"51",
          4497 => x"3f",
          4498 => x"ca",
          4499 => x"ac",
          4500 => x"2a",
          4501 => x"91",
          4502 => x"43",
          4503 => x"83",
          4504 => x"66",
          4505 => x"60",
          4506 => x"90",
          4507 => x"31",
          4508 => x"80",
          4509 => x"8a",
          4510 => x"56",
          4511 => x"26",
          4512 => x"77",
          4513 => x"81",
          4514 => x"74",
          4515 => x"38",
          4516 => x"55",
          4517 => x"83",
          4518 => x"81",
          4519 => x"80",
          4520 => x"38",
          4521 => x"55",
          4522 => x"5e",
          4523 => x"89",
          4524 => x"5a",
          4525 => x"09",
          4526 => x"e1",
          4527 => x"38",
          4528 => x"57",
          4529 => x"ba",
          4530 => x"5a",
          4531 => x"9d",
          4532 => x"26",
          4533 => x"ba",
          4534 => x"10",
          4535 => x"22",
          4536 => x"74",
          4537 => x"38",
          4538 => x"ee",
          4539 => x"66",
          4540 => x"f6",
          4541 => x"88",
          4542 => x"84",
          4543 => x"89",
          4544 => x"a0",
          4545 => x"91",
          4546 => x"fc",
          4547 => x"56",
          4548 => x"f0",
          4549 => x"80",
          4550 => x"d3",
          4551 => x"38",
          4552 => x"57",
          4553 => x"ba",
          4554 => x"5a",
          4555 => x"9d",
          4556 => x"26",
          4557 => x"ba",
          4558 => x"10",
          4559 => x"22",
          4560 => x"74",
          4561 => x"38",
          4562 => x"ee",
          4563 => x"66",
          4564 => x"96",
          4565 => x"88",
          4566 => x"05",
          4567 => x"88",
          4568 => x"26",
          4569 => x"0b",
          4570 => x"08",
          4571 => x"88",
          4572 => x"11",
          4573 => x"05",
          4574 => x"83",
          4575 => x"2a",
          4576 => x"a0",
          4577 => x"7d",
          4578 => x"69",
          4579 => x"05",
          4580 => x"72",
          4581 => x"5c",
          4582 => x"59",
          4583 => x"2e",
          4584 => x"89",
          4585 => x"60",
          4586 => x"84",
          4587 => x"5d",
          4588 => x"18",
          4589 => x"68",
          4590 => x"74",
          4591 => x"af",
          4592 => x"31",
          4593 => x"53",
          4594 => x"52",
          4595 => x"9a",
          4596 => x"88",
          4597 => x"83",
          4598 => x"06",
          4599 => x"ca",
          4600 => x"ff",
          4601 => x"dd",
          4602 => x"83",
          4603 => x"2a",
          4604 => x"be",
          4605 => x"39",
          4606 => x"09",
          4607 => x"c5",
          4608 => x"f5",
          4609 => x"88",
          4610 => x"38",
          4611 => x"79",
          4612 => x"80",
          4613 => x"38",
          4614 => x"96",
          4615 => x"06",
          4616 => x"2e",
          4617 => x"5e",
          4618 => x"91",
          4619 => x"9f",
          4620 => x"38",
          4621 => x"38",
          4622 => x"81",
          4623 => x"fc",
          4624 => x"ab",
          4625 => x"7d",
          4626 => x"81",
          4627 => x"7d",
          4628 => x"78",
          4629 => x"74",
          4630 => x"8e",
          4631 => x"9c",
          4632 => x"53",
          4633 => x"51",
          4634 => x"3f",
          4635 => x"b8",
          4636 => x"51",
          4637 => x"3f",
          4638 => x"8b",
          4639 => x"a1",
          4640 => x"8d",
          4641 => x"83",
          4642 => x"52",
          4643 => x"ff",
          4644 => x"81",
          4645 => x"34",
          4646 => x"70",
          4647 => x"2a",
          4648 => x"54",
          4649 => x"1b",
          4650 => x"88",
          4651 => x"74",
          4652 => x"26",
          4653 => x"83",
          4654 => x"52",
          4655 => x"ff",
          4656 => x"8a",
          4657 => x"a0",
          4658 => x"a1",
          4659 => x"0b",
          4660 => x"bf",
          4661 => x"51",
          4662 => x"3f",
          4663 => x"9a",
          4664 => x"a0",
          4665 => x"52",
          4666 => x"ff",
          4667 => x"7d",
          4668 => x"81",
          4669 => x"38",
          4670 => x"0a",
          4671 => x"1b",
          4672 => x"ce",
          4673 => x"a4",
          4674 => x"a0",
          4675 => x"52",
          4676 => x"ff",
          4677 => x"81",
          4678 => x"51",
          4679 => x"3f",
          4680 => x"1b",
          4681 => x"8c",
          4682 => x"0b",
          4683 => x"34",
          4684 => x"c2",
          4685 => x"53",
          4686 => x"52",
          4687 => x"51",
          4688 => x"88",
          4689 => x"a7",
          4690 => x"a0",
          4691 => x"83",
          4692 => x"52",
          4693 => x"ff",
          4694 => x"ff",
          4695 => x"1c",
          4696 => x"a6",
          4697 => x"53",
          4698 => x"52",
          4699 => x"ff",
          4700 => x"82",
          4701 => x"83",
          4702 => x"52",
          4703 => x"b4",
          4704 => x"60",
          4705 => x"7e",
          4706 => x"d7",
          4707 => x"91",
          4708 => x"83",
          4709 => x"83",
          4710 => x"06",
          4711 => x"75",
          4712 => x"05",
          4713 => x"7e",
          4714 => x"b7",
          4715 => x"53",
          4716 => x"51",
          4717 => x"3f",
          4718 => x"a4",
          4719 => x"51",
          4720 => x"3f",
          4721 => x"e4",
          4722 => x"e4",
          4723 => x"9f",
          4724 => x"18",
          4725 => x"1b",
          4726 => x"f6",
          4727 => x"83",
          4728 => x"ff",
          4729 => x"82",
          4730 => x"78",
          4731 => x"c4",
          4732 => x"60",
          4733 => x"7a",
          4734 => x"ff",
          4735 => x"75",
          4736 => x"53",
          4737 => x"51",
          4738 => x"3f",
          4739 => x"52",
          4740 => x"9f",
          4741 => x"56",
          4742 => x"83",
          4743 => x"06",
          4744 => x"52",
          4745 => x"9e",
          4746 => x"52",
          4747 => x"ff",
          4748 => x"f0",
          4749 => x"1b",
          4750 => x"87",
          4751 => x"55",
          4752 => x"83",
          4753 => x"74",
          4754 => x"ff",
          4755 => x"7c",
          4756 => x"74",
          4757 => x"38",
          4758 => x"54",
          4759 => x"52",
          4760 => x"99",
          4761 => x"ca",
          4762 => x"87",
          4763 => x"53",
          4764 => x"08",
          4765 => x"ff",
          4766 => x"76",
          4767 => x"31",
          4768 => x"cd",
          4769 => x"58",
          4770 => x"ff",
          4771 => x"55",
          4772 => x"83",
          4773 => x"61",
          4774 => x"26",
          4775 => x"57",
          4776 => x"53",
          4777 => x"51",
          4778 => x"3f",
          4779 => x"08",
          4780 => x"76",
          4781 => x"31",
          4782 => x"db",
          4783 => x"7d",
          4784 => x"38",
          4785 => x"83",
          4786 => x"8a",
          4787 => x"7d",
          4788 => x"38",
          4789 => x"81",
          4790 => x"80",
          4791 => x"80",
          4792 => x"7a",
          4793 => x"bc",
          4794 => x"d5",
          4795 => x"ff",
          4796 => x"83",
          4797 => x"77",
          4798 => x"0b",
          4799 => x"81",
          4800 => x"34",
          4801 => x"34",
          4802 => x"34",
          4803 => x"56",
          4804 => x"52",
          4805 => x"f4",
          4806 => x"0b",
          4807 => x"91",
          4808 => x"82",
          4809 => x"56",
          4810 => x"34",
          4811 => x"08",
          4812 => x"60",
          4813 => x"1b",
          4814 => x"96",
          4815 => x"83",
          4816 => x"ff",
          4817 => x"81",
          4818 => x"7a",
          4819 => x"ff",
          4820 => x"81",
          4821 => x"88",
          4822 => x"80",
          4823 => x"7e",
          4824 => x"e3",
          4825 => x"91",
          4826 => x"90",
          4827 => x"8e",
          4828 => x"81",
          4829 => x"91",
          4830 => x"56",
          4831 => x"88",
          4832 => x"0d",
          4833 => x"0d",
          4834 => x"93",
          4835 => x"38",
          4836 => x"91",
          4837 => x"52",
          4838 => x"91",
          4839 => x"81",
          4840 => x"bb",
          4841 => x"f9",
          4842 => x"f8",
          4843 => x"39",
          4844 => x"51",
          4845 => x"91",
          4846 => x"80",
          4847 => x"bc",
          4848 => x"dd",
          4849 => x"c0",
          4850 => x"39",
          4851 => x"51",
          4852 => x"91",
          4853 => x"80",
          4854 => x"bd",
          4855 => x"c1",
          4856 => x"98",
          4857 => x"91",
          4858 => x"b5",
          4859 => x"c8",
          4860 => x"91",
          4861 => x"a9",
          4862 => x"88",
          4863 => x"91",
          4864 => x"9d",
          4865 => x"bc",
          4866 => x"91",
          4867 => x"91",
          4868 => x"ec",
          4869 => x"91",
          4870 => x"85",
          4871 => x"90",
          4872 => x"fb",
          4873 => x"0d",
          4874 => x"0d",
          4875 => x"56",
          4876 => x"26",
          4877 => x"52",
          4878 => x"29",
          4879 => x"87",
          4880 => x"51",
          4881 => x"3f",
          4882 => x"08",
          4883 => x"fe",
          4884 => x"91",
          4885 => x"54",
          4886 => x"52",
          4887 => x"51",
          4888 => x"3f",
          4889 => x"04",
          4890 => x"7d",
          4891 => x"8c",
          4892 => x"05",
          4893 => x"15",
          4894 => x"5a",
          4895 => x"5c",
          4896 => x"bf",
          4897 => x"8c",
          4898 => x"bf",
          4899 => x"87",
          4900 => x"55",
          4901 => x"80",
          4902 => x"90",
          4903 => x"79",
          4904 => x"38",
          4905 => x"74",
          4906 => x"78",
          4907 => x"72",
          4908 => x"bf",
          4909 => x"8c",
          4910 => x"39",
          4911 => x"51",
          4912 => x"3f",
          4913 => x"80",
          4914 => x"16",
          4915 => x"27",
          4916 => x"08",
          4917 => x"c4",
          4918 => x"a7",
          4919 => x"91",
          4920 => x"ff",
          4921 => x"84",
          4922 => x"39",
          4923 => x"72",
          4924 => x"38",
          4925 => x"91",
          4926 => x"ff",
          4927 => x"89",
          4928 => x"ec",
          4929 => x"97",
          4930 => x"55",
          4931 => x"fa",
          4932 => x"80",
          4933 => x"f0",
          4934 => x"83",
          4935 => x"74",
          4936 => x"38",
          4937 => x"33",
          4938 => x"52",
          4939 => x"74",
          4940 => x"72",
          4941 => x"38",
          4942 => x"26",
          4943 => x"51",
          4944 => x"51",
          4945 => x"3f",
          4946 => x"d3",
          4947 => x"f4",
          4948 => x"cb",
          4949 => x"77",
          4950 => x"fe",
          4951 => x"91",
          4952 => x"98",
          4953 => x"2c",
          4954 => x"a0",
          4955 => x"06",
          4956 => x"fc",
          4957 => x"ca",
          4958 => x"2b",
          4959 => x"70",
          4960 => x"30",
          4961 => x"9f",
          4962 => x"56",
          4963 => x"9b",
          4964 => x"72",
          4965 => x"9b",
          4966 => x"06",
          4967 => x"53",
          4968 => x"1c",
          4969 => x"26",
          4970 => x"ff",
          4971 => x"ca",
          4972 => x"3d",
          4973 => x"3d",
          4974 => x"84",
          4975 => x"05",
          4976 => x"30",
          4977 => x"80",
          4978 => x"ff",
          4979 => x"51",
          4980 => x"5b",
          4981 => x"74",
          4982 => x"81",
          4983 => x"8c",
          4984 => x"57",
          4985 => x"91",
          4986 => x"56",
          4987 => x"08",
          4988 => x"ca",
          4989 => x"c0",
          4990 => x"91",
          4991 => x"59",
          4992 => x"05",
          4993 => x"53",
          4994 => x"51",
          4995 => x"91",
          4996 => x"56",
          4997 => x"08",
          4998 => x"55",
          4999 => x"89",
          5000 => x"75",
          5001 => x"d8",
          5002 => x"d8",
          5003 => x"e0",
          5004 => x"70",
          5005 => x"25",
          5006 => x"80",
          5007 => x"74",
          5008 => x"38",
          5009 => x"53",
          5010 => x"88",
          5011 => x"51",
          5012 => x"75",
          5013 => x"ca",
          5014 => x"3d",
          5015 => x"3d",
          5016 => x"84",
          5017 => x"33",
          5018 => x"57",
          5019 => x"52",
          5020 => x"c2",
          5021 => x"88",
          5022 => x"75",
          5023 => x"38",
          5024 => x"98",
          5025 => x"60",
          5026 => x"91",
          5027 => x"7e",
          5028 => x"77",
          5029 => x"88",
          5030 => x"39",
          5031 => x"91",
          5032 => x"89",
          5033 => x"fc",
          5034 => x"9b",
          5035 => x"c0",
          5036 => x"c0",
          5037 => x"ff",
          5038 => x"91",
          5039 => x"51",
          5040 => x"3f",
          5041 => x"54",
          5042 => x"53",
          5043 => x"33",
          5044 => x"a8",
          5045 => x"ab",
          5046 => x"2e",
          5047 => x"fe",
          5048 => x"3d",
          5049 => x"3d",
          5050 => x"96",
          5051 => x"ff",
          5052 => x"81",
          5053 => x"8c",
          5054 => x"c4",
          5055 => x"84",
          5056 => x"fe",
          5057 => x"72",
          5058 => x"81",
          5059 => x"71",
          5060 => x"38",
          5061 => x"f5",
          5062 => x"c0",
          5063 => x"f7",
          5064 => x"51",
          5065 => x"3f",
          5066 => x"70",
          5067 => x"52",
          5068 => x"95",
          5069 => x"fe",
          5070 => x"91",
          5071 => x"fe",
          5072 => x"80",
          5073 => x"bc",
          5074 => x"2a",
          5075 => x"51",
          5076 => x"2e",
          5077 => x"51",
          5078 => x"3f",
          5079 => x"51",
          5080 => x"3f",
          5081 => x"f5",
          5082 => x"84",
          5083 => x"06",
          5084 => x"80",
          5085 => x"81",
          5086 => x"88",
          5087 => x"98",
          5088 => x"80",
          5089 => x"fe",
          5090 => x"72",
          5091 => x"81",
          5092 => x"71",
          5093 => x"38",
          5094 => x"f4",
          5095 => x"c1",
          5096 => x"f6",
          5097 => x"51",
          5098 => x"3f",
          5099 => x"70",
          5100 => x"52",
          5101 => x"95",
          5102 => x"fe",
          5103 => x"91",
          5104 => x"fe",
          5105 => x"80",
          5106 => x"b8",
          5107 => x"2a",
          5108 => x"51",
          5109 => x"2e",
          5110 => x"51",
          5111 => x"3f",
          5112 => x"51",
          5113 => x"3f",
          5114 => x"f4",
          5115 => x"88",
          5116 => x"06",
          5117 => x"80",
          5118 => x"81",
          5119 => x"84",
          5120 => x"e8",
          5121 => x"fc",
          5122 => x"fe",
          5123 => x"fe",
          5124 => x"84",
          5125 => x"fa",
          5126 => x"70",
          5127 => x"55",
          5128 => x"2e",
          5129 => x"8e",
          5130 => x"0c",
          5131 => x"53",
          5132 => x"81",
          5133 => x"74",
          5134 => x"ff",
          5135 => x"53",
          5136 => x"83",
          5137 => x"74",
          5138 => x"38",
          5139 => x"75",
          5140 => x"53",
          5141 => x"09",
          5142 => x"38",
          5143 => x"81",
          5144 => x"80",
          5145 => x"29",
          5146 => x"05",
          5147 => x"70",
          5148 => x"fe",
          5149 => x"91",
          5150 => x"8b",
          5151 => x"33",
          5152 => x"2e",
          5153 => x"81",
          5154 => x"ff",
          5155 => x"95",
          5156 => x"38",
          5157 => x"91",
          5158 => x"88",
          5159 => x"cb",
          5160 => x"70",
          5161 => x"88",
          5162 => x"81",
          5163 => x"ff",
          5164 => x"91",
          5165 => x"81",
          5166 => x"78",
          5167 => x"81",
          5168 => x"91",
          5169 => x"99",
          5170 => x"59",
          5171 => x"3f",
          5172 => x"52",
          5173 => x"51",
          5174 => x"3f",
          5175 => x"08",
          5176 => x"38",
          5177 => x"51",
          5178 => x"81",
          5179 => x"91",
          5180 => x"fe",
          5181 => x"99",
          5182 => x"5a",
          5183 => x"80",
          5184 => x"fe",
          5185 => x"80",
          5186 => x"51",
          5187 => x"3f",
          5188 => x"f8",
          5189 => x"ff",
          5190 => x"88",
          5191 => x"70",
          5192 => x"59",
          5193 => x"2e",
          5194 => x"78",
          5195 => x"80",
          5196 => x"b0",
          5197 => x"38",
          5198 => x"aa",
          5199 => x"2e",
          5200 => x"78",
          5201 => x"38",
          5202 => x"ff",
          5203 => x"82",
          5204 => x"38",
          5205 => x"78",
          5206 => x"b8",
          5207 => x"2e",
          5208 => x"8e",
          5209 => x"bf",
          5210 => x"38",
          5211 => x"90",
          5212 => x"2e",
          5213 => x"78",
          5214 => x"fc",
          5215 => x"39",
          5216 => x"2e",
          5217 => x"78",
          5218 => x"88",
          5219 => x"b7",
          5220 => x"f8",
          5221 => x"38",
          5222 => x"24",
          5223 => x"80",
          5224 => x"cd",
          5225 => x"d1",
          5226 => x"78",
          5227 => x"8b",
          5228 => x"80",
          5229 => x"a8",
          5230 => x"39",
          5231 => x"2e",
          5232 => x"78",
          5233 => x"8c",
          5234 => x"fb",
          5235 => x"83",
          5236 => x"38",
          5237 => x"24",
          5238 => x"80",
          5239 => x"81",
          5240 => x"82",
          5241 => x"38",
          5242 => x"78",
          5243 => x"8d",
          5244 => x"81",
          5245 => x"f7",
          5246 => x"39",
          5247 => x"f4",
          5248 => x"f8",
          5249 => x"83",
          5250 => x"ca",
          5251 => x"38",
          5252 => x"51",
          5253 => x"b7",
          5254 => x"11",
          5255 => x"05",
          5256 => x"d4",
          5257 => x"88",
          5258 => x"88",
          5259 => x"25",
          5260 => x"43",
          5261 => x"05",
          5262 => x"80",
          5263 => x"51",
          5264 => x"3f",
          5265 => x"08",
          5266 => x"59",
          5267 => x"91",
          5268 => x"fe",
          5269 => x"81",
          5270 => x"39",
          5271 => x"51",
          5272 => x"b7",
          5273 => x"11",
          5274 => x"05",
          5275 => x"88",
          5276 => x"88",
          5277 => x"fc",
          5278 => x"53",
          5279 => x"80",
          5280 => x"51",
          5281 => x"3f",
          5282 => x"08",
          5283 => x"a0",
          5284 => x"39",
          5285 => x"f4",
          5286 => x"f8",
          5287 => x"82",
          5288 => x"ca",
          5289 => x"2e",
          5290 => x"89",
          5291 => x"38",
          5292 => x"f0",
          5293 => x"f8",
          5294 => x"82",
          5295 => x"ca",
          5296 => x"38",
          5297 => x"08",
          5298 => x"91",
          5299 => x"79",
          5300 => x"c5",
          5301 => x"cb",
          5302 => x"79",
          5303 => x"b4",
          5304 => x"b8",
          5305 => x"b5",
          5306 => x"ca",
          5307 => x"93",
          5308 => x"f8",
          5309 => x"a7",
          5310 => x"fb",
          5311 => x"3d",
          5312 => x"51",
          5313 => x"3f",
          5314 => x"08",
          5315 => x"f8",
          5316 => x"fe",
          5317 => x"81",
          5318 => x"88",
          5319 => x"51",
          5320 => x"80",
          5321 => x"3d",
          5322 => x"51",
          5323 => x"3f",
          5324 => x"08",
          5325 => x"f8",
          5326 => x"fe",
          5327 => x"91",
          5328 => x"b8",
          5329 => x"05",
          5330 => x"ea",
          5331 => x"ca",
          5332 => x"3d",
          5333 => x"52",
          5334 => x"bb",
          5335 => x"e4",
          5336 => x"bc",
          5337 => x"80",
          5338 => x"88",
          5339 => x"06",
          5340 => x"79",
          5341 => x"f5",
          5342 => x"ca",
          5343 => x"2e",
          5344 => x"91",
          5345 => x"51",
          5346 => x"fa",
          5347 => x"3d",
          5348 => x"53",
          5349 => x"51",
          5350 => x"3f",
          5351 => x"08",
          5352 => x"cb",
          5353 => x"fe",
          5354 => x"fe",
          5355 => x"ff",
          5356 => x"91",
          5357 => x"80",
          5358 => x"38",
          5359 => x"ec",
          5360 => x"f8",
          5361 => x"80",
          5362 => x"ca",
          5363 => x"38",
          5364 => x"08",
          5365 => x"ac",
          5366 => x"c3",
          5367 => x"5c",
          5368 => x"27",
          5369 => x"61",
          5370 => x"70",
          5371 => x"0c",
          5372 => x"f5",
          5373 => x"39",
          5374 => x"f4",
          5375 => x"f8",
          5376 => x"ff",
          5377 => x"ca",
          5378 => x"2e",
          5379 => x"b7",
          5380 => x"11",
          5381 => x"05",
          5382 => x"dc",
          5383 => x"88",
          5384 => x"f9",
          5385 => x"3d",
          5386 => x"53",
          5387 => x"51",
          5388 => x"3f",
          5389 => x"08",
          5390 => x"b3",
          5391 => x"b8",
          5392 => x"db",
          5393 => x"79",
          5394 => x"8c",
          5395 => x"79",
          5396 => x"5b",
          5397 => x"61",
          5398 => x"eb",
          5399 => x"fe",
          5400 => x"fe",
          5401 => x"fe",
          5402 => x"91",
          5403 => x"80",
          5404 => x"38",
          5405 => x"f0",
          5406 => x"f8",
          5407 => x"fe",
          5408 => x"ca",
          5409 => x"2e",
          5410 => x"b7",
          5411 => x"11",
          5412 => x"05",
          5413 => x"e0",
          5414 => x"88",
          5415 => x"f8",
          5416 => x"c3",
          5417 => x"f6",
          5418 => x"5a",
          5419 => x"a8",
          5420 => x"33",
          5421 => x"5a",
          5422 => x"2e",
          5423 => x"55",
          5424 => x"33",
          5425 => x"91",
          5426 => x"fe",
          5427 => x"81",
          5428 => x"05",
          5429 => x"39",
          5430 => x"51",
          5431 => x"b7",
          5432 => x"11",
          5433 => x"05",
          5434 => x"8c",
          5435 => x"88",
          5436 => x"38",
          5437 => x"33",
          5438 => x"2e",
          5439 => x"c6",
          5440 => x"b3",
          5441 => x"92",
          5442 => x"80",
          5443 => x"91",
          5444 => x"44",
          5445 => x"c7",
          5446 => x"78",
          5447 => x"c7",
          5448 => x"78",
          5449 => x"38",
          5450 => x"08",
          5451 => x"91",
          5452 => x"fc",
          5453 => x"b7",
          5454 => x"11",
          5455 => x"05",
          5456 => x"b4",
          5457 => x"88",
          5458 => x"38",
          5459 => x"33",
          5460 => x"2e",
          5461 => x"c6",
          5462 => x"b2",
          5463 => x"92",
          5464 => x"80",
          5465 => x"91",
          5466 => x"43",
          5467 => x"c7",
          5468 => x"78",
          5469 => x"c7",
          5470 => x"78",
          5471 => x"38",
          5472 => x"08",
          5473 => x"91",
          5474 => x"88",
          5475 => x"3d",
          5476 => x"53",
          5477 => x"51",
          5478 => x"3f",
          5479 => x"08",
          5480 => x"38",
          5481 => x"59",
          5482 => x"83",
          5483 => x"79",
          5484 => x"38",
          5485 => x"88",
          5486 => x"2e",
          5487 => x"42",
          5488 => x"51",
          5489 => x"3f",
          5490 => x"54",
          5491 => x"52",
          5492 => x"94",
          5493 => x"80",
          5494 => x"39",
          5495 => x"f4",
          5496 => x"f8",
          5497 => x"fc",
          5498 => x"ca",
          5499 => x"2e",
          5500 => x"b7",
          5501 => x"11",
          5502 => x"05",
          5503 => x"f8",
          5504 => x"88",
          5505 => x"a5",
          5506 => x"02",
          5507 => x"33",
          5508 => x"81",
          5509 => x"3d",
          5510 => x"53",
          5511 => x"51",
          5512 => x"3f",
          5513 => x"08",
          5514 => x"c3",
          5515 => x"33",
          5516 => x"c4",
          5517 => x"f9",
          5518 => x"f8",
          5519 => x"fe",
          5520 => x"79",
          5521 => x"59",
          5522 => x"f5",
          5523 => x"79",
          5524 => x"b7",
          5525 => x"11",
          5526 => x"05",
          5527 => x"98",
          5528 => x"88",
          5529 => x"91",
          5530 => x"02",
          5531 => x"33",
          5532 => x"81",
          5533 => x"b5",
          5534 => x"98",
          5535 => x"9f",
          5536 => x"39",
          5537 => x"e8",
          5538 => x"f8",
          5539 => x"fc",
          5540 => x"ca",
          5541 => x"2e",
          5542 => x"b7",
          5543 => x"11",
          5544 => x"05",
          5545 => x"c2",
          5546 => x"88",
          5547 => x"a6",
          5548 => x"02",
          5549 => x"79",
          5550 => x"5b",
          5551 => x"b7",
          5552 => x"11",
          5553 => x"05",
          5554 => x"9e",
          5555 => x"88",
          5556 => x"f4",
          5557 => x"70",
          5558 => x"91",
          5559 => x"fe",
          5560 => x"80",
          5561 => x"51",
          5562 => x"3f",
          5563 => x"33",
          5564 => x"2e",
          5565 => x"78",
          5566 => x"38",
          5567 => x"41",
          5568 => x"3d",
          5569 => x"53",
          5570 => x"51",
          5571 => x"3f",
          5572 => x"08",
          5573 => x"38",
          5574 => x"be",
          5575 => x"70",
          5576 => x"23",
          5577 => x"ae",
          5578 => x"98",
          5579 => x"ef",
          5580 => x"39",
          5581 => x"e8",
          5582 => x"f8",
          5583 => x"fb",
          5584 => x"ca",
          5585 => x"2e",
          5586 => x"b7",
          5587 => x"11",
          5588 => x"05",
          5589 => x"92",
          5590 => x"88",
          5591 => x"a1",
          5592 => x"71",
          5593 => x"84",
          5594 => x"3d",
          5595 => x"53",
          5596 => x"51",
          5597 => x"3f",
          5598 => x"08",
          5599 => x"ef",
          5600 => x"08",
          5601 => x"c4",
          5602 => x"f6",
          5603 => x"f8",
          5604 => x"fe",
          5605 => x"79",
          5606 => x"59",
          5607 => x"f2",
          5608 => x"79",
          5609 => x"b7",
          5610 => x"11",
          5611 => x"05",
          5612 => x"b6",
          5613 => x"88",
          5614 => x"99",
          5615 => x"60",
          5616 => x"ac",
          5617 => x"bb",
          5618 => x"71",
          5619 => x"84",
          5620 => x"ad",
          5621 => x"98",
          5622 => x"c3",
          5623 => x"39",
          5624 => x"51",
          5625 => x"3f",
          5626 => x"ef",
          5627 => x"ff",
          5628 => x"d0",
          5629 => x"a7",
          5630 => x"fe",
          5631 => x"f1",
          5632 => x"80",
          5633 => x"c0",
          5634 => x"84",
          5635 => x"87",
          5636 => x"0c",
          5637 => x"51",
          5638 => x"3f",
          5639 => x"91",
          5640 => x"fe",
          5641 => x"8c",
          5642 => x"87",
          5643 => x"0c",
          5644 => x"0b",
          5645 => x"94",
          5646 => x"39",
          5647 => x"f4",
          5648 => x"f8",
          5649 => x"f7",
          5650 => x"ca",
          5651 => x"2e",
          5652 => x"63",
          5653 => x"90",
          5654 => x"a7",
          5655 => x"78",
          5656 => x"fe",
          5657 => x"fe",
          5658 => x"fe",
          5659 => x"91",
          5660 => x"80",
          5661 => x"38",
          5662 => x"c5",
          5663 => x"f5",
          5664 => x"59",
          5665 => x"ca",
          5666 => x"91",
          5667 => x"80",
          5668 => x"38",
          5669 => x"08",
          5670 => x"c8",
          5671 => x"e3",
          5672 => x"39",
          5673 => x"51",
          5674 => x"3f",
          5675 => x"3f",
          5676 => x"91",
          5677 => x"fe",
          5678 => x"80",
          5679 => x"39",
          5680 => x"3f",
          5681 => x"64",
          5682 => x"59",
          5683 => x"f0",
          5684 => x"80",
          5685 => x"38",
          5686 => x"80",
          5687 => x"3d",
          5688 => x"51",
          5689 => x"3f",
          5690 => x"56",
          5691 => x"08",
          5692 => x"98",
          5693 => x"91",
          5694 => x"a3",
          5695 => x"5a",
          5696 => x"3f",
          5697 => x"58",
          5698 => x"57",
          5699 => x"81",
          5700 => x"05",
          5701 => x"91",
          5702 => x"91",
          5703 => x"79",
          5704 => x"3f",
          5705 => x"08",
          5706 => x"32",
          5707 => x"07",
          5708 => x"38",
          5709 => x"09",
          5710 => x"b3",
          5711 => x"ac",
          5712 => x"bf",
          5713 => x"39",
          5714 => x"80",
          5715 => x"bc",
          5716 => x"9b",
          5717 => x"98",
          5718 => x"9c",
          5719 => x"9c",
          5720 => x"e4",
          5721 => x"87",
          5722 => x"bc",
          5723 => x"94",
          5724 => x"c8",
          5725 => x"a7",
          5726 => x"e3",
          5727 => x"ea",
          5728 => x"ea",
          5729 => x"97",
          5730 => x"00",
          5731 => x"00",
          5732 => x"00",
          5733 => x"00",
          5734 => x"00",
          5735 => x"00",
          5736 => x"00",
          5737 => x"00",
          5738 => x"00",
          5739 => x"00",
          5740 => x"00",
          5741 => x"00",
          5742 => x"00",
          5743 => x"00",
          5744 => x"00",
          5745 => x"00",
          5746 => x"00",
          5747 => x"00",
          5748 => x"00",
          5749 => x"00",
          5750 => x"00",
          5751 => x"00",
          5752 => x"00",
          5753 => x"00",
          5754 => x"00",
          5755 => x"25",
          5756 => x"64",
          5757 => x"20",
          5758 => x"25",
          5759 => x"64",
          5760 => x"25",
          5761 => x"53",
          5762 => x"43",
          5763 => x"69",
          5764 => x"61",
          5765 => x"6e",
          5766 => x"20",
          5767 => x"6f",
          5768 => x"6f",
          5769 => x"6f",
          5770 => x"67",
          5771 => x"3a",
          5772 => x"76",
          5773 => x"73",
          5774 => x"70",
          5775 => x"65",
          5776 => x"64",
          5777 => x"20",
          5778 => x"49",
          5779 => x"20",
          5780 => x"4d",
          5781 => x"74",
          5782 => x"3d",
          5783 => x"58",
          5784 => x"69",
          5785 => x"25",
          5786 => x"29",
          5787 => x"20",
          5788 => x"42",
          5789 => x"20",
          5790 => x"61",
          5791 => x"25",
          5792 => x"2c",
          5793 => x"7a",
          5794 => x"30",
          5795 => x"2e",
          5796 => x"20",
          5797 => x"52",
          5798 => x"28",
          5799 => x"72",
          5800 => x"30",
          5801 => x"20",
          5802 => x"65",
          5803 => x"38",
          5804 => x"0a",
          5805 => x"20",
          5806 => x"49",
          5807 => x"4c",
          5808 => x"20",
          5809 => x"50",
          5810 => x"00",
          5811 => x"20",
          5812 => x"53",
          5813 => x"00",
          5814 => x"20",
          5815 => x"53",
          5816 => x"61",
          5817 => x"28",
          5818 => x"69",
          5819 => x"3d",
          5820 => x"58",
          5821 => x"00",
          5822 => x"20",
          5823 => x"49",
          5824 => x"52",
          5825 => x"54",
          5826 => x"4e",
          5827 => x"4c",
          5828 => x"0a",
          5829 => x"20",
          5830 => x"54",
          5831 => x"52",
          5832 => x"54",
          5833 => x"72",
          5834 => x"30",
          5835 => x"2e",
          5836 => x"41",
          5837 => x"65",
          5838 => x"73",
          5839 => x"20",
          5840 => x"43",
          5841 => x"52",
          5842 => x"74",
          5843 => x"63",
          5844 => x"20",
          5845 => x"72",
          5846 => x"20",
          5847 => x"30",
          5848 => x"00",
          5849 => x"20",
          5850 => x"43",
          5851 => x"4d",
          5852 => x"72",
          5853 => x"74",
          5854 => x"20",
          5855 => x"72",
          5856 => x"20",
          5857 => x"30",
          5858 => x"00",
          5859 => x"20",
          5860 => x"53",
          5861 => x"6b",
          5862 => x"61",
          5863 => x"41",
          5864 => x"65",
          5865 => x"20",
          5866 => x"20",
          5867 => x"30",
          5868 => x"00",
          5869 => x"20",
          5870 => x"5a",
          5871 => x"49",
          5872 => x"20",
          5873 => x"20",
          5874 => x"20",
          5875 => x"20",
          5876 => x"20",
          5877 => x"30",
          5878 => x"00",
          5879 => x"20",
          5880 => x"53",
          5881 => x"65",
          5882 => x"6c",
          5883 => x"20",
          5884 => x"71",
          5885 => x"20",
          5886 => x"20",
          5887 => x"30",
          5888 => x"00",
          5889 => x"53",
          5890 => x"6c",
          5891 => x"4d",
          5892 => x"75",
          5893 => x"46",
          5894 => x"00",
          5895 => x"45",
          5896 => x"45",
          5897 => x"69",
          5898 => x"55",
          5899 => x"6f",
          5900 => x"53",
          5901 => x"22",
          5902 => x"3a",
          5903 => x"3e",
          5904 => x"7c",
          5905 => x"46",
          5906 => x"46",
          5907 => x"32",
          5908 => x"eb",
          5909 => x"53",
          5910 => x"35",
          5911 => x"4e",
          5912 => x"41",
          5913 => x"20",
          5914 => x"41",
          5915 => x"20",
          5916 => x"4e",
          5917 => x"41",
          5918 => x"20",
          5919 => x"41",
          5920 => x"20",
          5921 => x"00",
          5922 => x"00",
          5923 => x"00",
          5924 => x"00",
          5925 => x"80",
          5926 => x"8e",
          5927 => x"45",
          5928 => x"49",
          5929 => x"90",
          5930 => x"99",
          5931 => x"59",
          5932 => x"9c",
          5933 => x"41",
          5934 => x"a5",
          5935 => x"a8",
          5936 => x"ac",
          5937 => x"b0",
          5938 => x"b4",
          5939 => x"b8",
          5940 => x"bc",
          5941 => x"c0",
          5942 => x"c4",
          5943 => x"c8",
          5944 => x"cc",
          5945 => x"d0",
          5946 => x"d4",
          5947 => x"d8",
          5948 => x"dc",
          5949 => x"e0",
          5950 => x"e4",
          5951 => x"e8",
          5952 => x"ec",
          5953 => x"f0",
          5954 => x"f4",
          5955 => x"f8",
          5956 => x"fc",
          5957 => x"2b",
          5958 => x"3d",
          5959 => x"5c",
          5960 => x"3c",
          5961 => x"7f",
          5962 => x"00",
          5963 => x"00",
          5964 => x"01",
          5965 => x"00",
          5966 => x"00",
          5967 => x"00",
          5968 => x"00",
          5969 => x"00",
          5970 => x"64",
          5971 => x"74",
          5972 => x"64",
          5973 => x"74",
          5974 => x"66",
          5975 => x"74",
          5976 => x"66",
          5977 => x"64",
          5978 => x"66",
          5979 => x"63",
          5980 => x"6d",
          5981 => x"61",
          5982 => x"6d",
          5983 => x"79",
          5984 => x"6d",
          5985 => x"66",
          5986 => x"6d",
          5987 => x"70",
          5988 => x"6d",
          5989 => x"6d",
          5990 => x"6d",
          5991 => x"68",
          5992 => x"68",
          5993 => x"68",
          5994 => x"68",
          5995 => x"63",
          5996 => x"00",
          5997 => x"6a",
          5998 => x"72",
          5999 => x"61",
          6000 => x"72",
          6001 => x"74",
          6002 => x"69",
          6003 => x"00",
          6004 => x"74",
          6005 => x"00",
          6006 => x"44",
          6007 => x"20",
          6008 => x"6f",
          6009 => x"49",
          6010 => x"72",
          6011 => x"20",
          6012 => x"6f",
          6013 => x"00",
          6014 => x"44",
          6015 => x"20",
          6016 => x"20",
          6017 => x"64",
          6018 => x"00",
          6019 => x"4e",
          6020 => x"69",
          6021 => x"66",
          6022 => x"64",
          6023 => x"4e",
          6024 => x"61",
          6025 => x"66",
          6026 => x"64",
          6027 => x"49",
          6028 => x"6c",
          6029 => x"66",
          6030 => x"6e",
          6031 => x"2e",
          6032 => x"41",
          6033 => x"73",
          6034 => x"65",
          6035 => x"64",
          6036 => x"46",
          6037 => x"20",
          6038 => x"65",
          6039 => x"20",
          6040 => x"73",
          6041 => x"0a",
          6042 => x"46",
          6043 => x"20",
          6044 => x"64",
          6045 => x"69",
          6046 => x"6c",
          6047 => x"0a",
          6048 => x"53",
          6049 => x"73",
          6050 => x"69",
          6051 => x"70",
          6052 => x"65",
          6053 => x"64",
          6054 => x"44",
          6055 => x"65",
          6056 => x"6d",
          6057 => x"20",
          6058 => x"69",
          6059 => x"6c",
          6060 => x"0a",
          6061 => x"44",
          6062 => x"20",
          6063 => x"20",
          6064 => x"62",
          6065 => x"2e",
          6066 => x"4e",
          6067 => x"6f",
          6068 => x"74",
          6069 => x"65",
          6070 => x"6c",
          6071 => x"73",
          6072 => x"20",
          6073 => x"6e",
          6074 => x"6e",
          6075 => x"73",
          6076 => x"00",
          6077 => x"46",
          6078 => x"61",
          6079 => x"62",
          6080 => x"65",
          6081 => x"00",
          6082 => x"54",
          6083 => x"6f",
          6084 => x"20",
          6085 => x"72",
          6086 => x"6f",
          6087 => x"61",
          6088 => x"6c",
          6089 => x"2e",
          6090 => x"46",
          6091 => x"20",
          6092 => x"6c",
          6093 => x"65",
          6094 => x"00",
          6095 => x"49",
          6096 => x"66",
          6097 => x"69",
          6098 => x"20",
          6099 => x"6f",
          6100 => x"0a",
          6101 => x"54",
          6102 => x"6d",
          6103 => x"20",
          6104 => x"6e",
          6105 => x"6c",
          6106 => x"0a",
          6107 => x"50",
          6108 => x"6d",
          6109 => x"72",
          6110 => x"6e",
          6111 => x"72",
          6112 => x"2e",
          6113 => x"53",
          6114 => x"65",
          6115 => x"0a",
          6116 => x"55",
          6117 => x"6f",
          6118 => x"65",
          6119 => x"72",
          6120 => x"0a",
          6121 => x"20",
          6122 => x"65",
          6123 => x"73",
          6124 => x"20",
          6125 => x"20",
          6126 => x"65",
          6127 => x"65",
          6128 => x"00",
          6129 => x"25",
          6130 => x"00",
          6131 => x"3a",
          6132 => x"25",
          6133 => x"00",
          6134 => x"20",
          6135 => x"20",
          6136 => x"00",
          6137 => x"25",
          6138 => x"00",
          6139 => x"20",
          6140 => x"20",
          6141 => x"7c",
          6142 => x"72",
          6143 => x"00",
          6144 => x"5a",
          6145 => x"41",
          6146 => x"0a",
          6147 => x"25",
          6148 => x"00",
          6149 => x"31",
          6150 => x"37",
          6151 => x"31",
          6152 => x"76",
          6153 => x"00",
          6154 => x"20",
          6155 => x"2c",
          6156 => x"76",
          6157 => x"32",
          6158 => x"25",
          6159 => x"73",
          6160 => x"0a",
          6161 => x"5a",
          6162 => x"41",
          6163 => x"74",
          6164 => x"75",
          6165 => x"48",
          6166 => x"6c",
          6167 => x"00",
          6168 => x"54",
          6169 => x"72",
          6170 => x"74",
          6171 => x"75",
          6172 => x"00",
          6173 => x"50",
          6174 => x"69",
          6175 => x"72",
          6176 => x"74",
          6177 => x"49",
          6178 => x"4c",
          6179 => x"20",
          6180 => x"65",
          6181 => x"70",
          6182 => x"49",
          6183 => x"4c",
          6184 => x"20",
          6185 => x"65",
          6186 => x"70",
          6187 => x"55",
          6188 => x"30",
          6189 => x"20",
          6190 => x"65",
          6191 => x"70",
          6192 => x"55",
          6193 => x"30",
          6194 => x"20",
          6195 => x"65",
          6196 => x"70",
          6197 => x"55",
          6198 => x"31",
          6199 => x"20",
          6200 => x"65",
          6201 => x"70",
          6202 => x"55",
          6203 => x"31",
          6204 => x"20",
          6205 => x"65",
          6206 => x"70",
          6207 => x"53",
          6208 => x"69",
          6209 => x"75",
          6210 => x"69",
          6211 => x"2e",
          6212 => x"00",
          6213 => x"45",
          6214 => x"6c",
          6215 => x"20",
          6216 => x"65",
          6217 => x"2e",
          6218 => x"30",
          6219 => x"46",
          6220 => x"65",
          6221 => x"6f",
          6222 => x"69",
          6223 => x"6c",
          6224 => x"20",
          6225 => x"63",
          6226 => x"20",
          6227 => x"70",
          6228 => x"73",
          6229 => x"6e",
          6230 => x"6d",
          6231 => x"61",
          6232 => x"2e",
          6233 => x"2a",
          6234 => x"42",
          6235 => x"64",
          6236 => x"20",
          6237 => x"0a",
          6238 => x"49",
          6239 => x"69",
          6240 => x"73",
          6241 => x"0a",
          6242 => x"46",
          6243 => x"65",
          6244 => x"6f",
          6245 => x"69",
          6246 => x"6c",
          6247 => x"2e",
          6248 => x"72",
          6249 => x"64",
          6250 => x"25",
          6251 => x"43",
          6252 => x"72",
          6253 => x"2e",
          6254 => x"43",
          6255 => x"69",
          6256 => x"2e",
          6257 => x"43",
          6258 => x"61",
          6259 => x"67",
          6260 => x"00",
          6261 => x"25",
          6262 => x"78",
          6263 => x"38",
          6264 => x"3e",
          6265 => x"6c",
          6266 => x"30",
          6267 => x"0a",
          6268 => x"44",
          6269 => x"20",
          6270 => x"6f",
          6271 => x"00",
          6272 => x"0a",
          6273 => x"70",
          6274 => x"65",
          6275 => x"25",
          6276 => x"20",
          6277 => x"58",
          6278 => x"3f",
          6279 => x"00",
          6280 => x"25",
          6281 => x"20",
          6282 => x"58",
          6283 => x"25",
          6284 => x"20",
          6285 => x"58",
          6286 => x"44",
          6287 => x"62",
          6288 => x"67",
          6289 => x"74",
          6290 => x"75",
          6291 => x"0a",
          6292 => x"45",
          6293 => x"6c",
          6294 => x"20",
          6295 => x"65",
          6296 => x"70",
          6297 => x"00",
          6298 => x"44",
          6299 => x"62",
          6300 => x"20",
          6301 => x"74",
          6302 => x"66",
          6303 => x"45",
          6304 => x"6c",
          6305 => x"20",
          6306 => x"74",
          6307 => x"66",
          6308 => x"45",
          6309 => x"75",
          6310 => x"67",
          6311 => x"64",
          6312 => x"20",
          6313 => x"78",
          6314 => x"2e",
          6315 => x"43",
          6316 => x"69",
          6317 => x"63",
          6318 => x"20",
          6319 => x"30",
          6320 => x"2e",
          6321 => x"00",
          6322 => x"43",
          6323 => x"20",
          6324 => x"75",
          6325 => x"64",
          6326 => x"64",
          6327 => x"25",
          6328 => x"0a",
          6329 => x"52",
          6330 => x"61",
          6331 => x"6e",
          6332 => x"70",
          6333 => x"63",
          6334 => x"6f",
          6335 => x"2e",
          6336 => x"43",
          6337 => x"20",
          6338 => x"6f",
          6339 => x"6e",
          6340 => x"2e",
          6341 => x"5a",
          6342 => x"62",
          6343 => x"25",
          6344 => x"25",
          6345 => x"73",
          6346 => x"00",
          6347 => x"42",
          6348 => x"63",
          6349 => x"61",
          6350 => x"0a",
          6351 => x"52",
          6352 => x"69",
          6353 => x"2e",
          6354 => x"45",
          6355 => x"6c",
          6356 => x"20",
          6357 => x"65",
          6358 => x"70",
          6359 => x"2e",
          6360 => x"00",
          6361 => x"00",
          6362 => x"00",
          6363 => x"00",
          6364 => x"00",
          6365 => x"00",
          6366 => x"00",
          6367 => x"00",
          6368 => x"00",
          6369 => x"00",
          6370 => x"00",
          6371 => x"05",
          6372 => x"00",
          6373 => x"01",
          6374 => x"80",
          6375 => x"01",
          6376 => x"00",
          6377 => x"01",
          6378 => x"00",
          6379 => x"01",
          6380 => x"00",
          6381 => x"00",
          6382 => x"00",
          6383 => x"01",
          6384 => x"00",
          6385 => x"00",
          6386 => x"00",
          6387 => x"01",
          6388 => x"00",
          6389 => x"00",
          6390 => x"00",
          6391 => x"01",
          6392 => x"00",
          6393 => x"00",
          6394 => x"00",
          6395 => x"01",
          6396 => x"00",
          6397 => x"00",
          6398 => x"00",
          6399 => x"01",
          6400 => x"00",
          6401 => x"00",
          6402 => x"00",
          6403 => x"01",
          6404 => x"00",
          6405 => x"00",
          6406 => x"00",
          6407 => x"01",
          6408 => x"00",
          6409 => x"00",
          6410 => x"00",
          6411 => x"01",
          6412 => x"00",
          6413 => x"00",
          6414 => x"00",
          6415 => x"01",
          6416 => x"00",
          6417 => x"00",
          6418 => x"00",
          6419 => x"01",
          6420 => x"00",
          6421 => x"00",
          6422 => x"00",
          6423 => x"01",
          6424 => x"00",
          6425 => x"00",
          6426 => x"00",
          6427 => x"01",
          6428 => x"00",
          6429 => x"00",
          6430 => x"00",
          6431 => x"01",
          6432 => x"00",
          6433 => x"00",
          6434 => x"00",
          6435 => x"01",
          6436 => x"00",
          6437 => x"00",
          6438 => x"00",
          6439 => x"01",
          6440 => x"00",
          6441 => x"00",
          6442 => x"00",
          6443 => x"01",
          6444 => x"00",
          6445 => x"00",
          6446 => x"00",
          6447 => x"01",
          6448 => x"00",
          6449 => x"00",
          6450 => x"00",
          6451 => x"01",
          6452 => x"00",
          6453 => x"00",
          6454 => x"00",
          6455 => x"01",
          6456 => x"00",
          6457 => x"00",
          6458 => x"00",
          6459 => x"01",
          6460 => x"00",
          6461 => x"00",
          6462 => x"00",
          6463 => x"01",
          6464 => x"00",
          6465 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
