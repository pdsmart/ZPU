-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87fa",
          2049 => x"f80d0b0b",
          2050 => x"0b93ed04",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"d1040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b93b4",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b82b7",
          2210 => x"ec738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93b90400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80d2",
          2219 => x"fe2d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80cd",
          2227 => x"fc2d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"96040b0b",
          2317 => x"0b8ca604",
          2318 => x"0b0b0b8c",
          2319 => x"b6040b0b",
          2320 => x"0b8cc604",
          2321 => x"0b0b0b8c",
          2322 => x"d6040b0b",
          2323 => x"0b8ce604",
          2324 => x"0b0b0b8c",
          2325 => x"f7040b0b",
          2326 => x"0b8d8804",
          2327 => x"0b0b0b8d",
          2328 => x"98040b0b",
          2329 => x"0b8da804",
          2330 => x"0b0b0b8d",
          2331 => x"b8040b0b",
          2332 => x"0b8dc904",
          2333 => x"0b0b0b8d",
          2334 => x"da040b0b",
          2335 => x"0b8deb04",
          2336 => x"0b0b0b8d",
          2337 => x"fc040b0b",
          2338 => x"0b8e8d04",
          2339 => x"0b0b0b8e",
          2340 => x"9e040b0b",
          2341 => x"0b8eaf04",
          2342 => x"0b0b0b8e",
          2343 => x"c0040b0b",
          2344 => x"0b8ed104",
          2345 => x"0b0b0b8e",
          2346 => x"e2040b0b",
          2347 => x"0b8ef304",
          2348 => x"0b0b0b8f",
          2349 => x"84040b0b",
          2350 => x"0b8f9504",
          2351 => x"0b0b0b8f",
          2352 => x"a6040b0b",
          2353 => x"0b8fb704",
          2354 => x"0b0b0b8f",
          2355 => x"c8040b0b",
          2356 => x"0b8fd904",
          2357 => x"0b0b0b8f",
          2358 => x"ea040b0b",
          2359 => x"0b8ffb04",
          2360 => x"0b0b0b90",
          2361 => x"8c040b0b",
          2362 => x"0b909d04",
          2363 => x"0b0b0b90",
          2364 => x"ae040b0b",
          2365 => x"0b90bf04",
          2366 => x"0b0b0b90",
          2367 => x"d0040b0b",
          2368 => x"0b90e104",
          2369 => x"0b0b0b90",
          2370 => x"f2040b0b",
          2371 => x"0b918304",
          2372 => x"0b0b0b91",
          2373 => x"94040b0b",
          2374 => x"0b91a504",
          2375 => x"0b0b0b91",
          2376 => x"b6040b0b",
          2377 => x"0b91c704",
          2378 => x"0b0b0b91",
          2379 => x"d8040b0b",
          2380 => x"0b91e904",
          2381 => x"0b0b0b91",
          2382 => x"fa040b0b",
          2383 => x"0b928b04",
          2384 => x"0b0b0b92",
          2385 => x"9c040b0b",
          2386 => x"0b92ad04",
          2387 => x"0b0b0b92",
          2388 => x"be040b0b",
          2389 => x"0b92cf04",
          2390 => x"0b0b0b92",
          2391 => x"e0040b0b",
          2392 => x"0b92f104",
          2393 => x"0b0b0b93",
          2394 => x"8204ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482e0a4",
          2434 => x"0c81818b",
          2435 => x"2d82e0a4",
          2436 => x"0880c080",
          2437 => x"900482e0",
          2438 => x"a40cb3e6",
          2439 => x"2d82e0a4",
          2440 => x"0880c080",
          2441 => x"900482e0",
          2442 => x"a40cb097",
          2443 => x"2d82e0a4",
          2444 => x"0880c080",
          2445 => x"900482e0",
          2446 => x"a40cafe1",
          2447 => x"2d82e0a4",
          2448 => x"0880c080",
          2449 => x"900482e0",
          2450 => x"a40c94e1",
          2451 => x"2d82e0a4",
          2452 => x"0880c080",
          2453 => x"900482e0",
          2454 => x"a40cb1f6",
          2455 => x"2d82e0a4",
          2456 => x"0880c080",
          2457 => x"900482e0",
          2458 => x"a40c80da",
          2459 => x"9f2d82e0",
          2460 => x"a40880c0",
          2461 => x"80900482",
          2462 => x"e0a40c80",
          2463 => x"d4ce2d82",
          2464 => x"e0a40880",
          2465 => x"c0809004",
          2466 => x"82e0a40c",
          2467 => x"948c2d82",
          2468 => x"e0a40880",
          2469 => x"c0809004",
          2470 => x"82e0a40c",
          2471 => x"96f42d82",
          2472 => x"e0a40880",
          2473 => x"c0809004",
          2474 => x"82e0a40c",
          2475 => x"98812d82",
          2476 => x"e0a40880",
          2477 => x"c0809004",
          2478 => x"82e0a40c",
          2479 => x"80e0e72d",
          2480 => x"82e0a408",
          2481 => x"80c08090",
          2482 => x"0482e0a4",
          2483 => x"0c80fff6",
          2484 => x"2d82e0a4",
          2485 => x"0880c080",
          2486 => x"900482e0",
          2487 => x"a40c8180",
          2488 => x"dd2d82e0",
          2489 => x"a40880c0",
          2490 => x"80900482",
          2491 => x"e0a40c80",
          2492 => x"fdb22d82",
          2493 => x"e0a40880",
          2494 => x"c0809004",
          2495 => x"82e0a40c",
          2496 => x"80fee52d",
          2497 => x"82e0a408",
          2498 => x"80c08090",
          2499 => x"0482e0a4",
          2500 => x"0c81f6a7",
          2501 => x"2d82e0a4",
          2502 => x"0880c080",
          2503 => x"900482e0",
          2504 => x"a40c8283",
          2505 => x"a72d82e0",
          2506 => x"a40880c0",
          2507 => x"80900482",
          2508 => x"e0a40c81",
          2509 => x"fb8c2d82",
          2510 => x"e0a40880",
          2511 => x"c0809004",
          2512 => x"82e0a40c",
          2513 => x"81fe8c2d",
          2514 => x"82e0a408",
          2515 => x"80c08090",
          2516 => x"0482e0a4",
          2517 => x"0c8288e5",
          2518 => x"2d82e0a4",
          2519 => x"0880c080",
          2520 => x"900482e0",
          2521 => x"a40c8291",
          2522 => x"ce2d82e0",
          2523 => x"a40880c0",
          2524 => x"80900482",
          2525 => x"e0a40c82",
          2526 => x"82842d82",
          2527 => x"e0a40880",
          2528 => x"c0809004",
          2529 => x"82e0a40c",
          2530 => x"828c882d",
          2531 => x"82e0a408",
          2532 => x"80c08090",
          2533 => x"0482e0a4",
          2534 => x"0c828da8",
          2535 => x"2d82e0a4",
          2536 => x"0880c080",
          2537 => x"900482e0",
          2538 => x"a40c828d",
          2539 => x"c72d82e0",
          2540 => x"a40880c0",
          2541 => x"80900482",
          2542 => x"e0a40c82",
          2543 => x"95bb2d82",
          2544 => x"e0a40880",
          2545 => x"c0809004",
          2546 => x"82e0a40c",
          2547 => x"82939d2d",
          2548 => x"82e0a408",
          2549 => x"80c08090",
          2550 => x"0482e0a4",
          2551 => x"0c829897",
          2552 => x"2d82e0a4",
          2553 => x"0880c080",
          2554 => x"900482e0",
          2555 => x"a40c828e",
          2556 => x"cd2d82e0",
          2557 => x"a40880c0",
          2558 => x"80900482",
          2559 => x"e0a40c82",
          2560 => x"9b9c2d82",
          2561 => x"e0a40880",
          2562 => x"c0809004",
          2563 => x"82e0a40c",
          2564 => x"829c9d2d",
          2565 => x"82e0a408",
          2566 => x"80c08090",
          2567 => x"0482e0a4",
          2568 => x"0c828487",
          2569 => x"2d82e0a4",
          2570 => x"0880c080",
          2571 => x"900482e0",
          2572 => x"a40c8283",
          2573 => x"e02d82e0",
          2574 => x"a40880c0",
          2575 => x"80900482",
          2576 => x"e0a40c82",
          2577 => x"858b2d82",
          2578 => x"e0a40880",
          2579 => x"c0809004",
          2580 => x"82e0a40c",
          2581 => x"828fa42d",
          2582 => x"82e0a408",
          2583 => x"80c08090",
          2584 => x"0482e0a4",
          2585 => x"0c829d8e",
          2586 => x"2d82e0a4",
          2587 => x"0880c080",
          2588 => x"900482e0",
          2589 => x"a40c829f",
          2590 => x"992d82e0",
          2591 => x"a40880c0",
          2592 => x"80900482",
          2593 => x"e0a40c82",
          2594 => x"a2a02d82",
          2595 => x"e0a40880",
          2596 => x"c0809004",
          2597 => x"82e0a40c",
          2598 => x"81f5c62d",
          2599 => x"82e0a408",
          2600 => x"80c08090",
          2601 => x"0482e0a4",
          2602 => x"0c82a58c",
          2603 => x"2d82e0a4",
          2604 => x"0880c080",
          2605 => x"900482e0",
          2606 => x"a40c82b4",
          2607 => x"e92d82e0",
          2608 => x"a40880c0",
          2609 => x"80900482",
          2610 => x"e0a40c82",
          2611 => x"b2d52d82",
          2612 => x"e0a40880",
          2613 => x"c0809004",
          2614 => x"82e0a40c",
          2615 => x"81b58b2d",
          2616 => x"82e0a408",
          2617 => x"80c08090",
          2618 => x"0482e0a4",
          2619 => x"0c81b6f5",
          2620 => x"2d82e0a4",
          2621 => x"0880c080",
          2622 => x"900482e0",
          2623 => x"a40c81b8",
          2624 => x"d92d82e0",
          2625 => x"a40880c0",
          2626 => x"80900482",
          2627 => x"e0a40c80",
          2628 => x"fbe42d82",
          2629 => x"e0a40880",
          2630 => x"c0809004",
          2631 => x"82e0a40c",
          2632 => x"80fd882d",
          2633 => x"82e0a408",
          2634 => x"80c08090",
          2635 => x"0482e0a4",
          2636 => x"0c818280",
          2637 => x"2d82e0a4",
          2638 => x"0880c080",
          2639 => x"900482e0",
          2640 => x"a40c80e0",
          2641 => x"ef2d82e0",
          2642 => x"a40880c0",
          2643 => x"80900482",
          2644 => x"e0a40c81",
          2645 => x"af9f2d82",
          2646 => x"e0a40880",
          2647 => x"c0809004",
          2648 => x"82e0a40c",
          2649 => x"81afc72d",
          2650 => x"82e0a408",
          2651 => x"80c08090",
          2652 => x"0482e0a4",
          2653 => x"0c81b3bf",
          2654 => x"2d82e0a4",
          2655 => x"0880c080",
          2656 => x"900482e0",
          2657 => x"a40c81ac",
          2658 => x"892d82e0",
          2659 => x"a40880c0",
          2660 => x"8090043c",
          2661 => x"04101010",
          2662 => x"10101010",
          2663 => x"10101010",
          2664 => x"10101010",
          2665 => x"10101010",
          2666 => x"10101010",
          2667 => x"10101010",
          2668 => x"10101010",
          2669 => x"53510400",
          2670 => x"007381ff",
          2671 => x"06738306",
          2672 => x"09810583",
          2673 => x"05101010",
          2674 => x"2b0772fc",
          2675 => x"060c5151",
          2676 => x"04727280",
          2677 => x"728106ff",
          2678 => x"05097206",
          2679 => x"05711052",
          2680 => x"720a100a",
          2681 => x"5372ed38",
          2682 => x"51515351",
          2683 => x"0482e098",
          2684 => x"7082fc84",
          2685 => x"278e3880",
          2686 => x"71708405",
          2687 => x"530c0b0b",
          2688 => x"0b93f004",
          2689 => x"8c815180",
          2690 => x"faa70400",
          2691 => x"82e0a408",
          2692 => x"0282e0a4",
          2693 => x"0cfb3d0d",
          2694 => x"82e0a408",
          2695 => x"8c057082",
          2696 => x"e0a408fc",
          2697 => x"050c82e0",
          2698 => x"a408fc05",
          2699 => x"085482e0",
          2700 => x"a4088805",
          2701 => x"085382fb",
          2702 => x"fc085254",
          2703 => x"849a3f82",
          2704 => x"e0980870",
          2705 => x"82e0a408",
          2706 => x"f8050c82",
          2707 => x"e0a408f8",
          2708 => x"05087082",
          2709 => x"e0980c51",
          2710 => x"54873d0d",
          2711 => x"82e0a40c",
          2712 => x"0482e0a4",
          2713 => x"080282e0",
          2714 => x"a40cfb3d",
          2715 => x"0d82e0a4",
          2716 => x"08900508",
          2717 => x"85113370",
          2718 => x"81327081",
          2719 => x"06515151",
          2720 => x"52718f38",
          2721 => x"800b82e0",
          2722 => x"a4088c05",
          2723 => x"08258338",
          2724 => x"8d39800b",
          2725 => x"82e0a408",
          2726 => x"f4050c81",
          2727 => x"c43982e0",
          2728 => x"a4088c05",
          2729 => x"08ff0582",
          2730 => x"e0a4088c",
          2731 => x"050c800b",
          2732 => x"82e0a408",
          2733 => x"f8050c82",
          2734 => x"e0a40888",
          2735 => x"050882e0",
          2736 => x"a408fc05",
          2737 => x"0c82e0a4",
          2738 => x"08f80508",
          2739 => x"8a2e80f6",
          2740 => x"38800b82",
          2741 => x"e0a4088c",
          2742 => x"05082580",
          2743 => x"e93882e0",
          2744 => x"a4089005",
          2745 => x"0851a090",
          2746 => x"3f82e098",
          2747 => x"087082e0",
          2748 => x"a408f805",
          2749 => x"0c5282e0",
          2750 => x"a408f805",
          2751 => x"08ff2e09",
          2752 => x"81068d38",
          2753 => x"800b82e0",
          2754 => x"a408f405",
          2755 => x"0c80d239",
          2756 => x"82e0a408",
          2757 => x"fc050882",
          2758 => x"e0a408f8",
          2759 => x"05085353",
          2760 => x"71733482",
          2761 => x"e0a4088c",
          2762 => x"0508ff05",
          2763 => x"82e0a408",
          2764 => x"8c050c82",
          2765 => x"e0a408fc",
          2766 => x"05088105",
          2767 => x"82e0a408",
          2768 => x"fc050cff",
          2769 => x"803982e0",
          2770 => x"a408fc05",
          2771 => x"08528072",
          2772 => x"3482e0a4",
          2773 => x"08880508",
          2774 => x"7082e0a4",
          2775 => x"08f4050c",
          2776 => x"5282e0a4",
          2777 => x"08f40508",
          2778 => x"82e0980c",
          2779 => x"873d0d82",
          2780 => x"e0a40c04",
          2781 => x"82e0a408",
          2782 => x"0282e0a4",
          2783 => x"0cf43d0d",
          2784 => x"860b82e0",
          2785 => x"a408e505",
          2786 => x"3482e0a4",
          2787 => x"08880508",
          2788 => x"82e0a408",
          2789 => x"e0050cfe",
          2790 => x"0a0b82e0",
          2791 => x"a408e805",
          2792 => x"0c82e0a4",
          2793 => x"08900570",
          2794 => x"82e0a408",
          2795 => x"fc050c82",
          2796 => x"e0a408fc",
          2797 => x"05085482",
          2798 => x"e0a4088c",
          2799 => x"05085382",
          2800 => x"e0a408e0",
          2801 => x"05705351",
          2802 => x"54818d3f",
          2803 => x"82e09808",
          2804 => x"7082e0a4",
          2805 => x"08dc050c",
          2806 => x"82e0a408",
          2807 => x"ec050882",
          2808 => x"e0a40888",
          2809 => x"05080551",
          2810 => x"54807434",
          2811 => x"82e0a408",
          2812 => x"dc050870",
          2813 => x"82e0980c",
          2814 => x"548e3d0d",
          2815 => x"82e0a40c",
          2816 => x"0482e0a4",
          2817 => x"080282e0",
          2818 => x"a40cfb3d",
          2819 => x"0d82e0a4",
          2820 => x"08900570",
          2821 => x"82e0a408",
          2822 => x"fc050c82",
          2823 => x"e0a408fc",
          2824 => x"05085482",
          2825 => x"e0a4088c",
          2826 => x"05085382",
          2827 => x"e0a40888",
          2828 => x"05085254",
          2829 => x"a33f82e0",
          2830 => x"98087082",
          2831 => x"e0a408f8",
          2832 => x"050c82e0",
          2833 => x"a408f805",
          2834 => x"087082e0",
          2835 => x"980c5154",
          2836 => x"873d0d82",
          2837 => x"e0a40c04",
          2838 => x"82e0a408",
          2839 => x"0282e0a4",
          2840 => x"0ced3d0d",
          2841 => x"800b82e0",
          2842 => x"a408e405",
          2843 => x"2382e0a4",
          2844 => x"08880508",
          2845 => x"53800b8c",
          2846 => x"140c82e0",
          2847 => x"a4088805",
          2848 => x"08851133",
          2849 => x"70812a70",
          2850 => x"81327081",
          2851 => x"06515151",
          2852 => x"51537280",
          2853 => x"2e8d38ff",
          2854 => x"0b82e0a4",
          2855 => x"08e0050c",
          2856 => x"96ac3982",
          2857 => x"e0a4088c",
          2858 => x"05085372",
          2859 => x"33537282",
          2860 => x"e0a408f8",
          2861 => x"05347281",
          2862 => x"ff065372",
          2863 => x"802e95fa",
          2864 => x"3882e0a4",
          2865 => x"088c0508",
          2866 => x"810582e0",
          2867 => x"a4088c05",
          2868 => x"0c82e0a4",
          2869 => x"08e40522",
          2870 => x"70810651",
          2871 => x"5372802e",
          2872 => x"958b3882",
          2873 => x"e0a408f8",
          2874 => x"053353af",
          2875 => x"732781fc",
          2876 => x"3882e0a4",
          2877 => x"08f80533",
          2878 => x"5372b926",
          2879 => x"81ee3882",
          2880 => x"e0a408f8",
          2881 => x"05335372",
          2882 => x"b02e0981",
          2883 => x"0680c538",
          2884 => x"82e0a408",
          2885 => x"e8053370",
          2886 => x"982b7098",
          2887 => x"2c515153",
          2888 => x"72b23882",
          2889 => x"e0a408e4",
          2890 => x"05227083",
          2891 => x"2a708132",
          2892 => x"70810651",
          2893 => x"51515372",
          2894 => x"802e9938",
          2895 => x"82e0a408",
          2896 => x"e4052270",
          2897 => x"82800751",
          2898 => x"537282e0",
          2899 => x"a408e405",
          2900 => x"23fed039",
          2901 => x"82e0a408",
          2902 => x"e8053370",
          2903 => x"982b7098",
          2904 => x"2c707083",
          2905 => x"2b721173",
          2906 => x"11515151",
          2907 => x"53515553",
          2908 => x"7282e0a4",
          2909 => x"08e80534",
          2910 => x"82e0a408",
          2911 => x"e8053354",
          2912 => x"82e0a408",
          2913 => x"f8053370",
          2914 => x"15d01151",
          2915 => x"51537282",
          2916 => x"e0a408e8",
          2917 => x"053482e0",
          2918 => x"a408e805",
          2919 => x"3370982b",
          2920 => x"70982c51",
          2921 => x"51537280",
          2922 => x"258b3880",
          2923 => x"ff0b82e0",
          2924 => x"a408e805",
          2925 => x"3482e0a4",
          2926 => x"08e40522",
          2927 => x"70832a70",
          2928 => x"81065151",
          2929 => x"5372fddb",
          2930 => x"3882e0a4",
          2931 => x"08e80533",
          2932 => x"70882b70",
          2933 => x"902b7090",
          2934 => x"2c70882c",
          2935 => x"51515151",
          2936 => x"537282e0",
          2937 => x"a408ec05",
          2938 => x"23fdb839",
          2939 => x"82e0a408",
          2940 => x"e4052270",
          2941 => x"832a7081",
          2942 => x"06515153",
          2943 => x"72802e9d",
          2944 => x"3882e0a4",
          2945 => x"08e80533",
          2946 => x"70982b70",
          2947 => x"982c5151",
          2948 => x"53728a38",
          2949 => x"810b82e0",
          2950 => x"a408e805",
          2951 => x"3482e0a4",
          2952 => x"08f80533",
          2953 => x"e01182e0",
          2954 => x"a408c405",
          2955 => x"0c5382e0",
          2956 => x"a408c405",
          2957 => x"0880d826",
          2958 => x"92943882",
          2959 => x"e0a408c4",
          2960 => x"05087082",
          2961 => x"2b82b9dc",
          2962 => x"11700851",
          2963 => x"51515372",
          2964 => x"0482e0a4",
          2965 => x"08e40522",
          2966 => x"70900751",
          2967 => x"537282e0",
          2968 => x"a408e405",
          2969 => x"2382e0a4",
          2970 => x"08e40522",
          2971 => x"70a00751",
          2972 => x"537282e0",
          2973 => x"a408e405",
          2974 => x"23fca839",
          2975 => x"82e0a408",
          2976 => x"e4052270",
          2977 => x"81800751",
          2978 => x"537282e0",
          2979 => x"a408e405",
          2980 => x"23fc9039",
          2981 => x"82e0a408",
          2982 => x"e4052270",
          2983 => x"80c00751",
          2984 => x"537282e0",
          2985 => x"a408e405",
          2986 => x"23fbf839",
          2987 => x"82e0a408",
          2988 => x"e4052270",
          2989 => x"88075153",
          2990 => x"7282e0a4",
          2991 => x"08e40523",
          2992 => x"800b82e0",
          2993 => x"a408e805",
          2994 => x"34fbd839",
          2995 => x"82e0a408",
          2996 => x"e4052270",
          2997 => x"84075153",
          2998 => x"7282e0a4",
          2999 => x"08e40523",
          3000 => x"fbc139bf",
          3001 => x"0b82e0a4",
          3002 => x"08fc0534",
          3003 => x"82e0a408",
          3004 => x"ec0522ff",
          3005 => x"11515372",
          3006 => x"82e0a408",
          3007 => x"ec052380",
          3008 => x"e30b82e0",
          3009 => x"a408f805",
          3010 => x"348da839",
          3011 => x"82e0a408",
          3012 => x"90050882",
          3013 => x"e0a40890",
          3014 => x"05088405",
          3015 => x"82e0a408",
          3016 => x"90050c70",
          3017 => x"08515372",
          3018 => x"82e0a408",
          3019 => x"fc053482",
          3020 => x"e0a408ec",
          3021 => x"0522ff11",
          3022 => x"51537282",
          3023 => x"e0a408ec",
          3024 => x"05238cef",
          3025 => x"3982e0a4",
          3026 => x"08900508",
          3027 => x"82e0a408",
          3028 => x"90050884",
          3029 => x"0582e0a4",
          3030 => x"0890050c",
          3031 => x"700882e0",
          3032 => x"a408fc05",
          3033 => x"0c82e0a4",
          3034 => x"08e40522",
          3035 => x"70832a70",
          3036 => x"81065151",
          3037 => x"51537280",
          3038 => x"2eab3882",
          3039 => x"e0a408e8",
          3040 => x"05337098",
          3041 => x"2b537298",
          3042 => x"2c5382e0",
          3043 => x"a408fc05",
          3044 => x"085253a4",
          3045 => x"833f82e0",
          3046 => x"98085372",
          3047 => x"82e0a408",
          3048 => x"f4052399",
          3049 => x"3982e0a4",
          3050 => x"08fc0508",
          3051 => x"519d8a3f",
          3052 => x"82e09808",
          3053 => x"537282e0",
          3054 => x"a408f405",
          3055 => x"2382e0a4",
          3056 => x"08ec0522",
          3057 => x"5382e0a4",
          3058 => x"08f40522",
          3059 => x"73713154",
          3060 => x"547282e0",
          3061 => x"a408ec05",
          3062 => x"238bd839",
          3063 => x"82e0a408",
          3064 => x"90050882",
          3065 => x"e0a40890",
          3066 => x"05088405",
          3067 => x"82e0a408",
          3068 => x"90050c70",
          3069 => x"0882e0a4",
          3070 => x"08fc050c",
          3071 => x"82e0a408",
          3072 => x"e4052270",
          3073 => x"832a7081",
          3074 => x"06515151",
          3075 => x"5372802e",
          3076 => x"ab3882e0",
          3077 => x"a408e805",
          3078 => x"3370982b",
          3079 => x"5372982c",
          3080 => x"5382e0a4",
          3081 => x"08fc0508",
          3082 => x"5253a2ec",
          3083 => x"3f82e098",
          3084 => x"08537282",
          3085 => x"e0a408f4",
          3086 => x"05239939",
          3087 => x"82e0a408",
          3088 => x"fc050851",
          3089 => x"9bf33f82",
          3090 => x"e0980853",
          3091 => x"7282e0a4",
          3092 => x"08f40523",
          3093 => x"82e0a408",
          3094 => x"ec052253",
          3095 => x"82e0a408",
          3096 => x"f4052273",
          3097 => x"71315454",
          3098 => x"7282e0a4",
          3099 => x"08ec0523",
          3100 => x"8ac13982",
          3101 => x"e0a408e4",
          3102 => x"05227082",
          3103 => x"2a708106",
          3104 => x"51515372",
          3105 => x"802ea438",
          3106 => x"82e0a408",
          3107 => x"90050882",
          3108 => x"e0a40890",
          3109 => x"05088405",
          3110 => x"82e0a408",
          3111 => x"90050c70",
          3112 => x"0882e0a4",
          3113 => x"08dc050c",
          3114 => x"53a23982",
          3115 => x"e0a40890",
          3116 => x"050882e0",
          3117 => x"a4089005",
          3118 => x"08840582",
          3119 => x"e0a40890",
          3120 => x"050c7008",
          3121 => x"82e0a408",
          3122 => x"dc050c53",
          3123 => x"82e0a408",
          3124 => x"dc050882",
          3125 => x"e0a408fc",
          3126 => x"050c82e0",
          3127 => x"a408fc05",
          3128 => x"088025a4",
          3129 => x"3882e0a4",
          3130 => x"08e40522",
          3131 => x"70820751",
          3132 => x"537282e0",
          3133 => x"a408e405",
          3134 => x"2382e0a4",
          3135 => x"08fc0508",
          3136 => x"3082e0a4",
          3137 => x"08fc050c",
          3138 => x"82e0a408",
          3139 => x"e4052270",
          3140 => x"ffbf0651",
          3141 => x"537282e0",
          3142 => x"a408e405",
          3143 => x"2381af39",
          3144 => x"880b82e0",
          3145 => x"a408f405",
          3146 => x"23a93982",
          3147 => x"e0a408e4",
          3148 => x"05227080",
          3149 => x"c0075153",
          3150 => x"7282e0a4",
          3151 => x"08e40523",
          3152 => x"80f80b82",
          3153 => x"e0a408f8",
          3154 => x"0534900b",
          3155 => x"82e0a408",
          3156 => x"f4052382",
          3157 => x"e0a408e4",
          3158 => x"05227082",
          3159 => x"2a708106",
          3160 => x"51515372",
          3161 => x"802ea438",
          3162 => x"82e0a408",
          3163 => x"90050882",
          3164 => x"e0a40890",
          3165 => x"05088405",
          3166 => x"82e0a408",
          3167 => x"90050c70",
          3168 => x"0882e0a4",
          3169 => x"08d8050c",
          3170 => x"53a23982",
          3171 => x"e0a40890",
          3172 => x"050882e0",
          3173 => x"a4089005",
          3174 => x"08840582",
          3175 => x"e0a40890",
          3176 => x"050c7008",
          3177 => x"82e0a408",
          3178 => x"d8050c53",
          3179 => x"82e0a408",
          3180 => x"d8050882",
          3181 => x"e0a408fc",
          3182 => x"050c82e0",
          3183 => x"a408e405",
          3184 => x"2270cf06",
          3185 => x"51537282",
          3186 => x"e0a408e4",
          3187 => x"052382e0",
          3188 => x"a80b82e0",
          3189 => x"a408f005",
          3190 => x"0c82e0a4",
          3191 => x"08f00508",
          3192 => x"82e0a408",
          3193 => x"f4052282",
          3194 => x"e0a408fc",
          3195 => x"05087155",
          3196 => x"70545654",
          3197 => x"55aaca3f",
          3198 => x"82e09808",
          3199 => x"53727534",
          3200 => x"82e0a408",
          3201 => x"f0050882",
          3202 => x"e0a408d4",
          3203 => x"050c82e0",
          3204 => x"a408f005",
          3205 => x"08703351",
          3206 => x"53897327",
          3207 => x"a43882e0",
          3208 => x"a408f005",
          3209 => x"08537233",
          3210 => x"5482e0a4",
          3211 => x"08f80533",
          3212 => x"7015df11",
          3213 => x"51515372",
          3214 => x"82e0a408",
          3215 => x"d0053497",
          3216 => x"3982e0a4",
          3217 => x"08f00508",
          3218 => x"537233b0",
          3219 => x"11515372",
          3220 => x"82e0a408",
          3221 => x"d0053482",
          3222 => x"e0a408d4",
          3223 => x"05085382",
          3224 => x"e0a408d0",
          3225 => x"05337334",
          3226 => x"82e0a408",
          3227 => x"f0050881",
          3228 => x"0582e0a4",
          3229 => x"08f0050c",
          3230 => x"82e0a408",
          3231 => x"f4052270",
          3232 => x"5382e0a4",
          3233 => x"08fc0508",
          3234 => x"5253a0c7",
          3235 => x"3f82e098",
          3236 => x"087082e0",
          3237 => x"a408fc05",
          3238 => x"0c5382e0",
          3239 => x"a408fc05",
          3240 => x"08802e84",
          3241 => x"38feb239",
          3242 => x"82e0a408",
          3243 => x"f0050882",
          3244 => x"e0a85455",
          3245 => x"72547470",
          3246 => x"75315153",
          3247 => x"7282e0a4",
          3248 => x"08fc0534",
          3249 => x"82e0a408",
          3250 => x"e4052270",
          3251 => x"b2065153",
          3252 => x"72802e94",
          3253 => x"3882e0a4",
          3254 => x"08ec0522",
          3255 => x"ff115153",
          3256 => x"7282e0a4",
          3257 => x"08ec0523",
          3258 => x"82e0a408",
          3259 => x"e4052270",
          3260 => x"862a7081",
          3261 => x"06515153",
          3262 => x"72802e80",
          3263 => x"e73882e0",
          3264 => x"a408ec05",
          3265 => x"2270902b",
          3266 => x"82e0a408",
          3267 => x"cc050c82",
          3268 => x"e0a408cc",
          3269 => x"0508902c",
          3270 => x"82e0a408",
          3271 => x"cc050c82",
          3272 => x"e0a408f4",
          3273 => x"05225153",
          3274 => x"72902e09",
          3275 => x"81069538",
          3276 => x"82e0a408",
          3277 => x"cc0508fe",
          3278 => x"05537282",
          3279 => x"e0a408c8",
          3280 => x"05239339",
          3281 => x"82e0a408",
          3282 => x"cc0508ff",
          3283 => x"05537282",
          3284 => x"e0a408c8",
          3285 => x"052382e0",
          3286 => x"a408c805",
          3287 => x"2282e0a4",
          3288 => x"08ec0523",
          3289 => x"82e0a408",
          3290 => x"e4052270",
          3291 => x"832a7081",
          3292 => x"06515153",
          3293 => x"72802e80",
          3294 => x"d03882e0",
          3295 => x"a408e805",
          3296 => x"3370982b",
          3297 => x"70982c82",
          3298 => x"e0a408fc",
          3299 => x"05335751",
          3300 => x"51537274",
          3301 => x"24973882",
          3302 => x"e0a408e4",
          3303 => x"052270f7",
          3304 => x"06515372",
          3305 => x"82e0a408",
          3306 => x"e405239d",
          3307 => x"3982e0a4",
          3308 => x"08e80533",
          3309 => x"5382e0a4",
          3310 => x"08fc0533",
          3311 => x"73713154",
          3312 => x"547282e0",
          3313 => x"a408e805",
          3314 => x"3482e0a4",
          3315 => x"08e40522",
          3316 => x"70832a70",
          3317 => x"81065151",
          3318 => x"5372802e",
          3319 => x"b13882e0",
          3320 => x"a408e805",
          3321 => x"3370882b",
          3322 => x"70902b70",
          3323 => x"902c7088",
          3324 => x"2c515151",
          3325 => x"51537254",
          3326 => x"82e0a408",
          3327 => x"ec052270",
          3328 => x"75315153",
          3329 => x"7282e0a4",
          3330 => x"08ec0523",
          3331 => x"af3982e0",
          3332 => x"a408fc05",
          3333 => x"3370882b",
          3334 => x"70902b70",
          3335 => x"902c7088",
          3336 => x"2c515151",
          3337 => x"51537254",
          3338 => x"82e0a408",
          3339 => x"ec052270",
          3340 => x"75315153",
          3341 => x"7282e0a4",
          3342 => x"08ec0523",
          3343 => x"82e0a408",
          3344 => x"e4052270",
          3345 => x"83800651",
          3346 => x"5372b038",
          3347 => x"82e0a408",
          3348 => x"ec0522ff",
          3349 => x"11545472",
          3350 => x"82e0a408",
          3351 => x"ec052373",
          3352 => x"902b7090",
          3353 => x"2c515380",
          3354 => x"73259038",
          3355 => x"82e0a408",
          3356 => x"88050852",
          3357 => x"a0518aee",
          3358 => x"3fd23982",
          3359 => x"e0a408e4",
          3360 => x"05227081",
          3361 => x"2a708106",
          3362 => x"51515372",
          3363 => x"802e9138",
          3364 => x"82e0a408",
          3365 => x"88050852",
          3366 => x"ad518aca",
          3367 => x"3f80c739",
          3368 => x"82e0a408",
          3369 => x"e4052270",
          3370 => x"842a7081",
          3371 => x"06515153",
          3372 => x"72802e90",
          3373 => x"3882e0a4",
          3374 => x"08880508",
          3375 => x"52ab518a",
          3376 => x"a53fa339",
          3377 => x"82e0a408",
          3378 => x"e4052270",
          3379 => x"852a7081",
          3380 => x"06515153",
          3381 => x"72802e8e",
          3382 => x"3882e0a4",
          3383 => x"08880508",
          3384 => x"52a0518a",
          3385 => x"813f82e0",
          3386 => x"a408e405",
          3387 => x"2270862a",
          3388 => x"70810651",
          3389 => x"51537280",
          3390 => x"2eb13882",
          3391 => x"e0a40888",
          3392 => x"050852b0",
          3393 => x"5189df3f",
          3394 => x"82e0a408",
          3395 => x"f4052253",
          3396 => x"72902e09",
          3397 => x"81069438",
          3398 => x"82e0a408",
          3399 => x"88050852",
          3400 => x"82e0a408",
          3401 => x"f8053351",
          3402 => x"89bc3f82",
          3403 => x"e0a408e4",
          3404 => x"05227088",
          3405 => x"2a708106",
          3406 => x"51515372",
          3407 => x"802eb038",
          3408 => x"82e0a408",
          3409 => x"ec0522ff",
          3410 => x"11545472",
          3411 => x"82e0a408",
          3412 => x"ec052373",
          3413 => x"902b7090",
          3414 => x"2c515380",
          3415 => x"73259038",
          3416 => x"82e0a408",
          3417 => x"88050852",
          3418 => x"b05188fa",
          3419 => x"3fd23982",
          3420 => x"e0a408e4",
          3421 => x"05227083",
          3422 => x"2a708106",
          3423 => x"51515372",
          3424 => x"802eb038",
          3425 => x"82e0a408",
          3426 => x"e80533ff",
          3427 => x"11545472",
          3428 => x"82e0a408",
          3429 => x"e8053473",
          3430 => x"982b7098",
          3431 => x"2c515380",
          3432 => x"73259038",
          3433 => x"82e0a408",
          3434 => x"88050852",
          3435 => x"b05188b6",
          3436 => x"3fd23982",
          3437 => x"e0a408e4",
          3438 => x"05227087",
          3439 => x"2a708106",
          3440 => x"51515372",
          3441 => x"b03882e0",
          3442 => x"a408ec05",
          3443 => x"22ff1154",
          3444 => x"547282e0",
          3445 => x"a408ec05",
          3446 => x"2373902b",
          3447 => x"70902c51",
          3448 => x"53807325",
          3449 => x"903882e0",
          3450 => x"a4088805",
          3451 => x"0852a051",
          3452 => x"87f43fd2",
          3453 => x"3982e0a4",
          3454 => x"08f80533",
          3455 => x"537280e3",
          3456 => x"2e098106",
          3457 => x"973882e0",
          3458 => x"a4088805",
          3459 => x"085282e0",
          3460 => x"a408fc05",
          3461 => x"335187ce",
          3462 => x"3f81ee39",
          3463 => x"82e0a408",
          3464 => x"f8053353",
          3465 => x"7280f32e",
          3466 => x"09810680",
          3467 => x"cb3882e0",
          3468 => x"a408f405",
          3469 => x"22ff1151",
          3470 => x"537282e0",
          3471 => x"a408f405",
          3472 => x"237283ff",
          3473 => x"ff065372",
          3474 => x"83ffff2e",
          3475 => x"81bb3882",
          3476 => x"e0a40888",
          3477 => x"05085282",
          3478 => x"e0a408fc",
          3479 => x"05087033",
          3480 => x"5282e0a4",
          3481 => x"08fc0508",
          3482 => x"810582e0",
          3483 => x"a408fc05",
          3484 => x"0c5386f2",
          3485 => x"3fffb739",
          3486 => x"82e0a408",
          3487 => x"f8053353",
          3488 => x"7280d32e",
          3489 => x"09810680",
          3490 => x"cb3882e0",
          3491 => x"a408f405",
          3492 => x"22ff1151",
          3493 => x"537282e0",
          3494 => x"a408f405",
          3495 => x"237283ff",
          3496 => x"ff065372",
          3497 => x"83ffff2e",
          3498 => x"80df3882",
          3499 => x"e0a40888",
          3500 => x"05085282",
          3501 => x"e0a408fc",
          3502 => x"05087033",
          3503 => x"525386a6",
          3504 => x"3f82e0a4",
          3505 => x"08fc0508",
          3506 => x"810582e0",
          3507 => x"a408fc05",
          3508 => x"0cffb739",
          3509 => x"82e0a408",
          3510 => x"f0050882",
          3511 => x"e0a82ea9",
          3512 => x"3882e0a4",
          3513 => x"08880508",
          3514 => x"5282e0a4",
          3515 => x"08f00508",
          3516 => x"ff0582e0",
          3517 => x"a408f005",
          3518 => x"0c82e0a4",
          3519 => x"08f00508",
          3520 => x"70335253",
          3521 => x"85e03fcc",
          3522 => x"3982e0a4",
          3523 => x"08e40522",
          3524 => x"70872a70",
          3525 => x"81065151",
          3526 => x"5372802e",
          3527 => x"80c33882",
          3528 => x"e0a408ec",
          3529 => x"0522ff11",
          3530 => x"54547282",
          3531 => x"e0a408ec",
          3532 => x"05237390",
          3533 => x"2b70902c",
          3534 => x"51538073",
          3535 => x"25a33882",
          3536 => x"e0a40888",
          3537 => x"050852a0",
          3538 => x"51859b3f",
          3539 => x"d23982e0",
          3540 => x"a4088805",
          3541 => x"085282e0",
          3542 => x"a408f805",
          3543 => x"33518586",
          3544 => x"3f800b82",
          3545 => x"e0a408e4",
          3546 => x"0523eab7",
          3547 => x"3982e0a4",
          3548 => x"08f80533",
          3549 => x"5372a52e",
          3550 => x"098106a8",
          3551 => x"38810b82",
          3552 => x"e0a408e4",
          3553 => x"0523800b",
          3554 => x"82e0a408",
          3555 => x"ec052380",
          3556 => x"0b82e0a4",
          3557 => x"08e80534",
          3558 => x"8a0b82e0",
          3559 => x"a408f405",
          3560 => x"23ea8039",
          3561 => x"82e0a408",
          3562 => x"88050852",
          3563 => x"82e0a408",
          3564 => x"f8053351",
          3565 => x"84b03fe9",
          3566 => x"ea3982e0",
          3567 => x"a4088805",
          3568 => x"088c1108",
          3569 => x"7082e0a4",
          3570 => x"08e0050c",
          3571 => x"515382e0",
          3572 => x"a408e005",
          3573 => x"0882e098",
          3574 => x"0c953d0d",
          3575 => x"82e0a40c",
          3576 => x"0482e0a4",
          3577 => x"080282e0",
          3578 => x"a40cfd3d",
          3579 => x"0d82fbf8",
          3580 => x"085382e0",
          3581 => x"a4088c05",
          3582 => x"085282e0",
          3583 => x"a4088805",
          3584 => x"0851e4dd",
          3585 => x"3f82e098",
          3586 => x"087082e0",
          3587 => x"980c5485",
          3588 => x"3d0d82e0",
          3589 => x"a40c0482",
          3590 => x"e0a40802",
          3591 => x"82e0a40c",
          3592 => x"fb3d0d80",
          3593 => x"0b82e0a4",
          3594 => x"08f8050c",
          3595 => x"82fbfc08",
          3596 => x"85113370",
          3597 => x"812a7081",
          3598 => x"32708106",
          3599 => x"51515151",
          3600 => x"5372802e",
          3601 => x"8d38ff0b",
          3602 => x"82e0a408",
          3603 => x"f4050c81",
          3604 => x"923982e0",
          3605 => x"a4088805",
          3606 => x"08537233",
          3607 => x"82e0a408",
          3608 => x"88050881",
          3609 => x"0582e0a4",
          3610 => x"0888050c",
          3611 => x"537282e0",
          3612 => x"a408fc05",
          3613 => x"347281ff",
          3614 => x"06537280",
          3615 => x"2eb03882",
          3616 => x"fbfc0882",
          3617 => x"fbfc0853",
          3618 => x"82e0a408",
          3619 => x"fc053352",
          3620 => x"90110851",
          3621 => x"53722d82",
          3622 => x"e0980853",
          3623 => x"72802eff",
          3624 => x"b138ff0b",
          3625 => x"82e0a408",
          3626 => x"f8050cff",
          3627 => x"a53982fb",
          3628 => x"fc0882fb",
          3629 => x"fc085353",
          3630 => x"8a519013",
          3631 => x"0853722d",
          3632 => x"82e09808",
          3633 => x"5372802e",
          3634 => x"8a38ff0b",
          3635 => x"82e0a408",
          3636 => x"f8050c82",
          3637 => x"e0a408f8",
          3638 => x"05087082",
          3639 => x"e0a408f4",
          3640 => x"050c5382",
          3641 => x"e0a408f4",
          3642 => x"050882e0",
          3643 => x"980c873d",
          3644 => x"0d82e0a4",
          3645 => x"0c0482e0",
          3646 => x"a4080282",
          3647 => x"e0a40cfb",
          3648 => x"3d0d800b",
          3649 => x"82e0a408",
          3650 => x"f8050c82",
          3651 => x"e0a4088c",
          3652 => x"05088511",
          3653 => x"3370812a",
          3654 => x"70813270",
          3655 => x"81065151",
          3656 => x"51515372",
          3657 => x"802e8d38",
          3658 => x"ff0b82e0",
          3659 => x"a408f405",
          3660 => x"0c80f339",
          3661 => x"82e0a408",
          3662 => x"88050853",
          3663 => x"723382e0",
          3664 => x"a4088805",
          3665 => x"08810582",
          3666 => x"e0a40888",
          3667 => x"050c5372",
          3668 => x"82e0a408",
          3669 => x"fc053472",
          3670 => x"81ff0653",
          3671 => x"72802eb6",
          3672 => x"3882e0a4",
          3673 => x"088c0508",
          3674 => x"82e0a408",
          3675 => x"8c050853",
          3676 => x"82e0a408",
          3677 => x"fc053352",
          3678 => x"90110851",
          3679 => x"53722d82",
          3680 => x"e0980853",
          3681 => x"72802eff",
          3682 => x"ab38ff0b",
          3683 => x"82e0a408",
          3684 => x"f8050cff",
          3685 => x"9f3982e0",
          3686 => x"a408f805",
          3687 => x"087082e0",
          3688 => x"a408f405",
          3689 => x"0c5382e0",
          3690 => x"a408f405",
          3691 => x"0882e098",
          3692 => x"0c873d0d",
          3693 => x"82e0a40c",
          3694 => x"0482e0a4",
          3695 => x"080282e0",
          3696 => x"a40cfe3d",
          3697 => x"0d82fbfc",
          3698 => x"085282e0",
          3699 => x"a4088805",
          3700 => x"0851933f",
          3701 => x"82e09808",
          3702 => x"7082e098",
          3703 => x"0c53843d",
          3704 => x"0d82e0a4",
          3705 => x"0c0482e0",
          3706 => x"a4080282",
          3707 => x"e0a40cfb",
          3708 => x"3d0d82e0",
          3709 => x"a4088c05",
          3710 => x"08851133",
          3711 => x"70812a70",
          3712 => x"81327081",
          3713 => x"06515151",
          3714 => x"51537280",
          3715 => x"2e8d38ff",
          3716 => x"0b82e0a4",
          3717 => x"08fc050c",
          3718 => x"81cb3982",
          3719 => x"e0a4088c",
          3720 => x"05088511",
          3721 => x"3370822a",
          3722 => x"70810651",
          3723 => x"51515372",
          3724 => x"802e80db",
          3725 => x"3882e0a4",
          3726 => x"088c0508",
          3727 => x"82e0a408",
          3728 => x"8c050854",
          3729 => x"548c1408",
          3730 => x"88140825",
          3731 => x"9f3882e0",
          3732 => x"a4088c05",
          3733 => x"08700870",
          3734 => x"82e0a408",
          3735 => x"88050852",
          3736 => x"57545472",
          3737 => x"75347308",
          3738 => x"8105740c",
          3739 => x"82e0a408",
          3740 => x"8c05088c",
          3741 => x"11088105",
          3742 => x"8c120c82",
          3743 => x"e0a40888",
          3744 => x"05087082",
          3745 => x"e0a408fc",
          3746 => x"050c5153",
          3747 => x"80d73982",
          3748 => x"e0a4088c",
          3749 => x"050882e0",
          3750 => x"a4088c05",
          3751 => x"085382e0",
          3752 => x"a4088805",
          3753 => x"087081ff",
          3754 => x"06539012",
          3755 => x"08515454",
          3756 => x"722d82e0",
          3757 => x"98085372",
          3758 => x"a33882e0",
          3759 => x"a4088c05",
          3760 => x"088c1108",
          3761 => x"81058c12",
          3762 => x"0c82e0a4",
          3763 => x"08880508",
          3764 => x"7082e0a4",
          3765 => x"08fc050c",
          3766 => x"51538a39",
          3767 => x"ff0b82e0",
          3768 => x"a408fc05",
          3769 => x"0c82e0a4",
          3770 => x"08fc0508",
          3771 => x"82e0980c",
          3772 => x"873d0d82",
          3773 => x"e0a40c04",
          3774 => x"82e0a408",
          3775 => x"0282e0a4",
          3776 => x"0cf93d0d",
          3777 => x"82e0a408",
          3778 => x"88050885",
          3779 => x"11337081",
          3780 => x"32708106",
          3781 => x"51515152",
          3782 => x"71802e8d",
          3783 => x"38ff0b82",
          3784 => x"e0a408f8",
          3785 => x"050c8394",
          3786 => x"3982e0a4",
          3787 => x"08880508",
          3788 => x"85113370",
          3789 => x"862a7081",
          3790 => x"06515151",
          3791 => x"5271802e",
          3792 => x"80c53882",
          3793 => x"e0a40888",
          3794 => x"050882e0",
          3795 => x"a4088805",
          3796 => x"08535385",
          3797 => x"123370ff",
          3798 => x"bf065152",
          3799 => x"71851434",
          3800 => x"82e0a408",
          3801 => x"8805088c",
          3802 => x"11088105",
          3803 => x"8c120c82",
          3804 => x"e0a40888",
          3805 => x"05088411",
          3806 => x"337082e0",
          3807 => x"a408f805",
          3808 => x"0c515152",
          3809 => x"82b63982",
          3810 => x"e0a40888",
          3811 => x"05088511",
          3812 => x"3370822a",
          3813 => x"70810651",
          3814 => x"51515271",
          3815 => x"802e80d7",
          3816 => x"3882e0a4",
          3817 => x"08880508",
          3818 => x"70087033",
          3819 => x"82e0a408",
          3820 => x"fc050c51",
          3821 => x"5282e0a4",
          3822 => x"08fc0508",
          3823 => x"a93882e0",
          3824 => x"a4088805",
          3825 => x"0882e0a4",
          3826 => x"08880508",
          3827 => x"53538512",
          3828 => x"3370a007",
          3829 => x"51527185",
          3830 => x"1434ff0b",
          3831 => x"82e0a408",
          3832 => x"f8050c81",
          3833 => x"d73982e0",
          3834 => x"a4088805",
          3835 => x"08700881",
          3836 => x"05710c52",
          3837 => x"81a13982",
          3838 => x"e0a40888",
          3839 => x"050882e0",
          3840 => x"a4088805",
          3841 => x"08529411",
          3842 => x"08515271",
          3843 => x"2d82e098",
          3844 => x"087082e0",
          3845 => x"a408fc05",
          3846 => x"0c5282e0",
          3847 => x"a408fc05",
          3848 => x"08802580",
          3849 => x"f23882e0",
          3850 => x"a4088805",
          3851 => x"0882e0a4",
          3852 => x"08f4050c",
          3853 => x"82e0a408",
          3854 => x"88050885",
          3855 => x"113382e0",
          3856 => x"a408f005",
          3857 => x"0c5282e0",
          3858 => x"a408fc05",
          3859 => x"08ff2e09",
          3860 => x"81069538",
          3861 => x"82e0a408",
          3862 => x"f0050890",
          3863 => x"07527182",
          3864 => x"e0a408ec",
          3865 => x"05349339",
          3866 => x"82e0a408",
          3867 => x"f00508a0",
          3868 => x"07527182",
          3869 => x"e0a408ec",
          3870 => x"053482e0",
          3871 => x"a408f405",
          3872 => x"085282e0",
          3873 => x"a408ec05",
          3874 => x"33851334",
          3875 => x"ff0b82e0",
          3876 => x"a408f805",
          3877 => x"0ca63982",
          3878 => x"e0a40888",
          3879 => x"05088c11",
          3880 => x"0881058c",
          3881 => x"120c82e0",
          3882 => x"a408fc05",
          3883 => x"087081ff",
          3884 => x"067082e0",
          3885 => x"a408f805",
          3886 => x"0c515152",
          3887 => x"82e0a408",
          3888 => x"f8050882",
          3889 => x"e0980c89",
          3890 => x"3d0d82e0",
          3891 => x"a40c0482",
          3892 => x"e0a40802",
          3893 => x"82e0a40c",
          3894 => x"fd3d0d82",
          3895 => x"e0a40888",
          3896 => x"050882e0",
          3897 => x"a408fc05",
          3898 => x"0c82e0a4",
          3899 => x"088c0508",
          3900 => x"82e0a408",
          3901 => x"f8050c82",
          3902 => x"e0a40890",
          3903 => x"0508802e",
          3904 => x"82a23882",
          3905 => x"e0a408f8",
          3906 => x"050882e0",
          3907 => x"a408fc05",
          3908 => x"082681ac",
          3909 => x"3882e0a4",
          3910 => x"08f80508",
          3911 => x"82e0a408",
          3912 => x"90050805",
          3913 => x"5182e0a4",
          3914 => x"08fc0508",
          3915 => x"71278190",
          3916 => x"3882e0a4",
          3917 => x"08fc0508",
          3918 => x"82e0a408",
          3919 => x"90050805",
          3920 => x"82e0a408",
          3921 => x"fc050c82",
          3922 => x"e0a408f8",
          3923 => x"050882e0",
          3924 => x"a4089005",
          3925 => x"080582e0",
          3926 => x"a408f805",
          3927 => x"0c82e0a4",
          3928 => x"08900508",
          3929 => x"810582e0",
          3930 => x"a4089005",
          3931 => x"0c82e0a4",
          3932 => x"08900508",
          3933 => x"ff0582e0",
          3934 => x"a4089005",
          3935 => x"0c82e0a4",
          3936 => x"08900508",
          3937 => x"802e819c",
          3938 => x"3882e0a4",
          3939 => x"08fc0508",
          3940 => x"ff0582e0",
          3941 => x"a408fc05",
          3942 => x"0c82e0a4",
          3943 => x"08f80508",
          3944 => x"ff0582e0",
          3945 => x"a408f805",
          3946 => x"0c82e0a4",
          3947 => x"08fc0508",
          3948 => x"82e0a408",
          3949 => x"f8050853",
          3950 => x"51713371",
          3951 => x"34ffae39",
          3952 => x"82e0a408",
          3953 => x"90050881",
          3954 => x"0582e0a4",
          3955 => x"0890050c",
          3956 => x"82e0a408",
          3957 => x"900508ff",
          3958 => x"0582e0a4",
          3959 => x"0890050c",
          3960 => x"82e0a408",
          3961 => x"90050880",
          3962 => x"2eba3882",
          3963 => x"e0a408f8",
          3964 => x"05085170",
          3965 => x"3382e0a4",
          3966 => x"08f80508",
          3967 => x"810582e0",
          3968 => x"a408f805",
          3969 => x"0c82e0a4",
          3970 => x"08fc0508",
          3971 => x"52527171",
          3972 => x"3482e0a4",
          3973 => x"08fc0508",
          3974 => x"810582e0",
          3975 => x"a408fc05",
          3976 => x"0cffad39",
          3977 => x"82e0a408",
          3978 => x"88050870",
          3979 => x"82e0980c",
          3980 => x"51853d0d",
          3981 => x"82e0a40c",
          3982 => x"0482e0a4",
          3983 => x"080282e0",
          3984 => x"a40cfe3d",
          3985 => x"0d82e0a4",
          3986 => x"08880508",
          3987 => x"82e0a408",
          3988 => x"fc050c82",
          3989 => x"e0a408fc",
          3990 => x"05085271",
          3991 => x"3382e0a4",
          3992 => x"08fc0508",
          3993 => x"810582e0",
          3994 => x"a408fc05",
          3995 => x"0c7081ff",
          3996 => x"06515170",
          3997 => x"802e8338",
          3998 => x"da3982e0",
          3999 => x"a408fc05",
          4000 => x"08ff0582",
          4001 => x"e0a408fc",
          4002 => x"050c82e0",
          4003 => x"a408fc05",
          4004 => x"0882e0a4",
          4005 => x"08880508",
          4006 => x"317082e0",
          4007 => x"980c5184",
          4008 => x"3d0d82e0",
          4009 => x"a40c0482",
          4010 => x"e0a40802",
          4011 => x"82e0a40c",
          4012 => x"fe3d0d82",
          4013 => x"e0a40888",
          4014 => x"050882e0",
          4015 => x"a408fc05",
          4016 => x"0c82e0a4",
          4017 => x"088c0508",
          4018 => x"52713382",
          4019 => x"e0a4088c",
          4020 => x"05088105",
          4021 => x"82e0a408",
          4022 => x"8c050c82",
          4023 => x"e0a408fc",
          4024 => x"05085351",
          4025 => x"70723482",
          4026 => x"e0a408fc",
          4027 => x"05088105",
          4028 => x"82e0a408",
          4029 => x"fc050c70",
          4030 => x"81ff0651",
          4031 => x"70802e84",
          4032 => x"38ffbe39",
          4033 => x"82e0a408",
          4034 => x"88050870",
          4035 => x"82e0980c",
          4036 => x"51843d0d",
          4037 => x"82e0a40c",
          4038 => x"0482e0a4",
          4039 => x"080282e0",
          4040 => x"a40cfd3d",
          4041 => x"0d82e0a4",
          4042 => x"08880508",
          4043 => x"82e0a408",
          4044 => x"fc050c82",
          4045 => x"e0a4088c",
          4046 => x"050882e0",
          4047 => x"a408f805",
          4048 => x"0c82e0a4",
          4049 => x"08900508",
          4050 => x"802e80e5",
          4051 => x"3882e0a4",
          4052 => x"08900508",
          4053 => x"810582e0",
          4054 => x"a4089005",
          4055 => x"0c82e0a4",
          4056 => x"08900508",
          4057 => x"ff0582e0",
          4058 => x"a4089005",
          4059 => x"0c82e0a4",
          4060 => x"08900508",
          4061 => x"802eba38",
          4062 => x"82e0a408",
          4063 => x"f8050851",
          4064 => x"703382e0",
          4065 => x"a408f805",
          4066 => x"08810582",
          4067 => x"e0a408f8",
          4068 => x"050c82e0",
          4069 => x"a408fc05",
          4070 => x"08525271",
          4071 => x"713482e0",
          4072 => x"a408fc05",
          4073 => x"08810582",
          4074 => x"e0a408fc",
          4075 => x"050cffad",
          4076 => x"3982e0a4",
          4077 => x"08880508",
          4078 => x"7082e098",
          4079 => x"0c51853d",
          4080 => x"0d82e0a4",
          4081 => x"0c0482e0",
          4082 => x"a4080282",
          4083 => x"e0a40cfd",
          4084 => x"3d0d82e0",
          4085 => x"a4089005",
          4086 => x"08802e81",
          4087 => x"f43882e0",
          4088 => x"a4088c05",
          4089 => x"08527133",
          4090 => x"82e0a408",
          4091 => x"8c050881",
          4092 => x"0582e0a4",
          4093 => x"088c050c",
          4094 => x"82e0a408",
          4095 => x"88050870",
          4096 => x"337281ff",
          4097 => x"06535454",
          4098 => x"5171712e",
          4099 => x"843880ce",
          4100 => x"3982e0a4",
          4101 => x"08880508",
          4102 => x"52713382",
          4103 => x"e0a40888",
          4104 => x"05088105",
          4105 => x"82e0a408",
          4106 => x"88050c70",
          4107 => x"81ff0651",
          4108 => x"51708d38",
          4109 => x"800b82e0",
          4110 => x"a408fc05",
          4111 => x"0c819b39",
          4112 => x"82e0a408",
          4113 => x"900508ff",
          4114 => x"0582e0a4",
          4115 => x"0890050c",
          4116 => x"82e0a408",
          4117 => x"90050880",
          4118 => x"2e8438ff",
          4119 => x"813982e0",
          4120 => x"a4089005",
          4121 => x"08802e80",
          4122 => x"e83882e0",
          4123 => x"a4088805",
          4124 => x"08703352",
          4125 => x"53708d38",
          4126 => x"ff0b82e0",
          4127 => x"a408fc05",
          4128 => x"0c80d739",
          4129 => x"82e0a408",
          4130 => x"8c0508ff",
          4131 => x"0582e0a4",
          4132 => x"088c050c",
          4133 => x"82e0a408",
          4134 => x"8c050870",
          4135 => x"33525270",
          4136 => x"8c38810b",
          4137 => x"82e0a408",
          4138 => x"fc050cae",
          4139 => x"3982e0a4",
          4140 => x"08880508",
          4141 => x"703382e0",
          4142 => x"a4088c05",
          4143 => x"08703372",
          4144 => x"71317082",
          4145 => x"e0a408fc",
          4146 => x"050c5355",
          4147 => x"5252538a",
          4148 => x"39800b82",
          4149 => x"e0a408fc",
          4150 => x"050c82e0",
          4151 => x"a408fc05",
          4152 => x"0882e098",
          4153 => x"0c853d0d",
          4154 => x"82e0a40c",
          4155 => x"0482e0a4",
          4156 => x"080282e0",
          4157 => x"a40cfa3d",
          4158 => x"0d82e0a4",
          4159 => x"088c0508",
          4160 => x"5282e0a4",
          4161 => x"08880508",
          4162 => x"51818d3f",
          4163 => x"82e09808",
          4164 => x"7082e0a4",
          4165 => x"08f8050c",
          4166 => x"82e0a408",
          4167 => x"f8050881",
          4168 => x"05705351",
          4169 => x"5480ecf7",
          4170 => x"3f82e098",
          4171 => x"087082e0",
          4172 => x"a408fc05",
          4173 => x"0c5482e0",
          4174 => x"a408fc05",
          4175 => x"088c3880",
          4176 => x"0b82e0a4",
          4177 => x"08f4050c",
          4178 => x"bc3982e0",
          4179 => x"a408fc05",
          4180 => x"0882e0a4",
          4181 => x"08f80508",
          4182 => x"05548074",
          4183 => x"3482e0a4",
          4184 => x"08f80508",
          4185 => x"5382e0a4",
          4186 => x"08880508",
          4187 => x"5282e0a4",
          4188 => x"08fc0508",
          4189 => x"51fba23f",
          4190 => x"82e09808",
          4191 => x"7082e0a4",
          4192 => x"08f4050c",
          4193 => x"5482e0a4",
          4194 => x"08f40508",
          4195 => x"82e0980c",
          4196 => x"883d0d82",
          4197 => x"e0a40c04",
          4198 => x"82e0a408",
          4199 => x"0282e0a4",
          4200 => x"0cfd3d0d",
          4201 => x"82e0a408",
          4202 => x"88050882",
          4203 => x"e0a408f8",
          4204 => x"050c82e0",
          4205 => x"a4088c05",
          4206 => x"088d3880",
          4207 => x"0b82e0a4",
          4208 => x"08fc050c",
          4209 => x"80ec3982",
          4210 => x"e0a408f8",
          4211 => x"05085271",
          4212 => x"3382e0a4",
          4213 => x"08f80508",
          4214 => x"810582e0",
          4215 => x"a408f805",
          4216 => x"0c7081ff",
          4217 => x"06515170",
          4218 => x"802e9f38",
          4219 => x"82e0a408",
          4220 => x"8c0508ff",
          4221 => x"0582e0a4",
          4222 => x"088c050c",
          4223 => x"82e0a408",
          4224 => x"8c0508ff",
          4225 => x"2e8438ff",
          4226 => x"be3982e0",
          4227 => x"a408f805",
          4228 => x"08ff0582",
          4229 => x"e0a408f8",
          4230 => x"050c82e0",
          4231 => x"a408f805",
          4232 => x"0882e0a4",
          4233 => x"08880508",
          4234 => x"317082e0",
          4235 => x"a408fc05",
          4236 => x"0c5182e0",
          4237 => x"a408fc05",
          4238 => x"0882e098",
          4239 => x"0c853d0d",
          4240 => x"82e0a40c",
          4241 => x"0482e0a4",
          4242 => x"080282e0",
          4243 => x"a40cfe3d",
          4244 => x"0d82e0a4",
          4245 => x"08880508",
          4246 => x"82e0a408",
          4247 => x"fc050c82",
          4248 => x"e0a40890",
          4249 => x"0508802e",
          4250 => x"80d43882",
          4251 => x"e0a40890",
          4252 => x"05088105",
          4253 => x"82e0a408",
          4254 => x"90050c82",
          4255 => x"e0a40890",
          4256 => x"0508ff05",
          4257 => x"82e0a408",
          4258 => x"90050c82",
          4259 => x"e0a40890",
          4260 => x"0508802e",
          4261 => x"a93882e0",
          4262 => x"a4088c05",
          4263 => x"08517082",
          4264 => x"e0a408fc",
          4265 => x"05085252",
          4266 => x"71713482",
          4267 => x"e0a408fc",
          4268 => x"05088105",
          4269 => x"82e0a408",
          4270 => x"fc050cff",
          4271 => x"be3982e0",
          4272 => x"a4088805",
          4273 => x"087082e0",
          4274 => x"980c5184",
          4275 => x"3d0d82e0",
          4276 => x"a40c0482",
          4277 => x"e0a40802",
          4278 => x"82e0a40c",
          4279 => x"fe3d0d82",
          4280 => x"e0a4088c",
          4281 => x"05085282",
          4282 => x"e0a40888",
          4283 => x"05085193",
          4284 => x"3f82e098",
          4285 => x"087082e0",
          4286 => x"980c5384",
          4287 => x"3d0d82e0",
          4288 => x"a40c0482",
          4289 => x"e0a40802",
          4290 => x"82e0a40c",
          4291 => x"f63d0da0",
          4292 => x"0b82e0a4",
          4293 => x"08fc050c",
          4294 => x"82e0a408",
          4295 => x"8c050880",
          4296 => x"2e9b3882",
          4297 => x"e0a4088c",
          4298 => x"05085183",
          4299 => x"fc3f82e0",
          4300 => x"98087082",
          4301 => x"e0a408e4",
          4302 => x"050c528f",
          4303 => x"3982e0a4",
          4304 => x"08fc0508",
          4305 => x"82e0a408",
          4306 => x"e4050c82",
          4307 => x"e0a40888",
          4308 => x"0508802e",
          4309 => x"a33882e0",
          4310 => x"a4088805",
          4311 => x"085183c9",
          4312 => x"3f82e098",
          4313 => x"0882e0a4",
          4314 => x"08e40508",
          4315 => x"713182e0",
          4316 => x"a408e005",
          4317 => x"0c529739",
          4318 => x"82e0a408",
          4319 => x"e4050882",
          4320 => x"e0a408fc",
          4321 => x"05083182",
          4322 => x"e0a408e0",
          4323 => x"050c82e0",
          4324 => x"a408e005",
          4325 => x"0882e0a4",
          4326 => x"08f8050c",
          4327 => x"82e0a408",
          4328 => x"fc0508ff",
          4329 => x"05527182",
          4330 => x"e0a408f8",
          4331 => x"0508278d",
          4332 => x"38800b82",
          4333 => x"e0a408e8",
          4334 => x"050c82da",
          4335 => x"3982e0a4",
          4336 => x"08fc0508",
          4337 => x"ff055271",
          4338 => x"82e0a408",
          4339 => x"f805082e",
          4340 => x"09810694",
          4341 => x"3882e0a4",
          4342 => x"08880508",
          4343 => x"7082e0a4",
          4344 => x"08e8050c",
          4345 => x"5282af39",
          4346 => x"82e0a408",
          4347 => x"f8050881",
          4348 => x"0582e0a4",
          4349 => x"08f8050c",
          4350 => x"82e0a408",
          4351 => x"88050882",
          4352 => x"e0a408f8",
          4353 => x"05082a82",
          4354 => x"e0a408f4",
          4355 => x"050c82e0",
          4356 => x"a408fc05",
          4357 => x"0882e0a4",
          4358 => x"08f80508",
          4359 => x"3182e0a4",
          4360 => x"08880508",
          4361 => x"712b82e0",
          4362 => x"a4088805",
          4363 => x"0c52800b",
          4364 => x"82e0a408",
          4365 => x"f0050c82",
          4366 => x"e0a408f8",
          4367 => x"0508802e",
          4368 => x"81ab3882",
          4369 => x"e0a408f4",
          4370 => x"05081082",
          4371 => x"e0a408fc",
          4372 => x"0508ff05",
          4373 => x"82e0a408",
          4374 => x"88050871",
          4375 => x"2a707307",
          4376 => x"82e0a408",
          4377 => x"f4050c82",
          4378 => x"e0a40888",
          4379 => x"05081070",
          4380 => x"82e0a408",
          4381 => x"f0050807",
          4382 => x"82e0a408",
          4383 => x"88050c82",
          4384 => x"e0a4088c",
          4385 => x"050882e0",
          4386 => x"a408f405",
          4387 => x"0831ff11",
          4388 => x"82e0a408",
          4389 => x"fc0508ff",
          4390 => x"0571712c",
          4391 => x"82e0a408",
          4392 => x"ec050c82",
          4393 => x"e0a408ec",
          4394 => x"05088106",
          4395 => x"82e0a408",
          4396 => x"f0050c82",
          4397 => x"e0a4088c",
          4398 => x"050882e0",
          4399 => x"a408ec05",
          4400 => x"080682e0",
          4401 => x"a408f405",
          4402 => x"08713182",
          4403 => x"e0a408f4",
          4404 => x"050c82e0",
          4405 => x"a408f805",
          4406 => x"08ff0582",
          4407 => x"e0a408f8",
          4408 => x"050c5152",
          4409 => x"55515151",
          4410 => x"5353fecb",
          4411 => x"3982e0a4",
          4412 => x"08880508",
          4413 => x"107082e0",
          4414 => x"a408f005",
          4415 => x"080782e0",
          4416 => x"a4088805",
          4417 => x"0c82e0a4",
          4418 => x"08880508",
          4419 => x"7082e0a4",
          4420 => x"08e8050c",
          4421 => x"515282e0",
          4422 => x"a408e805",
          4423 => x"0882e098",
          4424 => x"0c8c3d0d",
          4425 => x"82e0a40c",
          4426 => x"0482e0a4",
          4427 => x"080282e0",
          4428 => x"a40cf83d",
          4429 => x"0d82e0a4",
          4430 => x"08880508",
          4431 => x"82e0a408",
          4432 => x"fc050c82",
          4433 => x"e0a408fc",
          4434 => x"0508fc80",
          4435 => x"80065170",
          4436 => x"8c38900b",
          4437 => x"82e0a408",
          4438 => x"f0050c8a",
          4439 => x"39800b82",
          4440 => x"e0a408f0",
          4441 => x"050c82e0",
          4442 => x"a408f005",
          4443 => x"0882e0a4",
          4444 => x"08f8050c",
          4445 => x"900b82e0",
          4446 => x"a408f805",
          4447 => x"083182e0",
          4448 => x"a408fc05",
          4449 => x"08712a82",
          4450 => x"e0a408fc",
          4451 => x"050c82e0",
          4452 => x"a408f805",
          4453 => x"0882e0a4",
          4454 => x"08f4050c",
          4455 => x"82e0a408",
          4456 => x"fc050883",
          4457 => x"fe800651",
          4458 => x"51708c38",
          4459 => x"880b82e0",
          4460 => x"a408ec05",
          4461 => x"0c8a3980",
          4462 => x"0b82e0a4",
          4463 => x"08ec050c",
          4464 => x"82e0a408",
          4465 => x"ec050882",
          4466 => x"e0a408f8",
          4467 => x"050c880b",
          4468 => x"82e0a408",
          4469 => x"f8050831",
          4470 => x"82e0a408",
          4471 => x"fc050871",
          4472 => x"2a82e0a4",
          4473 => x"08fc050c",
          4474 => x"82e0a408",
          4475 => x"f4050882",
          4476 => x"e0a408f8",
          4477 => x"05080582",
          4478 => x"e0a408f4",
          4479 => x"050c82e0",
          4480 => x"a408fc05",
          4481 => x"0881f006",
          4482 => x"5151708c",
          4483 => x"38840b82",
          4484 => x"e0a408e8",
          4485 => x"050c8a39",
          4486 => x"800b82e0",
          4487 => x"a408e805",
          4488 => x"0c82e0a4",
          4489 => x"08e80508",
          4490 => x"82e0a408",
          4491 => x"f8050c84",
          4492 => x"0b82e0a4",
          4493 => x"08f80508",
          4494 => x"3182e0a4",
          4495 => x"08fc0508",
          4496 => x"712a82e0",
          4497 => x"a408fc05",
          4498 => x"0c82e0a4",
          4499 => x"08f40508",
          4500 => x"82e0a408",
          4501 => x"f8050805",
          4502 => x"82e0a408",
          4503 => x"f4050c82",
          4504 => x"e0a408fc",
          4505 => x"05088c06",
          4506 => x"5151708c",
          4507 => x"38820b82",
          4508 => x"e0a408e4",
          4509 => x"050c8a39",
          4510 => x"800b82e0",
          4511 => x"a408e405",
          4512 => x"0c82e0a4",
          4513 => x"08e40508",
          4514 => x"82e0a408",
          4515 => x"f8050c82",
          4516 => x"0b82e0a4",
          4517 => x"08f80508",
          4518 => x"3182e0a4",
          4519 => x"08fc0508",
          4520 => x"712a82e0",
          4521 => x"a408fc05",
          4522 => x"0c82e0a4",
          4523 => x"08f40508",
          4524 => x"82e0a408",
          4525 => x"f8050805",
          4526 => x"82e0a408",
          4527 => x"f4050c82",
          4528 => x"0b82e0a4",
          4529 => x"08fc0508",
          4530 => x"3182e0a4",
          4531 => x"08fc0508",
          4532 => x"812a7081",
          4533 => x"32708106",
          4534 => x"70307075",
          4535 => x"0682e0a4",
          4536 => x"08f40508",
          4537 => x"11707082",
          4538 => x"e0980c53",
          4539 => x"51555151",
          4540 => x"51525351",
          4541 => x"8a3d0d82",
          4542 => x"e0a40c04",
          4543 => x"82e0a408",
          4544 => x"0282e0a4",
          4545 => x"0cfe3d0d",
          4546 => x"82e0a408",
          4547 => x"8c050852",
          4548 => x"82e0a408",
          4549 => x"88050851",
          4550 => x"84e43f82",
          4551 => x"e0980870",
          4552 => x"82e0a408",
          4553 => x"8c050829",
          4554 => x"82e0a408",
          4555 => x"88050871",
          4556 => x"317082e0",
          4557 => x"980c5151",
          4558 => x"53843d0d",
          4559 => x"82e0a40c",
          4560 => x"0482e0a4",
          4561 => x"080282e0",
          4562 => x"a40cfe3d",
          4563 => x"0d82e0a4",
          4564 => x"088c0508",
          4565 => x"5282e0a4",
          4566 => x"08880508",
          4567 => x"51933f82",
          4568 => x"e0980870",
          4569 => x"82e0980c",
          4570 => x"53843d0d",
          4571 => x"82e0a40c",
          4572 => x"0482e0a4",
          4573 => x"080282e0",
          4574 => x"a40cf63d",
          4575 => x"0da00b82",
          4576 => x"e0a408fc",
          4577 => x"050c82e0",
          4578 => x"a4088c05",
          4579 => x"08802e9b",
          4580 => x"3882e0a4",
          4581 => x"088c0508",
          4582 => x"51fb8e3f",
          4583 => x"82e09808",
          4584 => x"7082e0a4",
          4585 => x"08e4050c",
          4586 => x"528f3982",
          4587 => x"e0a408fc",
          4588 => x"050882e0",
          4589 => x"a408e405",
          4590 => x"0c82e0a4",
          4591 => x"08880508",
          4592 => x"802ea338",
          4593 => x"82e0a408",
          4594 => x"88050851",
          4595 => x"fadb3f82",
          4596 => x"e0980882",
          4597 => x"e0a408e4",
          4598 => x"05087131",
          4599 => x"82e0a408",
          4600 => x"e0050c52",
          4601 => x"973982e0",
          4602 => x"a408e405",
          4603 => x"0882e0a4",
          4604 => x"08fc0508",
          4605 => x"3182e0a4",
          4606 => x"08e0050c",
          4607 => x"82e0a408",
          4608 => x"e0050882",
          4609 => x"e0a408f8",
          4610 => x"050c82e0",
          4611 => x"a408fc05",
          4612 => x"08ff0552",
          4613 => x"7182e0a4",
          4614 => x"08f80508",
          4615 => x"27943882",
          4616 => x"e0a40888",
          4617 => x"05087082",
          4618 => x"e0a408e8",
          4619 => x"050c5282",
          4620 => x"ba3982e0",
          4621 => x"a408fc05",
          4622 => x"08ff0552",
          4623 => x"7182e0a4",
          4624 => x"08f80508",
          4625 => x"2e098106",
          4626 => x"8d38800b",
          4627 => x"82e0a408",
          4628 => x"e8050c82",
          4629 => x"963982e0",
          4630 => x"a408f805",
          4631 => x"08810582",
          4632 => x"e0a408f8",
          4633 => x"050c82e0",
          4634 => x"a4088805",
          4635 => x"0882e0a4",
          4636 => x"08f80508",
          4637 => x"2a82e0a4",
          4638 => x"08f4050c",
          4639 => x"82e0a408",
          4640 => x"fc050882",
          4641 => x"e0a408f8",
          4642 => x"05083182",
          4643 => x"e0a40888",
          4644 => x"0508712b",
          4645 => x"82e0a408",
          4646 => x"88050c52",
          4647 => x"800b82e0",
          4648 => x"a408f005",
          4649 => x"0c82e0a4",
          4650 => x"08f80508",
          4651 => x"802e81ab",
          4652 => x"3882e0a4",
          4653 => x"08f40508",
          4654 => x"1082e0a4",
          4655 => x"08fc0508",
          4656 => x"ff0582e0",
          4657 => x"a4088805",
          4658 => x"08712a70",
          4659 => x"730782e0",
          4660 => x"a408f405",
          4661 => x"0c82e0a4",
          4662 => x"08880508",
          4663 => x"107082e0",
          4664 => x"a408f005",
          4665 => x"080782e0",
          4666 => x"a4088805",
          4667 => x"0c82e0a4",
          4668 => x"088c0508",
          4669 => x"82e0a408",
          4670 => x"f4050831",
          4671 => x"ff1182e0",
          4672 => x"a408fc05",
          4673 => x"08ff0571",
          4674 => x"712c82e0",
          4675 => x"a408ec05",
          4676 => x"0c82e0a4",
          4677 => x"08ec0508",
          4678 => x"810682e0",
          4679 => x"a408f005",
          4680 => x"0c82e0a4",
          4681 => x"088c0508",
          4682 => x"82e0a408",
          4683 => x"ec050806",
          4684 => x"82e0a408",
          4685 => x"f4050871",
          4686 => x"3182e0a4",
          4687 => x"08f4050c",
          4688 => x"82e0a408",
          4689 => x"f80508ff",
          4690 => x"0582e0a4",
          4691 => x"08f8050c",
          4692 => x"51525551",
          4693 => x"51515353",
          4694 => x"fecb3982",
          4695 => x"e0a408f4",
          4696 => x"05087082",
          4697 => x"e0a408e8",
          4698 => x"050c5282",
          4699 => x"e0a408e8",
          4700 => x"050882e0",
          4701 => x"980c8c3d",
          4702 => x"0d82e0a4",
          4703 => x"0c0482e0",
          4704 => x"a4080282",
          4705 => x"e0a40cfb",
          4706 => x"3d0d9f0b",
          4707 => x"82e0a408",
          4708 => x"fc050c82",
          4709 => x"e0a40888",
          4710 => x"050882e0",
          4711 => x"a408fc05",
          4712 => x"082c82e0",
          4713 => x"a408f805",
          4714 => x"0c82e0a4",
          4715 => x"088c0508",
          4716 => x"82e0a408",
          4717 => x"fc05082c",
          4718 => x"82e0a408",
          4719 => x"f4050c82",
          4720 => x"e0a40888",
          4721 => x"050882e0",
          4722 => x"a408f805",
          4723 => x"08327082",
          4724 => x"e0a408f8",
          4725 => x"05083182",
          4726 => x"e0a40888",
          4727 => x"050c82e0",
          4728 => x"a4088c05",
          4729 => x"0882e0a4",
          4730 => x"08f40508",
          4731 => x"327082e0",
          4732 => x"a408f405",
          4733 => x"083182e0",
          4734 => x"a4088c05",
          4735 => x"0c82e0a4",
          4736 => x"08f80508",
          4737 => x"82e0a408",
          4738 => x"f4050832",
          4739 => x"82e0a408",
          4740 => x"f8050c82",
          4741 => x"e0a4088c",
          4742 => x"05085482",
          4743 => x"e0a40888",
          4744 => x"05085351",
          4745 => x"53f1ac3f",
          4746 => x"82e09808",
          4747 => x"7082e0a4",
          4748 => x"08f80508",
          4749 => x"327082e0",
          4750 => x"a408f805",
          4751 => x"08317082",
          4752 => x"e0980c51",
          4753 => x"5153873d",
          4754 => x"0d82e0a4",
          4755 => x"0c0482e0",
          4756 => x"a4080282",
          4757 => x"e0a40cf7",
          4758 => x"3d0d800b",
          4759 => x"82e0a408",
          4760 => x"f0053482",
          4761 => x"e0a4088c",
          4762 => x"05085380",
          4763 => x"730c82e0",
          4764 => x"a4088805",
          4765 => x"08700851",
          4766 => x"53723353",
          4767 => x"7282e0a4",
          4768 => x"08f80534",
          4769 => x"7281ff06",
          4770 => x"5372a02e",
          4771 => x"09810691",
          4772 => x"3882e0a4",
          4773 => x"08880508",
          4774 => x"70088105",
          4775 => x"710c53ce",
          4776 => x"3982e0a4",
          4777 => x"08f80533",
          4778 => x"5372ad2e",
          4779 => x"098106a4",
          4780 => x"38810b82",
          4781 => x"e0a408f0",
          4782 => x"053482e0",
          4783 => x"a4088805",
          4784 => x"08700881",
          4785 => x"05710c70",
          4786 => x"08515372",
          4787 => x"3382e0a4",
          4788 => x"08f80534",
          4789 => x"82e0a408",
          4790 => x"f8053353",
          4791 => x"72b02e09",
          4792 => x"810681dc",
          4793 => x"3882e0a4",
          4794 => x"08880508",
          4795 => x"70088105",
          4796 => x"710c7008",
          4797 => x"51537233",
          4798 => x"82e0a408",
          4799 => x"f8053482",
          4800 => x"e0a408f8",
          4801 => x"053382e0",
          4802 => x"a408e805",
          4803 => x"0c82e0a4",
          4804 => x"08e80508",
          4805 => x"80e22eb6",
          4806 => x"3882e0a4",
          4807 => x"08e80508",
          4808 => x"80f82e84",
          4809 => x"3880cd39",
          4810 => x"900b82e0",
          4811 => x"a408f405",
          4812 => x"3482e0a4",
          4813 => x"08880508",
          4814 => x"70088105",
          4815 => x"710c7008",
          4816 => x"51537233",
          4817 => x"82e0a408",
          4818 => x"f8053481",
          4819 => x"a439820b",
          4820 => x"82e0a408",
          4821 => x"f4053482",
          4822 => x"e0a40888",
          4823 => x"05087008",
          4824 => x"8105710c",
          4825 => x"70085153",
          4826 => x"723382e0",
          4827 => x"a408f805",
          4828 => x"3480fe39",
          4829 => x"82e0a408",
          4830 => x"f8053353",
          4831 => x"72a0268d",
          4832 => x"38810b82",
          4833 => x"e0a408ec",
          4834 => x"050c8380",
          4835 => x"3982e0a4",
          4836 => x"08f80533",
          4837 => x"53af7327",
          4838 => x"903882e0",
          4839 => x"a408f805",
          4840 => x"335372b9",
          4841 => x"2683388d",
          4842 => x"39800b82",
          4843 => x"e0a408ec",
          4844 => x"050c82d8",
          4845 => x"39880b82",
          4846 => x"e0a408f4",
          4847 => x"0534b239",
          4848 => x"82e0a408",
          4849 => x"f8053353",
          4850 => x"af732790",
          4851 => x"3882e0a4",
          4852 => x"08f80533",
          4853 => x"5372b926",
          4854 => x"83388d39",
          4855 => x"800b82e0",
          4856 => x"a408ec05",
          4857 => x"0c82a539",
          4858 => x"8a0b82e0",
          4859 => x"a408f405",
          4860 => x"34800b82",
          4861 => x"e0a408fc",
          4862 => x"050c82e0",
          4863 => x"a408f805",
          4864 => x"3353a073",
          4865 => x"2781cf38",
          4866 => x"82e0a408",
          4867 => x"f8053353",
          4868 => x"80e07327",
          4869 => x"943882e0",
          4870 => x"a408f805",
          4871 => x"33e01151",
          4872 => x"537282e0",
          4873 => x"a408f805",
          4874 => x"3482e0a4",
          4875 => x"08f80533",
          4876 => x"d0115153",
          4877 => x"7282e0a4",
          4878 => x"08f80534",
          4879 => x"82e0a408",
          4880 => x"f8053353",
          4881 => x"907327ad",
          4882 => x"3882e0a4",
          4883 => x"08f80533",
          4884 => x"f9115153",
          4885 => x"7282e0a4",
          4886 => x"08f80534",
          4887 => x"82e0a408",
          4888 => x"f8053353",
          4889 => x"7289268d",
          4890 => x"38800b82",
          4891 => x"e0a408ec",
          4892 => x"050c8198",
          4893 => x"3982e0a4",
          4894 => x"08f80533",
          4895 => x"82e0a408",
          4896 => x"f4053354",
          4897 => x"54727426",
          4898 => x"8d38800b",
          4899 => x"82e0a408",
          4900 => x"ec050c80",
          4901 => x"f73982e0",
          4902 => x"a408f405",
          4903 => x"337082e0",
          4904 => x"a408fc05",
          4905 => x"082982e0",
          4906 => x"a408f805",
          4907 => x"33701282",
          4908 => x"e0a408fc",
          4909 => x"050c82e0",
          4910 => x"a4088805",
          4911 => x"08700881",
          4912 => x"05710c70",
          4913 => x"08515152",
          4914 => x"55537233",
          4915 => x"82e0a408",
          4916 => x"f80534fe",
          4917 => x"a53982e0",
          4918 => x"a408f005",
          4919 => x"33537280",
          4920 => x"2e903882",
          4921 => x"e0a408fc",
          4922 => x"05083082",
          4923 => x"e0a408fc",
          4924 => x"050c82e0",
          4925 => x"a4088c05",
          4926 => x"0882e0a4",
          4927 => x"08fc0508",
          4928 => x"710c5381",
          4929 => x"0b82e0a4",
          4930 => x"08ec050c",
          4931 => x"82e0a408",
          4932 => x"ec050882",
          4933 => x"e0980c8b",
          4934 => x"3d0d82e0",
          4935 => x"a40c0482",
          4936 => x"e0a40802",
          4937 => x"82e0a40c",
          4938 => x"f73d0d80",
          4939 => x"0b82e0a4",
          4940 => x"08f00534",
          4941 => x"82e0a408",
          4942 => x"8c050853",
          4943 => x"80730c82",
          4944 => x"e0a40888",
          4945 => x"05087008",
          4946 => x"51537233",
          4947 => x"537282e0",
          4948 => x"a408f805",
          4949 => x"347281ff",
          4950 => x"065372a0",
          4951 => x"2e098106",
          4952 => x"913882e0",
          4953 => x"a4088805",
          4954 => x"08700881",
          4955 => x"05710c53",
          4956 => x"ce3982e0",
          4957 => x"a408f805",
          4958 => x"335372ad",
          4959 => x"2e098106",
          4960 => x"a438810b",
          4961 => x"82e0a408",
          4962 => x"f0053482",
          4963 => x"e0a40888",
          4964 => x"05087008",
          4965 => x"8105710c",
          4966 => x"70085153",
          4967 => x"723382e0",
          4968 => x"a408f805",
          4969 => x"3482e0a4",
          4970 => x"08f80533",
          4971 => x"5372b02e",
          4972 => x"09810681",
          4973 => x"dc3882e0",
          4974 => x"a4088805",
          4975 => x"08700881",
          4976 => x"05710c70",
          4977 => x"08515372",
          4978 => x"3382e0a4",
          4979 => x"08f80534",
          4980 => x"82e0a408",
          4981 => x"f8053382",
          4982 => x"e0a408e8",
          4983 => x"050c82e0",
          4984 => x"a408e805",
          4985 => x"0880e22e",
          4986 => x"b63882e0",
          4987 => x"a408e805",
          4988 => x"0880f82e",
          4989 => x"843880cd",
          4990 => x"39900b82",
          4991 => x"e0a408f4",
          4992 => x"053482e0",
          4993 => x"a4088805",
          4994 => x"08700881",
          4995 => x"05710c70",
          4996 => x"08515372",
          4997 => x"3382e0a4",
          4998 => x"08f80534",
          4999 => x"81a43982",
          5000 => x"0b82e0a4",
          5001 => x"08f40534",
          5002 => x"82e0a408",
          5003 => x"88050870",
          5004 => x"08810571",
          5005 => x"0c700851",
          5006 => x"53723382",
          5007 => x"e0a408f8",
          5008 => x"053480fe",
          5009 => x"3982e0a4",
          5010 => x"08f80533",
          5011 => x"5372a026",
          5012 => x"8d38810b",
          5013 => x"82e0a408",
          5014 => x"ec050c83",
          5015 => x"803982e0",
          5016 => x"a408f805",
          5017 => x"3353af73",
          5018 => x"27903882",
          5019 => x"e0a408f8",
          5020 => x"05335372",
          5021 => x"b9268338",
          5022 => x"8d39800b",
          5023 => x"82e0a408",
          5024 => x"ec050c82",
          5025 => x"d839880b",
          5026 => x"82e0a408",
          5027 => x"f40534b2",
          5028 => x"3982e0a4",
          5029 => x"08f80533",
          5030 => x"53af7327",
          5031 => x"903882e0",
          5032 => x"a408f805",
          5033 => x"335372b9",
          5034 => x"2683388d",
          5035 => x"39800b82",
          5036 => x"e0a408ec",
          5037 => x"050c82a5",
          5038 => x"398a0b82",
          5039 => x"e0a408f4",
          5040 => x"0534800b",
          5041 => x"82e0a408",
          5042 => x"fc050c82",
          5043 => x"e0a408f8",
          5044 => x"053353a0",
          5045 => x"732781cf",
          5046 => x"3882e0a4",
          5047 => x"08f80533",
          5048 => x"5380e073",
          5049 => x"27943882",
          5050 => x"e0a408f8",
          5051 => x"0533e011",
          5052 => x"51537282",
          5053 => x"e0a408f8",
          5054 => x"053482e0",
          5055 => x"a408f805",
          5056 => x"33d01151",
          5057 => x"537282e0",
          5058 => x"a408f805",
          5059 => x"3482e0a4",
          5060 => x"08f80533",
          5061 => x"53907327",
          5062 => x"ad3882e0",
          5063 => x"a408f805",
          5064 => x"33f91151",
          5065 => x"537282e0",
          5066 => x"a408f805",
          5067 => x"3482e0a4",
          5068 => x"08f80533",
          5069 => x"53728926",
          5070 => x"8d38800b",
          5071 => x"82e0a408",
          5072 => x"ec050c81",
          5073 => x"983982e0",
          5074 => x"a408f805",
          5075 => x"3382e0a4",
          5076 => x"08f40533",
          5077 => x"54547274",
          5078 => x"268d3880",
          5079 => x"0b82e0a4",
          5080 => x"08ec050c",
          5081 => x"80f73982",
          5082 => x"e0a408f4",
          5083 => x"05337082",
          5084 => x"e0a408fc",
          5085 => x"05082982",
          5086 => x"e0a408f8",
          5087 => x"05337012",
          5088 => x"82e0a408",
          5089 => x"fc050c82",
          5090 => x"e0a40888",
          5091 => x"05087008",
          5092 => x"8105710c",
          5093 => x"70085151",
          5094 => x"52555372",
          5095 => x"3382e0a4",
          5096 => x"08f80534",
          5097 => x"fea53982",
          5098 => x"e0a408f0",
          5099 => x"05335372",
          5100 => x"802e9038",
          5101 => x"82e0a408",
          5102 => x"fc050830",
          5103 => x"82e0a408",
          5104 => x"fc050c82",
          5105 => x"e0a4088c",
          5106 => x"050882e0",
          5107 => x"a408fc05",
          5108 => x"08710c53",
          5109 => x"810b82e0",
          5110 => x"a408ec05",
          5111 => x"0c82e0a4",
          5112 => x"08ec0508",
          5113 => x"82e0980c",
          5114 => x"8b3d0d82",
          5115 => x"e0a40c04",
          5116 => x"f83d0d7a",
          5117 => x"70087056",
          5118 => x"56597480",
          5119 => x"2e80df38",
          5120 => x"8c397715",
          5121 => x"790c8516",
          5122 => x"335480d2",
          5123 => x"39743354",
          5124 => x"73a02e09",
          5125 => x"81068638",
          5126 => x"811555f1",
          5127 => x"39805776",
          5128 => x"902982db",
          5129 => x"a0057008",
          5130 => x"5256dc8d",
          5131 => x"3f82e098",
          5132 => x"0882e098",
          5133 => x"08547553",
          5134 => x"76085258",
          5135 => x"df883f82",
          5136 => x"e098088b",
          5137 => x"38841633",
          5138 => x"5473812e",
          5139 => x"ffb43881",
          5140 => x"177081ff",
          5141 => x"06585498",
          5142 => x"7727c438",
          5143 => x"ff547382",
          5144 => x"e0980c8a",
          5145 => x"3d0d0481",
          5146 => x"a00b82e0",
          5147 => x"980c04ff",
          5148 => x"3d0d7352",
          5149 => x"71932681",
          5150 => x"8e387184",
          5151 => x"2982b7fc",
          5152 => x"05527108",
          5153 => x"0482bde4",
          5154 => x"51818039",
          5155 => x"82bdf051",
          5156 => x"80f93982",
          5157 => x"be805180",
          5158 => x"f23982be",
          5159 => x"905180eb",
          5160 => x"3982bea0",
          5161 => x"5180e439",
          5162 => x"82beb051",
          5163 => x"80dd3982",
          5164 => x"bec45180",
          5165 => x"d63982be",
          5166 => x"d45180cf",
          5167 => x"3982beec",
          5168 => x"5180c839",
          5169 => x"82bf8451",
          5170 => x"80c13982",
          5171 => x"bf9c51bb",
          5172 => x"3982bfb8",
          5173 => x"51b53982",
          5174 => x"bfcc51af",
          5175 => x"3982bff4",
          5176 => x"51a93982",
          5177 => x"c08451a3",
          5178 => x"3982c0a4",
          5179 => x"519d3982",
          5180 => x"c0b45197",
          5181 => x"3982c0cc",
          5182 => x"51913982",
          5183 => x"c0e4518b",
          5184 => x"3982c0fc",
          5185 => x"51853982",
          5186 => x"c18851ce",
          5187 => x"8a3f833d",
          5188 => x"0d04fb3d",
          5189 => x"0d777956",
          5190 => x"567487e7",
          5191 => x"268a3874",
          5192 => x"527587e8",
          5193 => x"29519039",
          5194 => x"87e85274",
          5195 => x"51e3a43f",
          5196 => x"82e09808",
          5197 => x"527551e3",
          5198 => x"9a3f82e0",
          5199 => x"98085479",
          5200 => x"53755282",
          5201 => x"c19851ff",
          5202 => x"b1c23f87",
          5203 => x"3d0d04ec",
          5204 => x"3d0d6602",
          5205 => x"840580e3",
          5206 => x"05335b57",
          5207 => x"80687830",
          5208 => x"707a0773",
          5209 => x"25515759",
          5210 => x"59785677",
          5211 => x"87ff2683",
          5212 => x"38815674",
          5213 => x"76077081",
          5214 => x"ff065155",
          5215 => x"93567481",
          5216 => x"82388153",
          5217 => x"76528c3d",
          5218 => x"70525681",
          5219 => x"93993f82",
          5220 => x"e0980857",
          5221 => x"82e09808",
          5222 => x"b93882e0",
          5223 => x"980887c0",
          5224 => x"98880c82",
          5225 => x"e0980859",
          5226 => x"963dd405",
          5227 => x"54848053",
          5228 => x"77527551",
          5229 => x"8197d53f",
          5230 => x"82e09808",
          5231 => x"5782e098",
          5232 => x"0890387a",
          5233 => x"5574802e",
          5234 => x"89387419",
          5235 => x"75195959",
          5236 => x"d739963d",
          5237 => x"d8055181",
          5238 => x"9fcd3f76",
          5239 => x"30707807",
          5240 => x"80257b30",
          5241 => x"709f2a72",
          5242 => x"06515751",
          5243 => x"5674802e",
          5244 => x"903882c1",
          5245 => x"bc5387c0",
          5246 => x"98880852",
          5247 => x"7851fe92",
          5248 => x"3f765675",
          5249 => x"82e0980c",
          5250 => x"963d0d04",
          5251 => x"f83d0d7c",
          5252 => x"028405b7",
          5253 => x"05335859",
          5254 => x"ff588053",
          5255 => x"7b527a51",
          5256 => x"fead3f82",
          5257 => x"e09808a8",
          5258 => x"3876802e",
          5259 => x"88387681",
          5260 => x"2e9c389c",
          5261 => x"3982fbf8",
          5262 => x"56615560",
          5263 => x"5482e098",
          5264 => x"537f527e",
          5265 => x"51782d82",
          5266 => x"e0980858",
          5267 => x"83397804",
          5268 => x"7782e098",
          5269 => x"0c8a3d0d",
          5270 => x"04f33d0d",
          5271 => x"7f616302",
          5272 => x"8c0580cf",
          5273 => x"05337373",
          5274 => x"1568415f",
          5275 => x"5d5b5e5e",
          5276 => x"5e77a438",
          5277 => x"fbf13f82",
          5278 => x"e0980881",
          5279 => x"ff065388",
          5280 => x"5872a82e",
          5281 => x"92389058",
          5282 => x"7280d02e",
          5283 => x"8a388639",
          5284 => x"805382d2",
          5285 => x"39a0587a",
          5286 => x"5282c1c4",
          5287 => x"51ffaeec",
          5288 => x"3f82c1cc",
          5289 => x"51ffaee4",
          5290 => x"3f805574",
          5291 => x"78278180",
          5292 => x"387b902e",
          5293 => x"89387ba0",
          5294 => x"2ea73880",
          5295 => x"c6397419",
          5296 => x"53727a27",
          5297 => x"8e387222",
          5298 => x"5282c1d0",
          5299 => x"51ffaebc",
          5300 => x"3f893982",
          5301 => x"c1dc51ff",
          5302 => x"aeb23f82",
          5303 => x"155580c3",
          5304 => x"39741953",
          5305 => x"727a278e",
          5306 => x"38720852",
          5307 => x"82c1c451",
          5308 => x"ffae993f",
          5309 => x"893982c1",
          5310 => x"d851ffae",
          5311 => x"8f3f8415",
          5312 => x"55a13974",
          5313 => x"1953727a",
          5314 => x"278e3872",
          5315 => x"335282c1",
          5316 => x"e451ffad",
          5317 => x"f73f8939",
          5318 => x"82c1ec51",
          5319 => x"ffaded3f",
          5320 => x"81155582",
          5321 => x"fbfc0852",
          5322 => x"a051cdba",
          5323 => x"3ffefc39",
          5324 => x"82c1f051",
          5325 => x"ffadd53f",
          5326 => x"80557478",
          5327 => x"2780c638",
          5328 => x"74197033",
          5329 => x"55538056",
          5330 => x"727a2783",
          5331 => x"38815680",
          5332 => x"539f7427",
          5333 => x"83388153",
          5334 => x"75730670",
          5335 => x"81ff0651",
          5336 => x"5372802e",
          5337 => x"90387380",
          5338 => x"fe268a38",
          5339 => x"82fbfc08",
          5340 => x"52735188",
          5341 => x"3982fbfc",
          5342 => x"0852a051",
          5343 => x"cce83f81",
          5344 => x"1555ffb6",
          5345 => x"3982c1f4",
          5346 => x"51c98c3f",
          5347 => x"7719781c",
          5348 => x"5c598051",
          5349 => x"98e03f82",
          5350 => x"e0980898",
          5351 => x"2b70982c",
          5352 => x"515776a0",
          5353 => x"2e098106",
          5354 => x"ac388051",
          5355 => x"98c83f82",
          5356 => x"e0980898",
          5357 => x"2b70982c",
          5358 => x"70a03270",
          5359 => x"30729b32",
          5360 => x"70307072",
          5361 => x"07737507",
          5362 => x"06515858",
          5363 => x"59575157",
          5364 => x"807324d6",
          5365 => x"38769b2e",
          5366 => x"fdb6387c",
          5367 => x"1e537279",
          5368 => x"26fdb438",
          5369 => x"ff537282",
          5370 => x"e0980c8f",
          5371 => x"3d0d04fc",
          5372 => x"3d0d029b",
          5373 => x"0533558a",
          5374 => x"51cbbe3f",
          5375 => x"82c1f852",
          5376 => x"82c1fc51",
          5377 => x"ffac853f",
          5378 => x"82dee822",
          5379 => x"51a6d83f",
          5380 => x"82c28454",
          5381 => x"82c29053",
          5382 => x"82dee933",
          5383 => x"5282c298",
          5384 => x"51ffabe8",
          5385 => x"3f74802e",
          5386 => x"8438a289",
          5387 => x"3f863d0d",
          5388 => x"04fe3d0d",
          5389 => x"87c09680",
          5390 => x"0853a6f4",
          5391 => x"3f815199",
          5392 => x"bf3f82c2",
          5393 => x"b4519ad4",
          5394 => x"3f805199",
          5395 => x"b33f7281",
          5396 => x"2a708106",
          5397 => x"51527180",
          5398 => x"2e923881",
          5399 => x"5199a13f",
          5400 => x"82c2cc51",
          5401 => x"9ab63f80",
          5402 => x"5199953f",
          5403 => x"72822a70",
          5404 => x"81065152",
          5405 => x"71802e92",
          5406 => x"38815199",
          5407 => x"833f82c2",
          5408 => x"dc519a98",
          5409 => x"3f805198",
          5410 => x"f73f7283",
          5411 => x"2a708106",
          5412 => x"51527180",
          5413 => x"2e923881",
          5414 => x"5198e53f",
          5415 => x"82c2ec51",
          5416 => x"99fa3f80",
          5417 => x"5198d93f",
          5418 => x"72842a70",
          5419 => x"81065152",
          5420 => x"71802e92",
          5421 => x"38815198",
          5422 => x"c73f82c3",
          5423 => x"805199dc",
          5424 => x"3f805198",
          5425 => x"bb3f7285",
          5426 => x"2a708106",
          5427 => x"51527180",
          5428 => x"2e923881",
          5429 => x"5198a93f",
          5430 => x"82c39451",
          5431 => x"99be3f80",
          5432 => x"51989d3f",
          5433 => x"72862a70",
          5434 => x"81065152",
          5435 => x"71802e92",
          5436 => x"38815198",
          5437 => x"8b3f82c3",
          5438 => x"a85199a0",
          5439 => x"3f805197",
          5440 => x"ff3f7287",
          5441 => x"2a708106",
          5442 => x"51527180",
          5443 => x"2e923881",
          5444 => x"5197ed3f",
          5445 => x"82c3bc51",
          5446 => x"99823f80",
          5447 => x"5197e13f",
          5448 => x"72882a70",
          5449 => x"81065152",
          5450 => x"71802e92",
          5451 => x"38815197",
          5452 => x"cf3f82c3",
          5453 => x"d05198e4",
          5454 => x"3f805197",
          5455 => x"c33fa4f8",
          5456 => x"3f843d0d",
          5457 => x"04fb3d0d",
          5458 => x"77028405",
          5459 => x"a3053370",
          5460 => x"55565680",
          5461 => x"527551d9",
          5462 => x"ec3f0b0b",
          5463 => x"82db9c33",
          5464 => x"5473a938",
          5465 => x"815382c4",
          5466 => x"8c5282f7",
          5467 => x"a851818b",
          5468 => x"b63f82e0",
          5469 => x"98083070",
          5470 => x"82e09808",
          5471 => x"07802582",
          5472 => x"71315151",
          5473 => x"54730b0b",
          5474 => x"82db9c34",
          5475 => x"0b0b82db",
          5476 => x"9c335473",
          5477 => x"812e0981",
          5478 => x"06af3882",
          5479 => x"f7a85374",
          5480 => x"52755181",
          5481 => x"c7af3f82",
          5482 => x"e0980880",
          5483 => x"2e8b3882",
          5484 => x"e0980851",
          5485 => x"c4e13f91",
          5486 => x"3982f7a8",
          5487 => x"518197e7",
          5488 => x"3f820b0b",
          5489 => x"0b82db9c",
          5490 => x"340b0b82",
          5491 => x"db9c3354",
          5492 => x"73822e09",
          5493 => x"81068c38",
          5494 => x"82c49c53",
          5495 => x"74527551",
          5496 => x"aaf03f80",
          5497 => x"0b82e098",
          5498 => x"0c873d0d",
          5499 => x"04cd3d0d",
          5500 => x"8070415e",
          5501 => x"ff7e82f7",
          5502 => x"a40c5f81",
          5503 => x"527d5180",
          5504 => x"c88a3f82",
          5505 => x"e0980881",
          5506 => x"ff065978",
          5507 => x"7e2e0981",
          5508 => x"06a33897",
          5509 => x"3d598353",
          5510 => x"82c4a852",
          5511 => x"7851d1f9",
          5512 => x"3f7d5378",
          5513 => x"5282e1c4",
          5514 => x"5181899a",
          5515 => x"3f82e098",
          5516 => x"087e2e88",
          5517 => x"3882c4ac",
          5518 => x"518de539",
          5519 => x"8170415e",
          5520 => x"82c4e451",
          5521 => x"ffa7c53f",
          5522 => x"973d7047",
          5523 => x"5a80f852",
          5524 => x"7951fdf1",
          5525 => x"3fb53dff",
          5526 => x"840551f3",
          5527 => x"933f82e0",
          5528 => x"9808902b",
          5529 => x"70902c51",
          5530 => x"597880c2",
          5531 => x"2e87a538",
          5532 => x"7880c224",
          5533 => x"b23878bd",
          5534 => x"2e81d238",
          5535 => x"78bd2490",
          5536 => x"3878802e",
          5537 => x"ffba3878",
          5538 => x"bc2e80da",
          5539 => x"388adc39",
          5540 => x"7880c02e",
          5541 => x"83993878",
          5542 => x"80c02485",
          5543 => x"ce3878bf",
          5544 => x"2e828c38",
          5545 => x"8ac53978",
          5546 => x"80f92e89",
          5547 => x"df387880",
          5548 => x"f9249238",
          5549 => x"7880c32e",
          5550 => x"888d3878",
          5551 => x"80f82e89",
          5552 => x"a7388aa7",
          5553 => x"39788183",
          5554 => x"2e8a8d38",
          5555 => x"78818324",
          5556 => x"8b387881",
          5557 => x"822e89f1",
          5558 => x"388a9039",
          5559 => x"7881852e",
          5560 => x"8a83388a",
          5561 => x"8639b53d",
          5562 => x"ff801153",
          5563 => x"ff840551",
          5564 => x"ecad3f82",
          5565 => x"e0980880",
          5566 => x"2efec538",
          5567 => x"b53dfefc",
          5568 => x"1153ff84",
          5569 => x"0551ec97",
          5570 => x"3f82e098",
          5571 => x"08802efe",
          5572 => x"af38b53d",
          5573 => x"fef81153",
          5574 => x"ff840551",
          5575 => x"ec813f82",
          5576 => x"e0980886",
          5577 => x"3882e098",
          5578 => x"084382c4",
          5579 => x"e851ffa5",
          5580 => x"db3f6464",
          5581 => x"5c5a797b",
          5582 => x"2781ec38",
          5583 => x"6259787a",
          5584 => x"7084055c",
          5585 => x"0c7a7a26",
          5586 => x"f53881db",
          5587 => x"39b53dff",
          5588 => x"801153ff",
          5589 => x"840551eb",
          5590 => x"c63f82e0",
          5591 => x"9808802e",
          5592 => x"fdde38b5",
          5593 => x"3dfefc11",
          5594 => x"53ff8405",
          5595 => x"51ebb03f",
          5596 => x"82e09808",
          5597 => x"802efdc8",
          5598 => x"38b53dfe",
          5599 => x"f81153ff",
          5600 => x"840551eb",
          5601 => x"9a3f82e0",
          5602 => x"9808802e",
          5603 => x"fdb23882",
          5604 => x"c4f851ff",
          5605 => x"a4f63f64",
          5606 => x"5a796427",
          5607 => x"81893862",
          5608 => x"59797081",
          5609 => x"055b3379",
          5610 => x"34628105",
          5611 => x"43eb39b5",
          5612 => x"3dff8011",
          5613 => x"53ff8405",
          5614 => x"51eae43f",
          5615 => x"82e09808",
          5616 => x"802efcfc",
          5617 => x"38b53dfe",
          5618 => x"fc1153ff",
          5619 => x"840551ea",
          5620 => x"ce3f82e0",
          5621 => x"9808802e",
          5622 => x"fce638b5",
          5623 => x"3dfef811",
          5624 => x"53ff8405",
          5625 => x"51eab83f",
          5626 => x"82e09808",
          5627 => x"802efcd0",
          5628 => x"3882c584",
          5629 => x"51ffa494",
          5630 => x"3f645a79",
          5631 => x"6427a838",
          5632 => x"6270337b",
          5633 => x"335e5a5b",
          5634 => x"787c2e92",
          5635 => x"3878557a",
          5636 => x"54793353",
          5637 => x"795282c5",
          5638 => x"9451ffa3",
          5639 => x"ef3f811a",
          5640 => x"63810544",
          5641 => x"5ad5398a",
          5642 => x"51c38e3f",
          5643 => x"fc9239b5",
          5644 => x"3dff8011",
          5645 => x"53ff8405",
          5646 => x"51e9e43f",
          5647 => x"82e09808",
          5648 => x"80df3882",
          5649 => x"defc3359",
          5650 => x"78802e89",
          5651 => x"3882deb4",
          5652 => x"084580cd",
          5653 => x"3982defd",
          5654 => x"33597880",
          5655 => x"2e883882",
          5656 => x"debc0845",
          5657 => x"bc3982de",
          5658 => x"fe335978",
          5659 => x"802e8838",
          5660 => x"82dec408",
          5661 => x"45ab3982",
          5662 => x"deff3359",
          5663 => x"78802e88",
          5664 => x"3882decc",
          5665 => x"08459a39",
          5666 => x"82defa33",
          5667 => x"5978802e",
          5668 => x"883882de",
          5669 => x"d4084589",
          5670 => x"3982dee4",
          5671 => x"08fc8005",
          5672 => x"45b53dfe",
          5673 => x"fc1153ff",
          5674 => x"840551e8",
          5675 => x"f23f82e0",
          5676 => x"980880de",
          5677 => x"3882defc",
          5678 => x"33597880",
          5679 => x"2e893882",
          5680 => x"deb80844",
          5681 => x"80cc3982",
          5682 => x"defd3359",
          5683 => x"78802e88",
          5684 => x"3882dec0",
          5685 => x"0844bb39",
          5686 => x"82defe33",
          5687 => x"5978802e",
          5688 => x"883882de",
          5689 => x"c80844aa",
          5690 => x"3982deff",
          5691 => x"33597880",
          5692 => x"2e883882",
          5693 => x"ded00844",
          5694 => x"993982de",
          5695 => x"fa335978",
          5696 => x"802e8838",
          5697 => x"82ded808",
          5698 => x"44883982",
          5699 => x"dee40888",
          5700 => x"0544b53d",
          5701 => x"fef81153",
          5702 => x"ff840551",
          5703 => x"e8813f82",
          5704 => x"e0980880",
          5705 => x"2ea73880",
          5706 => x"635c5c7a",
          5707 => x"882e8338",
          5708 => x"815c7a90",
          5709 => x"32703070",
          5710 => x"72079f2a",
          5711 => x"707f0651",
          5712 => x"515a5a78",
          5713 => x"802e8838",
          5714 => x"7aa02e83",
          5715 => x"38884382",
          5716 => x"c5b051ff",
          5717 => x"bdc13f80",
          5718 => x"55645462",
          5719 => x"53635264",
          5720 => x"51f1f63f",
          5721 => x"82c5bc51",
          5722 => x"87b639b5",
          5723 => x"3dff8011",
          5724 => x"53ff8405",
          5725 => x"51e7a83f",
          5726 => x"82e09808",
          5727 => x"802ef9c0",
          5728 => x"38b53dfe",
          5729 => x"fc1153ff",
          5730 => x"840551e7",
          5731 => x"923f82e0",
          5732 => x"9808802e",
          5733 => x"a4386459",
          5734 => x"0280cf05",
          5735 => x"33793464",
          5736 => x"810545b5",
          5737 => x"3dfefc11",
          5738 => x"53ff8405",
          5739 => x"51e6f03f",
          5740 => x"82e09808",
          5741 => x"e138f988",
          5742 => x"39647033",
          5743 => x"545282c5",
          5744 => x"c851ffa0",
          5745 => x"c73f82fb",
          5746 => x"f8085380",
          5747 => x"f8527951",
          5748 => x"ffa18e3f",
          5749 => x"79467933",
          5750 => x"5978ae2e",
          5751 => x"f8e2389f",
          5752 => x"79279f38",
          5753 => x"b53dfefc",
          5754 => x"1153ff84",
          5755 => x"0551e6af",
          5756 => x"3f82e098",
          5757 => x"08802e91",
          5758 => x"38645902",
          5759 => x"80cf0533",
          5760 => x"79346481",
          5761 => x"0545ffb1",
          5762 => x"3982c5d4",
          5763 => x"51ffbc87",
          5764 => x"3fffa639",
          5765 => x"b53dfef4",
          5766 => x"1153ff84",
          5767 => x"0551e0ae",
          5768 => x"3f82e098",
          5769 => x"08802ef8",
          5770 => x"9738b53d",
          5771 => x"fef01153",
          5772 => x"ff840551",
          5773 => x"e0983f82",
          5774 => x"e0980880",
          5775 => x"2ea63861",
          5776 => x"590280c2",
          5777 => x"05227970",
          5778 => x"82055b23",
          5779 => x"7842b53d",
          5780 => x"fef01153",
          5781 => x"ff840551",
          5782 => x"dff43f82",
          5783 => x"e09808df",
          5784 => x"38f7dd39",
          5785 => x"61702254",
          5786 => x"5282c5d8",
          5787 => x"51ff9f9c",
          5788 => x"3f82fbf8",
          5789 => x"085380f8",
          5790 => x"527951ff",
          5791 => x"9fe33f79",
          5792 => x"46793359",
          5793 => x"78ae2ef7",
          5794 => x"b738789f",
          5795 => x"26873861",
          5796 => x"820542d0",
          5797 => x"39b53dfe",
          5798 => x"f01153ff",
          5799 => x"840551df",
          5800 => x"ad3f82e0",
          5801 => x"9808802e",
          5802 => x"93386159",
          5803 => x"0280c205",
          5804 => x"22797082",
          5805 => x"055b2378",
          5806 => x"42ffa939",
          5807 => x"82c5d451",
          5808 => x"ffbad43f",
          5809 => x"ff9e39b5",
          5810 => x"3dfef411",
          5811 => x"53ff8405",
          5812 => x"51defb3f",
          5813 => x"82e09808",
          5814 => x"802ef6e4",
          5815 => x"38b53dfe",
          5816 => x"f01153ff",
          5817 => x"840551de",
          5818 => x"e53f82e0",
          5819 => x"9808802e",
          5820 => x"a0386161",
          5821 => x"710c5961",
          5822 => x"840542b5",
          5823 => x"3dfef011",
          5824 => x"53ff8405",
          5825 => x"51dec73f",
          5826 => x"82e09808",
          5827 => x"e538f6b0",
          5828 => x"39617008",
          5829 => x"545282c5",
          5830 => x"e451ff9d",
          5831 => x"ef3f82fb",
          5832 => x"f8085380",
          5833 => x"f8527951",
          5834 => x"ff9eb63f",
          5835 => x"79467933",
          5836 => x"5978ae2e",
          5837 => x"f68a389f",
          5838 => x"79279b38",
          5839 => x"b53dfef0",
          5840 => x"1153ff84",
          5841 => x"0551de86",
          5842 => x"3f82e098",
          5843 => x"08802e8d",
          5844 => x"38616171",
          5845 => x"0c596184",
          5846 => x"0542ffb5",
          5847 => x"3982c5d4",
          5848 => x"51ffb9b3",
          5849 => x"3fffaa39",
          5850 => x"b53dff80",
          5851 => x"1153ff84",
          5852 => x"0551e3ab",
          5853 => x"3f82e098",
          5854 => x"08802ef5",
          5855 => x"c3386452",
          5856 => x"82c5f451",
          5857 => x"ff9d853f",
          5858 => x"64597804",
          5859 => x"b53dff80",
          5860 => x"1153ff84",
          5861 => x"0551e387",
          5862 => x"3f82e098",
          5863 => x"08802ef5",
          5864 => x"9f386452",
          5865 => x"82c69051",
          5866 => x"ff9ce13f",
          5867 => x"6459782d",
          5868 => x"82e09808",
          5869 => x"802ef588",
          5870 => x"3882e098",
          5871 => x"085282c6",
          5872 => x"ac51ff9c",
          5873 => x"c73ff4f8",
          5874 => x"3982c6c8",
          5875 => x"51ffb8c7",
          5876 => x"3fff9c99",
          5877 => x"3ff4e939",
          5878 => x"82c6e451",
          5879 => x"ffb8b83f",
          5880 => x"8059ffa6",
          5881 => x"3992ce3f",
          5882 => x"f4d63997",
          5883 => x"3d335978",
          5884 => x"802ef4cc",
          5885 => x"3880f852",
          5886 => x"7951c9f1",
          5887 => x"3f82e098",
          5888 => x"085d82e0",
          5889 => x"9808802e",
          5890 => x"82923882",
          5891 => x"e0980846",
          5892 => x"b53dff84",
          5893 => x"055183cc",
          5894 => x"3f82e098",
          5895 => x"08607f06",
          5896 => x"5a5c7880",
          5897 => x"2e81d238",
          5898 => x"82e09808",
          5899 => x"51c48a3f",
          5900 => x"82e09808",
          5901 => x"8f2681c1",
          5902 => x"38815b7a",
          5903 => x"822eb238",
          5904 => x"7a822489",
          5905 => x"387a812e",
          5906 => x"8c3880ca",
          5907 => x"397a832e",
          5908 => x"ad3880c2",
          5909 => x"3982c6f8",
          5910 => x"567b5582",
          5911 => x"c6fc5480",
          5912 => x"5382c780",
          5913 => x"52b53dff",
          5914 => x"b00551ff",
          5915 => x"9e863fb8",
          5916 => x"397b52b5",
          5917 => x"3dffb005",
          5918 => x"51c4ac3f",
          5919 => x"ab397b55",
          5920 => x"82c6fc54",
          5921 => x"805382c7",
          5922 => x"9052b53d",
          5923 => x"ffb00551",
          5924 => x"ff9de13f",
          5925 => x"93397b54",
          5926 => x"805382c7",
          5927 => x"9c52b53d",
          5928 => x"ffb00551",
          5929 => x"ff9dcd3f",
          5930 => x"82deb458",
          5931 => x"82e0c857",
          5932 => x"7c566555",
          5933 => x"80549080",
          5934 => x"0a539080",
          5935 => x"0a52b53d",
          5936 => x"ffb00551",
          5937 => x"eac63f82",
          5938 => x"e0980882",
          5939 => x"e0980809",
          5940 => x"70307072",
          5941 => x"07802551",
          5942 => x"5b5b5f80",
          5943 => x"5a7a8326",
          5944 => x"8338815a",
          5945 => x"787a0659",
          5946 => x"78802e8d",
          5947 => x"38811b70",
          5948 => x"81ff065c",
          5949 => x"597afec3",
          5950 => x"387f8132",
          5951 => x"7e813207",
          5952 => x"59788938",
          5953 => x"7eff2e09",
          5954 => x"81068938",
          5955 => x"82c7a451",
          5956 => x"ffb6843f",
          5957 => x"7c51b1f1",
          5958 => x"3ff2a539",
          5959 => x"82c7b451",
          5960 => x"ffb5f43f",
          5961 => x"f29a39f5",
          5962 => x"3d0d800b",
          5963 => x"82e0c834",
          5964 => x"87c0948c",
          5965 => x"70085455",
          5966 => x"87848052",
          5967 => x"7251cb93",
          5968 => x"3f82e098",
          5969 => x"08902b75",
          5970 => x"08555387",
          5971 => x"84805273",
          5972 => x"51cb803f",
          5973 => x"7282e098",
          5974 => x"0807750c",
          5975 => x"87c0949c",
          5976 => x"70085455",
          5977 => x"87848052",
          5978 => x"7251cae7",
          5979 => x"3f82e098",
          5980 => x"08902b75",
          5981 => x"08555387",
          5982 => x"84805273",
          5983 => x"51cad43f",
          5984 => x"7282e098",
          5985 => x"0807750c",
          5986 => x"8c80830b",
          5987 => x"87c09484",
          5988 => x"0c8c8083",
          5989 => x"0b87c094",
          5990 => x"940c8182",
          5991 => x"985a8185",
          5992 => x"845b8302",
          5993 => x"84059905",
          5994 => x"34805c82",
          5995 => x"fbf80b87",
          5996 => x"3d708813",
          5997 => x"0c70720c",
          5998 => x"82fbfc0c",
          5999 => x"548aaa3f",
          6000 => x"93ee3f82",
          6001 => x"c7e051ff",
          6002 => x"b4cd3f82",
          6003 => x"c7ec51ff",
          6004 => x"b4c53f80",
          6005 => x"e8b15193",
          6006 => x"d23f8151",
          6007 => x"ec913ff0",
          6008 => x"8c3f8004",
          6009 => x"fc3d0d76",
          6010 => x"70085455",
          6011 => x"80735254",
          6012 => x"72742e81",
          6013 => x"8a387233",
          6014 => x"5170a02e",
          6015 => x"09810686",
          6016 => x"38811353",
          6017 => x"f1397233",
          6018 => x"5170a22e",
          6019 => x"09810686",
          6020 => x"38811353",
          6021 => x"81547252",
          6022 => x"73812e09",
          6023 => x"81069f38",
          6024 => x"84398112",
          6025 => x"52807233",
          6026 => x"525470a2",
          6027 => x"2e833881",
          6028 => x"5470802e",
          6029 => x"9d3873ea",
          6030 => x"38983981",
          6031 => x"12528072",
          6032 => x"33525470",
          6033 => x"a02e8338",
          6034 => x"81547080",
          6035 => x"2e843873",
          6036 => x"ea388072",
          6037 => x"33525470",
          6038 => x"a02e0981",
          6039 => x"06833881",
          6040 => x"5470a232",
          6041 => x"70307080",
          6042 => x"25760751",
          6043 => x"51517080",
          6044 => x"2e883880",
          6045 => x"72708105",
          6046 => x"54347175",
          6047 => x"0c725170",
          6048 => x"82e0980c",
          6049 => x"863d0d04",
          6050 => x"fc3d0d76",
          6051 => x"53720880",
          6052 => x"2e913886",
          6053 => x"3dfc0552",
          6054 => x"7251d7b2",
          6055 => x"3f82e098",
          6056 => x"08853880",
          6057 => x"53833974",
          6058 => x"537282e0",
          6059 => x"980c863d",
          6060 => x"0d04fc3d",
          6061 => x"0d768211",
          6062 => x"33ff0552",
          6063 => x"53815270",
          6064 => x"8b268198",
          6065 => x"38831333",
          6066 => x"ff055182",
          6067 => x"52709e26",
          6068 => x"818a3884",
          6069 => x"13335183",
          6070 => x"52709726",
          6071 => x"80fe3885",
          6072 => x"13335184",
          6073 => x"5270bb26",
          6074 => x"80f23886",
          6075 => x"13335185",
          6076 => x"5270bb26",
          6077 => x"80e63888",
          6078 => x"13225586",
          6079 => x"527487e7",
          6080 => x"2680d938",
          6081 => x"8a132254",
          6082 => x"87527387",
          6083 => x"e72680cc",
          6084 => x"38810b87",
          6085 => x"c0989c0c",
          6086 => x"722287c0",
          6087 => x"98bc0c82",
          6088 => x"133387c0",
          6089 => x"98b80c83",
          6090 => x"133387c0",
          6091 => x"98b40c84",
          6092 => x"133387c0",
          6093 => x"98b00c85",
          6094 => x"133387c0",
          6095 => x"98ac0c86",
          6096 => x"133387c0",
          6097 => x"98a80c74",
          6098 => x"87c098a4",
          6099 => x"0c7387c0",
          6100 => x"98a00c80",
          6101 => x"0b87c098",
          6102 => x"9c0c8052",
          6103 => x"7182e098",
          6104 => x"0c863d0d",
          6105 => x"04f33d0d",
          6106 => x"7f5b87c0",
          6107 => x"989c5d81",
          6108 => x"7d0c87c0",
          6109 => x"98bc085e",
          6110 => x"7d7b2387",
          6111 => x"c098b808",
          6112 => x"5a79821c",
          6113 => x"3487c098",
          6114 => x"b4085a79",
          6115 => x"831c3487",
          6116 => x"c098b008",
          6117 => x"5a79841c",
          6118 => x"3487c098",
          6119 => x"ac085a79",
          6120 => x"851c3487",
          6121 => x"c098a808",
          6122 => x"5a79861c",
          6123 => x"3487c098",
          6124 => x"a4085c7b",
          6125 => x"881c2387",
          6126 => x"c098a008",
          6127 => x"5a798a1c",
          6128 => x"23807d0c",
          6129 => x"7983ffff",
          6130 => x"06597b83",
          6131 => x"ffff0658",
          6132 => x"861b3357",
          6133 => x"851b3356",
          6134 => x"841b3355",
          6135 => x"831b3354",
          6136 => x"821b3353",
          6137 => x"7d83ffff",
          6138 => x"065282c8",
          6139 => x"8451ff94",
          6140 => x"9b3f8f3d",
          6141 => x"0d04fd3d",
          6142 => x"0d029705",
          6143 => x"33538052",
          6144 => x"72812e09",
          6145 => x"81068338",
          6146 => x"72527283",
          6147 => x"32703070",
          6148 => x"80257407",
          6149 => x"51515170",
          6150 => x"802e8638",
          6151 => x"84973f84",
          6152 => x"3984f03f",
          6153 => x"82e09808",
          6154 => x"982b7098",
          6155 => x"2c515271",
          6156 => x"ff2e0981",
          6157 => x"069e3880",
          6158 => x"5472812e",
          6159 => x"09810683",
          6160 => x"38725472",
          6161 => x"83327030",
          6162 => x"70802576",
          6163 => x"07515151",
          6164 => x"70ffab38",
          6165 => x"7182e098",
          6166 => x"0c853d0d",
          6167 => x"04fd3d0d",
          6168 => x"80538354",
          6169 => x"72882b53",
          6170 => x"8151ff8a",
          6171 => x"3f82e098",
          6172 => x"08982b70",
          6173 => x"982c7407",
          6174 => x"ff165654",
          6175 => x"52738025",
          6176 => x"e3387282",
          6177 => x"e0980c85",
          6178 => x"3d0d04fb",
          6179 => x"3d0d029f",
          6180 => x"053382de",
          6181 => x"b0337081",
          6182 => x"ff065855",
          6183 => x"5587c094",
          6184 => x"84517580",
          6185 => x"2e863887",
          6186 => x"c0949451",
          6187 => x"70087096",
          6188 => x"2a708106",
          6189 => x"53545270",
          6190 => x"802e8c38",
          6191 => x"71912a70",
          6192 => x"81065151",
          6193 => x"70d73872",
          6194 => x"81327081",
          6195 => x"06515170",
          6196 => x"802e8d38",
          6197 => x"71932a70",
          6198 => x"81065151",
          6199 => x"70ffbe38",
          6200 => x"7381ff06",
          6201 => x"5187c094",
          6202 => x"80527080",
          6203 => x"2e863887",
          6204 => x"c0949052",
          6205 => x"74720c74",
          6206 => x"82e0980c",
          6207 => x"873d0d04",
          6208 => x"ff3d0d02",
          6209 => x"8f053370",
          6210 => x"30709f2a",
          6211 => x"51525270",
          6212 => x"82deb034",
          6213 => x"833d0d04",
          6214 => x"f93d0d02",
          6215 => x"a7053358",
          6216 => x"778a2e09",
          6217 => x"81068738",
          6218 => x"7a528d51",
          6219 => x"eb3f82de",
          6220 => x"b0337081",
          6221 => x"ff065856",
          6222 => x"87c09484",
          6223 => x"5376802e",
          6224 => x"863887c0",
          6225 => x"94945372",
          6226 => x"0870962a",
          6227 => x"70810655",
          6228 => x"56547280",
          6229 => x"2e8c3873",
          6230 => x"912a7081",
          6231 => x"06515372",
          6232 => x"d7387481",
          6233 => x"32708106",
          6234 => x"51537280",
          6235 => x"2e8d3873",
          6236 => x"932a7081",
          6237 => x"06515372",
          6238 => x"ffbe3875",
          6239 => x"81ff0653",
          6240 => x"87c09480",
          6241 => x"5472802e",
          6242 => x"863887c0",
          6243 => x"94905477",
          6244 => x"740c800b",
          6245 => x"82e0980c",
          6246 => x"893d0d04",
          6247 => x"f93d0d79",
          6248 => x"54807433",
          6249 => x"7081ff06",
          6250 => x"53535770",
          6251 => x"772e80fc",
          6252 => x"387181ff",
          6253 => x"06811582",
          6254 => x"deb03370",
          6255 => x"81ff0659",
          6256 => x"57555887",
          6257 => x"c0948451",
          6258 => x"75802e86",
          6259 => x"3887c094",
          6260 => x"94517008",
          6261 => x"70962a70",
          6262 => x"81065354",
          6263 => x"5270802e",
          6264 => x"8c387191",
          6265 => x"2a708106",
          6266 => x"515170d7",
          6267 => x"38728132",
          6268 => x"70810651",
          6269 => x"5170802e",
          6270 => x"8d387193",
          6271 => x"2a708106",
          6272 => x"515170ff",
          6273 => x"be387481",
          6274 => x"ff065187",
          6275 => x"c0948052",
          6276 => x"70802e86",
          6277 => x"3887c094",
          6278 => x"90527772",
          6279 => x"0c811774",
          6280 => x"337081ff",
          6281 => x"06535357",
          6282 => x"70ff8638",
          6283 => x"7682e098",
          6284 => x"0c893d0d",
          6285 => x"04fe3d0d",
          6286 => x"82deb033",
          6287 => x"7081ff06",
          6288 => x"545287c0",
          6289 => x"94845172",
          6290 => x"802e8638",
          6291 => x"87c09494",
          6292 => x"51700870",
          6293 => x"822a7081",
          6294 => x"06515151",
          6295 => x"70802ee2",
          6296 => x"387181ff",
          6297 => x"065187c0",
          6298 => x"94805270",
          6299 => x"802e8638",
          6300 => x"87c09490",
          6301 => x"52710870",
          6302 => x"81ff0682",
          6303 => x"e0980c51",
          6304 => x"843d0d04",
          6305 => x"ffaf3f82",
          6306 => x"e0980881",
          6307 => x"ff0682e0",
          6308 => x"980c04fe",
          6309 => x"3d0d82de",
          6310 => x"b0337081",
          6311 => x"ff065253",
          6312 => x"87c09484",
          6313 => x"5270802e",
          6314 => x"863887c0",
          6315 => x"94945271",
          6316 => x"0870822a",
          6317 => x"70810651",
          6318 => x"5151ff52",
          6319 => x"70802ea0",
          6320 => x"387281ff",
          6321 => x"065187c0",
          6322 => x"94805270",
          6323 => x"802e8638",
          6324 => x"87c09490",
          6325 => x"52710870",
          6326 => x"982b7098",
          6327 => x"2c515351",
          6328 => x"7182e098",
          6329 => x"0c843d0d",
          6330 => x"04ff3d0d",
          6331 => x"87c09e80",
          6332 => x"08709c2a",
          6333 => x"8a065151",
          6334 => x"70802e84",
          6335 => x"b43887c0",
          6336 => x"9ea40882",
          6337 => x"deb40c87",
          6338 => x"c09ea808",
          6339 => x"82deb80c",
          6340 => x"87c09e94",
          6341 => x"0882debc",
          6342 => x"0c87c09e",
          6343 => x"980882de",
          6344 => x"c00c87c0",
          6345 => x"9e9c0882",
          6346 => x"dec40c87",
          6347 => x"c09ea008",
          6348 => x"82dec80c",
          6349 => x"87c09eac",
          6350 => x"0882decc",
          6351 => x"0c87c09e",
          6352 => x"b00882de",
          6353 => x"d00c87c0",
          6354 => x"9eb40882",
          6355 => x"ded40c87",
          6356 => x"c09eb808",
          6357 => x"82ded80c",
          6358 => x"87c09ebc",
          6359 => x"0882dedc",
          6360 => x"0c87c09e",
          6361 => x"c00882de",
          6362 => x"e00c87c0",
          6363 => x"9ec40882",
          6364 => x"dee40c87",
          6365 => x"c09e8008",
          6366 => x"517082de",
          6367 => x"e82387c0",
          6368 => x"9e840882",
          6369 => x"deec0c87",
          6370 => x"c09e8808",
          6371 => x"82def00c",
          6372 => x"87c09e8c",
          6373 => x"0882def4",
          6374 => x"0c810b82",
          6375 => x"def83480",
          6376 => x"0b87c09e",
          6377 => x"90087084",
          6378 => x"800a0651",
          6379 => x"52527080",
          6380 => x"2e833881",
          6381 => x"527182de",
          6382 => x"f934800b",
          6383 => x"87c09e90",
          6384 => x"08708880",
          6385 => x"0a065152",
          6386 => x"5270802e",
          6387 => x"83388152",
          6388 => x"7182defa",
          6389 => x"34800b87",
          6390 => x"c09e9008",
          6391 => x"7090800a",
          6392 => x"06515252",
          6393 => x"70802e83",
          6394 => x"38815271",
          6395 => x"82defb34",
          6396 => x"800b87c0",
          6397 => x"9e900870",
          6398 => x"88808006",
          6399 => x"51525270",
          6400 => x"802e8338",
          6401 => x"81527182",
          6402 => x"defc3480",
          6403 => x"0b87c09e",
          6404 => x"900870a0",
          6405 => x"80800651",
          6406 => x"52527080",
          6407 => x"2e833881",
          6408 => x"527182de",
          6409 => x"fd34800b",
          6410 => x"87c09e90",
          6411 => x"08709080",
          6412 => x"80065152",
          6413 => x"5270802e",
          6414 => x"83388152",
          6415 => x"7182defe",
          6416 => x"34800b87",
          6417 => x"c09e9008",
          6418 => x"70848080",
          6419 => x"06515252",
          6420 => x"70802e83",
          6421 => x"38815271",
          6422 => x"82deff34",
          6423 => x"800b87c0",
          6424 => x"9e900870",
          6425 => x"82808006",
          6426 => x"51525270",
          6427 => x"802e8338",
          6428 => x"81527182",
          6429 => x"df803480",
          6430 => x"0b87c09e",
          6431 => x"90087081",
          6432 => x"80800651",
          6433 => x"52527080",
          6434 => x"2e833881",
          6435 => x"527182df",
          6436 => x"8134800b",
          6437 => x"87c09e90",
          6438 => x"087080c0",
          6439 => x"80065152",
          6440 => x"5270802e",
          6441 => x"83388152",
          6442 => x"7182df82",
          6443 => x"34800b87",
          6444 => x"c09e9008",
          6445 => x"70a08006",
          6446 => x"51525270",
          6447 => x"802e8338",
          6448 => x"81527182",
          6449 => x"df833487",
          6450 => x"c09e9008",
          6451 => x"70988006",
          6452 => x"708a2a51",
          6453 => x"51517082",
          6454 => x"df843480",
          6455 => x"0b87c09e",
          6456 => x"90087084",
          6457 => x"80065152",
          6458 => x"5270802e",
          6459 => x"83388152",
          6460 => x"7182df85",
          6461 => x"3487c09e",
          6462 => x"90087083",
          6463 => x"f0067084",
          6464 => x"2a515151",
          6465 => x"7082df86",
          6466 => x"34800b87",
          6467 => x"c09e9008",
          6468 => x"70880651",
          6469 => x"52527080",
          6470 => x"2e833881",
          6471 => x"527182df",
          6472 => x"873487c0",
          6473 => x"9e900870",
          6474 => x"87065151",
          6475 => x"7082df88",
          6476 => x"34833d0d",
          6477 => x"04fb3d0d",
          6478 => x"82c89c51",
          6479 => x"ff89cd3f",
          6480 => x"82def833",
          6481 => x"5473802e",
          6482 => x"893882c8",
          6483 => x"b051ff89",
          6484 => x"bb3f82c8",
          6485 => x"c451ffa5",
          6486 => x"be3f82de",
          6487 => x"fa335473",
          6488 => x"802e9438",
          6489 => x"82ded408",
          6490 => x"82ded808",
          6491 => x"11545282",
          6492 => x"c8dc51ff",
          6493 => x"89963f82",
          6494 => x"deff3354",
          6495 => x"73802e94",
          6496 => x"3882decc",
          6497 => x"0882ded0",
          6498 => x"08115452",
          6499 => x"82c8f851",
          6500 => x"ff88f93f",
          6501 => x"82defc33",
          6502 => x"5473802e",
          6503 => x"943882de",
          6504 => x"b40882de",
          6505 => x"b8081154",
          6506 => x"5282c994",
          6507 => x"51ff88dc",
          6508 => x"3f82defd",
          6509 => x"33547380",
          6510 => x"2e943882",
          6511 => x"debc0882",
          6512 => x"dec00811",
          6513 => x"545282c9",
          6514 => x"b051ff88",
          6515 => x"bf3f82de",
          6516 => x"fe335473",
          6517 => x"802e9438",
          6518 => x"82dec408",
          6519 => x"82dec808",
          6520 => x"11545282",
          6521 => x"c9cc51ff",
          6522 => x"88a23f82",
          6523 => x"df833354",
          6524 => x"73802e8e",
          6525 => x"3882df84",
          6526 => x"335282c9",
          6527 => x"e851ff88",
          6528 => x"8b3f82df",
          6529 => x"87335473",
          6530 => x"802e8e38",
          6531 => x"82df8833",
          6532 => x"5282ca88",
          6533 => x"51ff87f4",
          6534 => x"3f82df85",
          6535 => x"33547380",
          6536 => x"2e8e3882",
          6537 => x"df863352",
          6538 => x"82caa851",
          6539 => x"ff87dd3f",
          6540 => x"82def933",
          6541 => x"5473802e",
          6542 => x"893882ca",
          6543 => x"c851ffa3",
          6544 => x"d63f82de",
          6545 => x"fb335473",
          6546 => x"802e8938",
          6547 => x"82cadc51",
          6548 => x"ffa3c43f",
          6549 => x"82df8033",
          6550 => x"5473802e",
          6551 => x"893882ca",
          6552 => x"e851ffa3",
          6553 => x"b23f82df",
          6554 => x"81335473",
          6555 => x"802e8938",
          6556 => x"82caf451",
          6557 => x"ffa3a03f",
          6558 => x"82df8233",
          6559 => x"5473802e",
          6560 => x"893882ca",
          6561 => x"fc51ffa3",
          6562 => x"8e3f82cb",
          6563 => x"8451ffa3",
          6564 => x"863f82de",
          6565 => x"dc085282",
          6566 => x"cb9051ff",
          6567 => x"86ee3f82",
          6568 => x"dee00852",
          6569 => x"82cbb851",
          6570 => x"ff86e13f",
          6571 => x"82dee408",
          6572 => x"5282cbe0",
          6573 => x"51ff86d4",
          6574 => x"3f82cc88",
          6575 => x"51ffa2d7",
          6576 => x"3f82dee8",
          6577 => x"225282cc",
          6578 => x"9051ff86",
          6579 => x"bf3f82de",
          6580 => x"ec0856bd",
          6581 => x"84c05275",
          6582 => x"51ffb7f7",
          6583 => x"3f82e098",
          6584 => x"08bd84c0",
          6585 => x"29767131",
          6586 => x"545482e0",
          6587 => x"98085282",
          6588 => x"ccb851ff",
          6589 => x"86963f82",
          6590 => x"deff3354",
          6591 => x"73802eaa",
          6592 => x"3882def0",
          6593 => x"0856bd84",
          6594 => x"c0527551",
          6595 => x"ffb7c43f",
          6596 => x"82e09808",
          6597 => x"bd84c029",
          6598 => x"76713154",
          6599 => x"5482e098",
          6600 => x"085282cc",
          6601 => x"e451ff85",
          6602 => x"e33f82de",
          6603 => x"fa335473",
          6604 => x"802eaa38",
          6605 => x"82def408",
          6606 => x"56bd84c0",
          6607 => x"527551ff",
          6608 => x"b7913f82",
          6609 => x"e09808bd",
          6610 => x"84c02976",
          6611 => x"71315454",
          6612 => x"82e09808",
          6613 => x"5282cd90",
          6614 => x"51ff85b0",
          6615 => x"3f8a51ff",
          6616 => x"a4d73f87",
          6617 => x"3d0d04fe",
          6618 => x"3d0d0292",
          6619 => x"0533ff05",
          6620 => x"52718426",
          6621 => x"aa387184",
          6622 => x"2982b8cc",
          6623 => x"05527108",
          6624 => x"0482cdbc",
          6625 => x"519d3982",
          6626 => x"cdc45197",
          6627 => x"3982cdcc",
          6628 => x"51913982",
          6629 => x"cdd4518b",
          6630 => x"3982cdd8",
          6631 => x"51853982",
          6632 => x"cde051ff",
          6633 => x"84e63f84",
          6634 => x"3d0d0471",
          6635 => x"88800c04",
          6636 => x"800b87c0",
          6637 => x"96840c04",
          6638 => x"82df8c08",
          6639 => x"87c09684",
          6640 => x"0c04fd3d",
          6641 => x"0d76982b",
          6642 => x"70982c79",
          6643 => x"982b7098",
          6644 => x"2c721013",
          6645 => x"70822b51",
          6646 => x"53515451",
          6647 => x"51800b82",
          6648 => x"cdec1233",
          6649 => x"55537174",
          6650 => x"259c3882",
          6651 => x"cde81108",
          6652 => x"12028405",
          6653 => x"97053371",
          6654 => x"33525252",
          6655 => x"70722e09",
          6656 => x"81068338",
          6657 => x"81537282",
          6658 => x"e0980c85",
          6659 => x"3d0d04fb",
          6660 => x"3d0d7902",
          6661 => x"8405a305",
          6662 => x"33713355",
          6663 => x"56547280",
          6664 => x"2eb13882",
          6665 => x"fbfc0852",
          6666 => x"8851ffa3",
          6667 => x"b93f82fb",
          6668 => x"fc0852a0",
          6669 => x"51ffa3ae",
          6670 => x"3f82fbfc",
          6671 => x"08528851",
          6672 => x"ffa3a33f",
          6673 => x"7333ff05",
          6674 => x"53727434",
          6675 => x"7281ff06",
          6676 => x"53cc3977",
          6677 => x"51ff83b4",
          6678 => x"3f747434",
          6679 => x"873d0d04",
          6680 => x"f63d0d7c",
          6681 => x"028405b7",
          6682 => x"05330288",
          6683 => x"05bb0533",
          6684 => x"82dfe833",
          6685 => x"70842982",
          6686 => x"df900570",
          6687 => x"08515959",
          6688 => x"5a585974",
          6689 => x"802e8638",
          6690 => x"74519afd",
          6691 => x"3f82dfe8",
          6692 => x"33708429",
          6693 => x"82df9005",
          6694 => x"81197054",
          6695 => x"58565a9d",
          6696 => x"fe3f82e0",
          6697 => x"9808750c",
          6698 => x"82dfe833",
          6699 => x"70842982",
          6700 => x"df900570",
          6701 => x"0851565a",
          6702 => x"74802ea7",
          6703 => x"38755378",
          6704 => x"527451ff",
          6705 => x"acd33f82",
          6706 => x"dfe83381",
          6707 => x"05557482",
          6708 => x"dfe83474",
          6709 => x"81ff0655",
          6710 => x"93752787",
          6711 => x"38800b82",
          6712 => x"dfe83477",
          6713 => x"802eb638",
          6714 => x"82dfe408",
          6715 => x"5675802e",
          6716 => x"ac3882df",
          6717 => x"e0335574",
          6718 => x"a4388c3d",
          6719 => x"fc055476",
          6720 => x"53785275",
          6721 => x"5180ec84",
          6722 => x"3f82dfe4",
          6723 => x"08528a51",
          6724 => x"81a2d63f",
          6725 => x"82dfe408",
          6726 => x"5180efe8",
          6727 => x"3f8c3d0d",
          6728 => x"04fd3d0d",
          6729 => x"82df9053",
          6730 => x"93547208",
          6731 => x"5271802e",
          6732 => x"89387151",
          6733 => x"99d33f80",
          6734 => x"730cff14",
          6735 => x"84145454",
          6736 => x"738025e6",
          6737 => x"38800b82",
          6738 => x"dfe83482",
          6739 => x"dfe40852",
          6740 => x"71802e95",
          6741 => x"38715180",
          6742 => x"f0cd3f82",
          6743 => x"dfe40851",
          6744 => x"99a73f80",
          6745 => x"0b82dfe4",
          6746 => x"0c853d0d",
          6747 => x"04dc3d0d",
          6748 => x"81578052",
          6749 => x"82dfe408",
          6750 => x"5180f5e9",
          6751 => x"3f82e098",
          6752 => x"0880d338",
          6753 => x"82dfe408",
          6754 => x"5380f852",
          6755 => x"883d7052",
          6756 => x"56819fc1",
          6757 => x"3f82e098",
          6758 => x"08802eba",
          6759 => x"387551ff",
          6760 => x"a9973f82",
          6761 => x"e0980855",
          6762 => x"800b82e0",
          6763 => x"9808259d",
          6764 => x"3882e098",
          6765 => x"08ff0570",
          6766 => x"17555580",
          6767 => x"74347553",
          6768 => x"76528117",
          6769 => x"82d0dc52",
          6770 => x"57ff80c0",
          6771 => x"3f74ff2e",
          6772 => x"098106ff",
          6773 => x"af38a63d",
          6774 => x"0d04d93d",
          6775 => x"0daa3d08",
          6776 => x"ad3d085a",
          6777 => x"5a817058",
          6778 => x"58805282",
          6779 => x"dfe40851",
          6780 => x"80f4f23f",
          6781 => x"82e09808",
          6782 => x"819538ff",
          6783 => x"0b82dfe4",
          6784 => x"08545580",
          6785 => x"f8528b3d",
          6786 => x"70525681",
          6787 => x"9ec73f82",
          6788 => x"e0980880",
          6789 => x"2ea53875",
          6790 => x"51ffa89d",
          6791 => x"3f82e098",
          6792 => x"08811858",
          6793 => x"55800b82",
          6794 => x"e0980825",
          6795 => x"8e3882e0",
          6796 => x"9808ff05",
          6797 => x"70175555",
          6798 => x"80743474",
          6799 => x"09703070",
          6800 => x"72079f2a",
          6801 => x"51555578",
          6802 => x"772e8538",
          6803 => x"73ffac38",
          6804 => x"82dfe408",
          6805 => x"8c110853",
          6806 => x"5180f489",
          6807 => x"3f82e098",
          6808 => x"08802e89",
          6809 => x"3882d0e8",
          6810 => x"51feffa0",
          6811 => x"3f78772e",
          6812 => x"0981069b",
          6813 => x"38755279",
          6814 => x"51ffa8ab",
          6815 => x"3f7951ff",
          6816 => x"a7b73fab",
          6817 => x"3d085482",
          6818 => x"e0980874",
          6819 => x"34805877",
          6820 => x"82e0980c",
          6821 => x"a93d0d04",
          6822 => x"f63d0d7c",
          6823 => x"7e715c71",
          6824 => x"72335759",
          6825 => x"5a5873a0",
          6826 => x"2e098106",
          6827 => x"a2387833",
          6828 => x"78055677",
          6829 => x"76279838",
          6830 => x"8117705b",
          6831 => x"70713356",
          6832 => x"585573a0",
          6833 => x"2e098106",
          6834 => x"86387575",
          6835 => x"26ea3880",
          6836 => x"54738829",
          6837 => x"82dfec05",
          6838 => x"70085255",
          6839 => x"ffa6da3f",
          6840 => x"82e09808",
          6841 => x"53795274",
          6842 => x"0851ffa9",
          6843 => x"d93f82e0",
          6844 => x"980880c5",
          6845 => x"38841533",
          6846 => x"5574812e",
          6847 => x"88387482",
          6848 => x"2e8838b5",
          6849 => x"39fce63f",
          6850 => x"ac39811a",
          6851 => x"5a8c3dfc",
          6852 => x"1153f805",
          6853 => x"51c4883f",
          6854 => x"82e09808",
          6855 => x"802e9a38",
          6856 => x"ff1b5378",
          6857 => x"527751fd",
          6858 => x"b13f82e0",
          6859 => x"980881ff",
          6860 => x"06557485",
          6861 => x"38745491",
          6862 => x"39811470",
          6863 => x"81ff0651",
          6864 => x"54827427",
          6865 => x"ff8b3880",
          6866 => x"547382e0",
          6867 => x"980c8c3d",
          6868 => x"0d04d33d",
          6869 => x"0db03d08",
          6870 => x"b23d08b4",
          6871 => x"3d08595f",
          6872 => x"5a800baf",
          6873 => x"3d3482df",
          6874 => x"e83382df",
          6875 => x"e408555b",
          6876 => x"7381cb38",
          6877 => x"7382dfe0",
          6878 => x"33555573",
          6879 => x"83388155",
          6880 => x"76802e81",
          6881 => x"bc388170",
          6882 => x"76065556",
          6883 => x"73802e81",
          6884 => x"ad38a851",
          6885 => x"98893f82",
          6886 => x"e0980882",
          6887 => x"dfe40c82",
          6888 => x"e0980880",
          6889 => x"2e819238",
          6890 => x"93537652",
          6891 => x"82e09808",
          6892 => x"5180def3",
          6893 => x"3f82e098",
          6894 => x"08802e8c",
          6895 => x"3882d194",
          6896 => x"51ff98d3",
          6897 => x"3f80f739",
          6898 => x"82e09808",
          6899 => x"5b82dfe4",
          6900 => x"085380f8",
          6901 => x"52903d70",
          6902 => x"5254819a",
          6903 => x"f83f82e0",
          6904 => x"98085682",
          6905 => x"e0980874",
          6906 => x"2e098106",
          6907 => x"80d03882",
          6908 => x"e0980851",
          6909 => x"ffa4c23f",
          6910 => x"82e09808",
          6911 => x"55800b82",
          6912 => x"e0980825",
          6913 => x"a93882e0",
          6914 => x"9808ff05",
          6915 => x"70175555",
          6916 => x"80743480",
          6917 => x"537481ff",
          6918 => x"06527551",
          6919 => x"f8c23f81",
          6920 => x"1b7081ff",
          6921 => x"065c5493",
          6922 => x"7b278338",
          6923 => x"805b74ff",
          6924 => x"2e098106",
          6925 => x"ff973886",
          6926 => x"397582df",
          6927 => x"e034768c",
          6928 => x"3882dfe4",
          6929 => x"08802e84",
          6930 => x"38f9d63f",
          6931 => x"8f3d5d80",
          6932 => x"51e7a33f",
          6933 => x"82e09808",
          6934 => x"982b7098",
          6935 => x"2c515978",
          6936 => x"ff2eec38",
          6937 => x"7881ff06",
          6938 => x"82f7d433",
          6939 => x"70982b70",
          6940 => x"982c82f7",
          6941 => x"d0337098",
          6942 => x"2b70972c",
          6943 => x"71982c05",
          6944 => x"70842982",
          6945 => x"cde80570",
          6946 => x"08157033",
          6947 => x"51515151",
          6948 => x"59595159",
          6949 => x"5d588156",
          6950 => x"73782e80",
          6951 => x"e9387774",
          6952 => x"27b43874",
          6953 => x"81800a29",
          6954 => x"81ff0a05",
          6955 => x"70982c51",
          6956 => x"55807524",
          6957 => x"80ce3876",
          6958 => x"53745277",
          6959 => x"51f6833f",
          6960 => x"82e09808",
          6961 => x"81ff0654",
          6962 => x"73802ed7",
          6963 => x"387482f7",
          6964 => x"d0348156",
          6965 => x"b1397481",
          6966 => x"800a2981",
          6967 => x"800a0570",
          6968 => x"982c7081",
          6969 => x"ff065651",
          6970 => x"55739526",
          6971 => x"97387653",
          6972 => x"74527751",
          6973 => x"f5cc3f82",
          6974 => x"e0980881",
          6975 => x"ff065473",
          6976 => x"cc38d339",
          6977 => x"80567580",
          6978 => x"2e80ca38",
          6979 => x"811c5574",
          6980 => x"82f7d434",
          6981 => x"74982b70",
          6982 => x"982c82f7",
          6983 => x"d0337098",
          6984 => x"2b70982c",
          6985 => x"70101170",
          6986 => x"822b82cd",
          6987 => x"ec11335e",
          6988 => x"51515157",
          6989 => x"58515574",
          6990 => x"772e0981",
          6991 => x"06fe9038",
          6992 => x"82cdf014",
          6993 => x"087d0c80",
          6994 => x"0b82f7d4",
          6995 => x"34800b82",
          6996 => x"f7d03492",
          6997 => x"397582f7",
          6998 => x"d4347582",
          6999 => x"f7d03478",
          7000 => x"af3d3475",
          7001 => x"7d0c7e54",
          7002 => x"739526fd",
          7003 => x"df387384",
          7004 => x"2982b8e0",
          7005 => x"05547308",
          7006 => x"0482f7dc",
          7007 => x"3354737e",
          7008 => x"2efdc938",
          7009 => x"82f7d833",
          7010 => x"55737527",
          7011 => x"ab387498",
          7012 => x"2b70982c",
          7013 => x"51557375",
          7014 => x"249e3874",
          7015 => x"1a547333",
          7016 => x"81153474",
          7017 => x"81800a29",
          7018 => x"81ff0a05",
          7019 => x"70982c82",
          7020 => x"f7dc3356",
          7021 => x"5155df39",
          7022 => x"82f7dc33",
          7023 => x"81115654",
          7024 => x"7482f7dc",
          7025 => x"34731a54",
          7026 => x"ae3d3374",
          7027 => x"3482f7d8",
          7028 => x"3354737e",
          7029 => x"25893881",
          7030 => x"14547382",
          7031 => x"f7d83482",
          7032 => x"f7dc3370",
          7033 => x"81800a29",
          7034 => x"81ff0a05",
          7035 => x"70982c82",
          7036 => x"f7d8335a",
          7037 => x"51565674",
          7038 => x"7725a838",
          7039 => x"82fbfc08",
          7040 => x"52741a70",
          7041 => x"335254ff",
          7042 => x"97dc3f74",
          7043 => x"81800a29",
          7044 => x"81800a05",
          7045 => x"70982c82",
          7046 => x"f7d83356",
          7047 => x"51557375",
          7048 => x"24da3882",
          7049 => x"f7dc3370",
          7050 => x"982b7098",
          7051 => x"2c82f7d8",
          7052 => x"335a5156",
          7053 => x"56747725",
          7054 => x"fc923882",
          7055 => x"fbfc0852",
          7056 => x"8851ff97",
          7057 => x"a13f7481",
          7058 => x"800a2981",
          7059 => x"800a0570",
          7060 => x"982c82f7",
          7061 => x"d8335651",
          7062 => x"55737524",
          7063 => x"de38fbec",
          7064 => x"39837a34",
          7065 => x"800b811b",
          7066 => x"3482f7dc",
          7067 => x"53805282",
          7068 => x"c1b851f3",
          7069 => x"9a3f81fd",
          7070 => x"3982f7dc",
          7071 => x"337081ff",
          7072 => x"06555573",
          7073 => x"802efbc4",
          7074 => x"3882f7d8",
          7075 => x"33ff0554",
          7076 => x"7382f7d8",
          7077 => x"34ff1554",
          7078 => x"7382f7dc",
          7079 => x"3482fbfc",
          7080 => x"08528851",
          7081 => x"ff96bf3f",
          7082 => x"82f7dc33",
          7083 => x"70982b70",
          7084 => x"982c82f7",
          7085 => x"d8335751",
          7086 => x"56577474",
          7087 => x"25ad3874",
          7088 => x"1a548114",
          7089 => x"33743482",
          7090 => x"fbfc0852",
          7091 => x"733351ff",
          7092 => x"96943f74",
          7093 => x"81800a29",
          7094 => x"81800a05",
          7095 => x"70982c82",
          7096 => x"f7d83358",
          7097 => x"51557575",
          7098 => x"24d53882",
          7099 => x"fbfc0852",
          7100 => x"a051ff95",
          7101 => x"f13f82f7",
          7102 => x"dc337098",
          7103 => x"2b70982c",
          7104 => x"82f7d833",
          7105 => x"57515657",
          7106 => x"747424fa",
          7107 => x"bf3882fb",
          7108 => x"fc085288",
          7109 => x"51ff95ce",
          7110 => x"3f748180",
          7111 => x"0a298180",
          7112 => x"0a057098",
          7113 => x"2c82f7d8",
          7114 => x"33585155",
          7115 => x"757525de",
          7116 => x"38fa9939",
          7117 => x"82f7d833",
          7118 => x"7a055480",
          7119 => x"743482fb",
          7120 => x"fc08528a",
          7121 => x"51ff959e",
          7122 => x"3f82f7d8",
          7123 => x"527951f6",
          7124 => x"c73f82e0",
          7125 => x"980881ff",
          7126 => x"06547396",
          7127 => x"3882f7d8",
          7128 => x"33547380",
          7129 => x"2e8f3881",
          7130 => x"53735279",
          7131 => x"51f1f13f",
          7132 => x"8439807a",
          7133 => x"34800b82",
          7134 => x"f7dc3480",
          7135 => x"0b82f7d8",
          7136 => x"347982e0",
          7137 => x"980caf3d",
          7138 => x"0d0482f7",
          7139 => x"dc335473",
          7140 => x"802ef9b8",
          7141 => x"3882fbfc",
          7142 => x"08528851",
          7143 => x"ff94c73f",
          7144 => x"82f7dc33",
          7145 => x"ff055473",
          7146 => x"82f7dc34",
          7147 => x"7381ff06",
          7148 => x"54dd3982",
          7149 => x"f7dc3382",
          7150 => x"f7d83355",
          7151 => x"5573752e",
          7152 => x"f98a38ff",
          7153 => x"14547382",
          7154 => x"f7d83474",
          7155 => x"982b7098",
          7156 => x"2c7581ff",
          7157 => x"06565155",
          7158 => x"747425ad",
          7159 => x"38741a54",
          7160 => x"81143374",
          7161 => x"3482fbfc",
          7162 => x"08527333",
          7163 => x"51ff93f6",
          7164 => x"3f748180",
          7165 => x"0a298180",
          7166 => x"0a057098",
          7167 => x"2c82f7d8",
          7168 => x"33585155",
          7169 => x"757524d5",
          7170 => x"3882fbfc",
          7171 => x"0852a051",
          7172 => x"ff93d33f",
          7173 => x"82f7dc33",
          7174 => x"70982b70",
          7175 => x"982c82f7",
          7176 => x"d8335751",
          7177 => x"56577474",
          7178 => x"24f8a138",
          7179 => x"82fbfc08",
          7180 => x"528851ff",
          7181 => x"93b03f74",
          7182 => x"81800a29",
          7183 => x"81800a05",
          7184 => x"70982c82",
          7185 => x"f7d83358",
          7186 => x"51557575",
          7187 => x"25de38f7",
          7188 => x"fb3982f7",
          7189 => x"dc337081",
          7190 => x"ff0682f7",
          7191 => x"d8335956",
          7192 => x"54747727",
          7193 => x"f7e63882",
          7194 => x"fbfc0852",
          7195 => x"81145473",
          7196 => x"82f7dc34",
          7197 => x"741a7033",
          7198 => x"5254ff92",
          7199 => x"e93f82f7",
          7200 => x"dc337081",
          7201 => x"ff0682f7",
          7202 => x"d8335856",
          7203 => x"54757526",
          7204 => x"d638f7b8",
          7205 => x"3982f7dc",
          7206 => x"53805282",
          7207 => x"c1b851ee",
          7208 => x"ee3f800b",
          7209 => x"82f7dc34",
          7210 => x"800b82f7",
          7211 => x"d834f79c",
          7212 => x"397ab038",
          7213 => x"82dfdc08",
          7214 => x"5574802e",
          7215 => x"a6387451",
          7216 => x"ff9af63f",
          7217 => x"82e09808",
          7218 => x"82f7d834",
          7219 => x"82e09808",
          7220 => x"81ff0681",
          7221 => x"05537452",
          7222 => x"7951ff9c",
          7223 => x"bc3f935b",
          7224 => x"81c0397a",
          7225 => x"842982df",
          7226 => x"9005fc11",
          7227 => x"08565474",
          7228 => x"802ea738",
          7229 => x"7451ff9a",
          7230 => x"c03f82e0",
          7231 => x"980882f7",
          7232 => x"d83482e0",
          7233 => x"980881ff",
          7234 => x"06810553",
          7235 => x"74527951",
          7236 => x"ff9c863f",
          7237 => x"ff1b5480",
          7238 => x"fa397308",
          7239 => x"5574802e",
          7240 => x"f6aa3874",
          7241 => x"51ff9a91",
          7242 => x"3f99397a",
          7243 => x"932e0981",
          7244 => x"06ae3882",
          7245 => x"df900855",
          7246 => x"74802ea4",
          7247 => x"387451ff",
          7248 => x"99f73f82",
          7249 => x"e0980882",
          7250 => x"f7d83482",
          7251 => x"e0980881",
          7252 => x"ff068105",
          7253 => x"53745279",
          7254 => x"51ff9bbd",
          7255 => x"3f80c339",
          7256 => x"7a842982",
          7257 => x"df940570",
          7258 => x"08565474",
          7259 => x"802eab38",
          7260 => x"7451ff99",
          7261 => x"c43f82e0",
          7262 => x"980882f7",
          7263 => x"d83482e0",
          7264 => x"980881ff",
          7265 => x"06810553",
          7266 => x"74527951",
          7267 => x"ff9b8a3f",
          7268 => x"811b5473",
          7269 => x"81ff065b",
          7270 => x"89397482",
          7271 => x"f7d83474",
          7272 => x"7a3482f7",
          7273 => x"dc5382f7",
          7274 => x"d8335279",
          7275 => x"51ece03f",
          7276 => x"f59a3982",
          7277 => x"f7dc3370",
          7278 => x"81ff0682",
          7279 => x"f7d83359",
          7280 => x"56547477",
          7281 => x"27f58538",
          7282 => x"82fbfc08",
          7283 => x"52811454",
          7284 => x"7382f7dc",
          7285 => x"34741a70",
          7286 => x"335254ff",
          7287 => x"90883ff4",
          7288 => x"eb3982f7",
          7289 => x"dc335473",
          7290 => x"802ef4e0",
          7291 => x"3882fbfc",
          7292 => x"08528851",
          7293 => x"ff8fef3f",
          7294 => x"82f7dc33",
          7295 => x"ff055473",
          7296 => x"82f7dc34",
          7297 => x"f4c639f9",
          7298 => x"3d0d84fa",
          7299 => x"f40b82e0",
          7300 => x"880ca080",
          7301 => x"0b82e084",
          7302 => x"23828080",
          7303 => x"53805284",
          7304 => x"faf451ff",
          7305 => x"a09f3f82",
          7306 => x"e0880854",
          7307 => x"80587774",
          7308 => x"34815776",
          7309 => x"81153482",
          7310 => x"e0880854",
          7311 => x"77841534",
          7312 => x"76851534",
          7313 => x"82e08808",
          7314 => x"54778615",
          7315 => x"34768715",
          7316 => x"3482e088",
          7317 => x"0882e084",
          7318 => x"22ff05fe",
          7319 => x"80800770",
          7320 => x"83ffff06",
          7321 => x"70882a58",
          7322 => x"51555674",
          7323 => x"88173473",
          7324 => x"89173482",
          7325 => x"e0842270",
          7326 => x"882982e0",
          7327 => x"880805f8",
          7328 => x"11515555",
          7329 => x"77821534",
          7330 => x"76831534",
          7331 => x"893d0d04",
          7332 => x"ff3d0d73",
          7333 => x"52815184",
          7334 => x"72278f38",
          7335 => x"fb12832a",
          7336 => x"82117083",
          7337 => x"ffff0651",
          7338 => x"51517082",
          7339 => x"e0980c83",
          7340 => x"3d0d04f9",
          7341 => x"3d0d02a6",
          7342 => x"05220284",
          7343 => x"05aa0522",
          7344 => x"710582e0",
          7345 => x"88087183",
          7346 => x"2b711174",
          7347 => x"832b7311",
          7348 => x"70338112",
          7349 => x"3371882b",
          7350 => x"0702a405",
          7351 => x"ae052271",
          7352 => x"81ffff06",
          7353 => x"0770882a",
          7354 => x"53515259",
          7355 => x"545b5b57",
          7356 => x"53545571",
          7357 => x"77347081",
          7358 => x"183482e0",
          7359 => x"88081475",
          7360 => x"882a5254",
          7361 => x"70821534",
          7362 => x"74831534",
          7363 => x"82e08808",
          7364 => x"70177033",
          7365 => x"81123371",
          7366 => x"882b0770",
          7367 => x"832b8fff",
          7368 => x"f8065152",
          7369 => x"56527105",
          7370 => x"7383ffff",
          7371 => x"0670882a",
          7372 => x"54545171",
          7373 => x"82123472",
          7374 => x"81ff0653",
          7375 => x"72831234",
          7376 => x"82e08808",
          7377 => x"16567176",
          7378 => x"34728117",
          7379 => x"34893d0d",
          7380 => x"04fb3d0d",
          7381 => x"82e08808",
          7382 => x"0284059e",
          7383 => x"05227083",
          7384 => x"2b721186",
          7385 => x"11338712",
          7386 => x"33718b2b",
          7387 => x"71832b07",
          7388 => x"585b5952",
          7389 => x"55527205",
          7390 => x"84123385",
          7391 => x"13337188",
          7392 => x"2b077088",
          7393 => x"2a545656",
          7394 => x"52708413",
          7395 => x"34738513",
          7396 => x"3482e088",
          7397 => x"08701484",
          7398 => x"11338512",
          7399 => x"33718b2b",
          7400 => x"71832b07",
          7401 => x"56595752",
          7402 => x"72058612",
          7403 => x"33871333",
          7404 => x"71882b07",
          7405 => x"70882a54",
          7406 => x"56565270",
          7407 => x"86133473",
          7408 => x"87133482",
          7409 => x"e0880813",
          7410 => x"70338112",
          7411 => x"3371882b",
          7412 => x"077081ff",
          7413 => x"ff067088",
          7414 => x"2a535153",
          7415 => x"53537173",
          7416 => x"34708114",
          7417 => x"34873d0d",
          7418 => x"04fa3d0d",
          7419 => x"02a20522",
          7420 => x"82e08808",
          7421 => x"71832b71",
          7422 => x"11703381",
          7423 => x"12337188",
          7424 => x"2b077088",
          7425 => x"29157033",
          7426 => x"81123371",
          7427 => x"982b7190",
          7428 => x"2b07535f",
          7429 => x"5355525a",
          7430 => x"56575354",
          7431 => x"71802580",
          7432 => x"f6387251",
          7433 => x"feab3f82",
          7434 => x"e0880870",
          7435 => x"16703381",
          7436 => x"1233718b",
          7437 => x"2b71832b",
          7438 => x"07741170",
          7439 => x"33811233",
          7440 => x"71882b07",
          7441 => x"70832b8f",
          7442 => x"fff80651",
          7443 => x"52545153",
          7444 => x"5a585372",
          7445 => x"0574882a",
          7446 => x"54527282",
          7447 => x"13347383",
          7448 => x"133482e0",
          7449 => x"88087016",
          7450 => x"70338112",
          7451 => x"33718b2b",
          7452 => x"71832b07",
          7453 => x"56595755",
          7454 => x"72057033",
          7455 => x"81123371",
          7456 => x"882b0770",
          7457 => x"81ffff06",
          7458 => x"70882a57",
          7459 => x"51525852",
          7460 => x"72743471",
          7461 => x"81153488",
          7462 => x"3d0d04fb",
          7463 => x"3d0d82e0",
          7464 => x"88080284",
          7465 => x"059e0522",
          7466 => x"70832b72",
          7467 => x"11821133",
          7468 => x"83123371",
          7469 => x"8b2b7183",
          7470 => x"2b07595b",
          7471 => x"59525652",
          7472 => x"73057133",
          7473 => x"81133371",
          7474 => x"882b0702",
          7475 => x"8c05a205",
          7476 => x"22710770",
          7477 => x"882a5351",
          7478 => x"53535371",
          7479 => x"73347081",
          7480 => x"143482e0",
          7481 => x"88087015",
          7482 => x"70338112",
          7483 => x"33718b2b",
          7484 => x"71832b07",
          7485 => x"56595752",
          7486 => x"72058212",
          7487 => x"33831333",
          7488 => x"71882b07",
          7489 => x"70882a54",
          7490 => x"55565270",
          7491 => x"82133472",
          7492 => x"83133482",
          7493 => x"e0880814",
          7494 => x"82113383",
          7495 => x"12337188",
          7496 => x"2b0782e0",
          7497 => x"980c5254",
          7498 => x"873d0d04",
          7499 => x"f73d0d7b",
          7500 => x"82e08808",
          7501 => x"31832a70",
          7502 => x"83ffff06",
          7503 => x"70535753",
          7504 => x"fda73f82",
          7505 => x"e0880876",
          7506 => x"832b7111",
          7507 => x"82113383",
          7508 => x"1233718b",
          7509 => x"2b71832b",
          7510 => x"07751170",
          7511 => x"33811233",
          7512 => x"71982b71",
          7513 => x"902b0753",
          7514 => x"42405153",
          7515 => x"5b585559",
          7516 => x"54728025",
          7517 => x"8d388280",
          7518 => x"80527551",
          7519 => x"fe9d3f81",
          7520 => x"84398414",
          7521 => x"33851533",
          7522 => x"718b2b71",
          7523 => x"832b0776",
          7524 => x"1179882a",
          7525 => x"53515558",
          7526 => x"55768614",
          7527 => x"347581ff",
          7528 => x"06567587",
          7529 => x"143482e0",
          7530 => x"88087019",
          7531 => x"84123385",
          7532 => x"13337188",
          7533 => x"2b077088",
          7534 => x"2a54575b",
          7535 => x"56537284",
          7536 => x"16347385",
          7537 => x"163482e0",
          7538 => x"88081853",
          7539 => x"800b8614",
          7540 => x"34800b87",
          7541 => x"143482e0",
          7542 => x"88085376",
          7543 => x"84143475",
          7544 => x"85143482",
          7545 => x"e0880818",
          7546 => x"70338112",
          7547 => x"3371882b",
          7548 => x"07708280",
          7549 => x"80077088",
          7550 => x"2a535155",
          7551 => x"56547474",
          7552 => x"34728115",
          7553 => x"348b3d0d",
          7554 => x"04ff3d0d",
          7555 => x"735282e0",
          7556 => x"88088438",
          7557 => x"f7f13f71",
          7558 => x"802e8638",
          7559 => x"7151fe8c",
          7560 => x"3f833d0d",
          7561 => x"04f53d0d",
          7562 => x"807e5258",
          7563 => x"f8e23f82",
          7564 => x"e0980883",
          7565 => x"ffff0682",
          7566 => x"e0880884",
          7567 => x"11338512",
          7568 => x"3371882b",
          7569 => x"07705f59",
          7570 => x"56585a81",
          7571 => x"ffff5975",
          7572 => x"782e80cb",
          7573 => x"38758829",
          7574 => x"17703381",
          7575 => x"12337188",
          7576 => x"2b077081",
          7577 => x"ffff0679",
          7578 => x"317083ff",
          7579 => x"ff06707f",
          7580 => x"27525351",
          7581 => x"56595577",
          7582 => x"79278a38",
          7583 => x"73802e85",
          7584 => x"3875785a",
          7585 => x"5b841533",
          7586 => x"85163371",
          7587 => x"882b0757",
          7588 => x"5475c238",
          7589 => x"7881ffff",
          7590 => x"2e85387a",
          7591 => x"79595680",
          7592 => x"76832b82",
          7593 => x"e0880811",
          7594 => x"70338112",
          7595 => x"3371882b",
          7596 => x"077081ff",
          7597 => x"ff065152",
          7598 => x"5a565c55",
          7599 => x"73752e83",
          7600 => x"38815580",
          7601 => x"54797826",
          7602 => x"81cc3874",
          7603 => x"5474802e",
          7604 => x"81c43877",
          7605 => x"7a2e0981",
          7606 => x"06893875",
          7607 => x"51f8f23f",
          7608 => x"81ac3982",
          7609 => x"80805379",
          7610 => x"527551f7",
          7611 => x"c63f82e0",
          7612 => x"8808701c",
          7613 => x"86113387",
          7614 => x"1233718b",
          7615 => x"2b71832b",
          7616 => x"07535a5e",
          7617 => x"5574057a",
          7618 => x"177083ff",
          7619 => x"ff067088",
          7620 => x"2a5c5956",
          7621 => x"54788415",
          7622 => x"347681ff",
          7623 => x"06577685",
          7624 => x"153482e0",
          7625 => x"88087583",
          7626 => x"2b711172",
          7627 => x"1e861133",
          7628 => x"87123371",
          7629 => x"882b0770",
          7630 => x"882a535b",
          7631 => x"5e535a56",
          7632 => x"54738619",
          7633 => x"34758719",
          7634 => x"3482e088",
          7635 => x"08701c84",
          7636 => x"11338512",
          7637 => x"33718b2b",
          7638 => x"71832b07",
          7639 => x"535d5a55",
          7640 => x"74055478",
          7641 => x"86153476",
          7642 => x"87153482",
          7643 => x"e0880870",
          7644 => x"16711d84",
          7645 => x"11338512",
          7646 => x"3371882b",
          7647 => x"0770882a",
          7648 => x"535a5f52",
          7649 => x"56547384",
          7650 => x"16347585",
          7651 => x"163482e0",
          7652 => x"88081b84",
          7653 => x"05547382",
          7654 => x"e0980c8d",
          7655 => x"3d0d04fe",
          7656 => x"3d0d7452",
          7657 => x"82e08808",
          7658 => x"8438f4db",
          7659 => x"3f715371",
          7660 => x"802e8b38",
          7661 => x"7151fced",
          7662 => x"3f82e098",
          7663 => x"08537282",
          7664 => x"e0980c84",
          7665 => x"3d0d04ee",
          7666 => x"3d0d6466",
          7667 => x"405c8070",
          7668 => x"424082e0",
          7669 => x"8808602e",
          7670 => x"09810684",
          7671 => x"38f4a83f",
          7672 => x"7b8e387e",
          7673 => x"51ffb83f",
          7674 => x"82e09808",
          7675 => x"5483c739",
          7676 => x"7e8b387b",
          7677 => x"51fc923f",
          7678 => x"7e5483ba",
          7679 => x"397e51f5",
          7680 => x"8f3f82e0",
          7681 => x"980883ff",
          7682 => x"ff0682e0",
          7683 => x"88087d71",
          7684 => x"31832a70",
          7685 => x"83ffff06",
          7686 => x"70832b73",
          7687 => x"11703381",
          7688 => x"12337188",
          7689 => x"2b077075",
          7690 => x"317083ff",
          7691 => x"ff067088",
          7692 => x"29fc0573",
          7693 => x"88291a70",
          7694 => x"33811233",
          7695 => x"71882b07",
          7696 => x"70902b53",
          7697 => x"444e5348",
          7698 => x"41525c54",
          7699 => x"5b415c56",
          7700 => x"5b5b7380",
          7701 => x"258f3876",
          7702 => x"81ffff06",
          7703 => x"75317083",
          7704 => x"ffff0642",
          7705 => x"54821633",
          7706 => x"83173371",
          7707 => x"882b0770",
          7708 => x"88291c70",
          7709 => x"33811233",
          7710 => x"71982b71",
          7711 => x"902b0753",
          7712 => x"47455256",
          7713 => x"54738025",
          7714 => x"8b387875",
          7715 => x"317083ff",
          7716 => x"ff064154",
          7717 => x"777b2781",
          7718 => x"fe386018",
          7719 => x"54737b2e",
          7720 => x"0981068f",
          7721 => x"387851f6",
          7722 => x"c03f7a83",
          7723 => x"ffff0658",
          7724 => x"81e5397f",
          7725 => x"8e387a74",
          7726 => x"24893878",
          7727 => x"51f6aa3f",
          7728 => x"81a5397f",
          7729 => x"18557a75",
          7730 => x"2480c838",
          7731 => x"791d8211",
          7732 => x"33831233",
          7733 => x"71882b07",
          7734 => x"535754f4",
          7735 => x"f43f8052",
          7736 => x"7851f7b7",
          7737 => x"3f82e098",
          7738 => x"0883ffff",
          7739 => x"067e547c",
          7740 => x"5370832b",
          7741 => x"82e08808",
          7742 => x"11840553",
          7743 => x"5559ff87",
          7744 => x"ce3f82e0",
          7745 => x"88081484",
          7746 => x"057583ff",
          7747 => x"ff06595c",
          7748 => x"81853960",
          7749 => x"15547a74",
          7750 => x"2480d438",
          7751 => x"7851f5c9",
          7752 => x"3f82e088",
          7753 => x"081d8211",
          7754 => x"33831233",
          7755 => x"71882b07",
          7756 => x"534354f4",
          7757 => x"9c3f8052",
          7758 => x"7851f6df",
          7759 => x"3f82e098",
          7760 => x"0883ffff",
          7761 => x"067e547c",
          7762 => x"5370832b",
          7763 => x"82e08808",
          7764 => x"11840553",
          7765 => x"5559ff86",
          7766 => x"f63f82e0",
          7767 => x"88081484",
          7768 => x"05606205",
          7769 => x"19555c73",
          7770 => x"83ffff06",
          7771 => x"58a9397b",
          7772 => x"7f5254f9",
          7773 => x"b03f82e0",
          7774 => x"98085c82",
          7775 => x"e0980880",
          7776 => x"2e93387d",
          7777 => x"53735282",
          7778 => x"e0980851",
          7779 => x"ff8b8a3f",
          7780 => x"7351f798",
          7781 => x"3f7a587a",
          7782 => x"78279938",
          7783 => x"80537a52",
          7784 => x"7851f28f",
          7785 => x"3f7a1983",
          7786 => x"2b82e088",
          7787 => x"08058405",
          7788 => x"51f6f93f",
          7789 => x"7b547382",
          7790 => x"e0980c94",
          7791 => x"3d0d04fc",
          7792 => x"3d0d7777",
          7793 => x"29705254",
          7794 => x"fbd53f82",
          7795 => x"e0980855",
          7796 => x"82e09808",
          7797 => x"802e8e38",
          7798 => x"73538052",
          7799 => x"82e09808",
          7800 => x"51ff90e1",
          7801 => x"3f7482e0",
          7802 => x"980c863d",
          7803 => x"0d04ff3d",
          7804 => x"0d028f05",
          7805 => x"33518152",
          7806 => x"70722687",
          7807 => x"3882e094",
          7808 => x"11335271",
          7809 => x"82e0980c",
          7810 => x"833d0d04",
          7811 => x"fc3d0d02",
          7812 => x"9b053302",
          7813 => x"84059f05",
          7814 => x"33565383",
          7815 => x"51728126",
          7816 => x"80e03872",
          7817 => x"842b87c0",
          7818 => x"928c1153",
          7819 => x"51885474",
          7820 => x"802e8438",
          7821 => x"81885473",
          7822 => x"720c87c0",
          7823 => x"928c1151",
          7824 => x"81710c85",
          7825 => x"0b87c098",
          7826 => x"8c0c7052",
          7827 => x"71087082",
          7828 => x"06515170",
          7829 => x"802e8a38",
          7830 => x"87c0988c",
          7831 => x"085170ec",
          7832 => x"387108fc",
          7833 => x"80800652",
          7834 => x"71923887",
          7835 => x"c0988c08",
          7836 => x"5170802e",
          7837 => x"87387182",
          7838 => x"e0941434",
          7839 => x"82e09413",
          7840 => x"33517082",
          7841 => x"e0980c86",
          7842 => x"3d0d04f3",
          7843 => x"3d0d6062",
          7844 => x"64028c05",
          7845 => x"bf053357",
          7846 => x"40585b83",
          7847 => x"74525afe",
          7848 => x"cd3f82e0",
          7849 => x"98088106",
          7850 => x"7a545271",
          7851 => x"81be3871",
          7852 => x"7275842b",
          7853 => x"87c09280",
          7854 => x"1187c092",
          7855 => x"8c1287c0",
          7856 => x"92841341",
          7857 => x"5a40575a",
          7858 => x"58850b87",
          7859 => x"c0988c0c",
          7860 => x"767d0c84",
          7861 => x"760c7508",
          7862 => x"70852a70",
          7863 => x"81065153",
          7864 => x"5471802e",
          7865 => x"8e387b08",
          7866 => x"52717b70",
          7867 => x"81055d34",
          7868 => x"81195980",
          7869 => x"74a20653",
          7870 => x"5371732e",
          7871 => x"83388153",
          7872 => x"7883ff26",
          7873 => x"8f387280",
          7874 => x"2e8a3887",
          7875 => x"c0988c08",
          7876 => x"5271c338",
          7877 => x"87c0988c",
          7878 => x"08527180",
          7879 => x"2e873878",
          7880 => x"84802e99",
          7881 => x"3881760c",
          7882 => x"87c0928c",
          7883 => x"15537208",
          7884 => x"70820651",
          7885 => x"5271f738",
          7886 => x"ff1a5a8d",
          7887 => x"39848017",
          7888 => x"81197081",
          7889 => x"ff065a53",
          7890 => x"5779802e",
          7891 => x"903873fc",
          7892 => x"80800652",
          7893 => x"7187387d",
          7894 => x"7826feed",
          7895 => x"3873fc80",
          7896 => x"80065271",
          7897 => x"802e8338",
          7898 => x"81527153",
          7899 => x"7282e098",
          7900 => x"0c8f3d0d",
          7901 => x"04f33d0d",
          7902 => x"60626402",
          7903 => x"8c05bf05",
          7904 => x"33574058",
          7905 => x"5b835980",
          7906 => x"745258fc",
          7907 => x"e13f82e0",
          7908 => x"98088106",
          7909 => x"79545271",
          7910 => x"782e0981",
          7911 => x"0681b138",
          7912 => x"7774842b",
          7913 => x"87c09280",
          7914 => x"1187c092",
          7915 => x"8c1287c0",
          7916 => x"92841340",
          7917 => x"595f565a",
          7918 => x"850b87c0",
          7919 => x"988c0c76",
          7920 => x"7d0c8276",
          7921 => x"0c805875",
          7922 => x"0870842a",
          7923 => x"70810651",
          7924 => x"53547180",
          7925 => x"2e8c387a",
          7926 => x"7081055c",
          7927 => x"337c0c81",
          7928 => x"18587381",
          7929 => x"2a708106",
          7930 => x"51527180",
          7931 => x"2e8a3887",
          7932 => x"c0988c08",
          7933 => x"5271d038",
          7934 => x"87c0988c",
          7935 => x"08527180",
          7936 => x"2e873877",
          7937 => x"84802e99",
          7938 => x"3881760c",
          7939 => x"87c0928c",
          7940 => x"15537208",
          7941 => x"70820651",
          7942 => x"5271f738",
          7943 => x"ff19598d",
          7944 => x"39811a70",
          7945 => x"81ff0684",
          7946 => x"8019595b",
          7947 => x"5278802e",
          7948 => x"903873fc",
          7949 => x"80800652",
          7950 => x"7187387d",
          7951 => x"7a26fef8",
          7952 => x"3873fc80",
          7953 => x"80065271",
          7954 => x"802e8338",
          7955 => x"81527153",
          7956 => x"7282e098",
          7957 => x"0c8f3d0d",
          7958 => x"04fa3d0d",
          7959 => x"7a028405",
          7960 => x"a3053302",
          7961 => x"8805a705",
          7962 => x"33715454",
          7963 => x"5657fafe",
          7964 => x"3f82e098",
          7965 => x"08810653",
          7966 => x"83547280",
          7967 => x"fe38850b",
          7968 => x"87c0988c",
          7969 => x"0c815671",
          7970 => x"762e80dc",
          7971 => x"38717624",
          7972 => x"93387484",
          7973 => x"2b87c092",
          7974 => x"8c115454",
          7975 => x"71802e8d",
          7976 => x"3880d439",
          7977 => x"71832e80",
          7978 => x"c63880cb",
          7979 => x"39720870",
          7980 => x"812a7081",
          7981 => x"06515152",
          7982 => x"71802e8a",
          7983 => x"3887c098",
          7984 => x"8c085271",
          7985 => x"e83887c0",
          7986 => x"988c0852",
          7987 => x"71963881",
          7988 => x"730c87c0",
          7989 => x"928c1453",
          7990 => x"72087082",
          7991 => x"06515271",
          7992 => x"f7389639",
          7993 => x"80569239",
          7994 => x"88800a77",
          7995 => x"0c853981",
          7996 => x"80770c72",
          7997 => x"56833984",
          7998 => x"56755473",
          7999 => x"82e0980c",
          8000 => x"883d0d04",
          8001 => x"fe3d0d74",
          8002 => x"81113371",
          8003 => x"3371882b",
          8004 => x"0782e098",
          8005 => x"0c535184",
          8006 => x"3d0d04fd",
          8007 => x"3d0d7583",
          8008 => x"11338212",
          8009 => x"3371902b",
          8010 => x"71882b07",
          8011 => x"81143370",
          8012 => x"7207882b",
          8013 => x"75337107",
          8014 => x"82e0980c",
          8015 => x"52535456",
          8016 => x"5452853d",
          8017 => x"0d04ff3d",
          8018 => x"0d730284",
          8019 => x"05920522",
          8020 => x"52527072",
          8021 => x"70810554",
          8022 => x"3470882a",
          8023 => x"51707234",
          8024 => x"833d0d04",
          8025 => x"ff3d0d73",
          8026 => x"75525270",
          8027 => x"72708105",
          8028 => x"54347088",
          8029 => x"2a517072",
          8030 => x"70810554",
          8031 => x"3470882a",
          8032 => x"51707270",
          8033 => x"81055434",
          8034 => x"70882a51",
          8035 => x"70723483",
          8036 => x"3d0d04fe",
          8037 => x"3d0d7675",
          8038 => x"77545451",
          8039 => x"70802e92",
          8040 => x"38717081",
          8041 => x"05533373",
          8042 => x"70810555",
          8043 => x"34ff1151",
          8044 => x"eb39843d",
          8045 => x"0d04fe3d",
          8046 => x"0d757776",
          8047 => x"54525372",
          8048 => x"72708105",
          8049 => x"5434ff11",
          8050 => x"5170f438",
          8051 => x"843d0d04",
          8052 => x"fc3d0d78",
          8053 => x"77795656",
          8054 => x"53747081",
          8055 => x"05563374",
          8056 => x"70810556",
          8057 => x"33717131",
          8058 => x"ff165652",
          8059 => x"52527280",
          8060 => x"2e863871",
          8061 => x"802ee238",
          8062 => x"7182e098",
          8063 => x"0c863d0d",
          8064 => x"04fe3d0d",
          8065 => x"74765451",
          8066 => x"89397173",
          8067 => x"2e8a3881",
          8068 => x"11517033",
          8069 => x"5271f338",
          8070 => x"703382e0",
          8071 => x"980c843d",
          8072 => x"0d04800b",
          8073 => x"82e0980c",
          8074 => x"04fb3d0d",
          8075 => x"77700870",
          8076 => x"70810552",
          8077 => x"33705455",
          8078 => x"5556e73f",
          8079 => x"ff5582e0",
          8080 => x"9808a238",
          8081 => x"72802e98",
          8082 => x"3883b552",
          8083 => x"725180f9",
          8084 => x"a23f82e0",
          8085 => x"980883ff",
          8086 => x"ff065372",
          8087 => x"802e8638",
          8088 => x"73760c72",
          8089 => x"557482e0",
          8090 => x"980c873d",
          8091 => x"0d04f73d",
          8092 => x"0d7b5680",
          8093 => x"0b831733",
          8094 => x"565a747a",
          8095 => x"2e80d638",
          8096 => x"8154b416",
          8097 => x"0853b816",
          8098 => x"70538117",
          8099 => x"335259f9",
          8100 => x"e43f82e0",
          8101 => x"98087a2e",
          8102 => x"098106b7",
          8103 => x"3882e098",
          8104 => x"08831734",
          8105 => x"b4160870",
          8106 => x"a8180831",
          8107 => x"a0180859",
          8108 => x"56587477",
          8109 => x"279f3882",
          8110 => x"16335574",
          8111 => x"822e0981",
          8112 => x"06933881",
          8113 => x"54761853",
          8114 => x"78528116",
          8115 => x"3351f9a5",
          8116 => x"3f833981",
          8117 => x"5a7982e0",
          8118 => x"980c8b3d",
          8119 => x"0d04fa3d",
          8120 => x"0d787a56",
          8121 => x"56805774",
          8122 => x"b417082e",
          8123 => x"af387551",
          8124 => x"fefc3f82",
          8125 => x"e0980857",
          8126 => x"82e09808",
          8127 => x"9f388154",
          8128 => x"7453b816",
          8129 => x"52811633",
          8130 => x"51f7803f",
          8131 => x"82e09808",
          8132 => x"802e8538",
          8133 => x"ff558157",
          8134 => x"74b4170c",
          8135 => x"7682e098",
          8136 => x"0c883d0d",
          8137 => x"04f83d0d",
          8138 => x"7a705257",
          8139 => x"fec03f82",
          8140 => x"e0980858",
          8141 => x"82e09808",
          8142 => x"81913876",
          8143 => x"33557483",
          8144 => x"2e098106",
          8145 => x"80f03884",
          8146 => x"17335978",
          8147 => x"812e0981",
          8148 => x"0680e338",
          8149 => x"84805382",
          8150 => x"e0980852",
          8151 => x"b8177052",
          8152 => x"56fcd33f",
          8153 => x"82d4d552",
          8154 => x"84b61751",
          8155 => x"fbd83f84",
          8156 => x"8b85a4d2",
          8157 => x"527551fb",
          8158 => x"eb3f868a",
          8159 => x"85e4f252",
          8160 => x"849c1751",
          8161 => x"fbde3f94",
          8162 => x"17085284",
          8163 => x"a01751fb",
          8164 => x"d33f9017",
          8165 => x"085284a4",
          8166 => x"1751fbc8",
          8167 => x"3fa41708",
          8168 => x"810570b4",
          8169 => x"190c7955",
          8170 => x"53755281",
          8171 => x"173351f7",
          8172 => x"c43f7784",
          8173 => x"18348053",
          8174 => x"80528117",
          8175 => x"3351f999",
          8176 => x"3f82e098",
          8177 => x"08802e83",
          8178 => x"38815877",
          8179 => x"82e0980c",
          8180 => x"8a3d0d04",
          8181 => x"fb3d0d77",
          8182 => x"fe1a9c12",
          8183 => x"08fe0555",
          8184 => x"56548056",
          8185 => x"7473278d",
          8186 => x"388a1422",
          8187 => x"757129b0",
          8188 => x"16080557",
          8189 => x"537582e0",
          8190 => x"980c873d",
          8191 => x"0d04f93d",
          8192 => x"0d7a7a70",
          8193 => x"08565457",
          8194 => x"81772781",
          8195 => x"df38769c",
          8196 => x"15082781",
          8197 => x"d738ff74",
          8198 => x"33545872",
          8199 => x"822e80f5",
          8200 => x"38728224",
          8201 => x"89387281",
          8202 => x"2e8d3881",
          8203 => x"bf397283",
          8204 => x"2e818e38",
          8205 => x"81b63976",
          8206 => x"812a1770",
          8207 => x"892aa816",
          8208 => x"08055374",
          8209 => x"5255fd96",
          8210 => x"3f82e098",
          8211 => x"08819f38",
          8212 => x"7483ff06",
          8213 => x"14b81133",
          8214 => x"81177089",
          8215 => x"2aa81808",
          8216 => x"05557654",
          8217 => x"575753fc",
          8218 => x"f53f82e0",
          8219 => x"980880fe",
          8220 => x"387483ff",
          8221 => x"0614b811",
          8222 => x"3370882b",
          8223 => x"78077981",
          8224 => x"0671842a",
          8225 => x"5c525851",
          8226 => x"537280e2",
          8227 => x"38759fff",
          8228 => x"065880da",
          8229 => x"3976882a",
          8230 => x"a8150805",
          8231 => x"527351fc",
          8232 => x"bd3f82e0",
          8233 => x"980880c6",
          8234 => x"38761083",
          8235 => x"fe067405",
          8236 => x"b80551f8",
          8237 => x"cf3f82e0",
          8238 => x"980883ff",
          8239 => x"ff0658ae",
          8240 => x"3976872a",
          8241 => x"a8150805",
          8242 => x"527351fc",
          8243 => x"913f82e0",
          8244 => x"98089b38",
          8245 => x"76822b83",
          8246 => x"fc067405",
          8247 => x"b80551f8",
          8248 => x"ba3f82e0",
          8249 => x"9808f00a",
          8250 => x"06588339",
          8251 => x"81587782",
          8252 => x"e0980c89",
          8253 => x"3d0d04f8",
          8254 => x"3d0d7a7c",
          8255 => x"7e5a5856",
          8256 => x"82598177",
          8257 => x"27829e38",
          8258 => x"769c1708",
          8259 => x"27829638",
          8260 => x"75335372",
          8261 => x"792e819d",
          8262 => x"38727924",
          8263 => x"89387281",
          8264 => x"2e8d3882",
          8265 => x"80397283",
          8266 => x"2e81b838",
          8267 => x"81f73976",
          8268 => x"812a1770",
          8269 => x"892aa818",
          8270 => x"08055376",
          8271 => x"5255fb9e",
          8272 => x"3f82e098",
          8273 => x"085982e0",
          8274 => x"980881d9",
          8275 => x"387483ff",
          8276 => x"0616b805",
          8277 => x"81167881",
          8278 => x"06595654",
          8279 => x"77537680",
          8280 => x"2e8f3877",
          8281 => x"842b9ff0",
          8282 => x"0674338f",
          8283 => x"06710751",
          8284 => x"53727434",
          8285 => x"810b8317",
          8286 => x"3474892a",
          8287 => x"a8170805",
          8288 => x"527551fa",
          8289 => x"d93f82e0",
          8290 => x"98085982",
          8291 => x"e0980881",
          8292 => x"94387483",
          8293 => x"ff0616b8",
          8294 => x"0578842a",
          8295 => x"5454768f",
          8296 => x"3877882a",
          8297 => x"743381f0",
          8298 => x"06718f06",
          8299 => x"07515372",
          8300 => x"743480ec",
          8301 => x"3976882a",
          8302 => x"a8170805",
          8303 => x"527551fa",
          8304 => x"9d3f82e0",
          8305 => x"98085982",
          8306 => x"e0980880",
          8307 => x"d8387783",
          8308 => x"ffff0652",
          8309 => x"761083fe",
          8310 => x"067605b8",
          8311 => x"0551f6e6",
          8312 => x"3fbe3976",
          8313 => x"872aa817",
          8314 => x"08055275",
          8315 => x"51f9ef3f",
          8316 => x"82e09808",
          8317 => x"5982e098",
          8318 => x"08ab3877",
          8319 => x"f00a0677",
          8320 => x"822b83fc",
          8321 => x"067018b8",
          8322 => x"05705451",
          8323 => x"5454f68b",
          8324 => x"3f82e098",
          8325 => x"088f0a06",
          8326 => x"74075272",
          8327 => x"51f6c53f",
          8328 => x"810b8317",
          8329 => x"347882e0",
          8330 => x"980c8a3d",
          8331 => x"0d04f83d",
          8332 => x"0d7a7c7e",
          8333 => x"72085956",
          8334 => x"56598175",
          8335 => x"27a43874",
          8336 => x"9c170827",
          8337 => x"9d387380",
          8338 => x"2eaa38ff",
          8339 => x"53735275",
          8340 => x"51fda43f",
          8341 => x"82e09808",
          8342 => x"5482e098",
          8343 => x"0880f238",
          8344 => x"93398254",
          8345 => x"80eb3981",
          8346 => x"5480e639",
          8347 => x"82e09808",
          8348 => x"5480de39",
          8349 => x"74527851",
          8350 => x"fb843f82",
          8351 => x"e0980858",
          8352 => x"82e09808",
          8353 => x"802e80c7",
          8354 => x"3882e098",
          8355 => x"08812ed2",
          8356 => x"3882e098",
          8357 => x"08ff2ecf",
          8358 => x"38805374",
          8359 => x"527551fc",
          8360 => x"d63f82e0",
          8361 => x"9808c538",
          8362 => x"9c1608fe",
          8363 => x"11941808",
          8364 => x"57555774",
          8365 => x"74279038",
          8366 => x"81159417",
          8367 => x"0c841633",
          8368 => x"81075473",
          8369 => x"84173477",
          8370 => x"55767826",
          8371 => x"ffa63880",
          8372 => x"547382e0",
          8373 => x"980c8a3d",
          8374 => x"0d04f63d",
          8375 => x"0d7c7e71",
          8376 => x"08595b5b",
          8377 => x"79953890",
          8378 => x"17085877",
          8379 => x"802e8838",
          8380 => x"9c170878",
          8381 => x"26b23881",
          8382 => x"58ae3979",
          8383 => x"527a51f9",
          8384 => x"fd3f8155",
          8385 => x"7482e098",
          8386 => x"082782e0",
          8387 => x"3882e098",
          8388 => x"085582e0",
          8389 => x"9808ff2e",
          8390 => x"82d2389c",
          8391 => x"170882e0",
          8392 => x"98082682",
          8393 => x"c7387958",
          8394 => x"94170870",
          8395 => x"56547380",
          8396 => x"2e82b938",
          8397 => x"777a2e09",
          8398 => x"810680e2",
          8399 => x"38811a56",
          8400 => x"9c170876",
          8401 => x"26833882",
          8402 => x"5675527a",
          8403 => x"51f9af3f",
          8404 => x"805982e0",
          8405 => x"9808812e",
          8406 => x"09810686",
          8407 => x"3882e098",
          8408 => x"085982e0",
          8409 => x"98080970",
          8410 => x"30707207",
          8411 => x"8025707c",
          8412 => x"0782e098",
          8413 => x"08545151",
          8414 => x"55557381",
          8415 => x"ef3882e0",
          8416 => x"9808802e",
          8417 => x"95389017",
          8418 => x"08548174",
          8419 => x"27903873",
          8420 => x"9c180827",
          8421 => x"89387358",
          8422 => x"85397580",
          8423 => x"db387756",
          8424 => x"8116569c",
          8425 => x"17087626",
          8426 => x"89388256",
          8427 => x"75782681",
          8428 => x"ac387552",
          8429 => x"7a51f8c6",
          8430 => x"3f82e098",
          8431 => x"08802eb8",
          8432 => x"38805982",
          8433 => x"e0980881",
          8434 => x"2e098106",
          8435 => x"863882e0",
          8436 => x"98085982",
          8437 => x"e0980809",
          8438 => x"70307072",
          8439 => x"07802570",
          8440 => x"7c075151",
          8441 => x"55557380",
          8442 => x"f8387578",
          8443 => x"2e098106",
          8444 => x"ffae3873",
          8445 => x"5580f539",
          8446 => x"ff537552",
          8447 => x"7651f9f7",
          8448 => x"3f82e098",
          8449 => x"0882e098",
          8450 => x"08307082",
          8451 => x"e0980807",
          8452 => x"80255155",
          8453 => x"5579802e",
          8454 => x"94387380",
          8455 => x"2e8f3875",
          8456 => x"53795276",
          8457 => x"51f9d03f",
          8458 => x"82e09808",
          8459 => x"5574a538",
          8460 => x"7590180c",
          8461 => x"9c1708fe",
          8462 => x"05941808",
          8463 => x"56547474",
          8464 => x"268638ff",
          8465 => x"1594180c",
          8466 => x"84173381",
          8467 => x"07547384",
          8468 => x"18349739",
          8469 => x"ff567481",
          8470 => x"2e90388c",
          8471 => x"3980558c",
          8472 => x"3982e098",
          8473 => x"08558539",
          8474 => x"81567555",
          8475 => x"7482e098",
          8476 => x"0c8c3d0d",
          8477 => x"04f83d0d",
          8478 => x"7a705255",
          8479 => x"f3f03f82",
          8480 => x"e0980858",
          8481 => x"815682e0",
          8482 => x"980880d8",
          8483 => x"387b5274",
          8484 => x"51f6c13f",
          8485 => x"82e09808",
          8486 => x"82e09808",
          8487 => x"b4170c59",
          8488 => x"84805377",
          8489 => x"52b81570",
          8490 => x"5257f28a",
          8491 => x"3f775684",
          8492 => x"39811656",
          8493 => x"8a152258",
          8494 => x"75782797",
          8495 => x"38815475",
          8496 => x"19537652",
          8497 => x"81153351",
          8498 => x"edab3f82",
          8499 => x"e0980880",
          8500 => x"2edf388a",
          8501 => x"15227632",
          8502 => x"70307072",
          8503 => x"07709f2a",
          8504 => x"53515656",
          8505 => x"7582e098",
          8506 => x"0c8a3d0d",
          8507 => x"04f83d0d",
          8508 => x"7a7c7108",
          8509 => x"58565774",
          8510 => x"f0800a26",
          8511 => x"80f13874",
          8512 => x"9f065372",
          8513 => x"80e93874",
          8514 => x"90180c88",
          8515 => x"17085473",
          8516 => x"aa387533",
          8517 => x"53827327",
          8518 => x"8838ac16",
          8519 => x"0854739b",
          8520 => x"3874852a",
          8521 => x"53820b88",
          8522 => x"17225a58",
          8523 => x"72792780",
          8524 => x"fe38ac16",
          8525 => x"0898180c",
          8526 => x"80cd398a",
          8527 => x"16227089",
          8528 => x"2b545872",
          8529 => x"7526b238",
          8530 => x"73527651",
          8531 => x"f5b03f82",
          8532 => x"e0980854",
          8533 => x"82e09808",
          8534 => x"ff2ebd38",
          8535 => x"810b82e0",
          8536 => x"9808278b",
          8537 => x"389c1608",
          8538 => x"82e09808",
          8539 => x"26853882",
          8540 => x"58bd3974",
          8541 => x"733155cb",
          8542 => x"39735275",
          8543 => x"51f4d53f",
          8544 => x"82e09808",
          8545 => x"98180c73",
          8546 => x"94180c98",
          8547 => x"17085382",
          8548 => x"5872802e",
          8549 => x"9a388539",
          8550 => x"81589439",
          8551 => x"74892a13",
          8552 => x"98180c74",
          8553 => x"83ff0616",
          8554 => x"b8059c18",
          8555 => x"0c805877",
          8556 => x"82e0980c",
          8557 => x"8a3d0d04",
          8558 => x"f83d0d7a",
          8559 => x"70089012",
          8560 => x"08a00559",
          8561 => x"5754f080",
          8562 => x"0a772786",
          8563 => x"38800b98",
          8564 => x"150c9814",
          8565 => x"08538455",
          8566 => x"72802e81",
          8567 => x"cb387683",
          8568 => x"ff065877",
          8569 => x"81b53881",
          8570 => x"1398150c",
          8571 => x"94140855",
          8572 => x"74923876",
          8573 => x"852a8817",
          8574 => x"22565374",
          8575 => x"7326819b",
          8576 => x"3880c039",
          8577 => x"8a1622ff",
          8578 => x"0577892a",
          8579 => x"06537281",
          8580 => x"8a387452",
          8581 => x"7351f3e6",
          8582 => x"3f82e098",
          8583 => x"08538255",
          8584 => x"810b82e0",
          8585 => x"98082780",
          8586 => x"ff388155",
          8587 => x"82e09808",
          8588 => x"ff2e80f4",
          8589 => x"389c1608",
          8590 => x"82e09808",
          8591 => x"2680ca38",
          8592 => x"7b8a3877",
          8593 => x"98150c84",
          8594 => x"5580dd39",
          8595 => x"94140852",
          8596 => x"7351f986",
          8597 => x"3f82e098",
          8598 => x"08538755",
          8599 => x"82e09808",
          8600 => x"802e80c4",
          8601 => x"38825582",
          8602 => x"e0980881",
          8603 => x"2eba3881",
          8604 => x"5582e098",
          8605 => x"08ff2eb0",
          8606 => x"3882e098",
          8607 => x"08527551",
          8608 => x"fbf33f82",
          8609 => x"e09808a0",
          8610 => x"38729415",
          8611 => x"0c725275",
          8612 => x"51f2c13f",
          8613 => x"82e09808",
          8614 => x"98150c76",
          8615 => x"90150c77",
          8616 => x"16b8059c",
          8617 => x"150c8055",
          8618 => x"7482e098",
          8619 => x"0c8a3d0d",
          8620 => x"04f73d0d",
          8621 => x"7b7d7108",
          8622 => x"5b5b5780",
          8623 => x"527651fc",
          8624 => x"ac3f82e0",
          8625 => x"98085482",
          8626 => x"e0980880",
          8627 => x"ec3882e0",
          8628 => x"98085698",
          8629 => x"17085278",
          8630 => x"51f0833f",
          8631 => x"82e09808",
          8632 => x"5482e098",
          8633 => x"0880d238",
          8634 => x"82e09808",
          8635 => x"9c180870",
          8636 => x"33515458",
          8637 => x"7281e52e",
          8638 => x"09810683",
          8639 => x"38815882",
          8640 => x"e0980855",
          8641 => x"72833881",
          8642 => x"55777507",
          8643 => x"5372802e",
          8644 => x"8e388116",
          8645 => x"56757a2e",
          8646 => x"09810688",
          8647 => x"38a53982",
          8648 => x"e0980856",
          8649 => x"81527651",
          8650 => x"fd8e3f82",
          8651 => x"e0980854",
          8652 => x"82e09808",
          8653 => x"802eff9b",
          8654 => x"3873842e",
          8655 => x"09810683",
          8656 => x"38875473",
          8657 => x"82e0980c",
          8658 => x"8b3d0d04",
          8659 => x"fd3d0d76",
          8660 => x"9a115254",
          8661 => x"ebae3f82",
          8662 => x"e0980883",
          8663 => x"ffff0676",
          8664 => x"70335153",
          8665 => x"5371832e",
          8666 => x"09810690",
          8667 => x"38941451",
          8668 => x"eb923f82",
          8669 => x"e0980890",
          8670 => x"2b730753",
          8671 => x"7282e098",
          8672 => x"0c853d0d",
          8673 => x"04fc3d0d",
          8674 => x"77797083",
          8675 => x"ffff0654",
          8676 => x"9a125355",
          8677 => x"55ebaf3f",
          8678 => x"76703351",
          8679 => x"5372832e",
          8680 => x"0981068b",
          8681 => x"3873902a",
          8682 => x"52941551",
          8683 => x"eb983f86",
          8684 => x"3d0d04fd",
          8685 => x"3d0d7554",
          8686 => x"80518b53",
          8687 => x"70812a71",
          8688 => x"81802905",
          8689 => x"74708105",
          8690 => x"56337105",
          8691 => x"7081ff06",
          8692 => x"ff165651",
          8693 => x"515172e4",
          8694 => x"387082e0",
          8695 => x"980c853d",
          8696 => x"0d04f23d",
          8697 => x"0d606240",
          8698 => x"59847908",
          8699 => x"5f5b81ff",
          8700 => x"705d5d98",
          8701 => x"1908802e",
          8702 => x"83803898",
          8703 => x"1908527d",
          8704 => x"51eddb3f",
          8705 => x"82e09808",
          8706 => x"5b82e098",
          8707 => x"0882eb38",
          8708 => x"9c190870",
          8709 => x"33555573",
          8710 => x"8638845b",
          8711 => x"82dc398b",
          8712 => x"1533bf06",
          8713 => x"7081ff06",
          8714 => x"58537286",
          8715 => x"1a3482e0",
          8716 => x"98085673",
          8717 => x"81e52e09",
          8718 => x"81068338",
          8719 => x"815682e0",
          8720 => x"98085373",
          8721 => x"ae2e0981",
          8722 => x"06833881",
          8723 => x"53757307",
          8724 => x"53729938",
          8725 => x"82e09808",
          8726 => x"77df0654",
          8727 => x"5672882e",
          8728 => x"09810683",
          8729 => x"38815675",
          8730 => x"7f2e8738",
          8731 => x"81ff5c81",
          8732 => x"ef39768f",
          8733 => x"2e098106",
          8734 => x"81ca3873",
          8735 => x"862a7081",
          8736 => x"06515372",
          8737 => x"802e9238",
          8738 => x"8d153374",
          8739 => x"81bf0670",
          8740 => x"901c08ac",
          8741 => x"1d0c565d",
          8742 => x"5d737c2e",
          8743 => x"09810681",
          8744 => x"9c388d15",
          8745 => x"33537c73",
          8746 => x"2e098106",
          8747 => x"818f388c",
          8748 => x"1e089a16",
          8749 => x"525ae8cc",
          8750 => x"3f82e098",
          8751 => x"0883ffff",
          8752 => x"06537280",
          8753 => x"f8387433",
          8754 => x"7081bf06",
          8755 => x"8d29f305",
          8756 => x"5154817b",
          8757 => x"585882d2",
          8758 => x"a8173375",
          8759 => x"0551e8a4",
          8760 => x"3f82e098",
          8761 => x"0883ffff",
          8762 => x"06567780",
          8763 => x"2e963873",
          8764 => x"81fe2680",
          8765 => x"c8387310",
          8766 => x"1a765953",
          8767 => x"75732381",
          8768 => x"14548b39",
          8769 => x"7583ffff",
          8770 => x"2e098106",
          8771 => x"b0388117",
          8772 => x"578c7727",
          8773 => x"c1387433",
          8774 => x"70862a70",
          8775 => x"81065154",
          8776 => x"5572802e",
          8777 => x"8e387381",
          8778 => x"fe269238",
          8779 => x"73101a53",
          8780 => x"807323ff",
          8781 => x"1c7081ff",
          8782 => x"06515384",
          8783 => x"3981ff53",
          8784 => x"725c9d39",
          8785 => x"7b933874",
          8786 => x"51fce83f",
          8787 => x"82e09808",
          8788 => x"81ff0653",
          8789 => x"727d2ea7",
          8790 => x"38ff0bac",
          8791 => x"1a0ca039",
          8792 => x"80527851",
          8793 => x"f8d23f82",
          8794 => x"e098085b",
          8795 => x"82e09808",
          8796 => x"89389819",
          8797 => x"08fd8438",
          8798 => x"8639800b",
          8799 => x"981a0c7a",
          8800 => x"82e0980c",
          8801 => x"903d0d04",
          8802 => x"f23d0d60",
          8803 => x"70084059",
          8804 => x"80527851",
          8805 => x"f6d73f82",
          8806 => x"e0980858",
          8807 => x"82e09808",
          8808 => x"83a43881",
          8809 => x"ff705f5c",
          8810 => x"ff0bac1a",
          8811 => x"0c981908",
          8812 => x"527e51ea",
          8813 => x"a93f82e0",
          8814 => x"98085882",
          8815 => x"e0980883",
          8816 => x"85389c19",
          8817 => x"08703357",
          8818 => x"57758638",
          8819 => x"845882f6",
          8820 => x"398b1733",
          8821 => x"bf067081",
          8822 => x"ff065654",
          8823 => x"73861a34",
          8824 => x"7581e52e",
          8825 => x"82c33874",
          8826 => x"832a7081",
          8827 => x"06515474",
          8828 => x"8f2e8e38",
          8829 => x"7382b238",
          8830 => x"748f2e09",
          8831 => x"810681f7",
          8832 => x"38ab1933",
          8833 => x"70862a70",
          8834 => x"81065155",
          8835 => x"557382a1",
          8836 => x"3875862a",
          8837 => x"70810651",
          8838 => x"5473802e",
          8839 => x"92388d17",
          8840 => x"337681bf",
          8841 => x"0670901c",
          8842 => x"08ac1d0c",
          8843 => x"585d5e75",
          8844 => x"7c2e0981",
          8845 => x"0681b938",
          8846 => x"8d173356",
          8847 => x"7d762e09",
          8848 => x"810681ac",
          8849 => x"388c1f08",
          8850 => x"9a18525d",
          8851 => x"e5b63f82",
          8852 => x"e0980883",
          8853 => x"ffff0655",
          8854 => x"74819538",
          8855 => x"763370bf",
          8856 => x"068d29f3",
          8857 => x"05595681",
          8858 => x"755c5a82",
          8859 => x"d2a81b33",
          8860 => x"770551e5",
          8861 => x"8f3f82e0",
          8862 => x"980883ff",
          8863 => x"ff065679",
          8864 => x"802eb138",
          8865 => x"7781fe26",
          8866 => x"80e63875",
          8867 => x"5180e1a0",
          8868 => x"3f82e098",
          8869 => x"0878101e",
          8870 => x"70225355",
          8871 => x"81195955",
          8872 => x"80e18d3f",
          8873 => x"7482e098",
          8874 => x"082e0981",
          8875 => x"0680c138",
          8876 => x"755a8b39",
          8877 => x"7583ffff",
          8878 => x"2e098106",
          8879 => x"b338811b",
          8880 => x"5b8c7b27",
          8881 => x"ffa53876",
          8882 => x"3370862a",
          8883 => x"70810651",
          8884 => x"55577980",
          8885 => x"2e903873",
          8886 => x"802e8b38",
          8887 => x"77101d70",
          8888 => x"22515473",
          8889 => x"8b38ff1c",
          8890 => x"7081ff06",
          8891 => x"51548439",
          8892 => x"81ff5473",
          8893 => x"5cbb397b",
          8894 => x"93387651",
          8895 => x"f9b53f82",
          8896 => x"e0980881",
          8897 => x"ff065473",
          8898 => x"7e2ebb38",
          8899 => x"ab193381",
          8900 => x"06547395",
          8901 => x"388b53a0",
          8902 => x"19529c19",
          8903 => x"0851e5b0",
          8904 => x"3f82e098",
          8905 => x"08802e9e",
          8906 => x"3881ff5c",
          8907 => x"ff0bac1a",
          8908 => x"0c805278",
          8909 => x"51f5813f",
          8910 => x"82e09808",
          8911 => x"5882e098",
          8912 => x"08802efc",
          8913 => x"e8387782",
          8914 => x"e0980c90",
          8915 => x"3d0d04ee",
          8916 => x"3d0d6470",
          8917 => x"08ab1233",
          8918 => x"81a00656",
          8919 => x"5d5a8655",
          8920 => x"7385b538",
          8921 => x"738c1d08",
          8922 => x"70225656",
          8923 => x"5d73802e",
          8924 => x"8d38811d",
          8925 => x"70101670",
          8926 => x"2251555d",
          8927 => x"f0398c53",
          8928 => x"a01a7053",
          8929 => x"923d7053",
          8930 => x"5f59e487",
          8931 => x"3f0280cb",
          8932 => x"05338106",
          8933 => x"5473802e",
          8934 => x"82a83880",
          8935 => x"c00bab1b",
          8936 => x"34815b8c",
          8937 => x"1c087b56",
          8938 => x"588b537d",
          8939 => x"527851e3",
          8940 => x"e23f857b",
          8941 => x"2780c638",
          8942 => x"7a567722",
          8943 => x"7083ffff",
          8944 => x"06555573",
          8945 => x"802eb438",
          8946 => x"7483ffff",
          8947 => x"06821959",
          8948 => x"558f5774",
          8949 => x"81067610",
          8950 => x"0775812a",
          8951 => x"71902a70",
          8952 => x"81065156",
          8953 => x"56567380",
          8954 => x"2e873875",
          8955 => x"84a0a132",
          8956 => x"56ff1757",
          8957 => x"768025db",
          8958 => x"38c03975",
          8959 => x"55870284",
          8960 => x"05bf0557",
          8961 => x"5774b007",
          8962 => x"bf0654b9",
          8963 => x"74278438",
          8964 => x"87145473",
          8965 => x"7634ff16",
          8966 => x"ff187684",
          8967 => x"2a575856",
          8968 => x"74e33894",
          8969 => x"3dec0517",
          8970 => x"5480fe74",
          8971 => x"34807727",
          8972 => x"b5387833",
          8973 => x"5473a02e",
          8974 => x"ad387419",
          8975 => x"70335254",
          8976 => x"e3e03f82",
          8977 => x"e0980880",
          8978 => x"2e8c38ff",
          8979 => x"17547474",
          8980 => x"2e943881",
          8981 => x"15558115",
          8982 => x"55747727",
          8983 => x"89387419",
          8984 => x"70335154",
          8985 => x"d039943d",
          8986 => x"7705eb05",
          8987 => x"54781581",
          8988 => x"165658a0",
          8989 => x"56768726",
          8990 => x"8a388117",
          8991 => x"81157033",
          8992 => x"58555775",
          8993 => x"78348775",
          8994 => x"27e33879",
          8995 => x"51f9f93f",
          8996 => x"82e09808",
          8997 => x"8b38811b",
          8998 => x"5b80e37b",
          8999 => x"27fe8438",
          9000 => x"87557a80",
          9001 => x"e42e82f0",
          9002 => x"3882e098",
          9003 => x"085582e0",
          9004 => x"9808842e",
          9005 => x"09810682",
          9006 => x"df380280",
          9007 => x"cb0533ab",
          9008 => x"1b340280",
          9009 => x"cb053370",
          9010 => x"812a7081",
          9011 => x"0651555e",
          9012 => x"81597380",
          9013 => x"2e90388d",
          9014 => x"528c1d51",
          9015 => x"feebf43f",
          9016 => x"82e09808",
          9017 => x"19597852",
          9018 => x"7951f3c5",
          9019 => x"3f82e098",
          9020 => x"085782e0",
          9021 => x"9808829e",
          9022 => x"38ff1959",
          9023 => x"78802e81",
          9024 => x"d4387885",
          9025 => x"2b901b08",
          9026 => x"71315354",
          9027 => x"7951efdd",
          9028 => x"3f82e098",
          9029 => x"085782e0",
          9030 => x"980881fa",
          9031 => x"38a01a51",
          9032 => x"f5913f82",
          9033 => x"e0980881",
          9034 => x"ff065d98",
          9035 => x"1a08527b",
          9036 => x"51e3ab3f",
          9037 => x"82e09808",
          9038 => x"5782e098",
          9039 => x"0881d738",
          9040 => x"8c1c089c",
          9041 => x"1b087a81",
          9042 => x"ff065a57",
          9043 => x"5b7c8d17",
          9044 => x"348f0b8b",
          9045 => x"173482e0",
          9046 => x"98088c17",
          9047 => x"3482e098",
          9048 => x"08529a16",
          9049 => x"51dfdf3f",
          9050 => x"778d29f3",
          9051 => x"05775555",
          9052 => x"7383ffff",
          9053 => x"2e8b3874",
          9054 => x"101b7022",
          9055 => x"81175751",
          9056 => x"54735282",
          9057 => x"d2a81733",
          9058 => x"760551df",
          9059 => x"b93f7385",
          9060 => x"3883ffff",
          9061 => x"54811757",
          9062 => x"8c7727d4",
          9063 => x"387383ff",
          9064 => x"ff2e8b38",
          9065 => x"74101b70",
          9066 => x"22515473",
          9067 => x"86387780",
          9068 => x"c0075877",
          9069 => x"7634810b",
          9070 => x"831d3480",
          9071 => x"527951ef",
          9072 => x"f73f82e0",
          9073 => x"98085782",
          9074 => x"e0980880",
          9075 => x"c938ff19",
          9076 => x"5978fed7",
          9077 => x"38981a08",
          9078 => x"527b51e2",
          9079 => x"813f82e0",
          9080 => x"98085782",
          9081 => x"e09808ae",
          9082 => x"38a05382",
          9083 => x"e0980852",
          9084 => x"9c1a0851",
          9085 => x"dfc03f8b",
          9086 => x"53a01a52",
          9087 => x"9c1a0851",
          9088 => x"df913f9c",
          9089 => x"1a08ab1b",
          9090 => x"33980655",
          9091 => x"55738c16",
          9092 => x"34810b83",
          9093 => x"1d347655",
          9094 => x"7482e098",
          9095 => x"0c943d0d",
          9096 => x"04fa3d0d",
          9097 => x"78700890",
          9098 => x"1208ac13",
          9099 => x"08565957",
          9100 => x"5572ff2e",
          9101 => x"94387252",
          9102 => x"7451edb1",
          9103 => x"3f82e098",
          9104 => x"085482e0",
          9105 => x"980880c9",
          9106 => x"38981508",
          9107 => x"527551e1",
          9108 => x"8d3f82e0",
          9109 => x"98085482",
          9110 => x"e09808ab",
          9111 => x"389c1508",
          9112 => x"53e57334",
          9113 => x"810b8317",
          9114 => x"34901508",
          9115 => x"7727a238",
          9116 => x"82e09808",
          9117 => x"527451ee",
          9118 => x"bf3f82e0",
          9119 => x"98085482",
          9120 => x"e0980880",
          9121 => x"2ec33873",
          9122 => x"842e0981",
          9123 => x"06833882",
          9124 => x"547382e0",
          9125 => x"980c883d",
          9126 => x"0d04f43d",
          9127 => x"0d7e6071",
          9128 => x"085f595c",
          9129 => x"800b9619",
          9130 => x"34981c08",
          9131 => x"802e83e2",
          9132 => x"38ac1c08",
          9133 => x"ff2e81bb",
          9134 => x"38807071",
          9135 => x"7f8c0508",
          9136 => x"70225757",
          9137 => x"5b5c5772",
          9138 => x"772e819d",
          9139 => x"38781014",
          9140 => x"7022811b",
          9141 => x"5b56537a",
          9142 => x"973880d0",
          9143 => x"80157083",
          9144 => x"ffff0651",
          9145 => x"53728fff",
          9146 => x"26863874",
          9147 => x"5b80df39",
          9148 => x"76189611",
          9149 => x"81ff7931",
          9150 => x"585b5483",
          9151 => x"b5527a90",
          9152 => x"2b750751",
          9153 => x"80d7843f",
          9154 => x"82e09808",
          9155 => x"83ffff06",
          9156 => x"5581ff75",
          9157 => x"27953881",
          9158 => x"7627a538",
          9159 => x"74882a53",
          9160 => x"727a3474",
          9161 => x"97153482",
          9162 => x"559f3974",
          9163 => x"30763070",
          9164 => x"78078025",
          9165 => x"72802507",
          9166 => x"52545473",
          9167 => x"802e8538",
          9168 => x"80579a39",
          9169 => x"747a3481",
          9170 => x"55741757",
          9171 => x"805b8c1d",
          9172 => x"08791011",
          9173 => x"70225154",
          9174 => x"5472fef1",
          9175 => x"387a3070",
          9176 => x"80257030",
          9177 => x"79065951",
          9178 => x"53771794",
          9179 => x"0553800b",
          9180 => x"82143480",
          9181 => x"70891a58",
          9182 => x"5a579c1c",
          9183 => x"08197033",
          9184 => x"811b5b56",
          9185 => x"5374a02e",
          9186 => x"b7387485",
          9187 => x"2e098106",
          9188 => x"843881e5",
          9189 => x"55788932",
          9190 => x"70307072",
          9191 => x"07802551",
          9192 => x"5454768b",
          9193 => x"26903872",
          9194 => x"802e8b38",
          9195 => x"ae767081",
          9196 => x"05583481",
          9197 => x"17577476",
          9198 => x"70810558",
          9199 => x"34811757",
          9200 => x"8a7927ff",
          9201 => x"b5387717",
          9202 => x"88055380",
          9203 => x"0b811434",
          9204 => x"96183353",
          9205 => x"72818738",
          9206 => x"768b38bf",
          9207 => x"0b961934",
          9208 => x"815780e1",
          9209 => x"39727389",
          9210 => x"1a33555a",
          9211 => x"5772802e",
          9212 => x"80d33896",
          9213 => x"18891955",
          9214 => x"567333ff",
          9215 => x"bf115455",
          9216 => x"729926aa",
          9217 => x"389c1c08",
          9218 => x"8c113351",
          9219 => x"53887927",
          9220 => x"87387284",
          9221 => x"2a538539",
          9222 => x"72832a53",
          9223 => x"72810653",
          9224 => x"72802e8a",
          9225 => x"38a01570",
          9226 => x"83ffff06",
          9227 => x"56537476",
          9228 => x"70810558",
          9229 => x"34811981",
          9230 => x"15811971",
          9231 => x"33565955",
          9232 => x"5972ffb5",
          9233 => x"38771794",
          9234 => x"0553800b",
          9235 => x"8214349c",
          9236 => x"1c088c11",
          9237 => x"33515372",
          9238 => x"85387289",
          9239 => x"19349c1c",
          9240 => x"08538b13",
          9241 => x"33881934",
          9242 => x"9c1c089c",
          9243 => x"115253d9",
          9244 => x"aa3f82e0",
          9245 => x"9808780c",
          9246 => x"961351d9",
          9247 => x"873f82e0",
          9248 => x"98088619",
          9249 => x"23981351",
          9250 => x"d8fa3f82",
          9251 => x"e0980884",
          9252 => x"19238e3d",
          9253 => x"0d04f03d",
          9254 => x"0d627008",
          9255 => x"415e8064",
          9256 => x"70335155",
          9257 => x"5573af2e",
          9258 => x"83388155",
          9259 => x"7380dc2e",
          9260 => x"92387480",
          9261 => x"2e8d387f",
          9262 => x"98050888",
          9263 => x"1f0caa39",
          9264 => x"81154480",
          9265 => x"64703356",
          9266 => x"565673af",
          9267 => x"2e098106",
          9268 => x"83388156",
          9269 => x"7380dc32",
          9270 => x"70307080",
          9271 => x"25780751",
          9272 => x"515473dc",
          9273 => x"3873881f",
          9274 => x"0c637033",
          9275 => x"5154739f",
          9276 => x"269638ff",
          9277 => x"800bab1f",
          9278 => x"3480527d",
          9279 => x"51e7ee3f",
          9280 => x"82e09808",
          9281 => x"5687e139",
          9282 => x"63417d08",
          9283 => x"8c11085b",
          9284 => x"54805992",
          9285 => x"3dfc0551",
          9286 => x"da8f3f82",
          9287 => x"e09808ff",
          9288 => x"2e82b138",
          9289 => x"83ffff0b",
          9290 => x"82e09808",
          9291 => x"27923878",
          9292 => x"101a82e0",
          9293 => x"9808902a",
          9294 => x"55557375",
          9295 => x"23811959",
          9296 => x"82e09808",
          9297 => x"83ffff06",
          9298 => x"70af3270",
          9299 => x"309f7327",
          9300 => x"71802507",
          9301 => x"51515556",
          9302 => x"73b43875",
          9303 => x"80dc2eae",
          9304 => x"387580ff",
          9305 => x"26913875",
          9306 => x"5282d1c4",
          9307 => x"51d9923f",
          9308 => x"82e09808",
          9309 => x"81de3878",
          9310 => x"81fe2681",
          9311 => x"d7387810",
          9312 => x"1a547574",
          9313 => x"23811959",
          9314 => x"ff893981",
          9315 => x"15418061",
          9316 => x"70335656",
          9317 => x"5773af2e",
          9318 => x"09810683",
          9319 => x"38815773",
          9320 => x"80dc3270",
          9321 => x"30708025",
          9322 => x"79075151",
          9323 => x"5473dc38",
          9324 => x"74449f76",
          9325 => x"27822b57",
          9326 => x"78812e09",
          9327 => x"81068c38",
          9328 => x"79225473",
          9329 => x"ae2ea538",
          9330 => x"80d23978",
          9331 => x"822e0981",
          9332 => x"0680c938",
          9333 => x"821a2254",
          9334 => x"73ae2e09",
          9335 => x"810680c1",
          9336 => x"38792254",
          9337 => x"73ae2e09",
          9338 => x"8106b638",
          9339 => x"78101a54",
          9340 => x"80742380",
          9341 => x"0ba01f56",
          9342 => x"58ae5478",
          9343 => x"78268338",
          9344 => x"a0547375",
          9345 => x"70810557",
          9346 => x"34811858",
          9347 => x"8a7827e9",
          9348 => x"3876a007",
          9349 => x"5473ab1f",
          9350 => x"3484c439",
          9351 => x"78802ea8",
          9352 => x"3878101a",
          9353 => x"fe055574",
          9354 => x"22fe1671",
          9355 => x"72a03270",
          9356 => x"30709f2a",
          9357 => x"51515358",
          9358 => x"565475ae",
          9359 => x"2e843873",
          9360 => x"8738ff19",
          9361 => x"5978e038",
          9362 => x"78197a11",
          9363 => x"55568074",
          9364 => x"23788d38",
          9365 => x"86568590",
          9366 => x"39768307",
          9367 => x"57839939",
          9368 => x"807a2270",
          9369 => x"83ffff06",
          9370 => x"56565d73",
          9371 => x"a02e0981",
          9372 => x"06933881",
          9373 => x"1d70101b",
          9374 => x"70225155",
          9375 => x"5d73a02e",
          9376 => x"f2387c8f",
          9377 => x"387483ff",
          9378 => x"ff065473",
          9379 => x"ae2e0981",
          9380 => x"06853876",
          9381 => x"83075778",
          9382 => x"802eaa38",
          9383 => x"7916fe05",
          9384 => x"70225154",
          9385 => x"73ae2e9d",
          9386 => x"3878101a",
          9387 => x"fe0555ff",
          9388 => x"19597880",
          9389 => x"2e8f38fe",
          9390 => x"15702255",
          9391 => x"5573ae2e",
          9392 => x"098106eb",
          9393 => x"388b53a0",
          9394 => x"52a01e51",
          9395 => x"d5e83f80",
          9396 => x"70595c88",
          9397 => x"5f7c101a",
          9398 => x"7022811f",
          9399 => x"5f575475",
          9400 => x"802e8294",
          9401 => x"3875a02e",
          9402 => x"963875ae",
          9403 => x"32703070",
          9404 => x"80255151",
          9405 => x"547c792e",
          9406 => x"8c387380",
          9407 => x"2e893876",
          9408 => x"830757d1",
          9409 => x"39805473",
          9410 => x"5b7e7826",
          9411 => x"8338815b",
          9412 => x"7c793270",
          9413 => x"30707207",
          9414 => x"8025707e",
          9415 => x"07515155",
          9416 => x"5573802e",
          9417 => x"a6387e8b",
          9418 => x"2efeae38",
          9419 => x"7c792e8b",
          9420 => x"38768307",
          9421 => x"577c7926",
          9422 => x"81be3878",
          9423 => x"5d88588b",
          9424 => x"7c822b81",
          9425 => x"fc065d5f",
          9426 => x"ff8b3980",
          9427 => x"ff7627af",
          9428 => x"38768207",
          9429 => x"5783b552",
          9430 => x"755180ce",
          9431 => x"ae3f82e0",
          9432 => x"980883ff",
          9433 => x"ff067087",
          9434 => x"2a708106",
          9435 => x"51555673",
          9436 => x"802e8c38",
          9437 => x"7580ff06",
          9438 => x"82d2b811",
          9439 => x"33575481",
          9440 => x"ff7627a4",
          9441 => x"38ff1f54",
          9442 => x"7378268a",
          9443 => x"38768307",
          9444 => x"7f5957fe",
          9445 => x"c0397d18",
          9446 => x"a0057688",
          9447 => x"2a555573",
          9448 => x"75348118",
          9449 => x"5880c339",
          9450 => x"75802e92",
          9451 => x"38755282",
          9452 => x"d1d051d4",
          9453 => x"cc3f82e0",
          9454 => x"9808802e",
          9455 => x"8a3880df",
          9456 => x"77830758",
          9457 => x"56a439ff",
          9458 => x"bf165473",
          9459 => x"99268538",
          9460 => x"7b82075c",
          9461 => x"ff9f1654",
          9462 => x"7399268e",
          9463 => x"387b8107",
          9464 => x"e0177083",
          9465 => x"ffff0658",
          9466 => x"555c7d18",
          9467 => x"a0055475",
          9468 => x"74348118",
          9469 => x"58fdde39",
          9470 => x"a01e3354",
          9471 => x"7381e52e",
          9472 => x"09810686",
          9473 => x"38850ba0",
          9474 => x"1f347e88",
          9475 => x"2e098106",
          9476 => x"88387b82",
          9477 => x"2b81fc06",
          9478 => x"5c7b8c06",
          9479 => x"54738c2e",
          9480 => x"8d387b83",
          9481 => x"06547383",
          9482 => x"2e098106",
          9483 => x"85387682",
          9484 => x"07577681",
          9485 => x"2a708106",
          9486 => x"5154739f",
          9487 => x"387b8106",
          9488 => x"5473802e",
          9489 => x"85387690",
          9490 => x"07577b82",
          9491 => x"2a708106",
          9492 => x"51547380",
          9493 => x"2e853876",
          9494 => x"88075776",
          9495 => x"ab1f347d",
          9496 => x"51eaa53f",
          9497 => x"82e09808",
          9498 => x"ab1f3356",
          9499 => x"5682e098",
          9500 => x"08802ebe",
          9501 => x"3882e098",
          9502 => x"08842e09",
          9503 => x"810680e8",
          9504 => x"3874852a",
          9505 => x"70810676",
          9506 => x"822a5751",
          9507 => x"5473802e",
          9508 => x"96387481",
          9509 => x"06547380",
          9510 => x"2ef8ed38",
          9511 => x"ff800bab",
          9512 => x"1f348056",
          9513 => x"80c23974",
          9514 => x"81065473",
          9515 => x"bb388556",
          9516 => x"b7397482",
          9517 => x"2a708106",
          9518 => x"515473ac",
          9519 => x"38861e33",
          9520 => x"70842a70",
          9521 => x"81065155",
          9522 => x"5573802e",
          9523 => x"e138901e",
          9524 => x"0883ff06",
          9525 => x"6005b805",
          9526 => x"527f51e4",
          9527 => x"ef3f82e0",
          9528 => x"9808881f",
          9529 => x"0cf8a139",
          9530 => x"7582e098",
          9531 => x"0c923d0d",
          9532 => x"04f63d0d",
          9533 => x"7c5bff7b",
          9534 => x"08707173",
          9535 => x"55595c55",
          9536 => x"5973802e",
          9537 => x"81c63875",
          9538 => x"70810557",
          9539 => x"33709f26",
          9540 => x"525271ba",
          9541 => x"2e8d3870",
          9542 => x"ee3871ba",
          9543 => x"2e098106",
          9544 => x"81a53873",
          9545 => x"33d01170",
          9546 => x"81ff0651",
          9547 => x"52537089",
          9548 => x"26913882",
          9549 => x"147381ff",
          9550 => x"06d00556",
          9551 => x"5271762e",
          9552 => x"80f73880",
          9553 => x"0b82d298",
          9554 => x"59557708",
          9555 => x"7a555776",
          9556 => x"70810558",
          9557 => x"33747081",
          9558 => x"055633ff",
          9559 => x"9f125353",
          9560 => x"53709926",
          9561 => x"8938e013",
          9562 => x"7081ff06",
          9563 => x"5451ff9f",
          9564 => x"12517099",
          9565 => x"268938e0",
          9566 => x"127081ff",
          9567 => x"06535172",
          9568 => x"30709f2a",
          9569 => x"51517272",
          9570 => x"2e098106",
          9571 => x"853870ff",
          9572 => x"be387230",
          9573 => x"74773270",
          9574 => x"30707207",
          9575 => x"9f2a739f",
          9576 => x"2a075354",
          9577 => x"54517080",
          9578 => x"2e8f3881",
          9579 => x"15841959",
          9580 => x"55837525",
          9581 => x"ff94388b",
          9582 => x"39748324",
          9583 => x"86387476",
          9584 => x"7c0c5978",
          9585 => x"51863982",
          9586 => x"f7f43351",
          9587 => x"7082e098",
          9588 => x"0c8c3d0d",
          9589 => x"04fa3d0d",
          9590 => x"7856800b",
          9591 => x"831734ff",
          9592 => x"0bb4170c",
          9593 => x"79527551",
          9594 => x"d1f43f84",
          9595 => x"5582e098",
          9596 => x"08818038",
          9597 => x"84b61651",
          9598 => x"ce8a3f82",
          9599 => x"e0980883",
          9600 => x"ffff0654",
          9601 => x"83557382",
          9602 => x"d4d52e09",
          9603 => x"810680e3",
          9604 => x"38800bb8",
          9605 => x"17335657",
          9606 => x"7481e92e",
          9607 => x"09810683",
          9608 => x"38815774",
          9609 => x"81eb3270",
          9610 => x"30708025",
          9611 => x"79075151",
          9612 => x"54738a38",
          9613 => x"7481e82e",
          9614 => x"098106b5",
          9615 => x"38835382",
          9616 => x"d1d85280",
          9617 => x"ee1651cf",
          9618 => x"873f82e0",
          9619 => x"98085582",
          9620 => x"e0980880",
          9621 => x"2e9d3885",
          9622 => x"5382d1dc",
          9623 => x"52818a16",
          9624 => x"51ceed3f",
          9625 => x"82e09808",
          9626 => x"5582e098",
          9627 => x"08802e83",
          9628 => x"38825574",
          9629 => x"82e0980c",
          9630 => x"883d0d04",
          9631 => x"f23d0d61",
          9632 => x"02840580",
          9633 => x"cb053358",
          9634 => x"5580750c",
          9635 => x"6051fce1",
          9636 => x"3f82e098",
          9637 => x"08588b56",
          9638 => x"800b82e0",
          9639 => x"98082487",
          9640 => x"c73882e0",
          9641 => x"98088429",
          9642 => x"82f7e005",
          9643 => x"70085553",
          9644 => x"8c567380",
          9645 => x"2e87b138",
          9646 => x"73750c76",
          9647 => x"81fe0674",
          9648 => x"33545772",
          9649 => x"802eae38",
          9650 => x"81143351",
          9651 => x"c6a03f82",
          9652 => x"e0980881",
          9653 => x"ff067081",
          9654 => x"06545572",
          9655 => x"98387680",
          9656 => x"2e878338",
          9657 => x"74822a70",
          9658 => x"81065153",
          9659 => x"8a567286",
          9660 => x"f73886f2",
          9661 => x"39807434",
          9662 => x"77185982",
          9663 => x"e08c1933",
          9664 => x"81153481",
          9665 => x"52811433",
          9666 => x"51c6813f",
          9667 => x"82e09808",
          9668 => x"81ff0670",
          9669 => x"81065455",
          9670 => x"83567286",
          9671 => x"cb387680",
          9672 => x"2e8f3874",
          9673 => x"822a7081",
          9674 => x"0651538a",
          9675 => x"567286b8",
          9676 => x"38807053",
          9677 => x"74525bfd",
          9678 => x"9c3f82e0",
          9679 => x"980881ff",
          9680 => x"06577682",
          9681 => x"2e933876",
          9682 => x"8126819c",
          9683 => x"3882e08d",
          9684 => x"19335372",
          9685 => x"7b2e8190",
          9686 => x"388c3d74",
          9687 => x"56598356",
          9688 => x"83fa1533",
          9689 => x"70585372",
          9690 => x"802e8d38",
          9691 => x"83fe1551",
          9692 => x"cba93f82",
          9693 => x"e0980857",
          9694 => x"76797084",
          9695 => x"055b0cff",
          9696 => x"16901656",
          9697 => x"56758025",
          9698 => x"d7387718",
          9699 => x"82e08d11",
          9700 => x"33703070",
          9701 => x"9f2a7271",
          9702 => x"31953d71",
          9703 => x"842905f0",
          9704 => x"055a5351",
          9705 => x"55575974",
          9706 => x"085b8357",
          9707 => x"7a802e90",
          9708 => x"387a5273",
          9709 => x"51fc9e3f",
          9710 => x"82e09808",
          9711 => x"81ff0657",
          9712 => x"800b82e0",
          9713 => x"8d1a3354",
          9714 => x"5872782e",
          9715 => x"09810683",
          9716 => x"38815881",
          9717 => x"77279138",
          9718 => x"77802e8c",
          9719 => x"38811684",
          9720 => x"16565683",
          9721 => x"7627c038",
          9722 => x"81567684",
          9723 => x"2e84f938",
          9724 => x"8d567681",
          9725 => x"2684f138",
          9726 => x"80c31451",
          9727 => x"ca863f82",
          9728 => x"e0980883",
          9729 => x"ffff0653",
          9730 => x"7284802e",
          9731 => x"09810684",
          9732 => x"d73880ce",
          9733 => x"1451c9ec",
          9734 => x"3f82e098",
          9735 => x"0883ffff",
          9736 => x"0658778d",
          9737 => x"3880dc14",
          9738 => x"51c9f03f",
          9739 => x"82e09808",
          9740 => x"5877a015",
          9741 => x"0c80c814",
          9742 => x"33821534",
          9743 => x"80c81433",
          9744 => x"ff117081",
          9745 => x"ff065154",
          9746 => x"558d5672",
          9747 => x"81268498",
          9748 => x"387481ff",
          9749 => x"06787129",
          9750 => x"80c51633",
          9751 => x"52595372",
          9752 => x"8a152372",
          9753 => x"802e8b38",
          9754 => x"ff137306",
          9755 => x"5372802e",
          9756 => x"86388d56",
          9757 => x"83f23980",
          9758 => x"c91451c9",
          9759 => x"873f82e0",
          9760 => x"98085382",
          9761 => x"e0980888",
          9762 => x"1523728f",
          9763 => x"06578d56",
          9764 => x"7683d538",
          9765 => x"80cb1451",
          9766 => x"c8ea3f82",
          9767 => x"e0980883",
          9768 => x"ffff0655",
          9769 => x"748d3880",
          9770 => x"d81451c8",
          9771 => x"ee3f82e0",
          9772 => x"98085580",
          9773 => x"c61451c8",
          9774 => x"cb3f82e0",
          9775 => x"980883ff",
          9776 => x"ff06538d",
          9777 => x"5672802e",
          9778 => x"839e3888",
          9779 => x"14227814",
          9780 => x"71842a05",
          9781 => x"5a5a7875",
          9782 => x"26838d38",
          9783 => x"8a142252",
          9784 => x"74793151",
          9785 => x"fed3ec3f",
          9786 => x"82e09808",
          9787 => x"5582e098",
          9788 => x"08802e82",
          9789 => x"f33882e0",
          9790 => x"980880ff",
          9791 => x"fffff526",
          9792 => x"83388357",
          9793 => x"7483fff5",
          9794 => x"26833882",
          9795 => x"57749ff5",
          9796 => x"26853881",
          9797 => x"5789398d",
          9798 => x"5676802e",
          9799 => x"82ca3882",
          9800 => x"15709c16",
          9801 => x"0c7ba416",
          9802 => x"0c731c70",
          9803 => x"a8170c7a",
          9804 => x"1db0170c",
          9805 => x"54557683",
          9806 => x"2e098106",
          9807 => x"af3880e2",
          9808 => x"1451c7c0",
          9809 => x"3f82e098",
          9810 => x"0883ffff",
          9811 => x"06538d56",
          9812 => x"72829538",
          9813 => x"79829138",
          9814 => x"80e41451",
          9815 => x"c7bd3f82",
          9816 => x"e09808ac",
          9817 => x"150c7482",
          9818 => x"2b53a239",
          9819 => x"8d567980",
          9820 => x"2e81f538",
          9821 => x"7713ac15",
          9822 => x"0c741553",
          9823 => x"76822e8d",
          9824 => x"38741015",
          9825 => x"70812a76",
          9826 => x"81060551",
          9827 => x"5383ff13",
          9828 => x"892a538d",
          9829 => x"5672a015",
          9830 => x"082681cc",
          9831 => x"38ff0b94",
          9832 => x"150cff0b",
          9833 => x"90150cff",
          9834 => x"800b8415",
          9835 => x"3476832e",
          9836 => x"09810681",
          9837 => x"923880e8",
          9838 => x"1451c6c8",
          9839 => x"3f82e098",
          9840 => x"0883ffff",
          9841 => x"06537281",
          9842 => x"2e098106",
          9843 => x"80f93881",
          9844 => x"1b527351",
          9845 => x"ca883f82",
          9846 => x"e0980880",
          9847 => x"ea3882e0",
          9848 => x"98088415",
          9849 => x"3484b614",
          9850 => x"51c6993f",
          9851 => x"82e09808",
          9852 => x"83ffff06",
          9853 => x"537282d4",
          9854 => x"d52e0981",
          9855 => x"0680c838",
          9856 => x"b81451c6",
          9857 => x"963f82e0",
          9858 => x"9808848b",
          9859 => x"85a4d22e",
          9860 => x"098106b3",
          9861 => x"38849c14",
          9862 => x"51c6803f",
          9863 => x"82e09808",
          9864 => x"868a85e4",
          9865 => x"f22e0981",
          9866 => x"069d3884",
          9867 => x"a01451c5",
          9868 => x"ea3f82e0",
          9869 => x"98089415",
          9870 => x"0c84a414",
          9871 => x"51c5dc3f",
          9872 => x"82e09808",
          9873 => x"90150c76",
          9874 => x"743482f7",
          9875 => x"f0228105",
          9876 => x"537282f7",
          9877 => x"f0237286",
          9878 => x"152382f7",
          9879 => x"f80b8c15",
          9880 => x"0c800b98",
          9881 => x"150c8056",
          9882 => x"7582e098",
          9883 => x"0c903d0d",
          9884 => x"04fb3d0d",
          9885 => x"77548955",
          9886 => x"73802eba",
          9887 => x"38730853",
          9888 => x"72802eb2",
          9889 => x"38723352",
          9890 => x"71802eaa",
          9891 => x"38861322",
          9892 => x"84152257",
          9893 => x"5271762e",
          9894 => x"0981069a",
          9895 => x"38811333",
          9896 => x"51ffbeca",
          9897 => x"3f82e098",
          9898 => x"08810652",
          9899 => x"71883871",
          9900 => x"74085455",
          9901 => x"83398053",
          9902 => x"7873710c",
          9903 => x"527482e0",
          9904 => x"980c873d",
          9905 => x"0d04fa3d",
          9906 => x"0d02ab05",
          9907 => x"337a5889",
          9908 => x"3dfc0552",
          9909 => x"56f49a3f",
          9910 => x"8b54800b",
          9911 => x"82e09808",
          9912 => x"24bc3882",
          9913 => x"e0980884",
          9914 => x"2982f7e0",
          9915 => x"05700855",
          9916 => x"5573802e",
          9917 => x"84388074",
          9918 => x"34785473",
          9919 => x"802e8438",
          9920 => x"80743478",
          9921 => x"750c7554",
          9922 => x"75802e92",
          9923 => x"38805389",
          9924 => x"3d705384",
          9925 => x"0551f6e4",
          9926 => x"3f82e098",
          9927 => x"08547382",
          9928 => x"e0980c88",
          9929 => x"3d0d04ea",
          9930 => x"3d0d6802",
          9931 => x"840580eb",
          9932 => x"05335959",
          9933 => x"89547880",
          9934 => x"2e84c838",
          9935 => x"77bf0670",
          9936 => x"54993dcc",
          9937 => x"05539a3d",
          9938 => x"84055258",
          9939 => x"f6ae3f82",
          9940 => x"e0980855",
          9941 => x"82e09808",
          9942 => x"84a4387a",
          9943 => x"5c69528c",
          9944 => x"3d705256",
          9945 => x"eab03f82",
          9946 => x"e0980855",
          9947 => x"82e09808",
          9948 => x"92380280",
          9949 => x"d7053370",
          9950 => x"982b5557",
          9951 => x"73802583",
          9952 => x"38865577",
          9953 => x"9c065473",
          9954 => x"802e81ab",
          9955 => x"3874802e",
          9956 => x"95387484",
          9957 => x"2e098106",
          9958 => x"aa387551",
          9959 => x"dfb13f82",
          9960 => x"e0980855",
          9961 => x"9e3902b2",
          9962 => x"05339106",
          9963 => x"547381b8",
          9964 => x"3877822a",
          9965 => x"70810651",
          9966 => x"5473802e",
          9967 => x"8e388855",
          9968 => x"83bc3977",
          9969 => x"88075874",
          9970 => x"83b43877",
          9971 => x"832a7081",
          9972 => x"06515473",
          9973 => x"802e81af",
          9974 => x"3862527a",
          9975 => x"51d6ed3f",
          9976 => x"82e09808",
          9977 => x"568288b2",
          9978 => x"0a52628e",
          9979 => x"0551c2f4",
          9980 => x"3f6254a0",
          9981 => x"0b8b1534",
          9982 => x"80536252",
          9983 => x"7a51d785",
          9984 => x"3f805262",
          9985 => x"9c0551c2",
          9986 => x"db3f7a54",
          9987 => x"810b8315",
          9988 => x"3475802e",
          9989 => x"80f1387a",
          9990 => x"b4110851",
          9991 => x"54805375",
          9992 => x"52983dd0",
          9993 => x"0551cc86",
          9994 => x"3f82e098",
          9995 => x"085582e0",
          9996 => x"980882ca",
          9997 => x"38b73974",
          9998 => x"82c43802",
          9999 => x"b2053370",
         10000 => x"842a7081",
         10001 => x"06515556",
         10002 => x"73802e86",
         10003 => x"38845582",
         10004 => x"ad397781",
         10005 => x"2a708106",
         10006 => x"51547380",
         10007 => x"2ea93875",
         10008 => x"81065473",
         10009 => x"802ea038",
         10010 => x"87558292",
         10011 => x"3973527a",
         10012 => x"51c4eb3f",
         10013 => x"82e09808",
         10014 => x"7bff1890",
         10015 => x"120c5555",
         10016 => x"82e09808",
         10017 => x"81f83877",
         10018 => x"832a7081",
         10019 => x"06515473",
         10020 => x"802e8638",
         10021 => x"7780c007",
         10022 => x"587ab411",
         10023 => x"08a01b0c",
         10024 => x"63a41b0c",
         10025 => x"63537052",
         10026 => x"57d5a13f",
         10027 => x"82e09808",
         10028 => x"82e09808",
         10029 => x"881b0c63",
         10030 => x"9c05525a",
         10031 => x"c0dd3f82",
         10032 => x"e0980882",
         10033 => x"e098088c",
         10034 => x"1b0c777a",
         10035 => x"0c568617",
         10036 => x"22841a23",
         10037 => x"77901a34",
         10038 => x"800b911a",
         10039 => x"34800b9c",
         10040 => x"1a0c800b",
         10041 => x"941a0c77",
         10042 => x"852a7081",
         10043 => x"06515473",
         10044 => x"802e818d",
         10045 => x"3882e098",
         10046 => x"08802e81",
         10047 => x"843882e0",
         10048 => x"9808941a",
         10049 => x"0c8a1722",
         10050 => x"70892b7b",
         10051 => x"525957a8",
         10052 => x"39765278",
         10053 => x"51c5e73f",
         10054 => x"82e09808",
         10055 => x"5782e098",
         10056 => x"08812683",
         10057 => x"38825582",
         10058 => x"e09808ff",
         10059 => x"2e098106",
         10060 => x"83387955",
         10061 => x"75783156",
         10062 => x"74307076",
         10063 => x"07802551",
         10064 => x"54777627",
         10065 => x"8a388170",
         10066 => x"7506555a",
         10067 => x"73c33876",
         10068 => x"981a0c74",
         10069 => x"a9387583",
         10070 => x"ff065473",
         10071 => x"802ea238",
         10072 => x"76527a51",
         10073 => x"c4ee3f82",
         10074 => x"e0980885",
         10075 => x"3882558e",
         10076 => x"3975892a",
         10077 => x"82e09808",
         10078 => x"059c1a0c",
         10079 => x"84398079",
         10080 => x"0c745473",
         10081 => x"82e0980c",
         10082 => x"983d0d04",
         10083 => x"f23d0d60",
         10084 => x"63656440",
         10085 => x"405d5980",
         10086 => x"7e0c903d",
         10087 => x"fc055278",
         10088 => x"51f9ce3f",
         10089 => x"82e09808",
         10090 => x"5582e098",
         10091 => x"088a3891",
         10092 => x"19335574",
         10093 => x"802e8638",
         10094 => x"745682c7",
         10095 => x"39901933",
         10096 => x"81065587",
         10097 => x"5674802e",
         10098 => x"82b93895",
         10099 => x"39820b91",
         10100 => x"1a348256",
         10101 => x"82ad3981",
         10102 => x"0b911a34",
         10103 => x"815682a3",
         10104 => x"398c1908",
         10105 => x"941a0831",
         10106 => x"55747c27",
         10107 => x"8338745c",
         10108 => x"7b802e82",
         10109 => x"8c389419",
         10110 => x"087083ff",
         10111 => x"06565674",
         10112 => x"81b4387e",
         10113 => x"8a1122ff",
         10114 => x"0577892a",
         10115 => x"065b5579",
         10116 => x"a8387587",
         10117 => x"38881908",
         10118 => x"558f3998",
         10119 => x"19085278",
         10120 => x"51c3db3f",
         10121 => x"82e09808",
         10122 => x"55817527",
         10123 => x"ff9f3874",
         10124 => x"ff2effa3",
         10125 => x"3874981a",
         10126 => x"0c981908",
         10127 => x"527e51c3",
         10128 => x"933f82e0",
         10129 => x"9808802e",
         10130 => x"ff833882",
         10131 => x"e098081a",
         10132 => x"7c892a59",
         10133 => x"5777802e",
         10134 => x"80d83877",
         10135 => x"1a7f8a11",
         10136 => x"22585c55",
         10137 => x"75752785",
         10138 => x"38757a31",
         10139 => x"58775476",
         10140 => x"537c5281",
         10141 => x"1b3351ff",
         10142 => x"b8913f82",
         10143 => x"e09808fe",
         10144 => x"d6387e83",
         10145 => x"11335656",
         10146 => x"74802ea0",
         10147 => x"38b41608",
         10148 => x"77315574",
         10149 => x"78279538",
         10150 => x"848053b8",
         10151 => x"1652b416",
         10152 => x"08773189",
         10153 => x"2b7d0551",
         10154 => x"ffbde83f",
         10155 => x"77892b56",
         10156 => x"ba39769c",
         10157 => x"1a0c9419",
         10158 => x"0883ff06",
         10159 => x"84807131",
         10160 => x"57557b76",
         10161 => x"2783387b",
         10162 => x"569c1908",
         10163 => x"527e51c0",
         10164 => x"8d3f82e0",
         10165 => x"9808fdff",
         10166 => x"38755394",
         10167 => x"190883ff",
         10168 => x"061fb805",
         10169 => x"527c51ff",
         10170 => x"bda93f7b",
         10171 => x"76317e08",
         10172 => x"177f0c76",
         10173 => x"1e941b08",
         10174 => x"18941c0c",
         10175 => x"5e5cfdf0",
         10176 => x"39805675",
         10177 => x"82e0980c",
         10178 => x"903d0d04",
         10179 => x"f23d0d60",
         10180 => x"63656440",
         10181 => x"405d5880",
         10182 => x"7e0c903d",
         10183 => x"fc055277",
         10184 => x"51f6ce3f",
         10185 => x"82e09808",
         10186 => x"5582e098",
         10187 => x"088a3891",
         10188 => x"18335574",
         10189 => x"802e8638",
         10190 => x"745683bf",
         10191 => x"39901833",
         10192 => x"70812a70",
         10193 => x"81065156",
         10194 => x"56875674",
         10195 => x"802e83ab",
         10196 => x"38953982",
         10197 => x"0b911934",
         10198 => x"8256839f",
         10199 => x"39810b91",
         10200 => x"19348156",
         10201 => x"83953994",
         10202 => x"18087c11",
         10203 => x"56567476",
         10204 => x"27843875",
         10205 => x"095c7b80",
         10206 => x"2e82f338",
         10207 => x"94180870",
         10208 => x"83ff0656",
         10209 => x"56748282",
         10210 => x"387e8a11",
         10211 => x"22ff0577",
         10212 => x"892a065c",
         10213 => x"557abf38",
         10214 => x"758c3888",
         10215 => x"18085574",
         10216 => x"9c387a52",
         10217 => x"85399818",
         10218 => x"08527751",
         10219 => x"c6ac3f82",
         10220 => x"e0980855",
         10221 => x"82e09808",
         10222 => x"802e82b2",
         10223 => x"3874812e",
         10224 => x"ff913874",
         10225 => x"ff2eff95",
         10226 => x"38749819",
         10227 => x"0c881808",
         10228 => x"85387488",
         10229 => x"190c7e55",
         10230 => x"b415089c",
         10231 => x"19082e09",
         10232 => x"81068e38",
         10233 => x"7451ffbd",
         10234 => x"853f82e0",
         10235 => x"9808feed",
         10236 => x"38981808",
         10237 => x"527e51ff",
         10238 => x"bfda3f82",
         10239 => x"e0980880",
         10240 => x"2efed038",
         10241 => x"82e09808",
         10242 => x"1b7c892a",
         10243 => x"5a577880",
         10244 => x"2e80d738",
         10245 => x"781b7f8a",
         10246 => x"1122585b",
         10247 => x"55757527",
         10248 => x"8538757b",
         10249 => x"31597854",
         10250 => x"76537c52",
         10251 => x"811a3351",
         10252 => x"ffb6c23f",
         10253 => x"82e09808",
         10254 => x"fea3387e",
         10255 => x"b4110878",
         10256 => x"31565674",
         10257 => x"79279c38",
         10258 => x"848053b4",
         10259 => x"16087731",
         10260 => x"892b7d05",
         10261 => x"52b81651",
         10262 => x"ffbab83f",
         10263 => x"7e55800b",
         10264 => x"83163478",
         10265 => x"892b5680",
         10266 => x"de398c18",
         10267 => x"08941908",
         10268 => x"2694387e",
         10269 => x"51ffbbf6",
         10270 => x"3f82e098",
         10271 => x"08fdde38",
         10272 => x"7e77b412",
         10273 => x"0c55769c",
         10274 => x"190c9418",
         10275 => x"0883ff06",
         10276 => x"84807131",
         10277 => x"57557b76",
         10278 => x"2783387b",
         10279 => x"569c1808",
         10280 => x"527e51ff",
         10281 => x"bcb83f82",
         10282 => x"e09808fd",
         10283 => x"b0387553",
         10284 => x"7c529418",
         10285 => x"0883ff06",
         10286 => x"1fb80551",
         10287 => x"ffb9d43f",
         10288 => x"7e55810b",
         10289 => x"8316347b",
         10290 => x"76317e08",
         10291 => x"177f0c76",
         10292 => x"1e941a08",
         10293 => x"1870941c",
         10294 => x"0c8c1b08",
         10295 => x"58585e5c",
         10296 => x"74762783",
         10297 => x"38755574",
         10298 => x"8c190cfd",
         10299 => x"89399018",
         10300 => x"3380c007",
         10301 => x"55749019",
         10302 => x"34805675",
         10303 => x"82e0980c",
         10304 => x"903d0d04",
         10305 => x"f83d0d7a",
         10306 => x"8b3dfc05",
         10307 => x"53705256",
         10308 => x"f2df3f82",
         10309 => x"e0980857",
         10310 => x"82e09808",
         10311 => x"81803890",
         10312 => x"16337086",
         10313 => x"2a708106",
         10314 => x"51555573",
         10315 => x"802e80ee",
         10316 => x"38a01608",
         10317 => x"527851ff",
         10318 => x"bba43f82",
         10319 => x"e0980857",
         10320 => x"82e09808",
         10321 => x"80d838a4",
         10322 => x"16088b11",
         10323 => x"33a00755",
         10324 => x"55738b16",
         10325 => x"34881608",
         10326 => x"53745275",
         10327 => x"0851cca5",
         10328 => x"3f8c1608",
         10329 => x"529c1551",
         10330 => x"ffb7f93f",
         10331 => x"8288b20a",
         10332 => x"52961551",
         10333 => x"ffb7ed3f",
         10334 => x"76529215",
         10335 => x"51ffb7c6",
         10336 => x"3f785481",
         10337 => x"0b831534",
         10338 => x"7851ffbb",
         10339 => x"983f82e0",
         10340 => x"98089017",
         10341 => x"3381bf06",
         10342 => x"55577390",
         10343 => x"17347682",
         10344 => x"e0980c8a",
         10345 => x"3d0d04fc",
         10346 => x"3d0d7670",
         10347 => x"5254fed4",
         10348 => x"3f82e098",
         10349 => x"085382e0",
         10350 => x"98089c38",
         10351 => x"863dfc05",
         10352 => x"527351f1",
         10353 => x"ac3f82e0",
         10354 => x"98085382",
         10355 => x"e0980887",
         10356 => x"3882e098",
         10357 => x"08740c72",
         10358 => x"82e0980c",
         10359 => x"863d0d04",
         10360 => x"ff3d0d84",
         10361 => x"3d51e689",
         10362 => x"3f8b5280",
         10363 => x"0b82e098",
         10364 => x"08248b38",
         10365 => x"82e09808",
         10366 => x"82f7f434",
         10367 => x"80527182",
         10368 => x"e0980c83",
         10369 => x"3d0d04ee",
         10370 => x"3d0d8053",
         10371 => x"943dcc05",
         10372 => x"52953d51",
         10373 => x"e8e63f82",
         10374 => x"e0980855",
         10375 => x"82e09808",
         10376 => x"80e03876",
         10377 => x"58645294",
         10378 => x"3dd00551",
         10379 => x"dce83f82",
         10380 => x"e0980855",
         10381 => x"82e09808",
         10382 => x"bc380280",
         10383 => x"c7053370",
         10384 => x"982b5556",
         10385 => x"73802589",
         10386 => x"38767a98",
         10387 => x"120c54b2",
         10388 => x"3902a205",
         10389 => x"3370842a",
         10390 => x"70810651",
         10391 => x"55567380",
         10392 => x"2e9e3876",
         10393 => x"7f537052",
         10394 => x"54c9e13f",
         10395 => x"82e09808",
         10396 => x"98150c8e",
         10397 => x"3982e098",
         10398 => x"08842e09",
         10399 => x"81068338",
         10400 => x"85557482",
         10401 => x"e0980c94",
         10402 => x"3d0d04ff",
         10403 => x"a33d0d80",
         10404 => x"e13d0880",
         10405 => x"e13d085b",
         10406 => x"5b807a34",
         10407 => x"805380df",
         10408 => x"3dfdb405",
         10409 => x"5280e03d",
         10410 => x"51e7d13f",
         10411 => x"82e09808",
         10412 => x"5782e098",
         10413 => x"0883a138",
         10414 => x"7b80d43d",
         10415 => x"0c7a7c98",
         10416 => x"110880d8",
         10417 => x"3d0c5558",
         10418 => x"80d53d08",
         10419 => x"5473802e",
         10420 => x"828338a0",
         10421 => x"5280d33d",
         10422 => x"705255c4",
         10423 => x"903f82e0",
         10424 => x"98085782",
         10425 => x"e0980882",
         10426 => x"ef3880d9",
         10427 => x"3d08527b",
         10428 => x"51ffb7ea",
         10429 => x"3f82e098",
         10430 => x"085782e0",
         10431 => x"980882d8",
         10432 => x"3880da3d",
         10433 => x"08527b51",
         10434 => x"c8c23f82",
         10435 => x"e0980880",
         10436 => x"d63d0c76",
         10437 => x"527451c3",
         10438 => x"d43f82e0",
         10439 => x"98085782",
         10440 => x"e0980882",
         10441 => x"b3388052",
         10442 => x"7451c9b6",
         10443 => x"3f82e098",
         10444 => x"085782e0",
         10445 => x"9808a738",
         10446 => x"80da3d08",
         10447 => x"527b51c8",
         10448 => x"8b3f7382",
         10449 => x"e098082e",
         10450 => x"a6387652",
         10451 => x"7451c4e8",
         10452 => x"3f82e098",
         10453 => x"085782e0",
         10454 => x"9808802e",
         10455 => x"c9387684",
         10456 => x"2e098106",
         10457 => x"86388257",
         10458 => x"81ee3976",
         10459 => x"81ea3880",
         10460 => x"df3dfdb8",
         10461 => x"05527451",
         10462 => x"d6a03f76",
         10463 => x"933d7811",
         10464 => x"82113351",
         10465 => x"565a5673",
         10466 => x"802e9238",
         10467 => x"0280c605",
         10468 => x"55811681",
         10469 => x"16703356",
         10470 => x"565673f5",
         10471 => x"38811654",
         10472 => x"73782681",
         10473 => x"99387580",
         10474 => x"2e9c3878",
         10475 => x"16820555",
         10476 => x"ff1880e1",
         10477 => x"3d0811ff",
         10478 => x"18ff1858",
         10479 => x"58555874",
         10480 => x"33743475",
         10481 => x"eb38ff18",
         10482 => x"80e13d08",
         10483 => x"115558af",
         10484 => x"7434fdf4",
         10485 => x"39777b2e",
         10486 => x"0981068d",
         10487 => x"38ff1880",
         10488 => x"e13d0811",
         10489 => x"5558af74",
         10490 => x"34800b82",
         10491 => x"f7f43370",
         10492 => x"842982d2",
         10493 => x"98057008",
         10494 => x"7033525c",
         10495 => x"56565673",
         10496 => x"762e8d38",
         10497 => x"8116701a",
         10498 => x"70335155",
         10499 => x"5673f538",
         10500 => x"82165473",
         10501 => x"7826a738",
         10502 => x"80557476",
         10503 => x"27913874",
         10504 => x"19547333",
         10505 => x"7a708105",
         10506 => x"5c348115",
         10507 => x"55ec39ba",
         10508 => x"7a708105",
         10509 => x"5c3474ff",
         10510 => x"2e098106",
         10511 => x"85389157",
         10512 => x"973980e0",
         10513 => x"3d081881",
         10514 => x"19595473",
         10515 => x"337a7081",
         10516 => x"055c347a",
         10517 => x"7826eb38",
         10518 => x"807a3476",
         10519 => x"82e0980c",
         10520 => x"80df3d0d",
         10521 => x"04f73d0d",
         10522 => x"7b7d8d3d",
         10523 => x"fc055471",
         10524 => x"535755eb",
         10525 => x"fc3f82e0",
         10526 => x"98085382",
         10527 => x"e0980882",
         10528 => x"fe389115",
         10529 => x"33537282",
         10530 => x"f6388c15",
         10531 => x"08547376",
         10532 => x"27923890",
         10533 => x"15337081",
         10534 => x"2a708106",
         10535 => x"51545772",
         10536 => x"83387356",
         10537 => x"94150854",
         10538 => x"80709417",
         10539 => x"0c587578",
         10540 => x"2e829b38",
         10541 => x"798a1122",
         10542 => x"70892b59",
         10543 => x"51537378",
         10544 => x"2eb73876",
         10545 => x"52ff1651",
         10546 => x"febc883f",
         10547 => x"82e09808",
         10548 => x"ff157854",
         10549 => x"70535553",
         10550 => x"febbf83f",
         10551 => x"82e09808",
         10552 => x"73269638",
         10553 => x"76307075",
         10554 => x"06709418",
         10555 => x"0c777131",
         10556 => x"98180857",
         10557 => x"585153b2",
         10558 => x"39881508",
         10559 => x"5473a738",
         10560 => x"73527451",
         10561 => x"ffbbd33f",
         10562 => x"82e09808",
         10563 => x"5482e098",
         10564 => x"08812e81",
         10565 => x"9d3882e0",
         10566 => x"9808ff2e",
         10567 => x"819e3882",
         10568 => x"e0980888",
         10569 => x"160c7398",
         10570 => x"160c7380",
         10571 => x"2e819f38",
         10572 => x"76762780",
         10573 => x"de387577",
         10574 => x"31941608",
         10575 => x"1894170c",
         10576 => x"90163370",
         10577 => x"812a7081",
         10578 => x"0651555a",
         10579 => x"5672802e",
         10580 => x"9b387352",
         10581 => x"7451ffbb",
         10582 => x"813f82e0",
         10583 => x"98085482",
         10584 => x"e0980895",
         10585 => x"3882e098",
         10586 => x"0856a839",
         10587 => x"73527451",
         10588 => x"ffb58b3f",
         10589 => x"82e09808",
         10590 => x"5473ff2e",
         10591 => x"bf388174",
         10592 => x"27b03879",
         10593 => x"53739c14",
         10594 => x"0827a738",
         10595 => x"7398160c",
         10596 => x"ff9e3994",
         10597 => x"15081694",
         10598 => x"160c7583",
         10599 => x"ff065372",
         10600 => x"802eab38",
         10601 => x"73527951",
         10602 => x"ffb4a93f",
         10603 => x"82e09808",
         10604 => x"9438820b",
         10605 => x"91163482",
         10606 => x"5380c439",
         10607 => x"810b9116",
         10608 => x"348153bb",
         10609 => x"3975892a",
         10610 => x"82e09808",
         10611 => x"05589415",
         10612 => x"08548c15",
         10613 => x"08742790",
         10614 => x"38738c16",
         10615 => x"0c901533",
         10616 => x"80c00753",
         10617 => x"72901634",
         10618 => x"7383ff06",
         10619 => x"5372802e",
         10620 => x"8c38779c",
         10621 => x"16082e85",
         10622 => x"38779c16",
         10623 => x"0c805372",
         10624 => x"82e0980c",
         10625 => x"8b3d0d04",
         10626 => x"f93d0d79",
         10627 => x"56895475",
         10628 => x"802e818b",
         10629 => x"38805389",
         10630 => x"3dfc0552",
         10631 => x"8a3d8405",
         10632 => x"51e0d93f",
         10633 => x"82e09808",
         10634 => x"5582e098",
         10635 => x"0880eb38",
         10636 => x"77760c7a",
         10637 => x"527551d4",
         10638 => x"dd3f82e0",
         10639 => x"98085582",
         10640 => x"e0980880",
         10641 => x"c438ab16",
         10642 => x"3370982b",
         10643 => x"55578074",
         10644 => x"24a23886",
         10645 => x"16337084",
         10646 => x"2a708106",
         10647 => x"51555773",
         10648 => x"802eae38",
         10649 => x"9c160852",
         10650 => x"7751c1e0",
         10651 => x"3f82e098",
         10652 => x"0888170c",
         10653 => x"77548614",
         10654 => x"22841723",
         10655 => x"74527551",
         10656 => x"ffbcea3f",
         10657 => x"82e09808",
         10658 => x"5574842e",
         10659 => x"09810685",
         10660 => x"38855586",
         10661 => x"3974802e",
         10662 => x"84388076",
         10663 => x"0c745473",
         10664 => x"82e0980c",
         10665 => x"893d0d04",
         10666 => x"fc3d0d76",
         10667 => x"873dfc05",
         10668 => x"53705253",
         10669 => x"e7bb3f82",
         10670 => x"e0980887",
         10671 => x"3882e098",
         10672 => x"08730c86",
         10673 => x"3d0d04fb",
         10674 => x"3d0d7779",
         10675 => x"893dfc05",
         10676 => x"54715356",
         10677 => x"54e79a3f",
         10678 => x"82e09808",
         10679 => x"5382e098",
         10680 => x"0880e138",
         10681 => x"74943882",
         10682 => x"e0980852",
         10683 => x"7351ffbb",
         10684 => x"fc3f82e0",
         10685 => x"98085380",
         10686 => x"cb3982e0",
         10687 => x"98085273",
         10688 => x"51c1df3f",
         10689 => x"82e09808",
         10690 => x"5382e098",
         10691 => x"08842e09",
         10692 => x"81068538",
         10693 => x"80538739",
         10694 => x"82e09808",
         10695 => x"a7387452",
         10696 => x"7351cef6",
         10697 => x"3f725273",
         10698 => x"51ffbd8c",
         10699 => x"3f82e098",
         10700 => x"08843270",
         10701 => x"30707207",
         10702 => x"9f2c7082",
         10703 => x"e0980806",
         10704 => x"51515454",
         10705 => x"7282e098",
         10706 => x"0c873d0d",
         10707 => x"04ed3d0d",
         10708 => x"66578053",
         10709 => x"893d7053",
         10710 => x"973d5256",
         10711 => x"de9e3f82",
         10712 => x"e0980855",
         10713 => x"82e09808",
         10714 => x"b2386552",
         10715 => x"7551d2a6",
         10716 => x"3f82e098",
         10717 => x"085582e0",
         10718 => x"9808a038",
         10719 => x"0280cb05",
         10720 => x"3370982b",
         10721 => x"55587380",
         10722 => x"25853886",
         10723 => x"558d3976",
         10724 => x"802e8838",
         10725 => x"76527551",
         10726 => x"ce803f74",
         10727 => x"82e0980c",
         10728 => x"953d0d04",
         10729 => x"f03d0d63",
         10730 => x"65555c80",
         10731 => x"53923dec",
         10732 => x"0552933d",
         10733 => x"51ddc53f",
         10734 => x"82e09808",
         10735 => x"5b82e098",
         10736 => x"08828238",
         10737 => x"7c740c73",
         10738 => x"089c1108",
         10739 => x"fe119413",
         10740 => x"08595658",
         10741 => x"55757426",
         10742 => x"9138757c",
         10743 => x"0c81e639",
         10744 => x"815b81ce",
         10745 => x"39825b81",
         10746 => x"c93982e0",
         10747 => x"98087533",
         10748 => x"55597381",
         10749 => x"2e098106",
         10750 => x"80c03882",
         10751 => x"755f5776",
         10752 => x"52923df0",
         10753 => x"0551ffaf",
         10754 => x"f53f82e0",
         10755 => x"9808ff2e",
         10756 => x"cf3882e0",
         10757 => x"9808812e",
         10758 => x"cc3882e0",
         10759 => x"98083070",
         10760 => x"82e09808",
         10761 => x"0780257a",
         10762 => x"0581197f",
         10763 => x"53595a54",
         10764 => x"9c140877",
         10765 => x"26c93880",
         10766 => x"f939a815",
         10767 => x"0882e098",
         10768 => x"08575875",
         10769 => x"98387752",
         10770 => x"81187d52",
         10771 => x"58ffad8e",
         10772 => x"3f82e098",
         10773 => x"085b82e0",
         10774 => x"980880d6",
         10775 => x"387c7033",
         10776 => x"7712ff1a",
         10777 => x"5d525654",
         10778 => x"74822e09",
         10779 => x"81069e38",
         10780 => x"b81451ff",
         10781 => x"a98e3f82",
         10782 => x"e0980883",
         10783 => x"ffff0670",
         10784 => x"30708025",
         10785 => x"1b821959",
         10786 => x"5b51549b",
         10787 => x"39b81451",
         10788 => x"ffa9883f",
         10789 => x"82e09808",
         10790 => x"f00a0670",
         10791 => x"30708025",
         10792 => x"1b841959",
         10793 => x"5b515475",
         10794 => x"83ff067a",
         10795 => x"585679ff",
         10796 => x"9238787c",
         10797 => x"0c7c7994",
         10798 => x"120c8411",
         10799 => x"33810756",
         10800 => x"54748415",
         10801 => x"347a82e0",
         10802 => x"980c923d",
         10803 => x"0d04f93d",
         10804 => x"0d798a3d",
         10805 => x"fc055370",
         10806 => x"5257e395",
         10807 => x"3f82e098",
         10808 => x"085682e0",
         10809 => x"980881aa",
         10810 => x"38911733",
         10811 => x"567581a2",
         10812 => x"38901733",
         10813 => x"70812a70",
         10814 => x"81065155",
         10815 => x"55875573",
         10816 => x"802e8190",
         10817 => x"38941708",
         10818 => x"54738c18",
         10819 => x"08278182",
         10820 => x"38739c38",
         10821 => x"82e09808",
         10822 => x"53881708",
         10823 => x"527651ff",
         10824 => x"b28c3f82",
         10825 => x"e0980874",
         10826 => x"88190c56",
         10827 => x"80ca3998",
         10828 => x"17085276",
         10829 => x"51ffadc6",
         10830 => x"3f82e098",
         10831 => x"08ff2e09",
         10832 => x"81068338",
         10833 => x"815682e0",
         10834 => x"9808812e",
         10835 => x"09810685",
         10836 => x"388256a4",
         10837 => x"3975a138",
         10838 => x"775482e0",
         10839 => x"98089c15",
         10840 => x"08279538",
         10841 => x"98170853",
         10842 => x"82e09808",
         10843 => x"527651ff",
         10844 => x"b1bc3f82",
         10845 => x"e0980856",
         10846 => x"9417088c",
         10847 => x"180c9017",
         10848 => x"3380c007",
         10849 => x"54739018",
         10850 => x"3475802e",
         10851 => x"85387591",
         10852 => x"18347555",
         10853 => x"7482e098",
         10854 => x"0c893d0d",
         10855 => x"04e03d0d",
         10856 => x"8253a23d",
         10857 => x"ff9c0552",
         10858 => x"a33d51d9",
         10859 => x"cf3f82e0",
         10860 => x"98085582",
         10861 => x"e0980881",
         10862 => x"f9387846",
         10863 => x"a33d0852",
         10864 => x"963d7052",
         10865 => x"58cdcf3f",
         10866 => x"82e09808",
         10867 => x"5582e098",
         10868 => x"0881df38",
         10869 => x"0280ff05",
         10870 => x"3370852a",
         10871 => x"70810651",
         10872 => x"55568655",
         10873 => x"7381cb38",
         10874 => x"75982b54",
         10875 => x"80742481",
         10876 => x"c1380280",
         10877 => x"da053370",
         10878 => x"81065854",
         10879 => x"87557681",
         10880 => x"b1386c52",
         10881 => x"7851ffba",
         10882 => x"c33f82e0",
         10883 => x"98087484",
         10884 => x"2a708106",
         10885 => x"51555673",
         10886 => x"802e80d6",
         10887 => x"38785482",
         10888 => x"e0980898",
         10889 => x"15082e81",
         10890 => x"8938735a",
         10891 => x"82e09808",
         10892 => x"5c76528a",
         10893 => x"3d705254",
         10894 => x"ffb5b23f",
         10895 => x"82e09808",
         10896 => x"5582e098",
         10897 => x"0880eb38",
         10898 => x"82e09808",
         10899 => x"527351ff",
         10900 => x"bb903f82",
         10901 => x"e0980855",
         10902 => x"82e09808",
         10903 => x"86388755",
         10904 => x"80d03982",
         10905 => x"e0980884",
         10906 => x"2e883882",
         10907 => x"e0980880",
         10908 => x"c1387751",
         10909 => x"c7ab3f82",
         10910 => x"e0980882",
         10911 => x"e0980830",
         10912 => x"7082e098",
         10913 => x"08078025",
         10914 => x"51555575",
         10915 => x"802e9538",
         10916 => x"73802e90",
         10917 => x"38805375",
         10918 => x"527751ff",
         10919 => x"af903f82",
         10920 => x"e0980855",
         10921 => x"748c3878",
         10922 => x"51ffa8f9",
         10923 => x"3f82e098",
         10924 => x"08557482",
         10925 => x"e0980ca2",
         10926 => x"3d0d04e8",
         10927 => x"3d0d8253",
         10928 => x"9a3dffbc",
         10929 => x"05529b3d",
         10930 => x"51d7b13f",
         10931 => x"82e09808",
         10932 => x"5482e098",
         10933 => x"0882b738",
         10934 => x"785e6a52",
         10935 => x"8e3d7052",
         10936 => x"58cbb33f",
         10937 => x"82e09808",
         10938 => x"5482e098",
         10939 => x"08863888",
         10940 => x"54829b39",
         10941 => x"82e09808",
         10942 => x"842e0981",
         10943 => x"06828f38",
         10944 => x"0280df05",
         10945 => x"3370852a",
         10946 => x"81065155",
         10947 => x"86547481",
         10948 => x"fd38785a",
         10949 => x"74528a3d",
         10950 => x"705257ff",
         10951 => x"afbc3f82",
         10952 => x"e0980875",
         10953 => x"555682e0",
         10954 => x"98088338",
         10955 => x"875482e0",
         10956 => x"9808812e",
         10957 => x"09810683",
         10958 => x"38825482",
         10959 => x"e09808ff",
         10960 => x"2e098106",
         10961 => x"86388154",
         10962 => x"81ba3973",
         10963 => x"81b63882",
         10964 => x"e0980852",
         10965 => x"7851ffb2",
         10966 => x"9c3f82e0",
         10967 => x"98085482",
         10968 => x"e0980881",
         10969 => x"9f388b53",
         10970 => x"a052b819",
         10971 => x"51ffa4c6",
         10972 => x"3f7854ae",
         10973 => x"0bb81534",
         10974 => x"7854900b",
         10975 => x"80c31534",
         10976 => x"8288b20a",
         10977 => x"5280ce19",
         10978 => x"51ffa3d8",
         10979 => x"3f755378",
         10980 => x"b8115351",
         10981 => x"ffb7ee3f",
         10982 => x"a05378b8",
         10983 => x"115380d8",
         10984 => x"0551ffa3",
         10985 => x"ee3f7854",
         10986 => x"ae0b80d9",
         10987 => x"15347f53",
         10988 => x"7880d811",
         10989 => x"5351ffb7",
         10990 => x"cc3f7854",
         10991 => x"810b8315",
         10992 => x"347751ff",
         10993 => x"bf893f82",
         10994 => x"e0980854",
         10995 => x"82e09808",
         10996 => x"b3388288",
         10997 => x"b20a5264",
         10998 => x"960551ff",
         10999 => x"a3863f75",
         11000 => x"53645278",
         11001 => x"51ffb79d",
         11002 => x"3f645490",
         11003 => x"0b8b1534",
         11004 => x"7854810b",
         11005 => x"83153478",
         11006 => x"51ffa6a9",
         11007 => x"3f82e098",
         11008 => x"08548b39",
         11009 => x"80537552",
         11010 => x"7651ffac",
         11011 => x"a13f7382",
         11012 => x"e0980c9a",
         11013 => x"3d0d04d8",
         11014 => x"3d0dab3d",
         11015 => x"840551d1",
         11016 => x"d03f8253",
         11017 => x"aa3dfefc",
         11018 => x"0552ab3d",
         11019 => x"51d4cd3f",
         11020 => x"82e09808",
         11021 => x"5582e098",
         11022 => x"0882d838",
         11023 => x"784eab3d",
         11024 => x"08529e3d",
         11025 => x"705258c8",
         11026 => x"cd3f82e0",
         11027 => x"98085582",
         11028 => x"e0980882",
         11029 => x"be380281",
         11030 => x"9f053381",
         11031 => x"a0065486",
         11032 => x"557382af",
         11033 => x"38a053a5",
         11034 => x"3d0852aa",
         11035 => x"3dff8005",
         11036 => x"51ffa29f",
         11037 => x"3fb05377",
         11038 => x"52923d70",
         11039 => x"5254ffa2",
         11040 => x"923fac3d",
         11041 => x"08527351",
         11042 => x"c88c3f82",
         11043 => x"e0980855",
         11044 => x"82e09808",
         11045 => x"973863a1",
         11046 => x"3d082e09",
         11047 => x"81068838",
         11048 => x"65a33d08",
         11049 => x"2e923888",
         11050 => x"5581e839",
         11051 => x"82e09808",
         11052 => x"842e0981",
         11053 => x"0681bb38",
         11054 => x"7351ffbd",
         11055 => x"923f82e0",
         11056 => x"98085582",
         11057 => x"e0980881",
         11058 => x"ca386856",
         11059 => x"9353aa3d",
         11060 => x"ff8d0552",
         11061 => x"8d1651ff",
         11062 => x"a1b93f02",
         11063 => x"af05338b",
         11064 => x"17348b16",
         11065 => x"3370842a",
         11066 => x"70810651",
         11067 => x"55557389",
         11068 => x"3874a007",
         11069 => x"54738b17",
         11070 => x"34785481",
         11071 => x"0b831534",
         11072 => x"8b163370",
         11073 => x"842a7081",
         11074 => x"06515555",
         11075 => x"73802e80",
         11076 => x"e7386f64",
         11077 => x"2e80e138",
         11078 => x"75527851",
         11079 => x"ffb4ad3f",
         11080 => x"82e09808",
         11081 => x"527851ff",
         11082 => x"a5aa3f82",
         11083 => x"5582e098",
         11084 => x"08802e80",
         11085 => x"de3882e0",
         11086 => x"98085278",
         11087 => x"51ffa39e",
         11088 => x"3f82e098",
         11089 => x"087980d8",
         11090 => x"11585855",
         11091 => x"82e09808",
         11092 => x"80c13881",
         11093 => x"16335473",
         11094 => x"ae2e0981",
         11095 => x"069a3863",
         11096 => x"53755276",
         11097 => x"51ffb49d",
         11098 => x"3f785481",
         11099 => x"0b831534",
         11100 => x"873982e0",
         11101 => x"98089c38",
         11102 => x"7751c1a5",
         11103 => x"3f82e098",
         11104 => x"085582e0",
         11105 => x"98088c38",
         11106 => x"7851ffa3",
         11107 => x"983f82e0",
         11108 => x"98085574",
         11109 => x"82e0980c",
         11110 => x"aa3d0d04",
         11111 => x"ec3d0d02",
         11112 => x"80df0533",
         11113 => x"02840580",
         11114 => x"e3053357",
         11115 => x"57825396",
         11116 => x"3dcc0552",
         11117 => x"973d51d1",
         11118 => x"c33f82e0",
         11119 => x"98085582",
         11120 => x"e0980880",
         11121 => x"cf38785a",
         11122 => x"6652963d",
         11123 => x"d00551c5",
         11124 => x"c53f82e0",
         11125 => x"98085582",
         11126 => x"e09808b8",
         11127 => x"380280cf",
         11128 => x"053381a0",
         11129 => x"06548655",
         11130 => x"73aa3875",
         11131 => x"a7066171",
         11132 => x"098b1233",
         11133 => x"71067a74",
         11134 => x"06075157",
         11135 => x"5556748b",
         11136 => x"15347854",
         11137 => x"810b8315",
         11138 => x"347851ff",
         11139 => x"a2973f82",
         11140 => x"e0980855",
         11141 => x"7482e098",
         11142 => x"0c963d0d",
         11143 => x"04ee3d0d",
         11144 => x"65568253",
         11145 => x"943dcc05",
         11146 => x"52953d51",
         11147 => x"d0ce3f82",
         11148 => x"e0980855",
         11149 => x"82e09808",
         11150 => x"80cb3876",
         11151 => x"58645294",
         11152 => x"3dd00551",
         11153 => x"c4d03f82",
         11154 => x"e0980855",
         11155 => x"82e09808",
         11156 => x"b4380280",
         11157 => x"c7053381",
         11158 => x"a0065486",
         11159 => x"5573a638",
         11160 => x"84162286",
         11161 => x"17227190",
         11162 => x"2b075354",
         11163 => x"961f51ff",
         11164 => x"9df23f76",
         11165 => x"54810b83",
         11166 => x"15347651",
         11167 => x"ffa1a63f",
         11168 => x"82e09808",
         11169 => x"557482e0",
         11170 => x"980c943d",
         11171 => x"0d04e93d",
         11172 => x"0d6a6c5c",
         11173 => x"5a805399",
         11174 => x"3dcc0552",
         11175 => x"9a3d51cf",
         11176 => x"db3f82e0",
         11177 => x"980882e0",
         11178 => x"98083070",
         11179 => x"82e09808",
         11180 => x"07802551",
         11181 => x"55577980",
         11182 => x"2e818638",
         11183 => x"81707506",
         11184 => x"55557380",
         11185 => x"2e80fa38",
         11186 => x"7b5d805f",
         11187 => x"80528d3d",
         11188 => x"705254ff",
         11189 => x"ac973f82",
         11190 => x"e0980857",
         11191 => x"82e09808",
         11192 => x"80d23874",
         11193 => x"527351ff",
         11194 => x"b1f83f82",
         11195 => x"e0980857",
         11196 => x"82e09808",
         11197 => x"bf3882e0",
         11198 => x"980882e0",
         11199 => x"9808655b",
         11200 => x"59567818",
         11201 => x"81197b18",
         11202 => x"56595574",
         11203 => x"33743481",
         11204 => x"16568a78",
         11205 => x"27ec388b",
         11206 => x"56751a54",
         11207 => x"80743475",
         11208 => x"802e9e38",
         11209 => x"ff16701b",
         11210 => x"70335155",
         11211 => x"5673a02e",
         11212 => x"e8388e39",
         11213 => x"76842e09",
         11214 => x"81068638",
         11215 => x"807a3480",
         11216 => x"57763070",
         11217 => x"78078025",
         11218 => x"51547a80",
         11219 => x"2e80c138",
         11220 => x"73802ebc",
         11221 => x"387ba411",
         11222 => x"085351ff",
         11223 => x"9f803f82",
         11224 => x"e0980857",
         11225 => x"82e09808",
         11226 => x"a7387b70",
         11227 => x"33555580",
         11228 => x"c3567383",
         11229 => x"2e8b3880",
         11230 => x"e4567384",
         11231 => x"2e8338a7",
         11232 => x"567515b8",
         11233 => x"0551ff9b",
         11234 => x"923f82e0",
         11235 => x"98087b0c",
         11236 => x"7682e098",
         11237 => x"0c993d0d",
         11238 => x"04e63d0d",
         11239 => x"82539c3d",
         11240 => x"ffb40552",
         11241 => x"9d3d51cd",
         11242 => x"d33f82e0",
         11243 => x"980882e0",
         11244 => x"98085654",
         11245 => x"82e09808",
         11246 => x"82dd388b",
         11247 => x"53a0528a",
         11248 => x"3d705258",
         11249 => x"ff9bef3f",
         11250 => x"736d7033",
         11251 => x"5155569f",
         11252 => x"74278186",
         11253 => x"3877579d",
         11254 => x"3d51ff9c",
         11255 => x"cc3f82e0",
         11256 => x"980883ff",
         11257 => x"ff2680c4",
         11258 => x"3882e098",
         11259 => x"085196c0",
         11260 => x"3f83b552",
         11261 => x"82e09808",
         11262 => x"5195903f",
         11263 => x"82e09808",
         11264 => x"83ffff06",
         11265 => x"5574802e",
         11266 => x"a3387452",
         11267 => x"82d3b851",
         11268 => x"ff9bee3f",
         11269 => x"82e09808",
         11270 => x"933881ff",
         11271 => x"75278838",
         11272 => x"75892688",
         11273 => x"388b398a",
         11274 => x"76278638",
         11275 => x"865581e7",
         11276 => x"3981ff75",
         11277 => x"278f3874",
         11278 => x"882a5473",
         11279 => x"77708105",
         11280 => x"59348116",
         11281 => x"56747770",
         11282 => x"81055934",
         11283 => x"81166d70",
         11284 => x"33515556",
         11285 => x"739f26fe",
         11286 => x"fe388a3d",
         11287 => x"33548655",
         11288 => x"7381e52e",
         11289 => x"81b13875",
         11290 => x"802e9938",
         11291 => x"02a30555",
         11292 => x"75157033",
         11293 => x"515473a0",
         11294 => x"2e098106",
         11295 => x"8738ff16",
         11296 => x"5675ed38",
         11297 => x"78408042",
         11298 => x"8052903d",
         11299 => x"705255ff",
         11300 => x"a8db3f82",
         11301 => x"e0980854",
         11302 => x"82e09808",
         11303 => x"80f73881",
         11304 => x"527451ff",
         11305 => x"aebc3f82",
         11306 => x"e0980854",
         11307 => x"82e09808",
         11308 => x"8d387580",
         11309 => x"c4386654",
         11310 => x"e5743480",
         11311 => x"c63982e0",
         11312 => x"9808842e",
         11313 => x"09810680",
         11314 => x"cc388054",
         11315 => x"75742e80",
         11316 => x"c4388152",
         11317 => x"7451ffab",
         11318 => x"d83f82e0",
         11319 => x"98085482",
         11320 => x"e09808b1",
         11321 => x"38a05382",
         11322 => x"e0980852",
         11323 => x"6651ff99",
         11324 => x"c53f6654",
         11325 => x"880b8b15",
         11326 => x"348b5377",
         11327 => x"526651ff",
         11328 => x"99913f78",
         11329 => x"54810b83",
         11330 => x"15347851",
         11331 => x"ff9c963f",
         11332 => x"82e09808",
         11333 => x"54735574",
         11334 => x"82e0980c",
         11335 => x"9c3d0d04",
         11336 => x"f23d0d60",
         11337 => x"62028805",
         11338 => x"80cb0533",
         11339 => x"933dfc05",
         11340 => x"55725440",
         11341 => x"5e5ad2b9",
         11342 => x"3f82e098",
         11343 => x"085882e0",
         11344 => x"980882bd",
         11345 => x"38911a33",
         11346 => x"587782b5",
         11347 => x"387c802e",
         11348 => x"97388c1a",
         11349 => x"08597890",
         11350 => x"38901a33",
         11351 => x"70812a70",
         11352 => x"81065155",
         11353 => x"55739038",
         11354 => x"87548297",
         11355 => x"39825882",
         11356 => x"90398158",
         11357 => x"828b397e",
         11358 => x"8a112270",
         11359 => x"892b7055",
         11360 => x"7f545656",
         11361 => x"56fea2cb",
         11362 => x"3fff147d",
         11363 => x"06703070",
         11364 => x"72079f2a",
         11365 => x"82e09808",
         11366 => x"05901908",
         11367 => x"7c405a5d",
         11368 => x"55558177",
         11369 => x"2788389c",
         11370 => x"16087726",
         11371 => x"83388257",
         11372 => x"76775659",
         11373 => x"80567452",
         11374 => x"7951ff9c",
         11375 => x"c13f8115",
         11376 => x"7f55559c",
         11377 => x"14087526",
         11378 => x"83388255",
         11379 => x"82e09808",
         11380 => x"812eff99",
         11381 => x"3882e098",
         11382 => x"08ff2eff",
         11383 => x"953882e0",
         11384 => x"98088e38",
         11385 => x"81165675",
         11386 => x"7b2e0981",
         11387 => x"06873893",
         11388 => x"39745980",
         11389 => x"5674772e",
         11390 => x"098106ff",
         11391 => x"b9388758",
         11392 => x"80ff397d",
         11393 => x"802eba38",
         11394 => x"787b5555",
         11395 => x"7a802eb4",
         11396 => x"38811556",
         11397 => x"73812e09",
         11398 => x"81068338",
         11399 => x"ff567553",
         11400 => x"74527e51",
         11401 => x"ff9dd03f",
         11402 => x"82e09808",
         11403 => x"5882e098",
         11404 => x"0880ce38",
         11405 => x"748116ff",
         11406 => x"1656565c",
         11407 => x"73d33884",
         11408 => x"39ff195c",
         11409 => x"7e7c9012",
         11410 => x"0c557d80",
         11411 => x"2eb33878",
         11412 => x"881b0c7c",
         11413 => x"8c1b0c90",
         11414 => x"1a3380c0",
         11415 => x"07547390",
         11416 => x"1b349c15",
         11417 => x"08fe0594",
         11418 => x"16085754",
         11419 => x"75742691",
         11420 => x"38757b31",
         11421 => x"94160c84",
         11422 => x"15338107",
         11423 => x"54738416",
         11424 => x"34775473",
         11425 => x"82e0980c",
         11426 => x"903d0d04",
         11427 => x"e83d0d6c",
         11428 => x"6e028805",
         11429 => x"80ef0533",
         11430 => x"9e3d5445",
         11431 => x"5c59c4d1",
         11432 => x"3f8b5680",
         11433 => x"0b82e098",
         11434 => x"08248da0",
         11435 => x"3882e098",
         11436 => x"08842982",
         11437 => x"f7e00570",
         11438 => x"08515574",
         11439 => x"802e8438",
         11440 => x"80753482",
         11441 => x"e0980882",
         11442 => x"e0980805",
         11443 => x"82e08c11",
         11444 => x"3382e08d",
         11445 => x"12334741",
         11446 => x"5581527f",
         11447 => x"51ff8eac",
         11448 => x"3f82e098",
         11449 => x"0881ff06",
         11450 => x"70810656",
         11451 => x"57835674",
         11452 => x"8cda3876",
         11453 => x"822a7081",
         11454 => x"0651558a",
         11455 => x"56748ccc",
         11456 => x"389a3dfc",
         11457 => x"05538352",
         11458 => x"7f51ff92",
         11459 => x"cc3f82e0",
         11460 => x"98089938",
         11461 => x"68557480",
         11462 => x"2e923874",
         11463 => x"82808026",
         11464 => x"8b38ff15",
         11465 => x"75065574",
         11466 => x"802e8338",
         11467 => x"81497880",
         11468 => x"2e873884",
         11469 => x"80792692",
         11470 => x"38788180",
         11471 => x"0a268b38",
         11472 => x"ff197906",
         11473 => x"5574802e",
         11474 => x"86389356",
         11475 => x"8bfe3978",
         11476 => x"892a6f89",
         11477 => x"2a70892b",
         11478 => x"77594943",
         11479 => x"597a8338",
         11480 => x"81566130",
         11481 => x"70802577",
         11482 => x"07515591",
         11483 => x"56748bdc",
         11484 => x"3864802e",
         11485 => x"80e03881",
         11486 => x"5474537a",
         11487 => x"527f51ff",
         11488 => x"8e893f81",
         11489 => x"5682e098",
         11490 => x"088bc138",
         11491 => x"83fe1b51",
         11492 => x"ff92f13f",
         11493 => x"82e09808",
         11494 => x"83ffff06",
         11495 => x"558e5674",
         11496 => x"82d4d52e",
         11497 => x"0981068b",
         11498 => x"a3386490",
         11499 => x"291b83b2",
         11500 => x"11335657",
         11501 => x"74802e8b",
         11502 => x"933883b6",
         11503 => x"1751ff92",
         11504 => x"da3f82e0",
         11505 => x"980883ba",
         11506 => x"18525fff",
         11507 => x"92cd3f82",
         11508 => x"e0980848",
         11509 => x"b7399a3d",
         11510 => x"f8055381",
         11511 => x"527f51ff",
         11512 => x"90f73f81",
         11513 => x"5682e098",
         11514 => x"088ae138",
         11515 => x"62832a70",
         11516 => x"770682e0",
         11517 => x"98084151",
         11518 => x"55748338",
         11519 => x"bf5f6755",
         11520 => x"8e567e75",
         11521 => x"268ac538",
         11522 => x"747f3148",
         11523 => x"8e5680ff",
         11524 => x"68278ab8",
         11525 => x"38935678",
         11526 => x"8180268a",
         11527 => x"af386281",
         11528 => x"2a708106",
         11529 => x"56447480",
         11530 => x"2e953862",
         11531 => x"87065574",
         11532 => x"822e838d",
         11533 => x"38628106",
         11534 => x"5574802e",
         11535 => x"83833862",
         11536 => x"81065593",
         11537 => x"56825e74",
         11538 => x"802e8a80",
         11539 => x"38785a7d",
         11540 => x"832e0981",
         11541 => x"0680e138",
         11542 => x"78ae3867",
         11543 => x"912a5781",
         11544 => x"0b82d3dc",
         11545 => x"22565a74",
         11546 => x"802e9d38",
         11547 => x"74772698",
         11548 => x"3882d3dc",
         11549 => x"56791082",
         11550 => x"17702257",
         11551 => x"575a7480",
         11552 => x"2e863876",
         11553 => x"7527ee38",
         11554 => x"79526751",
         11555 => x"fe9cc43f",
         11556 => x"82e09808",
         11557 => x"84298487",
         11558 => x"0570892a",
         11559 => x"5e55a05c",
         11560 => x"800b82e0",
         11561 => x"9808fc80",
         11562 => x"8a055646",
         11563 => x"fdfff00a",
         11564 => x"752780ec",
         11565 => x"38898839",
         11566 => x"78ae3867",
         11567 => x"8c2a5781",
         11568 => x"0b82d3cc",
         11569 => x"22565a74",
         11570 => x"802e9d38",
         11571 => x"74772698",
         11572 => x"3882d3cc",
         11573 => x"56791082",
         11574 => x"17702257",
         11575 => x"575a7480",
         11576 => x"2e863876",
         11577 => x"7527ee38",
         11578 => x"79526751",
         11579 => x"fe9be43f",
         11580 => x"82e09808",
         11581 => x"10840557",
         11582 => x"82e09808",
         11583 => x"9ff52696",
         11584 => x"38810b82",
         11585 => x"e0980810",
         11586 => x"82e09808",
         11587 => x"05711172",
         11588 => x"2a830559",
         11589 => x"565e83ff",
         11590 => x"17892a5d",
         11591 => x"815ca046",
         11592 => x"7b1f7d11",
         11593 => x"67056a70",
         11594 => x"12ff0571",
         11595 => x"30707206",
         11596 => x"74315c52",
         11597 => x"59575941",
         11598 => x"7d832e09",
         11599 => x"81068938",
         11600 => x"761c6118",
         11601 => x"425c8439",
         11602 => x"761d5d79",
         11603 => x"90291870",
         11604 => x"60316958",
         11605 => x"51557476",
         11606 => x"2687e438",
         11607 => x"757c317d",
         11608 => x"317a5370",
         11609 => x"67315255",
         11610 => x"fe9ae83f",
         11611 => x"82e09808",
         11612 => x"587d832e",
         11613 => x"0981069b",
         11614 => x"3882e098",
         11615 => x"0883fff5",
         11616 => x"2680dd38",
         11617 => x"7887b838",
         11618 => x"79812a59",
         11619 => x"78fdbe38",
         11620 => x"87ad397d",
         11621 => x"822e0981",
         11622 => x"0680c538",
         11623 => x"83fff50b",
         11624 => x"82e09808",
         11625 => x"27a03878",
         11626 => x"8f38791a",
         11627 => x"557480c0",
         11628 => x"26863874",
         11629 => x"59fd9639",
         11630 => x"63810655",
         11631 => x"74802e8f",
         11632 => x"38835efd",
         11633 => x"883982e0",
         11634 => x"98089ff5",
         11635 => x"26923878",
         11636 => x"86ed3879",
         11637 => x"1a598180",
         11638 => x"7927fcf1",
         11639 => x"3886e039",
         11640 => x"80557d81",
         11641 => x"2e098106",
         11642 => x"83387d55",
         11643 => x"9ff57827",
         11644 => x"8b387481",
         11645 => x"06558e56",
         11646 => x"7486d138",
         11647 => x"84805380",
         11648 => x"527a51ff",
         11649 => x"8fb03f8b",
         11650 => x"5382d1e4",
         11651 => x"527a51ff",
         11652 => x"8f813f84",
         11653 => x"80528b1b",
         11654 => x"51ff8eaa",
         11655 => x"3f798d1c",
         11656 => x"347b83ff",
         11657 => x"ff06528e",
         11658 => x"1b51ff8e",
         11659 => x"993f810b",
         11660 => x"901c347d",
         11661 => x"83327030",
         11662 => x"70962a84",
         11663 => x"80065451",
         11664 => x"55911b51",
         11665 => x"ff8dff3f",
         11666 => x"67557483",
         11667 => x"ffff2690",
         11668 => x"387483ff",
         11669 => x"ff065293",
         11670 => x"1b51ff8d",
         11671 => x"e93f8a39",
         11672 => x"7452a01b",
         11673 => x"51ff8dfc",
         11674 => x"3ff80b95",
         11675 => x"1c34bf52",
         11676 => x"981b51ff",
         11677 => x"8dd03f81",
         11678 => x"ff529a1b",
         11679 => x"51ff8dc6",
         11680 => x"3f7e529c",
         11681 => x"1b51ff8d",
         11682 => x"db3f7d83",
         11683 => x"2e098106",
         11684 => x"80cb3882",
         11685 => x"88b20a52",
         11686 => x"80c31b51",
         11687 => x"ff8dc53f",
         11688 => x"7c52a41b",
         11689 => x"51ff8dbc",
         11690 => x"3f8252ac",
         11691 => x"1b51ff8d",
         11692 => x"b33f8152",
         11693 => x"b01b51ff",
         11694 => x"8d8c3f86",
         11695 => x"52b21b51",
         11696 => x"ff8d833f",
         11697 => x"ff800b80",
         11698 => x"c01c34a9",
         11699 => x"0b80c21c",
         11700 => x"34935382",
         11701 => x"d1f05280",
         11702 => x"c71b51ae",
         11703 => x"398288b2",
         11704 => x"0a52a71b",
         11705 => x"51ff8cfc",
         11706 => x"3f7c83ff",
         11707 => x"ff065296",
         11708 => x"1b51ff8c",
         11709 => x"d13fff80",
         11710 => x"0ba41c34",
         11711 => x"a90ba61c",
         11712 => x"34935382",
         11713 => x"d28452ab",
         11714 => x"1b51ff8d",
         11715 => x"863f82d4",
         11716 => x"d55283fe",
         11717 => x"1b705259",
         11718 => x"ff8cab3f",
         11719 => x"81547e53",
         11720 => x"7a527f51",
         11721 => x"ff88ce3f",
         11722 => x"815682e0",
         11723 => x"9808849c",
         11724 => x"387d832e",
         11725 => x"09810680",
         11726 => x"ec387554",
         11727 => x"861f537a",
         11728 => x"527f51ff",
         11729 => x"88af3f84",
         11730 => x"80538052",
         11731 => x"7a51ff8c",
         11732 => x"e53f848b",
         11733 => x"85a4d252",
         11734 => x"7a51ff8c",
         11735 => x"873f868a",
         11736 => x"85e4f252",
         11737 => x"83e41b51",
         11738 => x"ff8bf93f",
         11739 => x"ff185283",
         11740 => x"e81b51ff",
         11741 => x"8bee3f82",
         11742 => x"5283ec1b",
         11743 => x"51ff8be4",
         11744 => x"3f82d4d5",
         11745 => x"527851ff",
         11746 => x"8bbc3f75",
         11747 => x"54871f53",
         11748 => x"7a527f51",
         11749 => x"ff87de3f",
         11750 => x"7554751f",
         11751 => x"537a527f",
         11752 => x"51ff87d1",
         11753 => x"3f665380",
         11754 => x"527a51ff",
         11755 => x"8c883f60",
         11756 => x"5680587d",
         11757 => x"832e0981",
         11758 => x"069a38f8",
         11759 => x"527a51ff",
         11760 => x"8ba23fff",
         11761 => x"52841b51",
         11762 => x"ff8b993f",
         11763 => x"f00a5288",
         11764 => x"1b519139",
         11765 => x"87fffff8",
         11766 => x"557d812e",
         11767 => x"8338f855",
         11768 => x"74527a51",
         11769 => x"ff8afd3f",
         11770 => x"7c556157",
         11771 => x"74622683",
         11772 => x"38745776",
         11773 => x"5475537a",
         11774 => x"527f51ff",
         11775 => x"86f73f82",
         11776 => x"e0980882",
         11777 => x"be388480",
         11778 => x"5382e098",
         11779 => x"08527a51",
         11780 => x"ff8ba33f",
         11781 => x"76167578",
         11782 => x"31565674",
         11783 => x"cd388118",
         11784 => x"5877802e",
         11785 => x"ff8d3879",
         11786 => x"557d832e",
         11787 => x"83386555",
         11788 => x"61577462",
         11789 => x"26833874",
         11790 => x"57765475",
         11791 => x"537a527f",
         11792 => x"51ff86b1",
         11793 => x"3f82e098",
         11794 => x"0881f838",
         11795 => x"76167578",
         11796 => x"31565674",
         11797 => x"db388c57",
         11798 => x"7d832e93",
         11799 => x"38865767",
         11800 => x"83ffff26",
         11801 => x"8a388457",
         11802 => x"7d822e83",
         11803 => x"38815764",
         11804 => x"802eb238",
         11805 => x"81548053",
         11806 => x"7a527f51",
         11807 => x"ff848c3f",
         11808 => x"815682e0",
         11809 => x"980881c4",
         11810 => x"38649029",
         11811 => x"1b557683",
         11812 => x"b2163475",
         11813 => x"5482e098",
         11814 => x"08537a52",
         11815 => x"7f51ff85",
         11816 => x"d43f8181",
         11817 => x"3962832a",
         11818 => x"81065877",
         11819 => x"80fd3884",
         11820 => x"80537752",
         11821 => x"7a51ff89",
         11822 => x"fd3f82d4",
         11823 => x"d5527851",
         11824 => x"ff89833f",
         11825 => x"83be1b55",
         11826 => x"77753481",
         11827 => x"0b811634",
         11828 => x"810b8216",
         11829 => x"34778316",
         11830 => x"34768416",
         11831 => x"34671f56",
         11832 => x"80fdc152",
         11833 => x"7551fe93",
         11834 => x"ea3ffe0b",
         11835 => x"85163482",
         11836 => x"e0980882",
         11837 => x"2abf0756",
         11838 => x"75861634",
         11839 => x"82e09808",
         11840 => x"8716347e",
         11841 => x"5283c61b",
         11842 => x"51ff88d8",
         11843 => x"3f675283",
         11844 => x"ca1b51ff",
         11845 => x"88ce3f81",
         11846 => x"5477537a",
         11847 => x"527f51ff",
         11848 => x"84d33f81",
         11849 => x"5682e098",
         11850 => x"08a23880",
         11851 => x"5380527f",
         11852 => x"51ff86a5",
         11853 => x"3f815682",
         11854 => x"e0980890",
         11855 => x"3889398e",
         11856 => x"568a3981",
         11857 => x"56863982",
         11858 => x"e0980856",
         11859 => x"7582e098",
         11860 => x"0c9a3d0d",
         11861 => x"04f53d0d",
         11862 => x"7d605b59",
         11863 => x"807960ff",
         11864 => x"055a5757",
         11865 => x"767825b4",
         11866 => x"388d3df8",
         11867 => x"11555581",
         11868 => x"53fc1552",
         11869 => x"7951c894",
         11870 => x"3f7a812e",
         11871 => x"0981069c",
         11872 => x"388c3d33",
         11873 => x"55748d2e",
         11874 => x"db387476",
         11875 => x"70810558",
         11876 => x"34811757",
         11877 => x"748a2e09",
         11878 => x"8106c938",
         11879 => x"80763478",
         11880 => x"55768338",
         11881 => x"76557482",
         11882 => x"e0980c8d",
         11883 => x"3d0d04f7",
         11884 => x"3d0d7b02",
         11885 => x"8405b305",
         11886 => x"33595777",
         11887 => x"8a2e0981",
         11888 => x"0687388d",
         11889 => x"527651e7",
         11890 => x"3f841708",
         11891 => x"56807624",
         11892 => x"be388817",
         11893 => x"0877178c",
         11894 => x"05565977",
         11895 => x"75348116",
         11896 => x"56bb7625",
         11897 => x"a1388b3d",
         11898 => x"fc055475",
         11899 => x"538c1752",
         11900 => x"760851ca",
         11901 => x"973f7976",
         11902 => x"32703070",
         11903 => x"72079f2a",
         11904 => x"70305351",
         11905 => x"56567584",
         11906 => x"180c8119",
         11907 => x"88180c8b",
         11908 => x"3d0d04f9",
         11909 => x"3d0d7984",
         11910 => x"11085656",
         11911 => x"807524a7",
         11912 => x"38893dfc",
         11913 => x"05547453",
         11914 => x"8c165275",
         11915 => x"0851c9dc",
         11916 => x"3f82e098",
         11917 => x"08913884",
         11918 => x"1608782e",
         11919 => x"09810687",
         11920 => x"38881608",
         11921 => x"558339ff",
         11922 => x"557482e0",
         11923 => x"980c893d",
         11924 => x"0d04fd3d",
         11925 => x"0d755480",
         11926 => x"cc538052",
         11927 => x"7351ff86",
         11928 => x"d53f7674",
         11929 => x"0c853d0d",
         11930 => x"04ea3d0d",
         11931 => x"0280e305",
         11932 => x"336a5386",
         11933 => x"3d705354",
         11934 => x"54d83f73",
         11935 => x"527251fe",
         11936 => x"ae3f7251",
         11937 => x"ff8d3f98",
         11938 => x"3d0d04fd",
         11939 => x"3d0d7502",
         11940 => x"84059a05",
         11941 => x"22555380",
         11942 => x"527280ff",
         11943 => x"268a3872",
         11944 => x"83ffff06",
         11945 => x"5280c339",
         11946 => x"83ffff73",
         11947 => x"27517383",
         11948 => x"b52e0981",
         11949 => x"06b43870",
         11950 => x"802eaf38",
         11951 => x"82d3ec22",
         11952 => x"5172712e",
         11953 => x"9c388112",
         11954 => x"7083ffff",
         11955 => x"06535171",
         11956 => x"80ff268d",
         11957 => x"38711082",
         11958 => x"d3ec0570",
         11959 => x"225151e1",
         11960 => x"39818012",
         11961 => x"7081ff06",
         11962 => x"53517182",
         11963 => x"e0980c85",
         11964 => x"3d0d04fe",
         11965 => x"3d0d0292",
         11966 => x"05220284",
         11967 => x"05960522",
         11968 => x"53518053",
         11969 => x"7080ff26",
         11970 => x"85387053",
         11971 => x"9a397183",
         11972 => x"b52e0981",
         11973 => x"06913870",
         11974 => x"81ff268b",
         11975 => x"38701082",
         11976 => x"d1ec0570",
         11977 => x"22545172",
         11978 => x"82e0980c",
         11979 => x"843d0d04",
         11980 => x"fb3d0d77",
         11981 => x"517083ff",
         11982 => x"ff2681a7",
         11983 => x"387083ff",
         11984 => x"ff0682d5",
         11985 => x"ec57529f",
         11986 => x"ff722785",
         11987 => x"3882d9e0",
         11988 => x"56757082",
         11989 => x"05572270",
         11990 => x"30708025",
         11991 => x"72752607",
         11992 => x"51525570",
         11993 => x"80fb3875",
         11994 => x"70820557",
         11995 => x"2270882a",
         11996 => x"7181ff06",
         11997 => x"70185452",
         11998 => x"55537171",
         11999 => x"2580d738",
         12000 => x"73882680",
         12001 => x"dc387384",
         12002 => x"2982b9b8",
         12003 => x"05517008",
         12004 => x"04717531",
         12005 => x"10761170",
         12006 => x"22545151",
         12007 => x"80c33971",
         12008 => x"75318106",
         12009 => x"72713151",
         12010 => x"51a439f0",
         12011 => x"12519f39",
         12012 => x"e012519a",
         12013 => x"39d01251",
         12014 => x"9539e612",
         12015 => x"51903988",
         12016 => x"12518b39",
         12017 => x"ffb01251",
         12018 => x"8539c7a0",
         12019 => x"12517083",
         12020 => x"ffff0652",
         12021 => x"8c3973fe",
         12022 => x"f8387210",
         12023 => x"1656fef1",
         12024 => x"39715170",
         12025 => x"82e0980c",
         12026 => x"873d0d04",
         12027 => x"00ffffff",
         12028 => x"ff00ffff",
         12029 => x"ffff00ff",
         12030 => x"ffffff00",
         12031 => x"00003101",
         12032 => x"00003085",
         12033 => x"0000308c",
         12034 => x"00003093",
         12035 => x"0000309a",
         12036 => x"000030a1",
         12037 => x"000030a8",
         12038 => x"000030af",
         12039 => x"000030b6",
         12040 => x"000030bd",
         12041 => x"000030c4",
         12042 => x"000030cb",
         12043 => x"000030d1",
         12044 => x"000030d7",
         12045 => x"000030dd",
         12046 => x"000030e3",
         12047 => x"000030e9",
         12048 => x"000030ef",
         12049 => x"000030f5",
         12050 => x"000030fb",
         12051 => x"00004781",
         12052 => x"00004787",
         12053 => x"0000478d",
         12054 => x"00004793",
         12055 => x"00004799",
         12056 => x"00004d79",
         12057 => x"00004e79",
         12058 => x"00004f8a",
         12059 => x"000051e2",
         12060 => x"00004e61",
         12061 => x"00004c4c",
         12062 => x"00005052",
         12063 => x"000051b3",
         12064 => x"00005095",
         12065 => x"0000512b",
         12066 => x"000050b1",
         12067 => x"00004f34",
         12068 => x"00004c4c",
         12069 => x"00004f8a",
         12070 => x"00004fb3",
         12071 => x"00005052",
         12072 => x"00004c4c",
         12073 => x"00004c4c",
         12074 => x"000050b1",
         12075 => x"0000512b",
         12076 => x"000051b3",
         12077 => x"000051e2",
         12078 => x"00009b91",
         12079 => x"00009b9f",
         12080 => x"00009bab",
         12081 => x"00009bb0",
         12082 => x"00009bb5",
         12083 => x"00009bba",
         12084 => x"00009bbf",
         12085 => x"00009bc4",
         12086 => x"00009bca",
         12087 => x"00000e65",
         12088 => x"0000174e",
         12089 => x"0000174e",
         12090 => x"00000e94",
         12091 => x"0000174e",
         12092 => x"0000174e",
         12093 => x"0000174e",
         12094 => x"0000174e",
         12095 => x"0000174e",
         12096 => x"0000174e",
         12097 => x"0000174e",
         12098 => x"00000e51",
         12099 => x"0000174e",
         12100 => x"00000e7c",
         12101 => x"00000eac",
         12102 => x"0000174e",
         12103 => x"0000174e",
         12104 => x"0000174e",
         12105 => x"0000174e",
         12106 => x"0000174e",
         12107 => x"0000174e",
         12108 => x"0000174e",
         12109 => x"0000174e",
         12110 => x"0000174e",
         12111 => x"0000174e",
         12112 => x"0000174e",
         12113 => x"0000174e",
         12114 => x"0000174e",
         12115 => x"0000174e",
         12116 => x"0000174e",
         12117 => x"0000174e",
         12118 => x"0000174e",
         12119 => x"0000174e",
         12120 => x"0000174e",
         12121 => x"0000174e",
         12122 => x"0000174e",
         12123 => x"0000174e",
         12124 => x"0000174e",
         12125 => x"0000174e",
         12126 => x"0000174e",
         12127 => x"0000174e",
         12128 => x"0000174e",
         12129 => x"0000174e",
         12130 => x"0000174e",
         12131 => x"0000174e",
         12132 => x"0000174e",
         12133 => x"0000174e",
         12134 => x"0000174e",
         12135 => x"0000174e",
         12136 => x"0000174e",
         12137 => x"0000174e",
         12138 => x"00000fdc",
         12139 => x"0000174e",
         12140 => x"0000174e",
         12141 => x"0000174e",
         12142 => x"0000174e",
         12143 => x"0000114a",
         12144 => x"0000174e",
         12145 => x"0000174e",
         12146 => x"0000174e",
         12147 => x"0000174e",
         12148 => x"0000174e",
         12149 => x"0000174e",
         12150 => x"0000174e",
         12151 => x"0000174e",
         12152 => x"0000174e",
         12153 => x"0000174e",
         12154 => x"00000f0c",
         12155 => x"00001073",
         12156 => x"00000ee3",
         12157 => x"00000ee3",
         12158 => x"00000ee3",
         12159 => x"0000174e",
         12160 => x"00001073",
         12161 => x"0000174e",
         12162 => x"0000174e",
         12163 => x"00000ecc",
         12164 => x"0000174e",
         12165 => x"0000174e",
         12166 => x"00001120",
         12167 => x"0000112b",
         12168 => x"0000174e",
         12169 => x"0000174e",
         12170 => x"00000f45",
         12171 => x"0000174e",
         12172 => x"00001153",
         12173 => x"0000174e",
         12174 => x"0000174e",
         12175 => x"0000114a",
         12176 => x"64696e69",
         12177 => x"74000000",
         12178 => x"64696f63",
         12179 => x"746c0000",
         12180 => x"66696e69",
         12181 => x"74000000",
         12182 => x"666c6f61",
         12183 => x"64000000",
         12184 => x"66657865",
         12185 => x"63000000",
         12186 => x"6d636c65",
         12187 => x"61720000",
         12188 => x"6d636f70",
         12189 => x"79000000",
         12190 => x"6d646966",
         12191 => x"66000000",
         12192 => x"6d64756d",
         12193 => x"70000000",
         12194 => x"6d656200",
         12195 => x"6d656800",
         12196 => x"6d657700",
         12197 => x"68696400",
         12198 => x"68696500",
         12199 => x"68666400",
         12200 => x"68666500",
         12201 => x"63616c6c",
         12202 => x"00000000",
         12203 => x"6a6d7000",
         12204 => x"72657374",
         12205 => x"61727400",
         12206 => x"72657365",
         12207 => x"74000000",
         12208 => x"696e666f",
         12209 => x"00000000",
         12210 => x"74626173",
         12211 => x"69630000",
         12212 => x"6d626173",
         12213 => x"69630000",
         12214 => x"6b696c6f",
         12215 => x"00000000",
         12216 => x"65640000",
         12217 => x"4469736b",
         12218 => x"20457272",
         12219 => x"6f720000",
         12220 => x"496e7465",
         12221 => x"726e616c",
         12222 => x"20657272",
         12223 => x"6f722e00",
         12224 => x"4469736b",
         12225 => x"206e6f74",
         12226 => x"20726561",
         12227 => x"64792e00",
         12228 => x"4e6f2066",
         12229 => x"696c6520",
         12230 => x"666f756e",
         12231 => x"642e0000",
         12232 => x"4e6f2070",
         12233 => x"61746820",
         12234 => x"666f756e",
         12235 => x"642e0000",
         12236 => x"496e7661",
         12237 => x"6c696420",
         12238 => x"66696c65",
         12239 => x"6e616d65",
         12240 => x"2e000000",
         12241 => x"41636365",
         12242 => x"73732064",
         12243 => x"656e6965",
         12244 => x"642e0000",
         12245 => x"46696c65",
         12246 => x"20616c72",
         12247 => x"65616479",
         12248 => x"20657869",
         12249 => x"7374732e",
         12250 => x"00000000",
         12251 => x"46696c65",
         12252 => x"2068616e",
         12253 => x"646c6520",
         12254 => x"696e7661",
         12255 => x"6c69642e",
         12256 => x"00000000",
         12257 => x"53442069",
         12258 => x"73207772",
         12259 => x"69746520",
         12260 => x"70726f74",
         12261 => x"65637465",
         12262 => x"642e0000",
         12263 => x"44726976",
         12264 => x"65206e75",
         12265 => x"6d626572",
         12266 => x"20697320",
         12267 => x"696e7661",
         12268 => x"6c69642e",
         12269 => x"00000000",
         12270 => x"4469736b",
         12271 => x"206e6f74",
         12272 => x"20656e61",
         12273 => x"626c6564",
         12274 => x"2e000000",
         12275 => x"4e6f2063",
         12276 => x"6f6d7061",
         12277 => x"7469626c",
         12278 => x"65206669",
         12279 => x"6c657379",
         12280 => x"7374656d",
         12281 => x"20666f75",
         12282 => x"6e64206f",
         12283 => x"6e206469",
         12284 => x"736b2e00",
         12285 => x"466f726d",
         12286 => x"61742061",
         12287 => x"626f7274",
         12288 => x"65642e00",
         12289 => x"54696d65",
         12290 => x"6f75742c",
         12291 => x"206f7065",
         12292 => x"72617469",
         12293 => x"6f6e2063",
         12294 => x"616e6365",
         12295 => x"6c6c6564",
         12296 => x"2e000000",
         12297 => x"46696c65",
         12298 => x"20697320",
         12299 => x"6c6f636b",
         12300 => x"65642e00",
         12301 => x"496e7375",
         12302 => x"66666963",
         12303 => x"69656e74",
         12304 => x"206d656d",
         12305 => x"6f72792e",
         12306 => x"00000000",
         12307 => x"546f6f20",
         12308 => x"6d616e79",
         12309 => x"206f7065",
         12310 => x"6e206669",
         12311 => x"6c65732e",
         12312 => x"00000000",
         12313 => x"50617261",
         12314 => x"6d657465",
         12315 => x"72732069",
         12316 => x"6e636f72",
         12317 => x"72656374",
         12318 => x"2e000000",
         12319 => x"53756363",
         12320 => x"6573732e",
         12321 => x"00000000",
         12322 => x"556e6b6e",
         12323 => x"6f776e20",
         12324 => x"6572726f",
         12325 => x"722e0000",
         12326 => x"0a256c75",
         12327 => x"20627974",
         12328 => x"65732025",
         12329 => x"73206174",
         12330 => x"20256c75",
         12331 => x"20627974",
         12332 => x"65732f73",
         12333 => x"65632e0a",
         12334 => x"00000000",
         12335 => x"72656164",
         12336 => x"00000000",
         12337 => x"2530386c",
         12338 => x"58000000",
         12339 => x"3a202000",
         12340 => x"25303458",
         12341 => x"00000000",
         12342 => x"20202020",
         12343 => x"20202020",
         12344 => x"00000000",
         12345 => x"25303258",
         12346 => x"00000000",
         12347 => x"20200000",
         12348 => x"207c0000",
         12349 => x"7c000000",
         12350 => x"7a4f5300",
         12351 => x"2a2a2025",
         12352 => x"73202800",
         12353 => x"31312f31",
         12354 => x"322f3230",
         12355 => x"32300000",
         12356 => x"76312e31",
         12357 => x"63000000",
         12358 => x"205a5055",
         12359 => x"2c207265",
         12360 => x"76202530",
         12361 => x"32782920",
         12362 => x"25732025",
         12363 => x"73202a2a",
         12364 => x"0a0a0000",
         12365 => x"5a505520",
         12366 => x"496e7465",
         12367 => x"72727570",
         12368 => x"74204861",
         12369 => x"6e646c65",
         12370 => x"72000000",
         12371 => x"54696d65",
         12372 => x"7220696e",
         12373 => x"74657272",
         12374 => x"75707400",
         12375 => x"50533220",
         12376 => x"696e7465",
         12377 => x"72727570",
         12378 => x"74000000",
         12379 => x"494f4354",
         12380 => x"4c205244",
         12381 => x"20696e74",
         12382 => x"65727275",
         12383 => x"70740000",
         12384 => x"494f4354",
         12385 => x"4c205752",
         12386 => x"20696e74",
         12387 => x"65727275",
         12388 => x"70740000",
         12389 => x"55415254",
         12390 => x"30205258",
         12391 => x"20696e74",
         12392 => x"65727275",
         12393 => x"70740000",
         12394 => x"55415254",
         12395 => x"30205458",
         12396 => x"20696e74",
         12397 => x"65727275",
         12398 => x"70740000",
         12399 => x"55415254",
         12400 => x"31205258",
         12401 => x"20696e74",
         12402 => x"65727275",
         12403 => x"70740000",
         12404 => x"55415254",
         12405 => x"31205458",
         12406 => x"20696e74",
         12407 => x"65727275",
         12408 => x"70740000",
         12409 => x"53657474",
         12410 => x"696e6720",
         12411 => x"75702074",
         12412 => x"696d6572",
         12413 => x"2e2e2e00",
         12414 => x"456e6162",
         12415 => x"6c696e67",
         12416 => x"2074696d",
         12417 => x"65722e2e",
         12418 => x"2e000000",
         12419 => x"6175746f",
         12420 => x"65786563",
         12421 => x"2e626174",
         12422 => x"00000000",
         12423 => x"7a4f535f",
         12424 => x"7a70752e",
         12425 => x"68737400",
         12426 => x"303a0000",
         12427 => x"4661696c",
         12428 => x"65642074",
         12429 => x"6f20696e",
         12430 => x"69746961",
         12431 => x"6c697365",
         12432 => x"20736420",
         12433 => x"63617264",
         12434 => x"20302c20",
         12435 => x"706c6561",
         12436 => x"73652069",
         12437 => x"6e697420",
         12438 => x"6d616e75",
         12439 => x"616c6c79",
         12440 => x"2e000000",
         12441 => x"2a200000",
         12442 => x"436c6561",
         12443 => x"72696e67",
         12444 => x"2e2e2e2e",
         12445 => x"00000000",
         12446 => x"436f7079",
         12447 => x"696e672e",
         12448 => x"2e2e0000",
         12449 => x"436f6d70",
         12450 => x"6172696e",
         12451 => x"672e2e2e",
         12452 => x"00000000",
         12453 => x"2530386c",
         12454 => x"78282530",
         12455 => x"3878292d",
         12456 => x"3e253038",
         12457 => x"6c782825",
         12458 => x"30387829",
         12459 => x"0a000000",
         12460 => x"44756d70",
         12461 => x"204d656d",
         12462 => x"6f727900",
         12463 => x"0a436f6d",
         12464 => x"706c6574",
         12465 => x"652e0000",
         12466 => x"2530386c",
         12467 => x"58202530",
         12468 => x"32582d00",
         12469 => x"3f3f3f00",
         12470 => x"2530386c",
         12471 => x"58202530",
         12472 => x"34582d00",
         12473 => x"2530386c",
         12474 => x"58202530",
         12475 => x"386c582d",
         12476 => x"00000000",
         12477 => x"45786563",
         12478 => x"7574696e",
         12479 => x"6720636f",
         12480 => x"64652040",
         12481 => x"20253038",
         12482 => x"6c78202e",
         12483 => x"2e2e0a00",
         12484 => x"43616c6c",
         12485 => x"696e6720",
         12486 => x"636f6465",
         12487 => x"20402025",
         12488 => x"30386c78",
         12489 => x"202e2e2e",
         12490 => x"0a000000",
         12491 => x"43616c6c",
         12492 => x"20726574",
         12493 => x"75726e65",
         12494 => x"6420636f",
         12495 => x"64652028",
         12496 => x"2564292e",
         12497 => x"0a000000",
         12498 => x"52657374",
         12499 => x"61727469",
         12500 => x"6e672061",
         12501 => x"70706c69",
         12502 => x"63617469",
         12503 => x"6f6e2e2e",
         12504 => x"2e000000",
         12505 => x"436f6c64",
         12506 => x"20726562",
         12507 => x"6f6f7469",
         12508 => x"6e672e2e",
         12509 => x"2e000000",
         12510 => x"5a505500",
         12511 => x"62696e00",
         12512 => x"25643a5c",
         12513 => x"25735c25",
         12514 => x"732e2573",
         12515 => x"00000000",
         12516 => x"25643a5c",
         12517 => x"25735c25",
         12518 => x"73000000",
         12519 => x"25643a5c",
         12520 => x"25730000",
         12521 => x"42616420",
         12522 => x"636f6d6d",
         12523 => x"616e642e",
         12524 => x"00000000",
         12525 => x"4d656d6f",
         12526 => x"72792065",
         12527 => x"78686175",
         12528 => x"73746564",
         12529 => x"2c206361",
         12530 => x"6e6e6f74",
         12531 => x"2070726f",
         12532 => x"63657373",
         12533 => x"20636f6d",
         12534 => x"6d616e64",
         12535 => x"2e000000",
         12536 => x"52756e6e",
         12537 => x"696e672e",
         12538 => x"2e2e0000",
         12539 => x"456e6162",
         12540 => x"6c696e67",
         12541 => x"20696e74",
         12542 => x"65727275",
         12543 => x"7074732e",
         12544 => x"2e2e0000",
         12545 => x"25642f25",
         12546 => x"642f2564",
         12547 => x"2025643a",
         12548 => x"25643a25",
         12549 => x"642e2564",
         12550 => x"25640a00",
         12551 => x"536f4320",
         12552 => x"436f6e66",
         12553 => x"69677572",
         12554 => x"6174696f",
         12555 => x"6e000000",
         12556 => x"20286672",
         12557 => x"6f6d2053",
         12558 => x"6f432063",
         12559 => x"6f6e6669",
         12560 => x"67290000",
         12561 => x"3a0a4465",
         12562 => x"76696365",
         12563 => x"7320696d",
         12564 => x"706c656d",
         12565 => x"656e7465",
         12566 => x"643a0000",
         12567 => x"20202020",
         12568 => x"57422053",
         12569 => x"4452414d",
         12570 => x"20202825",
         12571 => x"3038583a",
         12572 => x"25303858",
         12573 => x"292e0a00",
         12574 => x"20202020",
         12575 => x"53445241",
         12576 => x"4d202020",
         12577 => x"20202825",
         12578 => x"3038583a",
         12579 => x"25303858",
         12580 => x"292e0a00",
         12581 => x"20202020",
         12582 => x"494e534e",
         12583 => x"20425241",
         12584 => x"4d202825",
         12585 => x"3038583a",
         12586 => x"25303858",
         12587 => x"292e0a00",
         12588 => x"20202020",
         12589 => x"4252414d",
         12590 => x"20202020",
         12591 => x"20202825",
         12592 => x"3038583a",
         12593 => x"25303858",
         12594 => x"292e0a00",
         12595 => x"20202020",
         12596 => x"52414d20",
         12597 => x"20202020",
         12598 => x"20202825",
         12599 => x"3038583a",
         12600 => x"25303858",
         12601 => x"292e0a00",
         12602 => x"20202020",
         12603 => x"53442043",
         12604 => x"41524420",
         12605 => x"20202844",
         12606 => x"65766963",
         12607 => x"6573203d",
         12608 => x"25303264",
         12609 => x"292e0a00",
         12610 => x"20202020",
         12611 => x"54494d45",
         12612 => x"52312020",
         12613 => x"20202854",
         12614 => x"696d6572",
         12615 => x"7320203d",
         12616 => x"25303264",
         12617 => x"292e0a00",
         12618 => x"20202020",
         12619 => x"494e5452",
         12620 => x"20435452",
         12621 => x"4c202843",
         12622 => x"68616e6e",
         12623 => x"656c733d",
         12624 => x"25303264",
         12625 => x"292e0a00",
         12626 => x"20202020",
         12627 => x"57495348",
         12628 => x"424f4e45",
         12629 => x"20425553",
         12630 => x"00000000",
         12631 => x"20202020",
         12632 => x"57422049",
         12633 => x"32430000",
         12634 => x"20202020",
         12635 => x"494f4354",
         12636 => x"4c000000",
         12637 => x"20202020",
         12638 => x"50533200",
         12639 => x"20202020",
         12640 => x"53504900",
         12641 => x"41646472",
         12642 => x"65737365",
         12643 => x"733a0000",
         12644 => x"20202020",
         12645 => x"43505520",
         12646 => x"52657365",
         12647 => x"74205665",
         12648 => x"63746f72",
         12649 => x"20416464",
         12650 => x"72657373",
         12651 => x"203d2025",
         12652 => x"3038580a",
         12653 => x"00000000",
         12654 => x"20202020",
         12655 => x"43505520",
         12656 => x"4d656d6f",
         12657 => x"72792053",
         12658 => x"74617274",
         12659 => x"20416464",
         12660 => x"72657373",
         12661 => x"203d2025",
         12662 => x"3038580a",
         12663 => x"00000000",
         12664 => x"20202020",
         12665 => x"53746163",
         12666 => x"6b205374",
         12667 => x"61727420",
         12668 => x"41646472",
         12669 => x"65737320",
         12670 => x"20202020",
         12671 => x"203d2025",
         12672 => x"3038580a",
         12673 => x"00000000",
         12674 => x"4d697363",
         12675 => x"3a000000",
         12676 => x"20202020",
         12677 => x"5a505520",
         12678 => x"49642020",
         12679 => x"20202020",
         12680 => x"20202020",
         12681 => x"20202020",
         12682 => x"20202020",
         12683 => x"203d2025",
         12684 => x"3034580a",
         12685 => x"00000000",
         12686 => x"20202020",
         12687 => x"53797374",
         12688 => x"656d2043",
         12689 => x"6c6f636b",
         12690 => x"20467265",
         12691 => x"71202020",
         12692 => x"20202020",
         12693 => x"203d2025",
         12694 => x"642e2530",
         12695 => x"34644d48",
         12696 => x"7a0a0000",
         12697 => x"20202020",
         12698 => x"53445241",
         12699 => x"4d20436c",
         12700 => x"6f636b20",
         12701 => x"46726571",
         12702 => x"20202020",
         12703 => x"20202020",
         12704 => x"203d2025",
         12705 => x"642e2530",
         12706 => x"34644d48",
         12707 => x"7a0a0000",
         12708 => x"20202020",
         12709 => x"57697368",
         12710 => x"626f6e65",
         12711 => x"20534452",
         12712 => x"414d2043",
         12713 => x"6c6f636b",
         12714 => x"20467265",
         12715 => x"713d2025",
         12716 => x"642e2530",
         12717 => x"34644d48",
         12718 => x"7a0a0000",
         12719 => x"536d616c",
         12720 => x"6c000000",
         12721 => x"4d656469",
         12722 => x"756d0000",
         12723 => x"466c6578",
         12724 => x"00000000",
         12725 => x"45564f00",
         12726 => x"45564f6d",
         12727 => x"00000000",
         12728 => x"556e6b6e",
         12729 => x"6f776e00",
         12730 => x"0000a844",
         12731 => x"01000000",
         12732 => x"00000002",
         12733 => x"0000a840",
         12734 => x"01000000",
         12735 => x"00000003",
         12736 => x"0000a83c",
         12737 => x"01000000",
         12738 => x"00000004",
         12739 => x"0000a838",
         12740 => x"01000000",
         12741 => x"00000005",
         12742 => x"0000a834",
         12743 => x"01000000",
         12744 => x"00000006",
         12745 => x"0000a830",
         12746 => x"01000000",
         12747 => x"00000007",
         12748 => x"0000a82c",
         12749 => x"01000000",
         12750 => x"00000001",
         12751 => x"0000a828",
         12752 => x"01000000",
         12753 => x"00000008",
         12754 => x"0000a824",
         12755 => x"01000000",
         12756 => x"0000000b",
         12757 => x"0000a820",
         12758 => x"01000000",
         12759 => x"00000009",
         12760 => x"0000a81c",
         12761 => x"01000000",
         12762 => x"0000000a",
         12763 => x"0000a818",
         12764 => x"04000000",
         12765 => x"0000000d",
         12766 => x"0000a814",
         12767 => x"04000000",
         12768 => x"0000000c",
         12769 => x"0000a810",
         12770 => x"04000000",
         12771 => x"0000000e",
         12772 => x"0000a80c",
         12773 => x"03000000",
         12774 => x"0000000f",
         12775 => x"0000a808",
         12776 => x"04000000",
         12777 => x"0000000f",
         12778 => x"0000a804",
         12779 => x"04000000",
         12780 => x"00000010",
         12781 => x"0000a800",
         12782 => x"04000000",
         12783 => x"00000011",
         12784 => x"0000a7fc",
         12785 => x"03000000",
         12786 => x"00000012",
         12787 => x"0000a7f8",
         12788 => x"03000000",
         12789 => x"00000013",
         12790 => x"0000a7f4",
         12791 => x"03000000",
         12792 => x"00000014",
         12793 => x"0000a7f0",
         12794 => x"03000000",
         12795 => x"00000015",
         12796 => x"1b5b4400",
         12797 => x"1b5b4300",
         12798 => x"1b5b4200",
         12799 => x"1b5b4100",
         12800 => x"1b5b367e",
         12801 => x"1b5b357e",
         12802 => x"1b5b347e",
         12803 => x"1b304600",
         12804 => x"1b5b337e",
         12805 => x"1b5b327e",
         12806 => x"1b5b317e",
         12807 => x"10000000",
         12808 => x"0e000000",
         12809 => x"0d000000",
         12810 => x"0b000000",
         12811 => x"08000000",
         12812 => x"06000000",
         12813 => x"05000000",
         12814 => x"04000000",
         12815 => x"03000000",
         12816 => x"02000000",
         12817 => x"01000000",
         12818 => x"68697374",
         12819 => x"6f727900",
         12820 => x"68697374",
         12821 => x"00000000",
         12822 => x"21000000",
         12823 => x"2530346c",
         12824 => x"75202025",
         12825 => x"730a0000",
         12826 => x"4661696c",
         12827 => x"65642074",
         12828 => x"6f207265",
         12829 => x"73657420",
         12830 => x"74686520",
         12831 => x"68697374",
         12832 => x"6f727920",
         12833 => x"66696c65",
         12834 => x"20746f20",
         12835 => x"454f462e",
         12836 => x"00000000",
         12837 => x"43616e6e",
         12838 => x"6f74206f",
         12839 => x"70656e2f",
         12840 => x"63726561",
         12841 => x"74652068",
         12842 => x"6973746f",
         12843 => x"72792066",
         12844 => x"696c652c",
         12845 => x"20646973",
         12846 => x"61626c69",
         12847 => x"6e672e00",
         12848 => x"53440000",
         12849 => x"222a3a3c",
         12850 => x"3e3f7c7f",
         12851 => x"00000000",
         12852 => x"2b2c3b3d",
         12853 => x"5b5d0000",
         12854 => x"46415400",
         12855 => x"46415433",
         12856 => x"32000000",
         12857 => x"ebfe904d",
         12858 => x"53444f53",
         12859 => x"352e3000",
         12860 => x"4e4f204e",
         12861 => x"414d4520",
         12862 => x"20202046",
         12863 => x"41543332",
         12864 => x"20202000",
         12865 => x"4e4f204e",
         12866 => x"414d4520",
         12867 => x"20202046",
         12868 => x"41542020",
         12869 => x"20202000",
         12870 => x"0000a8c0",
         12871 => x"00000000",
         12872 => x"00000000",
         12873 => x"00000000",
         12874 => x"01030507",
         12875 => x"090e1012",
         12876 => x"1416181c",
         12877 => x"1e000000",
         12878 => x"809a4541",
         12879 => x"8e418f80",
         12880 => x"45454549",
         12881 => x"49498e8f",
         12882 => x"9092924f",
         12883 => x"994f5555",
         12884 => x"59999a9b",
         12885 => x"9c9d9e9f",
         12886 => x"41494f55",
         12887 => x"a5a5a6a7",
         12888 => x"a8a9aaab",
         12889 => x"acadaeaf",
         12890 => x"b0b1b2b3",
         12891 => x"b4b5b6b7",
         12892 => x"b8b9babb",
         12893 => x"bcbdbebf",
         12894 => x"c0c1c2c3",
         12895 => x"c4c5c6c7",
         12896 => x"c8c9cacb",
         12897 => x"cccdcecf",
         12898 => x"d0d1d2d3",
         12899 => x"d4d5d6d7",
         12900 => x"d8d9dadb",
         12901 => x"dcdddedf",
         12902 => x"e0e1e2e3",
         12903 => x"e4e5e6e7",
         12904 => x"e8e9eaeb",
         12905 => x"ecedeeef",
         12906 => x"f0f1f2f3",
         12907 => x"f4f5f6f7",
         12908 => x"f8f9fafb",
         12909 => x"fcfdfeff",
         12910 => x"2b2e2c3b",
         12911 => x"3d5b5d2f",
         12912 => x"5c222a3a",
         12913 => x"3c3e3f7c",
         12914 => x"7f000000",
         12915 => x"00010004",
         12916 => x"00100040",
         12917 => x"01000200",
         12918 => x"00000000",
         12919 => x"00010002",
         12920 => x"00040008",
         12921 => x"00100020",
         12922 => x"00000000",
         12923 => x"00c700fc",
         12924 => x"00e900e2",
         12925 => x"00e400e0",
         12926 => x"00e500e7",
         12927 => x"00ea00eb",
         12928 => x"00e800ef",
         12929 => x"00ee00ec",
         12930 => x"00c400c5",
         12931 => x"00c900e6",
         12932 => x"00c600f4",
         12933 => x"00f600f2",
         12934 => x"00fb00f9",
         12935 => x"00ff00d6",
         12936 => x"00dc00a2",
         12937 => x"00a300a5",
         12938 => x"20a70192",
         12939 => x"00e100ed",
         12940 => x"00f300fa",
         12941 => x"00f100d1",
         12942 => x"00aa00ba",
         12943 => x"00bf2310",
         12944 => x"00ac00bd",
         12945 => x"00bc00a1",
         12946 => x"00ab00bb",
         12947 => x"25912592",
         12948 => x"25932502",
         12949 => x"25242561",
         12950 => x"25622556",
         12951 => x"25552563",
         12952 => x"25512557",
         12953 => x"255d255c",
         12954 => x"255b2510",
         12955 => x"25142534",
         12956 => x"252c251c",
         12957 => x"2500253c",
         12958 => x"255e255f",
         12959 => x"255a2554",
         12960 => x"25692566",
         12961 => x"25602550",
         12962 => x"256c2567",
         12963 => x"25682564",
         12964 => x"25652559",
         12965 => x"25582552",
         12966 => x"2553256b",
         12967 => x"256a2518",
         12968 => x"250c2588",
         12969 => x"2584258c",
         12970 => x"25902580",
         12971 => x"03b100df",
         12972 => x"039303c0",
         12973 => x"03a303c3",
         12974 => x"00b503c4",
         12975 => x"03a60398",
         12976 => x"03a903b4",
         12977 => x"221e03c6",
         12978 => x"03b52229",
         12979 => x"226100b1",
         12980 => x"22652264",
         12981 => x"23202321",
         12982 => x"00f72248",
         12983 => x"00b02219",
         12984 => x"00b7221a",
         12985 => x"207f00b2",
         12986 => x"25a000a0",
         12987 => x"0061031a",
         12988 => x"00e00317",
         12989 => x"00f80307",
         12990 => x"00ff0001",
         12991 => x"01780100",
         12992 => x"01300132",
         12993 => x"01060139",
         12994 => x"0110014a",
         12995 => x"012e0179",
         12996 => x"01060180",
         12997 => x"004d0243",
         12998 => x"01810182",
         12999 => x"01820184",
         13000 => x"01840186",
         13001 => x"01870187",
         13002 => x"0189018a",
         13003 => x"018b018b",
         13004 => x"018d018e",
         13005 => x"018f0190",
         13006 => x"01910191",
         13007 => x"01930194",
         13008 => x"01f60196",
         13009 => x"01970198",
         13010 => x"0198023d",
         13011 => x"019b019c",
         13012 => x"019d0220",
         13013 => x"019f01a0",
         13014 => x"01a001a2",
         13015 => x"01a201a4",
         13016 => x"01a401a6",
         13017 => x"01a701a7",
         13018 => x"01a901aa",
         13019 => x"01ab01ac",
         13020 => x"01ac01ae",
         13021 => x"01af01af",
         13022 => x"01b101b2",
         13023 => x"01b301b3",
         13024 => x"01b501b5",
         13025 => x"01b701b8",
         13026 => x"01b801ba",
         13027 => x"01bb01bc",
         13028 => x"01bc01be",
         13029 => x"01f701c0",
         13030 => x"01c101c2",
         13031 => x"01c301c4",
         13032 => x"01c501c4",
         13033 => x"01c701c8",
         13034 => x"01c701ca",
         13035 => x"01cb01ca",
         13036 => x"01cd0110",
         13037 => x"01dd0001",
         13038 => x"018e01de",
         13039 => x"011201f3",
         13040 => x"000301f1",
         13041 => x"01f401f4",
         13042 => x"01f80128",
         13043 => x"02220112",
         13044 => x"023a0009",
         13045 => x"2c65023b",
         13046 => x"023b023d",
         13047 => x"2c66023f",
         13048 => x"02400241",
         13049 => x"02410246",
         13050 => x"010a0253",
         13051 => x"00400181",
         13052 => x"01860255",
         13053 => x"0189018a",
         13054 => x"0258018f",
         13055 => x"025a0190",
         13056 => x"025c025d",
         13057 => x"025e025f",
         13058 => x"01930261",
         13059 => x"02620194",
         13060 => x"02640265",
         13061 => x"02660267",
         13062 => x"01970196",
         13063 => x"026a2c62",
         13064 => x"026c026d",
         13065 => x"026e019c",
         13066 => x"02700271",
         13067 => x"019d0273",
         13068 => x"0274019f",
         13069 => x"02760277",
         13070 => x"02780279",
         13071 => x"027a027b",
         13072 => x"027c2c64",
         13073 => x"027e027f",
         13074 => x"01a60281",
         13075 => x"028201a9",
         13076 => x"02840285",
         13077 => x"02860287",
         13078 => x"01ae0244",
         13079 => x"01b101b2",
         13080 => x"0245028d",
         13081 => x"028e028f",
         13082 => x"02900291",
         13083 => x"01b7037b",
         13084 => x"000303fd",
         13085 => x"03fe03ff",
         13086 => x"03ac0004",
         13087 => x"03860388",
         13088 => x"0389038a",
         13089 => x"03b10311",
         13090 => x"03c20002",
         13091 => x"03a303a3",
         13092 => x"03c40308",
         13093 => x"03cc0003",
         13094 => x"038c038e",
         13095 => x"038f03d8",
         13096 => x"011803f2",
         13097 => x"000a03f9",
         13098 => x"03f303f4",
         13099 => x"03f503f6",
         13100 => x"03f703f7",
         13101 => x"03f903fa",
         13102 => x"03fa0430",
         13103 => x"03200450",
         13104 => x"07100460",
         13105 => x"0122048a",
         13106 => x"013604c1",
         13107 => x"010e04cf",
         13108 => x"000104c0",
         13109 => x"04d00144",
         13110 => x"05610426",
         13111 => x"00000000",
         13112 => x"1d7d0001",
         13113 => x"2c631e00",
         13114 => x"01961ea0",
         13115 => x"015a1f00",
         13116 => x"06081f10",
         13117 => x"06061f20",
         13118 => x"06081f30",
         13119 => x"06081f40",
         13120 => x"06061f51",
         13121 => x"00071f59",
         13122 => x"1f521f5b",
         13123 => x"1f541f5d",
         13124 => x"1f561f5f",
         13125 => x"1f600608",
         13126 => x"1f70000e",
         13127 => x"1fba1fbb",
         13128 => x"1fc81fc9",
         13129 => x"1fca1fcb",
         13130 => x"1fda1fdb",
         13131 => x"1ff81ff9",
         13132 => x"1fea1feb",
         13133 => x"1ffa1ffb",
         13134 => x"1f800608",
         13135 => x"1f900608",
         13136 => x"1fa00608",
         13137 => x"1fb00004",
         13138 => x"1fb81fb9",
         13139 => x"1fb21fbc",
         13140 => x"1fcc0001",
         13141 => x"1fc31fd0",
         13142 => x"06021fe0",
         13143 => x"06021fe5",
         13144 => x"00011fec",
         13145 => x"1ff30001",
         13146 => x"1ffc214e",
         13147 => x"00012132",
         13148 => x"21700210",
         13149 => x"21840001",
         13150 => x"218324d0",
         13151 => x"051a2c30",
         13152 => x"042f2c60",
         13153 => x"01022c67",
         13154 => x"01062c75",
         13155 => x"01022c80",
         13156 => x"01642d00",
         13157 => x"0826ff41",
         13158 => x"031a0000",
         13159 => x"00000000",
         13160 => x"00009e40",
         13161 => x"01020100",
         13162 => x"00000000",
         13163 => x"00000000",
         13164 => x"00009e48",
         13165 => x"01040100",
         13166 => x"00000000",
         13167 => x"00000000",
         13168 => x"00009e50",
         13169 => x"01140300",
         13170 => x"00000000",
         13171 => x"00000000",
         13172 => x"00009e58",
         13173 => x"012b0300",
         13174 => x"00000000",
         13175 => x"00000000",
         13176 => x"00009e60",
         13177 => x"01300300",
         13178 => x"00000000",
         13179 => x"00000000",
         13180 => x"00009e68",
         13181 => x"013c0400",
         13182 => x"00000000",
         13183 => x"00000000",
         13184 => x"00009e70",
         13185 => x"013d0400",
         13186 => x"00000000",
         13187 => x"00000000",
         13188 => x"00009e78",
         13189 => x"013f0400",
         13190 => x"00000000",
         13191 => x"00000000",
         13192 => x"00009e80",
         13193 => x"01400400",
         13194 => x"00000000",
         13195 => x"00000000",
         13196 => x"00009e88",
         13197 => x"01410400",
         13198 => x"00000000",
         13199 => x"00000000",
         13200 => x"00009e8c",
         13201 => x"01420400",
         13202 => x"00000000",
         13203 => x"00000000",
         13204 => x"00009e90",
         13205 => x"01430400",
         13206 => x"00000000",
         13207 => x"00000000",
         13208 => x"00009e94",
         13209 => x"01500500",
         13210 => x"00000000",
         13211 => x"00000000",
         13212 => x"00009e98",
         13213 => x"01510500",
         13214 => x"00000000",
         13215 => x"00000000",
         13216 => x"00009e9c",
         13217 => x"01540500",
         13218 => x"00000000",
         13219 => x"00000000",
         13220 => x"00009ea0",
         13221 => x"01550500",
         13222 => x"00000000",
         13223 => x"00000000",
         13224 => x"00009ea4",
         13225 => x"01790700",
         13226 => x"00000000",
         13227 => x"00000000",
         13228 => x"00009eac",
         13229 => x"01780700",
         13230 => x"00000000",
         13231 => x"00000000",
         13232 => x"00009eb0",
         13233 => x"01820800",
         13234 => x"00000000",
         13235 => x"00000000",
         13236 => x"00009eb8",
         13237 => x"01830800",
         13238 => x"00000000",
         13239 => x"00000000",
         13240 => x"00009ec0",
         13241 => x"01850800",
         13242 => x"00000000",
         13243 => x"00000000",
         13244 => x"00009ec8",
         13245 => x"018c0900",
         13246 => x"00000000",
         13247 => x"00000000",
         13248 => x"00009ed0",
         13249 => x"018d0900",
         13250 => x"00000000",
         13251 => x"00000000",
         13252 => x"00009ed8",
         13253 => x"018e0900",
         13254 => x"00000000",
         13255 => x"00000000",
         13256 => x"00009ee0",
         13257 => x"018f0900",
         13258 => x"00000000",
         13259 => x"00000000",
         13260 => x"00000000",
         13261 => x"00000000",
         13262 => x"00007fff",
         13263 => x"00000000",
         13264 => x"00007fff",
         13265 => x"00010000",
         13266 => x"00007fff",
         13267 => x"00010000",
         13268 => x"00810000",
         13269 => x"01000000",
         13270 => x"017fffff",
         13271 => x"00000000",
         13272 => x"00000000",
         13273 => x"00007800",
         13274 => x"00000000",
         13275 => x"05f5e100",
         13276 => x"05f5e100",
         13277 => x"05f5e100",
         13278 => x"00000000",
         13279 => x"01010101",
         13280 => x"01010101",
         13281 => x"01011001",
         13282 => x"01000000",
         13283 => x"00000000",
         13284 => x"00000000",
         13285 => x"00000000",
         13286 => x"00000000",
         13287 => x"00000000",
         13288 => x"00000000",
         13289 => x"00000000",
         13290 => x"00000000",
         13291 => x"00000000",
         13292 => x"00000000",
         13293 => x"00000000",
         13294 => x"00000000",
         13295 => x"00000000",
         13296 => x"00000000",
         13297 => x"00000000",
         13298 => x"00000000",
         13299 => x"00000000",
         13300 => x"00000000",
         13301 => x"00000000",
         13302 => x"00000000",
         13303 => x"00000000",
         13304 => x"00000000",
         13305 => x"00000000",
         13306 => x"00000000",
         13307 => x"0000a848",
         13308 => x"01000000",
         13309 => x"0000a850",
         13310 => x"01000000",
         13311 => x"0000a858",
         13312 => x"02000000",
         13313 => x"00000000",
         13314 => x"00000000",
         13315 => x"00010002",
         13316 => x"00030004",
         13317 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

